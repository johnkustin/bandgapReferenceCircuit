magic
tech sky130A
magscale 1 2
timestamp 1620340193
<< nwell >>
rect -2813 -4398 2813 4364
<< pmoslvt >>
rect -2719 -4336 -2319 4264
rect -2261 -4336 -1861 4264
rect -1803 -4336 -1403 4264
rect -1345 -4336 -945 4264
rect -887 -4336 -487 4264
rect -429 -4336 -29 4264
rect 29 -4336 429 4264
rect 487 -4336 887 4264
rect 945 -4336 1345 4264
rect 1403 -4336 1803 4264
rect 1861 -4336 2261 4264
rect 2319 -4336 2719 4264
<< pdiff >>
rect -2777 4252 -2719 4264
rect -2777 -4324 -2765 4252
rect -2731 -4324 -2719 4252
rect -2777 -4336 -2719 -4324
rect -2319 4252 -2261 4264
rect -2319 -4324 -2307 4252
rect -2273 -4324 -2261 4252
rect -2319 -4336 -2261 -4324
rect -1861 4252 -1803 4264
rect -1861 -4324 -1849 4252
rect -1815 -4324 -1803 4252
rect -1861 -4336 -1803 -4324
rect -1403 4252 -1345 4264
rect -1403 -4324 -1391 4252
rect -1357 -4324 -1345 4252
rect -1403 -4336 -1345 -4324
rect -945 4252 -887 4264
rect -945 -4324 -933 4252
rect -899 -4324 -887 4252
rect -945 -4336 -887 -4324
rect -487 4252 -429 4264
rect -487 -4324 -475 4252
rect -441 -4324 -429 4252
rect -487 -4336 -429 -4324
rect -29 4252 29 4264
rect -29 -4324 -17 4252
rect 17 -4324 29 4252
rect -29 -4336 29 -4324
rect 429 4252 487 4264
rect 429 -4324 441 4252
rect 475 -4324 487 4252
rect 429 -4336 487 -4324
rect 887 4252 945 4264
rect 887 -4324 899 4252
rect 933 -4324 945 4252
rect 887 -4336 945 -4324
rect 1345 4252 1403 4264
rect 1345 -4324 1357 4252
rect 1391 -4324 1403 4252
rect 1345 -4336 1403 -4324
rect 1803 4252 1861 4264
rect 1803 -4324 1815 4252
rect 1849 -4324 1861 4252
rect 1803 -4336 1861 -4324
rect 2261 4252 2319 4264
rect 2261 -4324 2273 4252
rect 2307 -4324 2319 4252
rect 2261 -4336 2319 -4324
rect 2719 4252 2777 4264
rect 2719 -4324 2731 4252
rect 2765 -4324 2777 4252
rect 2719 -4336 2777 -4324
<< pdiffc >>
rect -2765 -4324 -2731 4252
rect -2307 -4324 -2273 4252
rect -1849 -4324 -1815 4252
rect -1391 -4324 -1357 4252
rect -933 -4324 -899 4252
rect -475 -4324 -441 4252
rect -17 -4324 17 4252
rect 441 -4324 475 4252
rect 899 -4324 933 4252
rect 1357 -4324 1391 4252
rect 1815 -4324 1849 4252
rect 2273 -4324 2307 4252
rect 2731 -4324 2765 4252
<< poly >>
rect -2719 4345 -2319 4361
rect -2719 4311 -2703 4345
rect -2335 4311 -2319 4345
rect -2719 4264 -2319 4311
rect -2261 4345 -1861 4361
rect -2261 4311 -2245 4345
rect -1877 4311 -1861 4345
rect -2261 4264 -1861 4311
rect -1803 4345 -1403 4361
rect -1803 4311 -1787 4345
rect -1419 4311 -1403 4345
rect -1803 4264 -1403 4311
rect -1345 4345 -945 4361
rect -1345 4311 -1329 4345
rect -961 4311 -945 4345
rect -1345 4264 -945 4311
rect -887 4345 -487 4361
rect -887 4311 -871 4345
rect -503 4311 -487 4345
rect -887 4264 -487 4311
rect -429 4345 -29 4361
rect -429 4311 -413 4345
rect -45 4311 -29 4345
rect -429 4264 -29 4311
rect 29 4345 429 4361
rect 29 4311 45 4345
rect 413 4311 429 4345
rect 29 4264 429 4311
rect 487 4345 887 4361
rect 487 4311 503 4345
rect 871 4311 887 4345
rect 487 4264 887 4311
rect 945 4345 1345 4361
rect 945 4311 961 4345
rect 1329 4311 1345 4345
rect 945 4264 1345 4311
rect 1403 4345 1803 4361
rect 1403 4311 1419 4345
rect 1787 4311 1803 4345
rect 1403 4264 1803 4311
rect 1861 4345 2261 4361
rect 1861 4311 1877 4345
rect 2245 4311 2261 4345
rect 1861 4264 2261 4311
rect 2319 4345 2719 4361
rect 2319 4311 2335 4345
rect 2703 4311 2719 4345
rect 2319 4264 2719 4311
rect -2719 -4362 -2319 -4336
rect -2261 -4362 -1861 -4336
rect -1803 -4362 -1403 -4336
rect -1345 -4362 -945 -4336
rect -887 -4362 -487 -4336
rect -429 -4362 -29 -4336
rect 29 -4362 429 -4336
rect 487 -4362 887 -4336
rect 945 -4362 1345 -4336
rect 1403 -4362 1803 -4336
rect 1861 -4362 2261 -4336
rect 2319 -4362 2719 -4336
<< polycont >>
rect -2703 4311 -2335 4345
rect -2245 4311 -1877 4345
rect -1787 4311 -1419 4345
rect -1329 4311 -961 4345
rect -871 4311 -503 4345
rect -413 4311 -45 4345
rect 45 4311 413 4345
rect 503 4311 871 4345
rect 961 4311 1329 4345
rect 1419 4311 1787 4345
rect 1877 4311 2245 4345
rect 2335 4311 2703 4345
<< locali >>
rect -2719 4311 -2703 4345
rect -2335 4311 -2319 4345
rect -2261 4311 -2245 4345
rect -1877 4311 -1861 4345
rect -1803 4311 -1787 4345
rect -1419 4311 -1403 4345
rect -1345 4311 -1329 4345
rect -961 4311 -945 4345
rect -887 4311 -871 4345
rect -503 4311 -487 4345
rect -429 4311 -413 4345
rect -45 4311 -29 4345
rect 29 4311 45 4345
rect 413 4311 429 4345
rect 487 4311 503 4345
rect 871 4311 887 4345
rect 945 4311 961 4345
rect 1329 4311 1345 4345
rect 1403 4311 1419 4345
rect 1787 4311 1803 4345
rect 1861 4311 1877 4345
rect 2245 4311 2261 4345
rect 2319 4311 2335 4345
rect 2703 4311 2719 4345
rect -2765 4252 -2731 4268
rect -2765 -4340 -2731 -4324
rect -2307 4252 -2273 4268
rect -2307 -4340 -2273 -4324
rect -1849 4252 -1815 4268
rect -1849 -4340 -1815 -4324
rect -1391 4252 -1357 4268
rect -1391 -4340 -1357 -4324
rect -933 4252 -899 4268
rect -933 -4340 -899 -4324
rect -475 4252 -441 4268
rect -475 -4340 -441 -4324
rect -17 4252 17 4268
rect -17 -4340 17 -4324
rect 441 4252 475 4268
rect 441 -4340 475 -4324
rect 899 4252 933 4268
rect 899 -4340 933 -4324
rect 1357 4252 1391 4268
rect 1357 -4340 1391 -4324
rect 1815 4252 1849 4268
rect 1815 -4340 1849 -4324
rect 2273 4252 2307 4268
rect 2273 -4340 2307 -4324
rect 2731 4252 2765 4268
rect 2731 -4340 2765 -4324
<< viali >>
rect -2611 4311 -2427 4345
rect -2153 4311 -1969 4345
rect -1695 4311 -1511 4345
rect -1237 4311 -1053 4345
rect -779 4311 -595 4345
rect -321 4311 -137 4345
rect 137 4311 321 4345
rect 595 4311 779 4345
rect 1053 4311 1237 4345
rect 1511 4311 1695 4345
rect 1969 4311 2153 4345
rect 2427 4311 2611 4345
rect -2765 -4324 -2731 4252
rect -2307 -4324 -2273 4252
rect -1849 -4324 -1815 4252
rect -1391 -4324 -1357 4252
rect -933 -4324 -899 4252
rect -475 -4324 -441 4252
rect -17 -4324 17 4252
rect 441 -4324 475 4252
rect 899 -4324 933 4252
rect 1357 -4324 1391 4252
rect 1815 -4324 1849 4252
rect 2273 -4324 2307 4252
rect 2731 -4324 2765 4252
<< metal1 >>
rect -2623 4345 -2415 4351
rect -2623 4311 -2611 4345
rect -2427 4311 -2415 4345
rect -2623 4305 -2415 4311
rect -2165 4345 -1957 4351
rect -2165 4311 -2153 4345
rect -1969 4311 -1957 4345
rect -2165 4305 -1957 4311
rect -1707 4345 -1499 4351
rect -1707 4311 -1695 4345
rect -1511 4311 -1499 4345
rect -1707 4305 -1499 4311
rect -1249 4345 -1041 4351
rect -1249 4311 -1237 4345
rect -1053 4311 -1041 4345
rect -1249 4305 -1041 4311
rect -791 4345 -583 4351
rect -791 4311 -779 4345
rect -595 4311 -583 4345
rect -791 4305 -583 4311
rect -333 4345 -125 4351
rect -333 4311 -321 4345
rect -137 4311 -125 4345
rect -333 4305 -125 4311
rect 125 4345 333 4351
rect 125 4311 137 4345
rect 321 4311 333 4345
rect 125 4305 333 4311
rect 583 4345 791 4351
rect 583 4311 595 4345
rect 779 4311 791 4345
rect 583 4305 791 4311
rect 1041 4345 1249 4351
rect 1041 4311 1053 4345
rect 1237 4311 1249 4345
rect 1041 4305 1249 4311
rect 1499 4345 1707 4351
rect 1499 4311 1511 4345
rect 1695 4311 1707 4345
rect 1499 4305 1707 4311
rect 1957 4345 2165 4351
rect 1957 4311 1969 4345
rect 2153 4311 2165 4345
rect 1957 4305 2165 4311
rect 2415 4345 2623 4351
rect 2415 4311 2427 4345
rect 2611 4311 2623 4345
rect 2415 4305 2623 4311
rect -2771 4252 -2725 4264
rect -2771 -4324 -2765 4252
rect -2731 -4324 -2725 4252
rect -2771 -4336 -2725 -4324
rect -2313 4252 -2267 4264
rect -2313 -4324 -2307 4252
rect -2273 -4324 -2267 4252
rect -2313 -4336 -2267 -4324
rect -1855 4252 -1809 4264
rect -1855 -4324 -1849 4252
rect -1815 -4324 -1809 4252
rect -1855 -4336 -1809 -4324
rect -1397 4252 -1351 4264
rect -1397 -4324 -1391 4252
rect -1357 -4324 -1351 4252
rect -1397 -4336 -1351 -4324
rect -939 4252 -893 4264
rect -939 -4324 -933 4252
rect -899 -4324 -893 4252
rect -939 -4336 -893 -4324
rect -481 4252 -435 4264
rect -481 -4324 -475 4252
rect -441 -4324 -435 4252
rect -481 -4336 -435 -4324
rect -23 4252 23 4264
rect -23 -4324 -17 4252
rect 17 -4324 23 4252
rect -23 -4336 23 -4324
rect 435 4252 481 4264
rect 435 -4324 441 4252
rect 475 -4324 481 4252
rect 435 -4336 481 -4324
rect 893 4252 939 4264
rect 893 -4324 899 4252
rect 933 -4324 939 4252
rect 893 -4336 939 -4324
rect 1351 4252 1397 4264
rect 1351 -4324 1357 4252
rect 1391 -4324 1397 4252
rect 1351 -4336 1397 -4324
rect 1809 4252 1855 4264
rect 1809 -4324 1815 4252
rect 1849 -4324 1855 4252
rect 1809 -4336 1855 -4324
rect 2267 4252 2313 4264
rect 2267 -4324 2273 4252
rect 2307 -4324 2313 4252
rect 2267 -4336 2313 -4324
rect 2725 4252 2771 4264
rect 2725 -4324 2731 4252
rect 2765 -4324 2771 4252
rect 2725 -4336 2771 -4324
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 43 l 2 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 50 viadrn 100 viasrc 100
string library sky130
<< end >>
