magic
tech sky130A
magscale 1 2
timestamp 1620316209
<< nwell >>
rect -294 -364 294 364
<< pmoslvt >>
rect -200 64 200 264
rect -200 -264 200 -64
<< pdiff >>
rect -258 252 -200 264
rect -258 76 -246 252
rect -212 76 -200 252
rect -258 64 -200 76
rect 200 252 258 264
rect 200 76 212 252
rect 246 76 258 252
rect 200 64 258 76
rect -258 -76 -200 -64
rect -258 -252 -246 -76
rect -212 -252 -200 -76
rect -258 -264 -200 -252
rect 200 -76 258 -64
rect 200 -252 212 -76
rect 246 -252 258 -76
rect 200 -264 258 -252
<< pdiffc >>
rect -246 76 -212 252
rect 212 76 246 252
rect -246 -252 -212 -76
rect 212 -252 246 -76
<< poly >>
rect -200 345 200 361
rect -200 311 -184 345
rect 184 311 200 345
rect -200 264 200 311
rect -200 17 200 64
rect -200 -17 -184 17
rect 184 -17 200 17
rect -200 -64 200 -17
rect -200 -311 200 -264
rect -200 -345 -184 -311
rect 184 -345 200 -311
rect -200 -361 200 -345
<< polycont >>
rect -184 311 184 345
rect -184 -17 184 17
rect -184 -345 184 -311
<< locali >>
rect -200 311 -184 345
rect 184 311 200 345
rect -246 252 -212 268
rect -246 60 -212 76
rect 212 252 246 268
rect 212 60 246 76
rect -200 -17 -184 17
rect 184 -17 200 17
rect -246 -76 -212 -60
rect -246 -268 -212 -252
rect 212 -76 246 -60
rect 212 -268 246 -252
rect -200 -345 -184 -311
rect 184 -345 200 -311
<< viali >>
rect -184 311 184 345
rect -246 76 -212 252
rect 212 76 246 252
rect -184 -17 184 17
rect -246 -252 -212 -76
rect 212 -252 246 -76
rect -184 -345 184 -311
<< metal1 >>
rect -196 345 196 351
rect -196 311 -184 345
rect 184 311 196 345
rect -196 305 196 311
rect -252 252 -206 264
rect -252 76 -246 252
rect -212 76 -206 252
rect -252 64 -206 76
rect 206 252 252 264
rect 206 76 212 252
rect 246 76 252 252
rect 206 64 252 76
rect -196 17 196 23
rect -196 -17 -184 17
rect 184 -17 196 17
rect -196 -23 196 -17
rect -252 -76 -206 -64
rect -252 -252 -246 -76
rect -212 -252 -206 -76
rect -252 -264 -206 -252
rect 206 -76 252 -64
rect 206 -252 212 -76
rect 246 -252 252 -76
rect 206 -264 252 -252
rect -196 -311 196 -305
rect -196 -345 -184 -311
rect 184 -345 196 -311
rect -196 -351 196 -345
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 1 l 2 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
