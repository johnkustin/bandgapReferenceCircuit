magic
tech sky130A
magscale 1 2
timestamp 1620596302
<< nwell >>
rect -900 -200 20 7700
rect 4700 -200 5700 7700
rect 10300 -200 11200 7700
rect 15900 -200 16800 7700
<< nsubdiff >>
rect -800 7200 -200 7400
rect -800 200 -600 7200
rect -400 200 -200 7200
rect -800 0 -200 200
rect 4800 7200 5400 7400
rect 4800 200 5000 7200
rect 5200 200 5400 7200
rect 4800 0 5400 200
rect 10400 7200 11000 7400
rect 10400 200 10600 7200
rect 10800 200 11000 7200
rect 10400 0 11000 200
rect 16000 7200 16600 7400
rect 16000 200 16200 7200
rect 16400 200 16600 7200
rect 16000 0 16600 200
<< nsubdiffcont >>
rect -600 200 -400 7200
rect 5000 200 5200 7200
rect 10600 200 10800 7200
rect 16200 200 16400 7200
<< locali >>
rect -800 8200 -200 8300
rect -800 8100 -700 8200
rect -300 8100 -200 8200
rect -800 7200 -200 8100
rect -800 200 -600 7200
rect -400 200 -200 7200
rect -800 0 -200 200
rect 4800 8200 5400 8300
rect 4800 8100 4900 8200
rect 5300 8100 5400 8200
rect 4800 7200 5400 8100
rect 4800 200 5000 7200
rect 5200 200 5400 7200
rect 4800 0 5400 200
rect 10400 8200 11000 8300
rect 10400 8100 10500 8200
rect 10900 8100 11000 8200
rect 10400 7200 11000 8100
rect 10400 200 10600 7200
rect 10800 200 11000 7200
rect 10400 0 11000 200
rect 16000 8200 16600 8300
rect 16000 8100 16100 8200
rect 16500 8100 16600 8200
rect 16000 7200 16600 8100
rect 16000 200 16200 7200
rect 16400 200 16600 7200
rect 16000 0 16600 200
<< viali >>
rect -700 8100 -300 8200
rect 4900 8100 5300 8200
rect 10500 8100 10900 8200
rect 16100 8100 16500 8200
<< metal1 >>
rect -800 8200 -200 8300
rect -800 8100 -700 8200
rect -300 8100 -200 8200
rect -800 8000 -200 8100
rect 4800 8200 5400 8300
rect 4800 8100 4900 8200
rect 5300 8100 5400 8200
rect 460 8060 580 8080
rect 460 7980 480 8060
rect 560 7980 580 8060
rect 460 7960 580 7980
rect 1380 8060 1500 8080
rect 1380 7980 1400 8060
rect 1480 7980 1500 8060
rect 1380 7960 1500 7980
rect 2300 8060 2420 8080
rect 2300 7980 2320 8060
rect 2400 7980 2420 8060
rect 2300 7960 2420 7980
rect 3220 8060 3340 8080
rect 3220 7980 3240 8060
rect 3320 7980 3340 8060
rect 3220 7960 3340 7980
rect 4140 8060 4260 8080
rect 4140 7980 4160 8060
rect 4240 7980 4260 8060
rect 4800 8000 5400 8100
rect 10400 8200 11000 8300
rect 10400 8100 10500 8200
rect 10900 8100 11000 8200
rect 6060 8060 6180 8080
rect 4140 7960 4260 7980
rect 6060 7980 6080 8060
rect 6160 7980 6180 8060
rect 6060 7960 6180 7980
rect 6980 8060 7100 8080
rect 6980 7980 7000 8060
rect 7080 7980 7100 8060
rect 6980 7960 7100 7980
rect 7900 8060 8020 8080
rect 7900 7980 7920 8060
rect 8000 7980 8020 8060
rect 7900 7960 8020 7980
rect 8820 8060 8940 8080
rect 8820 7980 8840 8060
rect 8920 7980 8940 8060
rect 8820 7960 8940 7980
rect 9740 8060 9860 8080
rect 9740 7980 9760 8060
rect 9840 7980 9860 8060
rect 10400 8000 11000 8100
rect 16000 8200 16600 8300
rect 16000 8100 16100 8200
rect 16500 8100 16600 8200
rect 11660 8060 11780 8080
rect 9740 7960 9860 7980
rect 11660 7980 11680 8060
rect 11760 7980 11780 8060
rect 11660 7960 11780 7980
rect 12580 8060 12700 8080
rect 12580 7980 12600 8060
rect 12680 7980 12700 8060
rect 12580 7960 12700 7980
rect 13500 8060 13620 8080
rect 13500 7980 13520 8060
rect 13600 7980 13620 8060
rect 13500 7960 13620 7980
rect 14420 8060 14540 8080
rect 14420 7980 14440 8060
rect 14520 7980 14540 8060
rect 14420 7960 14540 7980
rect 15340 8060 15460 8080
rect 15340 7980 15360 8060
rect 15440 7980 15460 8060
rect 16000 8000 16600 8100
rect 15340 7960 15460 7980
rect 200 7900 380 7920
rect 200 7780 220 7900
rect 360 7780 380 7900
rect 200 7640 380 7780
rect 500 7580 540 7960
rect 660 7900 840 7920
rect 660 7780 680 7900
rect 820 7780 840 7900
rect 660 7640 840 7780
rect 1120 7900 1300 7920
rect 1120 7780 1140 7900
rect 1280 7780 1300 7900
rect 1120 7640 1300 7780
rect 1420 7580 1460 7960
rect 1580 7900 1760 7920
rect 1580 7780 1600 7900
rect 1740 7780 1760 7900
rect 1580 7640 1760 7780
rect 2040 7900 2220 7920
rect 2040 7780 2060 7900
rect 2200 7780 2220 7900
rect 2040 7640 2220 7780
rect 2340 7580 2380 7960
rect 2500 7900 2680 7920
rect 2500 7780 2520 7900
rect 2660 7780 2680 7900
rect 2500 7640 2680 7780
rect 2960 7900 3140 7920
rect 2960 7780 2980 7900
rect 3120 7780 3140 7900
rect 2960 7640 3140 7780
rect 3240 7580 3280 7960
rect 3420 7900 3600 7920
rect 3420 7780 3440 7900
rect 3580 7780 3600 7900
rect 3420 7640 3600 7780
rect 3880 7900 4060 7920
rect 3880 7780 3900 7900
rect 4040 7780 4060 7900
rect 3880 7640 4060 7780
rect 4160 7580 4200 7960
rect 4340 7900 4520 7920
rect 4340 7780 4360 7900
rect 4500 7780 4520 7900
rect 4340 7640 4520 7780
rect 5800 7900 5980 7920
rect 5800 7780 5820 7900
rect 5960 7780 5980 7900
rect 5800 7640 5980 7780
rect 6100 7580 6140 7960
rect 6260 7900 6440 7920
rect 6260 7780 6280 7900
rect 6420 7780 6440 7900
rect 6260 7640 6440 7780
rect 6720 7900 6900 7920
rect 6720 7780 6740 7900
rect 6880 7780 6900 7900
rect 6720 7640 6900 7780
rect 7020 7580 7060 7960
rect 7180 7900 7360 7920
rect 7180 7780 7200 7900
rect 7340 7780 7360 7900
rect 7180 7640 7360 7780
rect 7640 7900 7820 7920
rect 7640 7780 7660 7900
rect 7800 7780 7820 7900
rect 7640 7640 7820 7780
rect 7940 7580 7980 7960
rect 8100 7900 8280 7920
rect 8100 7780 8120 7900
rect 8260 7780 8280 7900
rect 8100 7640 8280 7780
rect 8560 7900 8740 7920
rect 8560 7780 8580 7900
rect 8720 7780 8740 7900
rect 8560 7640 8740 7780
rect 8840 7580 8880 7960
rect 9020 7900 9200 7920
rect 9020 7780 9040 7900
rect 9180 7780 9200 7900
rect 9020 7640 9200 7780
rect 9480 7900 9660 7920
rect 9480 7780 9500 7900
rect 9640 7780 9660 7900
rect 9480 7640 9660 7780
rect 9760 7580 9800 7960
rect 9940 7900 10120 7920
rect 9940 7780 9960 7900
rect 10100 7780 10120 7900
rect 9940 7640 10120 7780
rect 11400 7900 11580 7920
rect 11400 7780 11420 7900
rect 11560 7780 11580 7900
rect 11400 7640 11580 7780
rect 11700 7580 11740 7960
rect 11860 7900 12040 7920
rect 11860 7780 11880 7900
rect 12020 7780 12040 7900
rect 11860 7640 12040 7780
rect 12320 7900 12500 7920
rect 12320 7780 12340 7900
rect 12480 7780 12500 7900
rect 12320 7640 12500 7780
rect 12620 7580 12660 7960
rect 12780 7900 12960 7920
rect 12780 7780 12800 7900
rect 12940 7780 12960 7900
rect 12780 7640 12960 7780
rect 13240 7900 13420 7920
rect 13240 7780 13260 7900
rect 13400 7780 13420 7900
rect 13240 7640 13420 7780
rect 13540 7580 13580 7960
rect 13700 7900 13880 7920
rect 13700 7780 13720 7900
rect 13860 7780 13880 7900
rect 13700 7640 13880 7780
rect 14160 7900 14340 7920
rect 14160 7780 14180 7900
rect 14320 7780 14340 7900
rect 14160 7640 14340 7780
rect 14440 7580 14480 7960
rect 14620 7900 14800 7920
rect 14620 7780 14640 7900
rect 14780 7780 14800 7900
rect 14620 7640 14800 7780
rect 15080 7900 15260 7920
rect 15080 7780 15100 7900
rect 15240 7780 15260 7900
rect 15080 7640 15260 7780
rect 15360 7580 15400 7960
rect 15540 7900 15720 7920
rect 15540 7780 15560 7900
rect 15700 7780 15720 7900
rect 15540 7640 15720 7780
rect 40 -200 80 -100
rect 960 -180 1000 -120
rect 0 -760 240 -200
rect 920 -420 1040 -180
rect 1880 -200 1920 -100
rect 2780 -200 2840 -120
rect 3700 -200 3760 -100
rect 4620 -200 4680 -100
rect 5640 -200 5680 -120
rect 6560 -200 6600 -120
rect 7480 -200 7520 -100
rect 8400 -200 8440 -100
rect 9300 -200 9360 -100
rect 10220 -200 10280 -100
rect 11240 -200 11280 -100
rect 12160 -200 12200 -100
rect 13080 -200 13120 -100
rect 13980 -200 14040 -100
rect 14900 -200 14960 -120
rect 15820 -200 15860 -120
rect 1840 -220 1960 -200
rect 1840 -300 1860 -220
rect 1940 -300 1960 -220
rect 1840 -340 1960 -300
rect 920 -460 1080 -420
rect 920 -620 940 -460
rect 1060 -620 1080 -460
rect 920 -640 1080 -620
rect 0 -820 260 -760
rect 0 -1160 40 -820
rect 220 -1160 260 -820
rect 0 -1200 260 -1160
rect 2700 -820 2960 -200
rect 3640 -440 3800 -200
rect 4600 -220 4720 -200
rect 4600 -300 4620 -220
rect 4700 -300 4720 -220
rect 4600 -340 4720 -300
rect 3640 -600 3660 -440
rect 3780 -600 3800 -440
rect 3640 -620 3800 -600
rect 2700 -1160 2740 -820
rect 2920 -1160 2960 -820
rect 2700 -1180 2960 -1160
rect 5560 -820 5820 -200
rect 6480 -460 6680 -200
rect 7440 -220 7560 -200
rect 7440 -300 7460 -220
rect 7540 -300 7560 -220
rect 7440 -340 7560 -300
rect 6480 -620 6520 -460
rect 6660 -620 6680 -460
rect 6480 -660 6680 -620
rect 5560 -1160 5600 -820
rect 5780 -1160 5820 -820
rect 5560 -1180 5820 -1160
rect 8260 -820 8520 -200
rect 9220 -440 9420 -200
rect 10180 -220 10300 -200
rect 10180 -300 10200 -220
rect 10280 -300 10300 -220
rect 10180 -340 10300 -300
rect 9220 -640 9240 -440
rect 9400 -640 9420 -440
rect 9220 -660 9420 -640
rect 8260 -1160 8300 -820
rect 8480 -1160 8520 -820
rect 8260 -1180 8520 -1160
rect 11120 -820 11380 -200
rect 12080 -440 12280 -200
rect 13040 -220 13160 -200
rect 13040 -300 13060 -220
rect 13140 -300 13160 -220
rect 13040 -340 13160 -300
rect 12080 -640 12100 -440
rect 12260 -640 12280 -440
rect 12080 -660 12280 -640
rect 11120 -1160 11160 -820
rect 11340 -1160 11380 -820
rect 11120 -1180 11380 -1160
rect 13860 -800 14140 -200
rect 14820 -460 15040 -200
rect 15780 -300 15800 -200
rect 15900 -300 15920 -200
rect 15780 -340 15920 -300
rect 14820 -620 14860 -460
rect 15000 -620 15040 -460
rect 14820 -660 15040 -620
rect 13860 -1160 13880 -800
rect 14120 -1160 14140 -800
rect 13860 -1180 14140 -1160
<< via1 >>
rect -700 8100 -300 8200
rect 4900 8100 5300 8200
rect 480 7980 560 8060
rect 1400 7980 1480 8060
rect 2320 7980 2400 8060
rect 3240 7980 3320 8060
rect 4160 7980 4240 8060
rect 10500 8100 10900 8200
rect 6080 7980 6160 8060
rect 7000 7980 7080 8060
rect 7920 7980 8000 8060
rect 8840 7980 8920 8060
rect 9760 7980 9840 8060
rect 16100 8100 16500 8200
rect 11680 7980 11760 8060
rect 12600 7980 12680 8060
rect 13520 7980 13600 8060
rect 14440 7980 14520 8060
rect 15360 7980 15440 8060
rect 220 7780 360 7900
rect 680 7780 820 7900
rect 1140 7780 1280 7900
rect 1600 7780 1740 7900
rect 2060 7780 2200 7900
rect 2520 7780 2660 7900
rect 2980 7780 3120 7900
rect 3440 7780 3580 7900
rect 3900 7780 4040 7900
rect 4360 7780 4500 7900
rect 5820 7780 5960 7900
rect 6280 7780 6420 7900
rect 6740 7780 6880 7900
rect 7200 7780 7340 7900
rect 7660 7780 7800 7900
rect 8120 7780 8260 7900
rect 8580 7780 8720 7900
rect 9040 7780 9180 7900
rect 9500 7780 9640 7900
rect 9960 7780 10100 7900
rect 11420 7780 11560 7900
rect 11880 7780 12020 7900
rect 12340 7780 12480 7900
rect 12800 7780 12940 7900
rect 13260 7780 13400 7900
rect 13720 7780 13860 7900
rect 14180 7780 14320 7900
rect 14640 7780 14780 7900
rect 15100 7780 15240 7900
rect 15560 7780 15700 7900
rect 1860 -300 1940 -220
rect 940 -620 1060 -460
rect 40 -1160 220 -820
rect 4620 -300 4700 -220
rect 3660 -600 3780 -440
rect 2740 -1160 2920 -820
rect 7460 -300 7540 -220
rect 6520 -620 6660 -460
rect 5600 -1160 5780 -820
rect 10200 -300 10280 -220
rect 9240 -640 9400 -440
rect 8300 -1160 8480 -820
rect 13060 -300 13140 -220
rect 12100 -640 12260 -440
rect 11160 -1160 11340 -820
rect 15800 -300 15900 -200
rect 14860 -620 15000 -460
rect 13880 -1160 14120 -800
<< metal2 >>
rect -800 8200 -200 8300
rect -800 8100 -700 8200
rect -300 8100 -200 8200
rect -800 8000 -200 8100
rect 4800 8200 5400 8300
rect 4800 8100 4900 8200
rect 5300 8100 5400 8200
rect 460 8060 580 8080
rect 460 7980 480 8060
rect 560 7980 580 8060
rect 460 7960 580 7980
rect 1380 8060 1500 8080
rect 1380 7980 1400 8060
rect 1480 7980 1500 8060
rect 1380 7960 1500 7980
rect 2300 8060 2420 8080
rect 2300 7980 2320 8060
rect 2400 7980 2420 8060
rect 2300 7960 2420 7980
rect 3220 8060 3340 8080
rect 3220 7980 3240 8060
rect 3320 7980 3340 8060
rect 3220 7960 3340 7980
rect 4140 8060 4260 8080
rect 4140 7980 4160 8060
rect 4240 7980 4260 8060
rect 4800 8000 5400 8100
rect 10400 8200 11000 8300
rect 10400 8100 10500 8200
rect 10900 8100 11000 8200
rect 6060 8060 6180 8080
rect 4140 7960 4260 7980
rect 6060 7980 6080 8060
rect 6160 7980 6180 8060
rect 6060 7960 6180 7980
rect 6980 8060 7100 8080
rect 6980 7980 7000 8060
rect 7080 7980 7100 8060
rect 6980 7960 7100 7980
rect 7900 8060 8020 8080
rect 7900 7980 7920 8060
rect 8000 7980 8020 8060
rect 7900 7960 8020 7980
rect 8820 8060 8940 8080
rect 8820 7980 8840 8060
rect 8920 7980 8940 8060
rect 8820 7960 8940 7980
rect 9740 8060 9860 8080
rect 9740 7980 9760 8060
rect 9840 7980 9860 8060
rect 10400 8000 11000 8100
rect 16000 8200 16600 8300
rect 16000 8100 16100 8200
rect 16500 8100 16600 8200
rect 11660 8060 11780 8080
rect 9740 7960 9860 7980
rect 11660 7980 11680 8060
rect 11760 7980 11780 8060
rect 11660 7960 11780 7980
rect 12580 8060 12700 8080
rect 12580 7980 12600 8060
rect 12680 7980 12700 8060
rect 12580 7960 12700 7980
rect 13500 8060 13620 8080
rect 13500 7980 13520 8060
rect 13600 7980 13620 8060
rect 13500 7960 13620 7980
rect 14420 8060 14540 8080
rect 14420 7980 14440 8060
rect 14520 7980 14540 8060
rect 14420 7960 14540 7980
rect 15340 8060 15460 8080
rect 15340 7980 15360 8060
rect 15440 7980 15460 8060
rect 16000 8000 16600 8100
rect 15340 7960 15460 7980
rect 200 7900 15720 7920
rect 200 7780 220 7900
rect 360 7780 680 7900
rect 820 7780 1140 7900
rect 1280 7780 1600 7900
rect 1740 7780 2060 7900
rect 2200 7780 2520 7900
rect 2660 7780 2980 7900
rect 3120 7780 3440 7900
rect 3580 7780 3900 7900
rect 4040 7780 4360 7900
rect 4500 7780 5820 7900
rect 5960 7780 6280 7900
rect 6420 7780 6740 7900
rect 6880 7780 7200 7900
rect 7340 7780 7660 7900
rect 7800 7780 8120 7900
rect 8260 7780 8580 7900
rect 8720 7780 9040 7900
rect 9180 7780 9500 7900
rect 9640 7780 9960 7900
rect 10100 7780 11420 7900
rect 11560 7780 11880 7900
rect 12020 7780 12340 7900
rect 12480 7780 12800 7900
rect 12940 7780 13260 7900
rect 13400 7780 13720 7900
rect 13860 7780 14180 7900
rect 14320 7780 14640 7900
rect 14780 7780 15100 7900
rect 15240 7780 15560 7900
rect 15700 7780 15720 7900
rect 200 7760 15720 7780
rect 1800 -220 15800 -200
rect 1800 -300 1860 -220
rect 1940 -300 4620 -220
rect 4700 -300 7460 -220
rect 7540 -300 10200 -220
rect 10280 -300 13060 -220
rect 13140 -300 15800 -220
rect 15900 -300 15920 -200
rect 1800 -340 15920 -300
rect 900 -440 15100 -400
rect 900 -460 3660 -440
rect 900 -620 940 -460
rect 1060 -600 3660 -460
rect 3780 -460 9240 -440
rect 3780 -600 6520 -460
rect 1060 -620 6520 -600
rect 6660 -620 9240 -460
rect 900 -640 9240 -620
rect 9400 -640 12100 -440
rect 12260 -460 15100 -440
rect 12260 -620 14860 -460
rect 15000 -620 15100 -460
rect 12260 -640 15100 -620
rect 900 -700 15100 -640
rect 0 -820 13880 -800
rect 0 -1160 40 -820
rect 220 -1160 2740 -820
rect 2920 -1160 5600 -820
rect 5780 -1160 8300 -820
rect 8480 -1160 11160 -820
rect 11340 -1160 13880 -820
rect 14120 -1160 14180 -800
rect 0 -1200 14180 -1160
<< via2 >>
rect -700 8100 -300 8200
rect 4900 8100 5300 8200
rect 480 7980 560 8060
rect 1400 7980 1480 8060
rect 2320 7980 2400 8060
rect 3240 7980 3320 8060
rect 4160 7980 4240 8060
rect 10500 8100 10900 8200
rect 6080 7980 6160 8060
rect 7000 7980 7080 8060
rect 7920 7980 8000 8060
rect 8840 7980 8920 8060
rect 9760 7980 9840 8060
rect 16100 8100 16500 8200
rect 11680 7980 11760 8060
rect 12600 7980 12680 8060
rect 13520 7980 13600 8060
rect 14440 7980 14520 8060
rect 15360 7980 15440 8060
<< metal3 >>
rect -800 8280 -200 8300
rect 4800 8280 5400 8300
rect 10400 8280 11000 8300
rect 15340 8280 16600 8300
rect -800 8200 16600 8280
rect -800 8100 -700 8200
rect -300 8100 4900 8200
rect 5300 8100 10500 8200
rect 10900 8100 16100 8200
rect 16500 8100 16600 8200
rect -800 8060 16600 8100
rect -800 7980 480 8060
rect 560 7980 1400 8060
rect 1480 7980 2320 8060
rect 2400 7980 3240 8060
rect 3320 7980 4160 8060
rect 4240 7980 6080 8060
rect 6160 7980 7000 8060
rect 7080 7980 7920 8060
rect 8000 7980 8840 8060
rect 8920 7980 9760 8060
rect 9840 7980 11680 8060
rect 11760 7980 12600 8060
rect 12680 7980 13520 8060
rect 13600 7980 14440 8060
rect 14520 7980 15360 8060
rect 15440 7980 16600 8060
rect -800 7960 16600 7980
use sky130_fd_pr__pfet_01v8_lvt_8QZ6MX  sky130_fd_pr__pfet_01v8_lvt_8QZ6MX_0
timestamp 1620594042
transform 1 0 2355 0 1 3768
box -2355 -3968 2355 3934
use sky130_fd_pr__pfet_01v8_lvt_8QZ6MX  sky130_fd_pr__pfet_01v8_lvt_8QZ6MX_2
timestamp 1620594042
transform 1 0 13555 0 1 3768
box -2355 -3968 2355 3934
use sky130_fd_pr__pfet_01v8_lvt_8QZ6MX  sky130_fd_pr__pfet_01v8_lvt_8QZ6MX_1
timestamp 1620594042
transform 1 0 7955 0 1 3768
box -2355 -3968 2355 3934
<< labels >>
flabel space 960 -140 1000 -100 1 FreeSans 800 0 0 0 m2
flabel metal1 1880 -140 1920 -100 1 FreeSans 800 0 0 0 m3
rlabel via1 272 7840 318 7884 1 Vgate
port 1 n
rlabel metal2 13862 -1108 13996 -990 1 Va
port 3 n
rlabel metal2 14808 -610 14942 -492 1 Vb
port 4 n
rlabel metal3 994 8122 1128 8240 1 VDD!
port 0 n
flabel metal1 40 -140 80 -100 1 FreeSans 2 0 0 0 m4
flabel metal1 40 -140 80 -100 1 FreeSans 800 0 0 0 m1
rlabel metal2 15766 -334 15900 -216 1 Vbg
port 2 n
<< end >>
