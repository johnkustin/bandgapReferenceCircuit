magic
tech sky130A
magscale 1 2
timestamp 1620883575
<< psubdiff >>
rect 7484 8216 7590 8232
rect 7484 6600 7500 8216
rect 7574 6600 7590 8216
rect 7484 6584 7590 6600
<< psubdiffcont >>
rect 7500 6600 7574 8216
<< xpolycontact >>
rect 10102 6600 10172 7032
rect 10902 6600 10972 7032
rect 12102 6600 12172 7032
rect 12902 6600 12972 7032
rect 13702 6600 13772 7032
rect 14502 6600 14572 7032
<< locali >>
rect 7484 8216 7590 8232
rect 7484 6600 7500 8216
rect 7574 6600 7590 8216
rect 7484 6584 7590 6600
rect 8400 -5000 8600 5300
rect 9500 -5000 9900 5200
rect 10800 -5000 11200 5200
rect 12100 -5000 12500 5200
rect 13300 -5000 13800 5300
rect 14600 -5000 14800 5300
<< viali >>
rect 7518 7801 7556 8198
rect 7518 6618 7556 7015
rect 10118 6618 10156 7015
rect 10918 6618 10956 7015
rect 12118 6618 12156 7015
rect 12918 6618 12956 7015
rect 13718 6618 13756 7015
rect 14518 6618 14556 7015
<< metal1 >>
rect 13288 8328 13388 8348
rect 13288 8268 13308 8328
rect 13368 8268 13388 8328
rect 13288 8248 13388 8268
rect 7512 8198 7772 8216
rect 7512 7801 7518 8198
rect 7556 7801 7772 8198
rect 7512 7784 7772 7801
rect 8102 8196 8172 8216
rect 8102 8144 8108 8196
rect 8160 8144 8172 8196
rect 8102 7784 8172 8144
rect 8502 7864 8572 8216
rect 8502 7812 8508 7864
rect 8560 7812 8572 7864
rect 8502 7784 8572 7812
rect 8902 8196 8972 8216
rect 8902 8144 8908 8196
rect 8960 8144 8972 8196
rect 8902 7784 8972 8144
rect 9302 7864 9372 8216
rect 9302 7812 9308 7864
rect 9360 7812 9372 7864
rect 9302 7784 9372 7812
rect 9702 8196 9772 8216
rect 9702 8144 9708 8196
rect 9760 8144 9772 8196
rect 9702 7784 9772 8144
rect 10102 7864 10172 8216
rect 10102 7812 10108 7864
rect 10160 7812 10172 7864
rect 10102 7784 10172 7812
rect 10502 8196 10572 8216
rect 10502 8144 10508 8196
rect 10560 8144 10572 8196
rect 10502 7784 10572 8144
rect 10902 7864 10972 8216
rect 10902 7812 10908 7864
rect 10960 7812 10972 7864
rect 10902 7784 10972 7812
rect 8502 7448 8572 7468
rect 8502 7396 8510 7448
rect 8562 7396 8572 7448
rect 7512 7015 7772 7032
rect 7512 6618 7518 7015
rect 7556 6618 7772 7015
rect 7512 6600 7772 6618
rect 8102 5900 8172 7032
rect 8502 6492 8572 7396
rect 11302 7448 11372 8216
rect 11702 8196 11772 8216
rect 11702 8144 11708 8196
rect 11760 8144 11772 8196
rect 11702 7784 11772 8144
rect 12102 7864 12172 8216
rect 12102 7812 12108 7864
rect 12160 7812 12172 7864
rect 12102 7784 12172 7812
rect 12502 8196 12572 8216
rect 12502 8144 12508 8196
rect 12560 8144 12572 8196
rect 12502 7784 12572 8144
rect 12902 7864 12972 8216
rect 12902 7812 12908 7864
rect 12960 7812 12972 7864
rect 12902 7784 12972 7812
rect 13302 7784 13372 8248
rect 13702 7864 13772 8216
rect 13702 7812 13708 7864
rect 13760 7812 13772 7864
rect 13702 7784 13772 7812
rect 14102 8196 14172 8216
rect 14102 8144 14108 8196
rect 14160 8144 14172 8196
rect 14102 7784 14172 8144
rect 14502 7864 14572 8216
rect 14502 7812 14508 7864
rect 14560 7812 14572 7864
rect 14502 7784 14572 7812
rect 11302 7396 11308 7448
rect 11360 7396 11372 7448
rect 11302 7368 11372 7396
rect 8902 6680 8972 7032
rect 8902 6628 8908 6680
rect 8960 6628 8972 6680
rect 8902 6600 8972 6628
rect 9302 7012 9372 7032
rect 9302 6960 9308 7012
rect 9360 6960 9372 7012
rect 9302 6600 9372 6960
rect 9702 6680 9772 7032
rect 9702 6628 9708 6680
rect 9760 6628 9772 6680
rect 9702 6600 9772 6628
rect 10102 7015 10172 7032
rect 10102 7012 10118 7015
rect 10156 7012 10172 7015
rect 10102 6960 10108 7012
rect 10160 6960 10172 7012
rect 10102 6618 10118 6960
rect 10156 6618 10172 6960
rect 10102 6600 10172 6618
rect 10502 6680 10572 7032
rect 10502 6628 10508 6680
rect 10560 6628 10572 6680
rect 10502 6600 10572 6628
rect 10902 7015 10972 7032
rect 10902 7012 10918 7015
rect 10956 7012 10972 7015
rect 10902 6960 10908 7012
rect 10960 6960 10972 7012
rect 10902 6618 10918 6960
rect 10956 6618 10972 6960
rect 10902 6600 10972 6618
rect 11302 6500 11372 7032
rect 11702 6680 11772 7032
rect 11702 6628 11708 6680
rect 11760 6628 11772 6680
rect 11702 6600 11772 6628
rect 12102 7015 12172 7032
rect 12102 7012 12118 7015
rect 12156 7012 12172 7015
rect 12102 6960 12108 7012
rect 12160 6960 12172 7012
rect 12102 6618 12118 6960
rect 12156 6618 12172 6960
rect 12102 6600 12172 6618
rect 12502 6680 12572 7032
rect 12502 6628 12508 6680
rect 12560 6628 12572 6680
rect 12502 6600 12572 6628
rect 12902 7015 12972 7032
rect 12902 7012 12918 7015
rect 12956 7012 12972 7015
rect 12902 6960 12908 7012
rect 12960 6960 12972 7012
rect 12902 6618 12918 6960
rect 12956 6618 12972 6960
rect 12902 6600 12972 6618
rect 13302 6680 13372 7032
rect 13302 6628 13308 6680
rect 13360 6628 13372 6680
rect 13302 6600 13372 6628
rect 13702 7015 13772 7032
rect 13702 6618 13718 7015
rect 13756 6832 13772 7015
rect 14102 6832 14172 7032
rect 13756 6732 14172 6832
rect 13756 6618 13772 6732
rect 13702 6600 13772 6618
rect 14102 6568 14172 6732
rect 14502 7015 14572 7032
rect 14502 7012 14518 7015
rect 14556 7012 14572 7015
rect 14502 6960 14508 7012
rect 14560 6960 14572 7012
rect 14502 6618 14518 6960
rect 14556 6618 14572 6960
rect 14502 6600 14572 6618
rect 14088 6548 14188 6568
rect 8444 6486 8630 6492
rect 8444 6300 8450 6486
rect 8624 6300 8630 6486
rect 8444 6294 8630 6300
rect 8102 5686 9400 5900
rect 8102 5500 8450 5686
rect 8624 5500 9400 5686
rect 8102 4300 9400 5500
rect 11000 5000 11700 6500
rect 14088 6488 14108 6548
rect 14168 6488 14188 6548
rect 14088 6468 14188 6488
rect 10000 3700 14600 5000
rect 8700 -4700 14600 3700
<< via1 >>
rect 13308 8268 13368 8328
rect 8108 8144 8160 8196
rect 8508 7812 8560 7864
rect 8908 8144 8960 8196
rect 9308 7812 9360 7864
rect 9708 8144 9760 8196
rect 10108 7812 10160 7864
rect 10508 8144 10560 8196
rect 10908 7812 10960 7864
rect 8510 7396 8562 7448
rect 11708 8144 11760 8196
rect 12108 7812 12160 7864
rect 12508 8144 12560 8196
rect 12908 7812 12960 7864
rect 13708 7812 13760 7864
rect 14108 8144 14160 8196
rect 14508 7812 14560 7864
rect 11308 7396 11360 7448
rect 8908 6628 8960 6680
rect 9308 6960 9360 7012
rect 9708 6628 9760 6680
rect 10108 6960 10118 7012
rect 10118 6960 10156 7012
rect 10156 6960 10160 7012
rect 10508 6628 10560 6680
rect 10908 6960 10918 7012
rect 10918 6960 10956 7012
rect 10956 6960 10960 7012
rect 11708 6628 11760 6680
rect 12108 6960 12118 7012
rect 12118 6960 12156 7012
rect 12156 6960 12160 7012
rect 12508 6628 12560 6680
rect 12908 6960 12918 7012
rect 12918 6960 12956 7012
rect 12956 6960 12960 7012
rect 13308 6628 13360 6680
rect 14508 6960 14518 7012
rect 14518 6960 14556 7012
rect 14556 6960 14560 7012
rect 8450 6300 8624 6486
rect 8450 5500 8624 5686
rect 14108 6488 14168 6548
<< metal2 >>
rect 13288 8328 14900 8348
rect 13288 8268 13308 8328
rect 13368 8268 14900 8328
rect 13288 8248 14900 8268
rect 8090 8196 8990 8216
rect 8090 8144 8108 8196
rect 8160 8144 8908 8196
rect 8960 8144 8990 8196
rect 8090 8116 8990 8144
rect 9690 8196 10590 8216
rect 9690 8144 9708 8196
rect 9760 8144 10508 8196
rect 10560 8144 10590 8196
rect 9690 8116 10590 8144
rect 11690 8196 14190 8216
rect 11690 8144 11708 8196
rect 11760 8144 12508 8196
rect 12560 8144 14108 8196
rect 14160 8144 14190 8196
rect 11690 8116 14190 8144
rect 8490 7864 9390 7884
rect 8490 7812 8508 7864
rect 8560 7812 9308 7864
rect 9360 7812 9390 7864
rect 8490 7784 9390 7812
rect 10090 7864 10990 7884
rect 10090 7812 10108 7864
rect 10160 7812 10908 7864
rect 10960 7812 10990 7864
rect 10090 7784 10990 7812
rect 12090 7864 13790 7884
rect 12090 7812 12108 7864
rect 12160 7812 12908 7864
rect 12960 7812 13708 7864
rect 13760 7812 13790 7864
rect 12090 7784 13790 7812
rect 14490 7864 14900 7884
rect 14490 7812 14508 7864
rect 14560 7812 14900 7864
rect 14490 7784 14900 7812
rect 8500 7448 11390 7468
rect 8500 7396 8510 7448
rect 8562 7396 11308 7448
rect 11360 7396 11390 7448
rect 8500 7368 11390 7396
rect 9290 7012 10190 7032
rect 9290 6960 9308 7012
rect 9360 6960 10108 7012
rect 10160 6960 10190 7012
rect 9290 6932 10190 6960
rect 10890 7012 12190 7032
rect 10890 6960 10908 7012
rect 10960 6960 12108 7012
rect 12160 6960 12190 7012
rect 10890 6932 12190 6960
rect 12890 7012 14590 7032
rect 12890 6960 12908 7012
rect 12960 6960 14508 7012
rect 14560 6960 14590 7012
rect 12890 6932 14590 6960
rect 8890 6680 9790 6700
rect 8890 6628 8908 6680
rect 8960 6628 9708 6680
rect 9760 6628 9790 6680
rect 8890 6600 9790 6628
rect 10490 6680 11790 6700
rect 10490 6628 10508 6680
rect 10560 6628 11708 6680
rect 11760 6628 11790 6680
rect 10490 6600 11790 6628
rect 12490 6680 13390 6700
rect 12490 6628 12508 6680
rect 12560 6628 13308 6680
rect 13360 6628 13390 6680
rect 12490 6600 13390 6628
rect 14088 6548 14900 6568
rect 8444 6486 8630 6492
rect 8444 6300 8450 6486
rect 8624 6300 8630 6486
rect 14088 6488 14108 6548
rect 14168 6488 14900 6548
rect 14088 6468 14900 6488
rect 8444 6294 8630 6300
rect 8444 5686 8630 5692
rect 8444 5500 8450 5686
rect 8624 5500 8630 5686
rect 8444 5494 8630 5500
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_0
timestamp 1620883575
transform 1 0 8137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_1
timestamp 1620883575
transform 1 0 8537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_4
timestamp 1620883575
transform 1 0 9737 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_3
timestamp 1620883575
transform 1 0 9337 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_2
timestamp 1620883575
transform 1 0 8937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_7
timestamp 1620883575
transform 1 0 10937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_6
timestamp 1620883575
transform 1 0 10537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_5
timestamp 1620883575
transform 1 0 10137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_8
timestamp 1620883575
transform 1 0 11337 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_12
timestamp 1620883575
transform 1 0 12937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_11
timestamp 1620883575
transform 1 0 12537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_10
timestamp 1620883575
transform 1 0 12137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_9
timestamp 1620883575
transform 1 0 11737 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_13
timestamp 1620883575
transform 1 0 13337 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_16
timestamp 1620883575
transform 1 0 14537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_15
timestamp 1620883575
transform 1 0 14137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_14
timestamp 1620883575
transform 1 0 13737 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 7 1288
timestamp 1620883575
transform 1 0 8374 0 1 -5042
box 26 26 1314 1314
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_18
timestamp 1620883575
transform 1 0 14937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_17
timestamp 1620883575
transform 1 0 7737 0 1 7408
box -37 -808 37 808
<< labels >>
flabel metal1 11240 5360 11440 5580 1 FreeSans 800 0 0 0 Vbneg
flabel metal1 8700 5500 9000 5800 1 FreeSans 1600 0 0 0 Va
port 1 n
flabel via1 8458 6304 8606 6468 1 FreeSans 1600 0 0 0 Vb
port 0 n
<< end >>
