magic
tech sky130A
magscale 1 2
timestamp 1620316209
<< nwell >>
rect -396 -13247 396 13247
<< pmoslvt >>
rect -200 4428 200 13028
rect -200 -4300 200 4300
rect -200 -13028 200 -4428
<< pdiff >>
rect -258 13016 -200 13028
rect -258 4440 -246 13016
rect -212 4440 -200 13016
rect -258 4428 -200 4440
rect 200 13016 258 13028
rect 200 4440 212 13016
rect 246 4440 258 13016
rect 200 4428 258 4440
rect -258 4288 -200 4300
rect -258 -4288 -246 4288
rect -212 -4288 -200 4288
rect -258 -4300 -200 -4288
rect 200 4288 258 4300
rect 200 -4288 212 4288
rect 246 -4288 258 4288
rect 200 -4300 258 -4288
rect -258 -4440 -200 -4428
rect -258 -13016 -246 -4440
rect -212 -13016 -200 -4440
rect -258 -13028 -200 -13016
rect 200 -4440 258 -4428
rect 200 -13016 212 -4440
rect 246 -13016 258 -4440
rect 200 -13028 258 -13016
<< pdiffc >>
rect -246 4440 -212 13016
rect 212 4440 246 13016
rect -246 -4288 -212 4288
rect 212 -4288 246 4288
rect -246 -13016 -212 -4440
rect 212 -13016 246 -4440
<< nsubdiff >>
rect -360 13177 -264 13211
rect 264 13177 360 13211
rect -360 13115 -326 13177
rect 326 13115 360 13177
rect -360 -13177 -326 -13115
rect 326 -13177 360 -13115
rect -360 -13211 -264 -13177
rect 264 -13211 360 -13177
<< nsubdiffcont >>
rect -264 13177 264 13211
rect -360 -13115 -326 13115
rect 326 -13115 360 13115
rect -264 -13211 264 -13177
<< poly >>
rect -200 13109 200 13125
rect -200 13075 -184 13109
rect 184 13075 200 13109
rect -200 13028 200 13075
rect -200 4381 200 4428
rect -200 4347 -184 4381
rect 184 4347 200 4381
rect -200 4300 200 4347
rect -200 -4347 200 -4300
rect -200 -4381 -184 -4347
rect 184 -4381 200 -4347
rect -200 -4428 200 -4381
rect -200 -13075 200 -13028
rect -200 -13109 -184 -13075
rect 184 -13109 200 -13075
rect -200 -13125 200 -13109
<< polycont >>
rect -184 13075 184 13109
rect -184 4347 184 4381
rect -184 -4381 184 -4347
rect -184 -13109 184 -13075
<< locali >>
rect -360 13177 -264 13211
rect 264 13177 360 13211
rect -360 13115 -326 13177
rect 326 13115 360 13177
rect -200 13075 -184 13109
rect 184 13075 200 13109
rect -246 13016 -212 13032
rect -246 4424 -212 4440
rect 212 13016 246 13032
rect 212 4424 246 4440
rect -200 4347 -184 4381
rect 184 4347 200 4381
rect -246 4288 -212 4304
rect -246 -4304 -212 -4288
rect 212 4288 246 4304
rect 212 -4304 246 -4288
rect -200 -4381 -184 -4347
rect 184 -4381 200 -4347
rect -246 -4440 -212 -4424
rect -246 -13032 -212 -13016
rect 212 -4440 246 -4424
rect 212 -13032 246 -13016
rect -200 -13109 -184 -13075
rect 184 -13109 200 -13075
rect -360 -13177 -326 -13115
rect 326 -13177 360 -13115
rect -360 -13211 -264 -13177
rect 264 -13211 360 -13177
<< viali >>
rect -184 13075 184 13109
rect -246 4440 -212 13016
rect 212 4440 246 13016
rect -184 4347 184 4381
rect -246 -4288 -212 4288
rect 212 -4288 246 4288
rect -184 -4381 184 -4347
rect -246 -13016 -212 -4440
rect 212 -13016 246 -4440
rect -184 -13109 184 -13075
<< metal1 >>
rect -196 13109 196 13115
rect -196 13075 -184 13109
rect 184 13075 196 13109
rect -196 13069 196 13075
rect -252 13016 -206 13028
rect -252 4440 -246 13016
rect -212 4440 -206 13016
rect -252 4428 -206 4440
rect 206 13016 252 13028
rect 206 4440 212 13016
rect 246 4440 252 13016
rect 206 4428 252 4440
rect -196 4381 196 4387
rect -196 4347 -184 4381
rect 184 4347 196 4381
rect -196 4341 196 4347
rect -252 4288 -206 4300
rect -252 -4288 -246 4288
rect -212 -4288 -206 4288
rect -252 -4300 -206 -4288
rect 206 4288 252 4300
rect 206 -4288 212 4288
rect 246 -4288 252 4288
rect 206 -4300 252 -4288
rect -196 -4347 196 -4341
rect -196 -4381 -184 -4347
rect 184 -4381 196 -4347
rect -196 -4387 196 -4381
rect -252 -4440 -206 -4428
rect -252 -13016 -246 -4440
rect -212 -13016 -206 -4440
rect -252 -13028 -206 -13016
rect 206 -4440 252 -4428
rect 206 -13016 212 -4440
rect 246 -13016 252 -4440
rect 206 -13028 252 -13016
rect -196 -13075 196 -13069
rect -196 -13109 -184 -13075
rect 184 -13109 196 -13075
rect -196 -13115 196 -13109
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -343 -13194 343 13194
string parameters w 43 l 2 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
