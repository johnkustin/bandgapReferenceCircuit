magic
tech sky130A
magscale 1 2
timestamp 1621192096
<< nwell >>
rect -3090 5156 6438 5762
rect -3090 5148 5106 5156
rect -3090 2420 -2290 5148
rect -1774 2420 5106 5148
rect 5622 2420 6438 5156
<< psubdiff >>
rect -1174 1720 -974 1820
rect -1174 120 -1124 1720
rect -1024 120 -974 1720
rect -1174 20 -974 120
rect 4326 1720 4526 1820
rect 4326 120 4376 1720
rect 4476 120 4526 1720
rect 4326 20 4526 120
<< nsubdiff >>
rect 542 5566 3084 5616
rect 542 5466 642 5566
rect 2984 5466 3084 5566
rect 542 5416 3084 5466
rect -2990 4962 -2790 5062
rect -2990 2620 -2940 4962
rect -2840 2620 -2790 4962
rect -2990 2520 -2790 2620
rect 6138 4962 6338 5062
rect 6138 2620 6188 4962
rect 6288 2620 6338 4962
rect 6138 2520 6338 2620
<< psubdiffcont >>
rect -1124 120 -1024 1720
rect 4376 120 4476 1720
<< nsubdiffcont >>
rect 642 5466 2984 5566
rect -2940 2620 -2840 4962
rect 6188 2620 6288 4962
<< locali >>
rect 630 5566 3000 5582
rect 630 5466 642 5566
rect 2984 5466 3000 5566
rect 630 5450 3000 5466
rect -2956 4962 -2824 4978
rect -2956 2620 -2940 4962
rect -2840 2620 -2824 4962
rect -2956 2608 -2824 2620
rect 6172 4962 6304 4978
rect 6172 2620 6188 4962
rect 6288 2620 6304 4962
rect 6172 2608 6304 2620
rect -1140 1720 -1008 1736
rect -1140 120 -1124 1720
rect -1024 120 -1008 1720
rect -1140 104 -1008 120
rect 4360 1720 4492 1736
rect 4360 120 4376 1720
rect 4476 120 4492 1720
rect 4360 104 4492 120
<< viali >>
rect 642 5466 2984 5566
rect -2940 2620 -2840 4962
rect 6188 2620 6288 4962
rect -1124 120 -1024 1718
rect 4376 120 4476 1718
<< metal1 >>
rect 630 5566 3084 5582
rect -1744 5514 -1672 5524
rect -1744 5410 -1734 5514
rect -1682 5410 -1672 5514
rect -1744 5400 -1672 5410
rect -1172 5514 -1100 5524
rect -1172 5410 -1162 5514
rect -1110 5410 -1100 5514
rect -1172 5400 -1100 5410
rect -600 5514 -528 5524
rect -600 5410 -590 5514
rect -538 5410 -528 5514
rect 630 5466 642 5566
rect 2984 5466 3084 5566
rect 630 5450 3084 5466
rect 3404 5514 3476 5524
rect -600 5400 -528 5410
rect 3404 5410 3414 5514
rect 3466 5410 3476 5514
rect 3404 5400 3476 5410
rect 3976 5514 4048 5524
rect 3976 5410 3986 5514
rect 4038 5410 4048 5514
rect 3976 5400 4048 5410
rect 4548 5514 4620 5524
rect 4548 5410 4558 5514
rect 4610 5410 4620 5514
rect 4548 5400 4620 5410
rect -2956 5314 -2824 5324
rect -2956 5210 -2930 5314
rect -2878 5210 -2824 5314
rect -2956 4962 -2824 5210
rect -2318 5314 -2246 5324
rect -2318 5210 -2308 5314
rect -2256 5210 -2246 5314
rect -2318 5200 -2246 5210
rect -1860 5314 -1788 5324
rect -1860 5210 -1850 5314
rect -1798 5210 -1788 5314
rect -1860 5200 -1788 5210
rect -2956 2620 -2940 4962
rect -2840 2620 -2824 4962
rect -2956 2608 -2824 2620
rect -2304 2480 -2258 5200
rect -1846 2480 -1800 5200
rect -1730 2520 -1688 5400
rect -1284 5314 -1212 5324
rect -1284 5210 -1274 5314
rect -1222 5210 -1212 5314
rect -1284 5200 -1212 5210
rect -1268 2536 -1234 5200
rect -1158 2520 -1116 5400
rect -712 5314 -640 5324
rect -712 5210 -702 5314
rect -650 5210 -640 5314
rect -712 5200 -640 5210
rect -696 2536 -654 5200
rect -586 2520 -544 5400
rect -140 5314 -68 5324
rect -140 5210 -130 5314
rect -78 5210 -68 5314
rect -140 5200 -68 5210
rect 432 5314 504 5324
rect 432 5210 442 5314
rect 494 5210 504 5314
rect 432 5200 504 5210
rect 1004 5314 1076 5324
rect 1004 5210 1014 5314
rect 1066 5210 1076 5314
rect 1004 5200 1076 5210
rect 1576 5314 1648 5324
rect 1576 5210 1586 5314
rect 1638 5210 1648 5314
rect 1576 5200 1648 5210
rect 2148 5314 2220 5324
rect 2148 5210 2158 5314
rect 2210 5210 2220 5314
rect 2148 5200 2220 5210
rect 2720 5314 2792 5324
rect 2720 5210 2730 5314
rect 2782 5210 2792 5314
rect 2720 5200 2792 5210
rect 3292 5314 3360 5324
rect 3292 5210 3302 5314
rect 3354 5210 3360 5314
rect 3292 5200 3360 5210
rect -124 2536 -74 5200
rect 448 2536 490 5200
rect 1020 2536 1062 5200
rect -2304 2432 -1800 2480
rect -1584 2386 -1376 2480
rect -1584 2132 -1458 2386
rect -1406 2132 -1376 2386
rect -1584 2126 -1376 2132
rect -1024 2386 -816 2480
rect -1024 2132 -898 2386
rect -846 2132 -816 2386
rect -1024 2126 -816 2132
rect -464 2386 -256 2480
rect -464 2132 -338 2386
rect -286 2132 -256 2386
rect -464 2126 -256 2132
rect -2 2478 32 2536
rect 1592 2532 1626 5200
rect 2164 2532 2198 5200
rect 2736 2532 2770 5200
rect 3308 2532 3342 5200
rect 134 2480 354 2490
rect 134 2478 140 2480
rect -2 2438 140 2478
rect -1140 1718 -1008 1736
rect -1140 120 -1124 1718
rect -1024 120 -1008 1718
rect -1140 104 -1008 120
rect -1130 76 -1016 104
rect -578 76 -532 1902
rect -120 76 -74 1902
rect -2 1896 32 2438
rect 134 2422 140 2438
rect 348 2478 354 2480
rect 348 2442 444 2478
rect 348 2422 354 2442
rect 134 2420 354 2422
rect 570 2392 604 2532
rect 706 2484 926 2490
rect 706 2426 712 2484
rect 920 2426 926 2484
rect 706 2420 926 2426
rect 1142 2474 1176 2532
rect 1278 2480 1498 2486
rect 1278 2474 1284 2480
rect 1142 2438 1284 2474
rect 556 2386 620 2392
rect 556 2132 562 2386
rect 614 2132 620 2386
rect 556 2126 620 2132
rect 432 2086 504 2096
rect 432 1982 442 2086
rect 494 1982 504 2086
rect 432 1972 504 1982
rect 458 120 492 1972
rect 570 1896 604 2126
rect 1004 2086 1076 2096
rect 1004 1982 1014 2086
rect 1066 1982 1076 2086
rect 1004 1972 1076 1982
rect 1030 120 1064 1972
rect 1142 1896 1176 2438
rect 1278 2422 1284 2438
rect 1492 2474 1498 2480
rect 1492 2438 1588 2474
rect 1492 2422 1498 2438
rect 1278 2416 1498 2422
rect 1714 2392 1748 2532
rect 1850 2480 2070 2486
rect 1850 2422 1856 2480
rect 2064 2422 2070 2480
rect 1850 2416 2070 2422
rect 2286 2474 2320 2532
rect 2422 2480 2642 2486
rect 2422 2474 2428 2480
rect 2286 2438 2428 2474
rect 1700 2386 1764 2392
rect 1700 2132 1706 2386
rect 1758 2132 1764 2386
rect 1700 2126 1764 2132
rect 1576 2086 1648 2096
rect 1576 1982 1586 2086
rect 1638 1982 1648 2086
rect 1576 1972 1648 1982
rect 1602 120 1636 1972
rect 1714 1896 1748 2126
rect 2148 2086 2220 2096
rect 2148 1982 2158 2086
rect 2210 1982 2220 2086
rect 2148 1972 2220 1982
rect 2174 120 2208 1972
rect 2286 1896 2320 2438
rect 2422 2422 2428 2438
rect 2636 2474 2642 2480
rect 2636 2438 2732 2474
rect 2636 2422 2642 2438
rect 2422 2416 2642 2422
rect 2858 2392 2892 2532
rect 3418 2520 3460 5400
rect 3864 5314 3932 5324
rect 3864 5210 3874 5314
rect 3926 5210 3932 5314
rect 3864 5200 3932 5210
rect 3880 2532 3914 5200
rect 3990 2520 4032 5400
rect 4436 5314 4504 5324
rect 4436 5210 4446 5314
rect 4498 5210 4504 5314
rect 4436 5200 4504 5210
rect 4452 2532 4486 5200
rect 4562 2520 4604 5400
rect 5008 5314 5076 5324
rect 5008 5210 5018 5314
rect 5070 5210 5076 5314
rect 5008 5200 5076 5210
rect 5118 5314 5190 5324
rect 5118 5210 5128 5314
rect 5180 5210 5190 5314
rect 5118 5200 5190 5210
rect 5576 5314 5648 5324
rect 5576 5210 5586 5314
rect 5638 5210 5648 5314
rect 5576 5200 5648 5210
rect 6172 5314 6304 5324
rect 6172 5210 6198 5314
rect 6250 5210 6304 5314
rect 5024 2532 5058 5200
rect 5132 5088 5178 5200
rect 2994 2480 3214 2486
rect 5132 2480 5178 2532
rect 5590 2480 5636 5200
rect 6172 4962 6304 5210
rect 6172 2620 6188 4962
rect 6288 2620 6304 4962
rect 6172 2608 6304 2620
rect 2994 2422 3000 2480
rect 3208 2422 3214 2480
rect 2994 2416 3214 2422
rect 2844 2386 2908 2392
rect 2844 2132 2850 2386
rect 2902 2132 2908 2386
rect 2844 2126 2908 2132
rect 3564 2386 3772 2480
rect 3564 2132 3650 2386
rect 3702 2132 3772 2386
rect 3564 2126 3772 2132
rect 4124 2386 4332 2480
rect 4124 2132 4210 2386
rect 4262 2132 4332 2386
rect 4124 2126 4332 2132
rect 4684 2386 4892 2480
rect 5132 2432 5636 2480
rect 4684 2132 4770 2386
rect 4822 2132 4892 2386
rect 4684 2126 4892 2132
rect 2720 2086 2792 2096
rect 2720 1982 2730 2086
rect 2782 1982 2792 2086
rect 2720 1972 2792 1982
rect 2746 120 2780 1972
rect 2858 1896 2892 2126
rect 3292 2086 3364 2096
rect 3292 1982 3302 2086
rect 3354 1982 3364 2086
rect 3292 1972 3364 1982
rect 3318 120 3352 1972
rect -1130 30 -74 76
rect 3426 76 3472 1902
rect 4360 1718 4492 1736
rect 4360 120 4376 1718
rect 4476 120 4492 1718
rect 3884 76 3930 120
rect 4360 104 4492 120
rect 4368 76 4482 104
rect 154 -30 338 70
rect 154 -84 174 -30
rect 318 -84 338 -30
rect 154 -104 338 -84
rect 726 -170 910 56
rect 1298 -30 1482 30
rect 1298 -84 1318 -30
rect 1462 -84 1482 -30
rect 1298 -104 1482 -84
rect 726 -224 746 -170
rect 890 -224 910 -170
rect 726 -244 910 -224
rect 1870 -170 2054 56
rect 2442 -30 2626 30
rect 2442 -84 2462 -30
rect 2606 -84 2626 -30
rect 2442 -104 2626 -84
rect 1870 -224 1890 -170
rect 2034 -224 2054 -170
rect 1870 -244 2054 -224
rect 3014 -170 3198 56
rect 3426 30 4482 76
rect 3014 -224 3034 -170
rect 3178 -224 3198 -170
rect 3014 -244 3198 -224
<< via1 >>
rect -1734 5410 -1682 5514
rect -1162 5410 -1110 5514
rect -590 5410 -538 5514
rect 3414 5410 3466 5514
rect 3986 5410 4038 5514
rect 4558 5410 4610 5514
rect -2930 5210 -2878 5314
rect -2308 5210 -2256 5314
rect -1850 5210 -1798 5314
rect -1274 5210 -1222 5314
rect -702 5210 -650 5314
rect -130 5210 -78 5314
rect 442 5210 494 5314
rect 1014 5210 1066 5314
rect 1586 5210 1638 5314
rect 2158 5210 2210 5314
rect 2730 5210 2782 5314
rect 3302 5210 3354 5314
rect -1458 2132 -1406 2386
rect -898 2132 -846 2386
rect -338 2132 -286 2386
rect 140 2422 348 2480
rect 712 2426 920 2484
rect 562 2132 614 2386
rect 442 1982 494 2086
rect 1014 1982 1066 2086
rect 1284 2422 1492 2480
rect 1856 2422 2064 2480
rect 1706 2132 1758 2386
rect 1586 1982 1638 2086
rect 2158 1982 2210 2086
rect 2428 2422 2636 2480
rect 3874 5210 3926 5314
rect 4446 5210 4498 5314
rect 5018 5210 5070 5314
rect 5128 5210 5180 5314
rect 5586 5210 5638 5314
rect 6198 5210 6250 5314
rect 3000 2422 3208 2480
rect 2850 2132 2902 2386
rect 3650 2132 3702 2386
rect 4210 2132 4262 2386
rect 4770 2132 4822 2386
rect 2730 1982 2782 2086
rect 3302 1982 3354 2086
rect 174 -84 318 -30
rect 1318 -84 1462 -30
rect 746 -224 890 -170
rect 2462 -84 2606 -30
rect 1890 -224 2034 -170
rect 3034 -224 3178 -170
<< metal2 >>
rect -1744 5514 4620 5524
rect -1744 5410 -1734 5514
rect -1682 5410 -1162 5514
rect -1110 5410 -590 5514
rect -538 5410 3414 5514
rect 3466 5410 3986 5514
rect 4038 5410 4558 5514
rect 4610 5410 4620 5514
rect -1744 5400 4620 5410
rect -2956 5314 6304 5324
rect -2956 5210 -2930 5314
rect -2878 5210 -2308 5314
rect -2256 5210 -1850 5314
rect -1798 5210 -1274 5314
rect -1222 5210 -702 5314
rect -650 5210 -130 5314
rect -78 5210 442 5314
rect 494 5210 1014 5314
rect 1066 5210 1586 5314
rect 1638 5210 2158 5314
rect 2210 5210 2730 5314
rect 2782 5210 3302 5314
rect 3354 5210 3874 5314
rect 3926 5210 4446 5314
rect 4498 5210 5018 5314
rect 5070 5210 5128 5314
rect 5180 5210 5586 5314
rect 5638 5210 6198 5314
rect 6250 5210 6304 5314
rect -2956 5200 6304 5210
rect 134 2486 1180 2490
rect 134 2484 3214 2486
rect 134 2480 712 2484
rect 134 2422 140 2480
rect 348 2426 712 2480
rect 920 2480 3214 2484
rect 920 2426 1284 2480
rect 348 2422 1284 2426
rect 1492 2422 1856 2480
rect 2064 2422 2428 2480
rect 2636 2422 3000 2480
rect 3208 2422 3214 2480
rect 134 2420 3214 2422
rect -1740 2386 5144 2392
rect -1740 2132 -1458 2386
rect -1406 2132 -898 2386
rect -846 2132 -338 2386
rect -286 2132 562 2386
rect 614 2132 1706 2386
rect 1758 2132 2850 2386
rect 2902 2132 3650 2386
rect 3702 2132 4210 2386
rect 4262 2132 4770 2386
rect 4822 2132 5144 2386
rect -1740 2126 5144 2132
rect 432 2096 842 2098
rect 432 2086 3364 2096
rect 432 1982 442 2086
rect 494 1982 1014 2086
rect 1066 1982 1586 2086
rect 1638 1982 2158 2086
rect 2210 1982 2730 2086
rect 2782 1982 3302 2086
rect 3354 1982 3364 2086
rect 432 1972 3364 1982
rect 154 -30 2626 -24
rect 154 -84 174 -30
rect 318 -84 1318 -30
rect 1462 -84 2462 -30
rect 2606 -84 2626 -30
rect 154 -104 2626 -84
rect 726 -170 3198 -164
rect 726 -224 746 -170
rect 890 -224 1890 -170
rect 2034 -224 3034 -170
rect 3178 -224 3198 -170
rect 726 -244 3198 -224
use sky130_fd_pr__pfet_01v8_lvt_654NJ6  sky130_fd_pr__pfet_01v8_lvt_654NJ6_0
timestamp 1620881708
transform 1 0 1666 0 1 3774
box -4012 -1354 4012 1388
use sky130_fd_pr__nfet_01v8_lvt_VQR4RW  sky130_fd_pr__nfet_01v8_lvt_VQR4RW_0
timestamp 1620881708
transform 1 0 1676 0 1 977
box -2260 -957 2260 957
<< labels >>
flabel metal2 1750 5200 1766 5324 1 FreeSans 800 0 0 0 VDD!
port 0 n
flabel metal2 2404 1972 2420 2096 1 FreeSans 800 0 0 0 Vq
port 6 n
flabel metal2 2346 -244 2362 -164 1 FreeSans 800 0 0 0 Va
port 3 n
flabel metal2 1574 -104 1590 -24 1 FreeSans 800 0 0 0 Vb
port 5 n
flabel metal2 3080 2126 3174 2392 1 FreeSans 800 0 0 0 Vgate
port 1 n
flabel metal2 1356 2126 1450 2392 1 FreeSans 800 0 0 0 Vgate
port 1 n
flabel metal1 -2 2286 32 2378 1 FreeSans 800 0 0 0 vg
flabel metal2 4098 5400 4120 5524 1 FreeSans 800 0 0 0 Vx
port 2 n
flabel psubdiffcont -1124 120 -1024 1720 1 FreeSans 800 0 0 0 GND!
port 4 n
flabel psubdiff 4326 20 4526 120 1 FreeSans 800 180 0 0 GND!
<< end >>
