magic
tech sky130A
magscale 1 2
timestamp 1621288169
<< psubdiff >>
rect -21540 25036 -10308 25060
rect -21540 24270 -21516 25036
rect -10332 24270 -10308 25036
rect -21540 24246 -10308 24270
rect -17906 9382 -11406 9406
rect -17906 9050 -17882 9382
rect -11430 9050 -11406 9382
rect -17906 9026 -11406 9050
<< psubdiffcont >>
rect -21516 24270 -10332 25036
rect -17882 9050 -11430 9382
<< locali >>
rect -17898 9388 -11414 9398
rect -17898 9044 -17888 9388
rect -11424 9044 -11414 9388
rect -17898 9034 -11414 9044
<< viali >>
rect -21532 25036 -10316 25052
rect -21532 24270 -21516 25036
rect -21516 24270 -10332 25036
rect -10332 24270 -10316 25036
rect -21532 24254 -10316 24270
rect -17888 9382 -11424 9388
rect -17888 9050 -17882 9382
rect -17882 9050 -11430 9382
rect -11430 9050 -11424 9382
rect -17888 9044 -11424 9050
<< metal1 >>
rect -21552 25066 -10296 25072
rect -21552 24240 -21546 25066
rect -10302 24240 -10296 25066
rect -21552 24234 -10296 24240
rect -8104 15426 -7556 16438
rect 9804 13500 10508 15196
rect -2890 12808 10508 13500
rect 9278 12640 10226 12646
rect 9278 12122 9286 12640
rect 10220 12122 10226 12640
rect -8390 11860 -6390 11902
rect -8390 11410 -8384 11860
rect -6396 11410 -6390 11860
rect -9908 11104 -9776 11110
rect -9908 10690 -9902 11104
rect -9782 10690 -9776 11104
rect -8390 10996 -6390 11410
rect 5310 11860 7310 11902
rect 5310 11410 5316 11860
rect 7304 11410 7310 11860
rect 5310 10996 7310 11410
rect -10364 10398 -10232 10684
rect -10364 10106 -10358 10398
rect -10238 10106 -10232 10398
rect -17900 9388 -11412 9400
rect -17900 9044 -17888 9388
rect -11424 9044 -11412 9388
rect -17900 8832 -11412 9044
rect -19254 8502 -17208 8710
rect -17894 8038 -11418 8394
rect -18930 5002 -18724 5008
rect -18930 4944 -18924 5002
rect -18730 4944 -18724 5002
rect -18930 1358 -18724 4944
rect -17894 4282 -17686 8038
rect -11626 4282 -11418 8038
rect -10364 6866 -10232 10106
rect -9908 7006 -9776 10690
rect -5690 9502 -3690 10408
rect 2610 9502 4610 10408
rect -9908 6926 -9902 7006
rect -9782 6926 -9776 7006
rect -9908 6920 -9776 6926
rect -10364 6786 -10358 6866
rect -10248 6786 -10232 6866
rect -10364 6780 -10232 6786
rect -9496 4630 -9016 4636
rect -9496 4376 -9490 4630
rect -9022 4376 -9016 4630
rect -9496 1536 -9016 4376
rect 9278 2220 10226 12122
rect 11440 10396 12144 15196
rect 11440 10108 11448 10396
rect 12138 10108 12144 10396
rect 11440 10102 12144 10108
rect -9496 1388 -9490 1536
rect -9022 1388 -9016 1536
rect -9496 1382 -9016 1388
rect -18930 1244 -18924 1358
rect -18730 1244 -18724 1358
rect -18930 1238 -18724 1244
<< via1 >>
rect -21546 25052 -10302 25066
rect -21546 24254 -21532 25052
rect -21532 24254 -10316 25052
rect -10316 24254 -10302 25052
rect -21546 24240 -10302 24254
rect 9286 12122 10220 12640
rect -8384 11410 -6396 11860
rect -9902 10690 -9782 11104
rect 5316 11410 7304 11860
rect -10358 10106 -10238 10398
rect -18924 4944 -18730 5002
rect -9902 6926 -9782 7006
rect -10358 6786 -10248 6866
rect -9490 4376 -9022 4630
rect 10628 11410 11320 11860
rect 11448 10108 12138 10396
rect -9490 1388 -9022 1536
rect -18924 1244 -18730 1358
<< metal2 >>
rect -21561 25072 -10287 25081
rect -21561 24234 -21552 25072
rect -10296 24234 -10287 25072
rect -21561 24225 -10287 24234
rect 5714 12646 6416 14640
rect 5714 12640 10226 12646
rect 5714 12122 9286 12640
rect 10220 12122 10226 12640
rect 5714 12116 10226 12122
rect -9906 11860 11340 11868
rect -9906 11786 -8384 11860
rect -6396 11786 5316 11860
rect 7304 11786 10628 11860
rect -9906 11110 -9252 11786
rect 11320 11410 11340 11860
rect -9908 11104 -9252 11110
rect -9908 10690 -9902 11104
rect -9782 10802 -9252 11104
rect 11070 10802 11340 11410
rect -9782 10690 11340 10802
rect -9908 10686 11340 10690
rect -9908 10684 -9776 10686
rect -10364 10398 12144 10402
rect -10364 10106 -10358 10398
rect -10238 10396 12144 10398
rect -10238 10108 11448 10396
rect 12138 10108 12144 10396
rect -10238 10106 12144 10108
rect -10364 9802 12144 10106
rect -14276 6926 -9902 7006
rect -9782 6926 -9776 7006
rect -14848 6786 -10358 6866
rect -10248 6786 -10242 6866
rect -19536 5002 -18724 5008
rect -19536 4944 -18924 5002
rect -18730 4944 -18724 5002
rect -19536 4938 -18724 4944
rect -21317 4664 -12946 4798
rect -18620 4630 -17980 4636
rect -11488 4630 -9016 4636
rect -18620 4629 -17981 4630
rect -18620 4377 -18600 4629
rect -18000 4377 -17981 4629
rect -18620 4376 -17981 4377
rect -11488 4629 -9490 4630
rect -11488 4377 -10109 4629
rect -9509 4377 -9490 4629
rect -11488 4376 -9490 4377
rect -9022 4376 -9016 4630
rect -18620 4370 -17980 4376
rect -11488 4370 -9016 4376
rect -19268 1438 -19266 1562
rect -10006 1438 -10002 1562
rect -9496 1536 -8010 1542
rect -9496 1388 -9490 1536
rect -9022 1388 -8010 1536
rect -9496 1382 -8010 1388
rect -18930 1362 -18724 1364
rect -18930 1358 -17838 1362
rect -18930 1244 -18924 1358
rect -18730 1244 -17838 1358
rect -18930 1238 -17838 1244
rect -9504 1324 8454 1334
rect -9504 1006 -9494 1324
rect 8444 1006 8454 1324
rect -9504 998 8454 1006
<< via2 >>
rect -21552 25066 -10296 25072
rect -21552 24240 -21546 25066
rect -21546 24240 -10302 25066
rect -10302 24240 -10296 25066
rect -21552 24234 -10296 24240
rect -9252 11410 -8384 11786
rect -8384 11410 -6396 11786
rect -6396 11410 5316 11786
rect 5316 11410 7304 11786
rect 7304 11410 10628 11786
rect 10628 11410 11070 11786
rect -9252 10802 11070 11410
rect -18600 4377 -18000 4629
rect -10109 4377 -9509 4629
rect -19258 1442 -10012 1556
rect -9494 1006 8444 1324
<< metal3 >>
rect -21567 25081 -10281 25087
rect -21567 24225 -21561 25081
rect -10287 24225 -10281 25081
rect -21567 24219 -10281 24225
rect -18620 4643 -17980 4649
rect -18620 4363 -18614 4643
rect -17986 4363 -17980 4643
rect -18620 4357 -17980 4363
rect -17888 1562 -10718 16666
rect -9257 11786 11075 11791
rect -9257 10802 -9252 11786
rect 11070 10802 11075 11786
rect -9257 10797 11075 10802
rect -10129 4643 -9489 4649
rect -10129 4363 -10123 4643
rect -9495 4363 -9489 4643
rect -10129 4357 -9489 4363
rect -19266 1556 8465 1562
rect -19266 1442 -19258 1556
rect -10012 1442 8465 1556
rect -20266 1324 8465 1442
rect -20266 1006 -9494 1324
rect 8444 1006 8465 1324
rect -20266 1000 8465 1006
rect -17888 966 -10718 1000
<< via3 >>
rect -21561 25072 -10287 25081
rect -21561 24234 -21552 25072
rect -21552 24234 -10296 25072
rect -10296 24234 -10287 25072
rect -21561 24225 -10287 24234
rect -18614 4629 -17986 4643
rect -18614 4377 -18600 4629
rect -18600 4377 -18000 4629
rect -18000 4377 -17986 4629
rect -18614 4363 -17986 4377
rect -9246 10808 11064 11780
rect -10123 4629 -9495 4643
rect -10123 4377 -10109 4629
rect -10109 4377 -9509 4629
rect -9509 4377 -9495 4629
rect -10123 4363 -9495 4377
<< metal4 >>
rect -21578 25081 -10252 25118
rect -21578 24225 -21561 25081
rect -10287 24225 -10252 25081
rect -21578 16956 -10252 24225
rect -21532 16950 -10252 16956
rect -17788 9698 -17388 16566
rect -17068 9698 -16668 16566
rect -16348 9698 -15948 16566
rect -15628 9698 -15228 16566
rect -14908 9698 -14508 16566
rect -14188 9698 -13788 16566
rect -13468 9698 -13068 16566
rect -12748 9698 -12348 16566
rect -12028 9698 -11628 16566
rect -11317 16166 -10908 16566
rect -11308 9706 -10908 16166
rect -9247 11780 11065 11781
rect -9247 10808 -9246 11780
rect 11064 10808 11065 11780
rect -9247 10807 11065 10808
rect -11308 9698 -10888 9706
rect -17788 9691 -10888 9698
rect -18614 4645 -9482 9691
rect -18616 4643 -9482 4645
rect -18616 4363 -18614 4643
rect -17986 4363 -10123 4643
rect -9495 4363 -9482 4643
rect -18616 4361 -9482 4363
rect -18614 4360 -9482 4361
<< via4 >>
rect -9246 10808 11064 11780
<< metal5 >>
rect -21532 23950 11082 24225
rect -21532 11780 11238 23950
rect -21532 10808 -9246 11780
rect 11064 10808 11238 11780
rect -21532 10748 11238 10808
rect -9246 10710 11238 10748
use bandgapcorev3  bandgapcorev3_0
timestamp 1621287318
transform 0 1 30186 -1 0 28802
box 5270 -39968 26884 -11302
use amplifier  amplifier_0
timestamp 1621270775
transform 1 0 -16310 0 -1 6762
box -3090 -244 6438 5762
use currentmirror  currentmirror_0
timestamp 1621270775
transform 1 0 -8490 0 -1 9302
box -1748 -4198 17156 8302
use sky130_fd_pr__nfet_01v8_lvt_5FLLME  sky130_fd_pr__nfet_01v8_lvt_5FLLME_0
timestamp 1621270775
transform 0 1 -14507 -1 0 8606
box -258 -2757 258 2757
use sky130_fd_pr__cap_mim_m3_1_LZDD7Y  sky130_fd_pr__cap_mim_m3_1_LZDD7Y_0
timestamp 1621270775
transform 1 0 -14303 0 1 13216
box -3585 -3450 3585 3450
use sky130_fd_pr__cap_mim_m3_2_MZ9F78  sky130_fd_pr__cap_mim_m3_2_MZ9F78_0
timestamp 1621277573
transform 1 0 -15978 0 1 20456
box -5600 -3500 5600 3500
use ampcurrentsource  ampcurrentsource_0
timestamp 1621278611
transform 1 0 -21372 0 1 5166
box -960 -438 2860 694
<< labels >>
flabel metal1 -19254 8502 -18792 8700 1 FreeSans 1600 0 0 0 porst
port 2 n
flabel metal1 -2858 12824 1810 13500 1 FreeSans 1600 0 0 0 Vbg
port 1 n
flabel metal3 -20266 1000 -19556 1422 1 FreeSans 1600 0 0 0 VDD!
<< end >>
