magic
tech sky130A
timestamp 1621277573
<< error_p >>
rect -1798 1495 -1688 1725
rect -2800 1425 -2403 1495
rect -2238 1425 -1688 1495
rect -1678 1495 -1568 1725
rect -1237 1495 -1127 1725
rect -1678 1425 -1127 1495
rect -1117 1495 -1007 1725
rect -676 1495 -566 1725
rect -1117 1425 -566 1495
rect -556 1495 -446 1725
rect -115 1495 -5 1725
rect -556 1425 -5 1495
rect 5 1495 115 1725
rect 446 1495 556 1725
rect 5 1425 556 1495
rect 566 1495 676 1725
rect 1007 1495 1117 1725
rect 566 1425 1117 1495
rect 1127 1495 1237 1725
rect 1568 1495 1678 1725
rect 1127 1425 1678 1495
rect 1688 1495 1798 1725
rect 2129 1495 2239 1725
rect 1688 1425 2239 1495
rect 2249 1495 2359 1725
rect 2249 1425 2800 1495
rect -2800 1305 -2403 1375
rect -2238 1305 -1688 1375
rect -1798 1145 -1688 1305
rect -2800 1075 -2403 1145
rect -2238 1075 -1688 1145
rect -1678 1305 -1127 1375
rect -1678 1145 -1568 1305
rect -1237 1145 -1127 1305
rect -1678 1075 -1127 1145
rect -1117 1305 -566 1375
rect -1117 1145 -1007 1305
rect -676 1145 -566 1305
rect -1117 1075 -566 1145
rect -556 1305 -5 1375
rect -556 1145 -446 1305
rect -115 1145 -5 1305
rect -556 1075 -5 1145
rect 5 1305 556 1375
rect 5 1145 115 1305
rect 446 1145 556 1305
rect 5 1075 556 1145
rect 566 1305 1117 1375
rect 566 1145 676 1305
rect 1007 1145 1117 1305
rect 566 1075 1117 1145
rect 1127 1305 1678 1375
rect 1127 1145 1237 1305
rect 1568 1145 1678 1305
rect 1127 1075 1678 1145
rect 1688 1305 2239 1375
rect 1688 1145 1798 1305
rect 2129 1145 2239 1305
rect 1688 1075 2239 1145
rect 2249 1305 2800 1375
rect 2249 1145 2359 1305
rect 2249 1075 2800 1145
rect -2800 955 -2403 1025
rect -2238 955 -1688 1025
rect -1798 795 -1688 955
rect -2800 725 -2403 795
rect -2238 725 -1688 795
rect -1678 955 -1127 1025
rect -1678 795 -1568 955
rect -1237 795 -1127 955
rect -1678 725 -1127 795
rect -1117 955 -566 1025
rect -1117 795 -1007 955
rect -676 795 -566 955
rect -1117 725 -566 795
rect -556 955 -5 1025
rect -556 795 -446 955
rect -115 795 -5 955
rect -556 725 -5 795
rect 5 955 556 1025
rect 5 795 115 955
rect 446 795 556 955
rect 5 725 556 795
rect 566 955 1117 1025
rect 566 795 676 955
rect 1007 795 1117 955
rect 566 725 1117 795
rect 1127 955 1678 1025
rect 1127 795 1237 955
rect 1568 795 1678 955
rect 1127 725 1678 795
rect 1688 955 2239 1025
rect 1688 795 1798 955
rect 2129 795 2239 955
rect 1688 725 2239 795
rect 2249 955 2800 1025
rect 2249 795 2359 955
rect 2249 725 2800 795
rect -2800 605 -2403 675
rect -2238 605 -1688 675
rect -1798 445 -1688 605
rect -2800 375 -2403 445
rect -2238 375 -1688 445
rect -1678 605 -1127 675
rect -1678 445 -1568 605
rect -1237 445 -1127 605
rect -1678 375 -1127 445
rect -1117 605 -566 675
rect -1117 445 -1007 605
rect -676 445 -566 605
rect -1117 375 -566 445
rect -556 605 -5 675
rect -556 445 -446 605
rect -115 445 -5 605
rect -556 375 -5 445
rect 5 605 556 675
rect 5 445 115 605
rect 446 445 556 605
rect 5 375 556 445
rect 566 605 1117 675
rect 566 445 676 605
rect 1007 445 1117 605
rect 566 375 1117 445
rect 1127 605 1678 675
rect 1127 445 1237 605
rect 1568 445 1678 605
rect 1127 375 1678 445
rect 1688 605 2239 675
rect 1688 445 1798 605
rect 2129 445 2239 605
rect 1688 375 2239 445
rect 2249 605 2800 675
rect 2249 445 2359 605
rect 2249 375 2800 445
rect -2800 255 -2403 325
rect -2238 255 -1688 325
rect -1798 95 -1688 255
rect -2800 25 -2403 95
rect -2238 25 -1688 95
rect -1678 255 -1127 325
rect -1678 95 -1568 255
rect -1237 95 -1127 255
rect -1678 25 -1127 95
rect -1117 255 -566 325
rect -1117 95 -1007 255
rect -676 95 -566 255
rect -1117 25 -566 95
rect -556 255 -5 325
rect -556 95 -446 255
rect -115 95 -5 255
rect -556 25 -5 95
rect 5 255 556 325
rect 5 95 115 255
rect 446 95 556 255
rect 5 25 556 95
rect 566 255 1117 325
rect 566 95 676 255
rect 1007 95 1117 255
rect 566 25 1117 95
rect 1127 255 1678 325
rect 1127 95 1237 255
rect 1568 95 1678 255
rect 1127 25 1678 95
rect 1688 255 2239 325
rect 1688 95 1798 255
rect 2129 95 2239 255
rect 1688 25 2239 95
rect 2249 255 2800 325
rect 2249 95 2359 255
rect 2249 25 2800 95
rect -2800 -95 -2403 -25
rect -2238 -95 -1688 -25
rect -1798 -255 -1688 -95
rect -2800 -325 -2403 -255
rect -2238 -325 -1688 -255
rect -1678 -95 -1127 -25
rect -1678 -255 -1568 -95
rect -1237 -255 -1127 -95
rect -1678 -325 -1127 -255
rect -1117 -95 -566 -25
rect -1117 -255 -1007 -95
rect -676 -255 -566 -95
rect -1117 -325 -566 -255
rect -556 -95 -5 -25
rect -556 -255 -446 -95
rect -115 -255 -5 -95
rect -556 -325 -5 -255
rect 5 -95 556 -25
rect 5 -255 115 -95
rect 446 -255 556 -95
rect 5 -325 556 -255
rect 566 -95 1117 -25
rect 566 -255 676 -95
rect 1007 -255 1117 -95
rect 566 -325 1117 -255
rect 1127 -95 1678 -25
rect 1127 -255 1237 -95
rect 1568 -255 1678 -95
rect 1127 -325 1678 -255
rect 1688 -95 2239 -25
rect 1688 -255 1798 -95
rect 2129 -255 2239 -95
rect 1688 -325 2239 -255
rect 2249 -95 2800 -25
rect 2249 -255 2359 -95
rect 2249 -325 2800 -255
rect -2800 -445 -2403 -375
rect -2238 -445 -1688 -375
rect -1798 -605 -1688 -445
rect -2800 -675 -2403 -605
rect -2238 -675 -1688 -605
rect -1678 -445 -1127 -375
rect -1678 -605 -1568 -445
rect -1237 -605 -1127 -445
rect -1678 -675 -1127 -605
rect -1117 -445 -566 -375
rect -1117 -605 -1007 -445
rect -676 -605 -566 -445
rect -1117 -675 -566 -605
rect -556 -445 -5 -375
rect -556 -605 -446 -445
rect -115 -605 -5 -445
rect -556 -675 -5 -605
rect 5 -445 556 -375
rect 5 -605 115 -445
rect 446 -605 556 -445
rect 5 -675 556 -605
rect 566 -445 1117 -375
rect 566 -605 676 -445
rect 1007 -605 1117 -445
rect 566 -675 1117 -605
rect 1127 -445 1678 -375
rect 1127 -605 1237 -445
rect 1568 -605 1678 -445
rect 1127 -675 1678 -605
rect 1688 -445 2239 -375
rect 1688 -605 1798 -445
rect 2129 -605 2239 -445
rect 1688 -675 2239 -605
rect 2249 -445 2800 -375
rect 2249 -605 2359 -445
rect 2249 -675 2800 -605
rect -2800 -795 -2403 -725
rect -2238 -795 -1688 -725
rect -1798 -955 -1688 -795
rect -2800 -1025 -2403 -955
rect -2238 -1025 -1688 -955
rect -1678 -795 -1127 -725
rect -1678 -955 -1568 -795
rect -1237 -955 -1127 -795
rect -1678 -1025 -1127 -955
rect -1117 -795 -566 -725
rect -1117 -955 -1007 -795
rect -676 -955 -566 -795
rect -1117 -1025 -566 -955
rect -556 -795 -5 -725
rect -556 -955 -446 -795
rect -115 -955 -5 -795
rect -556 -1025 -5 -955
rect 5 -795 556 -725
rect 5 -955 115 -795
rect 446 -955 556 -795
rect 5 -1025 556 -955
rect 566 -795 1117 -725
rect 566 -955 676 -795
rect 1007 -955 1117 -795
rect 566 -1025 1117 -955
rect 1127 -795 1678 -725
rect 1127 -955 1237 -795
rect 1568 -955 1678 -795
rect 1127 -1025 1678 -955
rect 1688 -795 2239 -725
rect 1688 -955 1798 -795
rect 2129 -955 2239 -795
rect 1688 -1025 2239 -955
rect 2249 -795 2800 -725
rect 2249 -955 2359 -795
rect 2249 -1025 2800 -955
rect -2800 -1145 -2403 -1075
rect -2238 -1145 -1688 -1075
rect -1798 -1305 -1688 -1145
rect -2800 -1375 -2403 -1305
rect -2238 -1375 -1688 -1305
rect -1678 -1145 -1127 -1075
rect -1678 -1305 -1568 -1145
rect -1237 -1305 -1127 -1145
rect -1678 -1375 -1127 -1305
rect -1117 -1145 -566 -1075
rect -1117 -1305 -1007 -1145
rect -676 -1305 -566 -1145
rect -1117 -1375 -566 -1305
rect -556 -1145 -5 -1075
rect -556 -1305 -446 -1145
rect -115 -1305 -5 -1145
rect -556 -1375 -5 -1305
rect 5 -1145 556 -1075
rect 5 -1305 115 -1145
rect 446 -1305 556 -1145
rect 5 -1375 556 -1305
rect 566 -1145 1117 -1075
rect 566 -1305 676 -1145
rect 1007 -1305 1117 -1145
rect 566 -1375 1117 -1305
rect 1127 -1145 1678 -1075
rect 1127 -1305 1237 -1145
rect 1568 -1305 1678 -1145
rect 1127 -1375 1678 -1305
rect 1688 -1145 2239 -1075
rect 1688 -1305 1798 -1145
rect 2129 -1305 2239 -1145
rect 1688 -1375 2239 -1305
rect 2249 -1145 2800 -1075
rect 2249 -1305 2359 -1145
rect 2249 -1375 2800 -1305
rect -2800 -1495 -2403 -1425
rect -2238 -1495 -1688 -1425
rect -1798 -1725 -1688 -1495
rect -1678 -1495 -1127 -1425
rect -1678 -1725 -1568 -1495
rect -1237 -1725 -1127 -1495
rect -1117 -1495 -566 -1425
rect -1117 -1725 -1007 -1495
rect -676 -1725 -566 -1495
rect -556 -1495 -5 -1425
rect -556 -1725 -446 -1495
rect -115 -1725 -5 -1495
rect 5 -1495 556 -1425
rect 5 -1725 115 -1495
rect 446 -1725 556 -1495
rect 566 -1495 1117 -1425
rect 566 -1725 676 -1495
rect 1007 -1725 1117 -1495
rect 1127 -1495 1678 -1425
rect 1127 -1725 1237 -1495
rect 1568 -1725 1678 -1495
rect 1688 -1495 2239 -1425
rect 1688 -1725 1798 -1495
rect 2129 -1725 2239 -1495
rect 2249 -1495 2800 -1425
rect 2249 -1725 2359 -1495
<< metal4 >>
rect -2800 1425 -2403 1725
rect -2238 1425 -1688 1725
rect -1678 1425 -1127 1725
rect -1117 1425 -566 1725
rect -556 1425 -5 1725
rect 5 1425 556 1725
rect 566 1425 1117 1725
rect 1127 1425 1678 1725
rect 1688 1425 2239 1725
rect 2249 1425 2800 1725
rect -2800 1075 -2403 1375
rect -2238 1075 -1688 1375
rect -1678 1075 -1127 1375
rect -1117 1075 -566 1375
rect -556 1075 -5 1375
rect 5 1075 556 1375
rect 566 1075 1117 1375
rect 1127 1075 1678 1375
rect 1688 1075 2239 1375
rect 2249 1075 2800 1375
rect -2800 725 -2403 1025
rect -2238 725 -1688 1025
rect -1678 725 -1127 1025
rect -1117 725 -566 1025
rect -556 725 -5 1025
rect 5 725 556 1025
rect 566 725 1117 1025
rect 1127 725 1678 1025
rect 1688 725 2239 1025
rect 2249 725 2800 1025
rect -2800 375 -2403 675
rect -2238 375 -1688 675
rect -1678 375 -1127 675
rect -1117 375 -566 675
rect -556 375 -5 675
rect 5 375 556 675
rect 566 375 1117 675
rect 1127 375 1678 675
rect 1688 375 2239 675
rect 2249 375 2800 675
rect -2800 25 -2403 325
rect -2238 25 -1688 325
rect -1678 25 -1127 325
rect -1117 25 -566 325
rect -556 25 -5 325
rect 5 25 556 325
rect 566 25 1117 325
rect 1127 25 1678 325
rect 1688 25 2239 325
rect 2249 25 2800 325
rect -2800 -325 -2403 -25
rect -2238 -325 -1688 -25
rect -1678 -325 -1127 -25
rect -1117 -325 -566 -25
rect -556 -325 -5 -25
rect 5 -325 556 -25
rect 566 -325 1117 -25
rect 1127 -325 1678 -25
rect 1688 -325 2239 -25
rect 2249 -325 2800 -25
rect -2800 -675 -2403 -375
rect -2238 -675 -1688 -375
rect -1678 -675 -1127 -375
rect -1117 -675 -566 -375
rect -556 -675 -5 -375
rect 5 -675 556 -375
rect 566 -675 1117 -375
rect 1127 -675 1678 -375
rect 1688 -675 2239 -375
rect 2249 -675 2800 -375
rect -2800 -1025 -2403 -725
rect -2238 -1025 -1688 -725
rect -1678 -1025 -1127 -725
rect -1117 -1025 -566 -725
rect -556 -1025 -5 -725
rect 5 -1025 556 -725
rect 566 -1025 1117 -725
rect 1127 -1025 1678 -725
rect 1688 -1025 2239 -725
rect 2249 -1025 2800 -725
rect -2800 -1375 -2403 -1075
rect -2238 -1375 -1688 -1075
rect -1678 -1375 -1127 -1075
rect -1117 -1375 -566 -1075
rect -556 -1375 -5 -1075
rect 5 -1375 556 -1075
rect 566 -1375 1117 -1075
rect 1127 -1375 1678 -1075
rect 1688 -1375 2239 -1075
rect 2249 -1375 2800 -1075
rect -2800 -1725 -2403 -1425
rect -2238 -1725 -1688 -1425
rect -1678 -1725 -1127 -1425
rect -1117 -1725 -566 -1425
rect -556 -1725 -5 -1425
rect 5 -1725 556 -1425
rect 566 -1725 1117 -1425
rect 1127 -1725 1678 -1425
rect 1688 -1725 2239 -1425
rect 2249 -1725 2800 -1425
<< mimcap2 >>
rect -2750 1655 -2550 1675
rect -2750 1495 -2730 1655
rect -2570 1495 -2550 1655
rect -2750 1475 -2550 1495
rect -2189 1475 -1989 1675
rect -1628 1475 -1428 1675
rect -1067 1475 -867 1675
rect -506 1475 -306 1675
rect 55 1475 255 1675
rect 616 1475 816 1675
rect 1177 1475 1377 1675
rect 1738 1475 1938 1675
rect 2299 1475 2499 1675
rect -2750 1305 -2550 1325
rect -2750 1145 -2730 1305
rect -2570 1145 -2550 1305
rect -2750 1125 -2550 1145
rect -2189 1125 -1989 1325
rect -1628 1125 -1428 1325
rect -1067 1125 -867 1325
rect -506 1125 -306 1325
rect 55 1125 255 1325
rect 616 1125 816 1325
rect 1177 1125 1377 1325
rect 1738 1125 1938 1325
rect 2299 1125 2499 1325
rect -2750 955 -2550 975
rect -2750 795 -2730 955
rect -2570 795 -2550 955
rect -2750 775 -2550 795
rect -2189 775 -1989 975
rect -1628 775 -1428 975
rect -1067 775 -867 975
rect -506 775 -306 975
rect 55 775 255 975
rect 616 775 816 975
rect 1177 775 1377 975
rect 1738 775 1938 975
rect 2299 775 2499 975
rect -2750 605 -2550 625
rect -2750 445 -2730 605
rect -2570 445 -2550 605
rect -2750 425 -2550 445
rect -2189 425 -1989 625
rect -1628 425 -1428 625
rect -1067 425 -867 625
rect -506 425 -306 625
rect 55 425 255 625
rect 616 425 816 625
rect 1177 425 1377 625
rect 1738 425 1938 625
rect 2299 425 2499 625
rect -2750 255 -2550 275
rect -2750 95 -2730 255
rect -2570 95 -2550 255
rect -2750 75 -2550 95
rect -2189 75 -1989 275
rect -1628 75 -1428 275
rect -1067 75 -867 275
rect -506 75 -306 275
rect 55 75 255 275
rect 616 75 816 275
rect 1177 75 1377 275
rect 1738 75 1938 275
rect 2299 75 2499 275
rect -2750 -95 -2550 -75
rect -2750 -255 -2730 -95
rect -2570 -255 -2550 -95
rect -2750 -275 -2550 -255
rect -2189 -275 -1989 -75
rect -1628 -275 -1428 -75
rect -1067 -275 -867 -75
rect -506 -275 -306 -75
rect 55 -275 255 -75
rect 616 -275 816 -75
rect 1177 -275 1377 -75
rect 1738 -275 1938 -75
rect 2299 -275 2499 -75
rect -2750 -445 -2550 -425
rect -2750 -605 -2730 -445
rect -2570 -605 -2550 -445
rect -2750 -625 -2550 -605
rect -2189 -625 -1989 -425
rect -1628 -625 -1428 -425
rect -1067 -625 -867 -425
rect -506 -625 -306 -425
rect 55 -625 255 -425
rect 616 -625 816 -425
rect 1177 -625 1377 -425
rect 1738 -625 1938 -425
rect 2299 -625 2499 -425
rect -2750 -795 -2550 -775
rect -2750 -955 -2730 -795
rect -2570 -955 -2550 -795
rect -2750 -975 -2550 -955
rect -2189 -975 -1989 -775
rect -1628 -975 -1428 -775
rect -1067 -975 -867 -775
rect -506 -975 -306 -775
rect 55 -975 255 -775
rect 616 -975 816 -775
rect 1177 -975 1377 -775
rect 1738 -975 1938 -775
rect 2299 -975 2499 -775
rect -2750 -1145 -2550 -1125
rect -2750 -1305 -2730 -1145
rect -2570 -1305 -2550 -1145
rect -2750 -1325 -2550 -1305
rect -2189 -1325 -1989 -1125
rect -1628 -1325 -1428 -1125
rect -1067 -1325 -867 -1125
rect -506 -1325 -306 -1125
rect 55 -1325 255 -1125
rect 616 -1325 816 -1125
rect 1177 -1325 1377 -1125
rect 1738 -1325 1938 -1125
rect 2299 -1325 2499 -1125
rect -2750 -1495 -2550 -1475
rect -2750 -1655 -2730 -1495
rect -2570 -1655 -2550 -1495
rect -2750 -1675 -2550 -1655
rect -2189 -1675 -1989 -1475
rect -1628 -1675 -1428 -1475
rect -1067 -1675 -867 -1475
rect -506 -1675 -306 -1475
rect 55 -1675 255 -1475
rect 616 -1675 816 -1475
rect 1177 -1675 1377 -1475
rect 1738 -1675 1938 -1475
rect 2299 -1675 2499 -1475
<< mimcap2contact >>
rect -2730 1495 -2570 1655
rect -2730 1145 -2570 1305
rect -2730 795 -2570 955
rect -2730 445 -2570 605
rect -2730 95 -2570 255
rect -2730 -255 -2570 -95
rect -2730 -605 -2570 -445
rect -2730 -955 -2570 -795
rect -2730 -1305 -2570 -1145
rect -2730 -1655 -2570 -1495
<< metal5 >>
rect -2730 1667 -2410 1750
rect -2742 1655 -2410 1667
rect -2742 1495 -2730 1655
rect -2570 1495 -2410 1655
rect -2742 1483 -2410 1495
rect -2730 1317 -2410 1483
rect -2742 1305 -2410 1317
rect -2742 1145 -2730 1305
rect -2570 1145 -2410 1305
rect -2742 1133 -2410 1145
rect -2730 967 -2410 1133
rect -2742 955 -2410 967
rect -2742 795 -2730 955
rect -2570 795 -2410 955
rect -2742 783 -2410 795
rect -2730 617 -2410 783
rect -2742 605 -2410 617
rect -2742 445 -2730 605
rect -2570 445 -2410 605
rect -2742 433 -2410 445
rect -2730 267 -2410 433
rect -2742 255 -2410 267
rect -2742 95 -2730 255
rect -2570 95 -2410 255
rect -2742 83 -2410 95
rect -2730 -83 -2410 83
rect -2742 -95 -2410 -83
rect -2742 -255 -2730 -95
rect -2570 -255 -2410 -95
rect -2742 -267 -2410 -255
rect -2730 -433 -2410 -267
rect -2742 -445 -2410 -433
rect -2742 -605 -2730 -445
rect -2570 -605 -2410 -445
rect -2742 -617 -2410 -605
rect -2730 -783 -2410 -617
rect -2742 -795 -2410 -783
rect -2742 -955 -2730 -795
rect -2570 -955 -2410 -795
rect -2742 -967 -2410 -955
rect -2730 -1133 -2410 -967
rect -2742 -1145 -2410 -1133
rect -2742 -1305 -2730 -1145
rect -2570 -1305 -2410 -1145
rect -2742 -1317 -2410 -1305
rect -2730 -1483 -2410 -1317
rect -2742 -1495 -2410 -1483
rect -2742 -1655 -2730 -1495
rect -2570 -1655 -2410 -1495
rect -2742 -1667 -2410 -1655
rect -2730 -1750 -2410 -1667
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX 2249 1425 2549 1725
string parameters w 2.00 l 2.00 val 5.36 carea 1.00 cperi 0.17 nx 10 ny 10 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
