magic
tech sky130A
magscale 1 2
timestamp 1622134248
<< psubdiff >>
rect 298846 617944 298856 624600
rect 343126 617944 343136 624600
<< locali >>
rect 298846 617944 298880 624600
rect 343126 617944 343160 624600
<< viali >>
rect 298876 642594 298976 642694
rect 299100 642594 299200 642694
rect 299324 642594 299424 642694
rect 299548 642594 299648 642694
rect 299772 642594 299872 642694
rect 299996 642594 300096 642694
rect 300220 642594 300320 642694
rect 300444 642594 300544 642694
rect 300668 642594 300768 642694
rect 300892 642594 300992 642694
rect 301116 642594 301216 642694
rect 301340 642594 301440 642694
rect 301564 642594 301664 642694
rect 301788 642594 301888 642694
rect 302012 642594 302112 642694
rect 302236 642594 302336 642694
rect 302460 642594 302560 642694
rect 302684 642594 302784 642694
rect 302908 642594 303008 642694
rect 303132 642594 303232 642694
rect 303356 642594 303456 642694
rect 303580 642594 303680 642694
rect 303804 642594 303904 642694
rect 304028 642594 304128 642694
rect 304252 642594 304352 642694
rect 304476 642594 304576 642694
rect 304700 642594 304800 642694
rect 304924 642594 305024 642694
rect 305148 642594 305248 642694
rect 305372 642594 305472 642694
rect 309346 642594 309446 642694
rect 309570 642594 309670 642694
rect 309794 642594 309894 642694
rect 310018 642594 310118 642694
rect 310242 642594 310342 642694
rect 310466 642594 310566 642694
rect 310690 642594 310790 642694
rect 310914 642594 311014 642694
rect 311138 642594 311238 642694
rect 311362 642594 311462 642694
rect 311586 642594 311686 642694
rect 311810 642594 311910 642694
rect 312034 642594 312134 642694
rect 312258 642594 312358 642694
rect 312482 642594 312582 642694
rect 312706 642594 312806 642694
rect 312930 642594 313030 642694
rect 313154 642594 313254 642694
rect 313378 642594 313478 642694
rect 313602 642594 313702 642694
rect 313826 642594 313926 642694
rect 314050 642594 314150 642694
rect 314274 642594 314374 642694
rect 314498 642594 314598 642694
rect 314722 642594 314822 642694
rect 314946 642594 315046 642694
rect 315170 642594 315270 642694
rect 315394 642594 315494 642694
rect 315618 642594 315718 642694
rect 315842 642594 315942 642694
rect 335616 642614 335716 642714
rect 335840 642614 335940 642714
rect 336064 642614 336164 642714
rect 336288 642614 336388 642714
rect 336512 642614 336612 642714
rect 336736 642614 336836 642714
rect 336960 642614 337060 642714
rect 337184 642614 337284 642714
rect 337408 642614 337508 642714
rect 337632 642614 337732 642714
rect 337856 642614 337956 642714
rect 338080 642614 338180 642714
rect 338304 642614 338404 642714
rect 338528 642614 338628 642714
rect 338752 642614 338852 642714
rect 338976 642614 339076 642714
rect 339200 642614 339300 642714
rect 339424 642614 339524 642714
rect 339648 642614 339748 642714
rect 339872 642614 339972 642714
rect 340096 642614 340196 642714
rect 340320 642614 340420 642714
rect 340544 642614 340644 642714
rect 340768 642614 340868 642714
rect 340992 642614 341092 642714
rect 341216 642614 341316 642714
rect 341440 642614 341540 642714
rect 341664 642614 341764 642714
rect 341888 642614 341988 642714
rect 342112 642614 342212 642714
rect 298876 642370 298976 642470
rect 299100 642370 299200 642470
rect 299324 642370 299424 642470
rect 299548 642370 299648 642470
rect 299772 642370 299872 642470
rect 299996 642370 300096 642470
rect 300220 642370 300320 642470
rect 300444 642370 300544 642470
rect 300668 642370 300768 642470
rect 300892 642370 300992 642470
rect 301116 642370 301216 642470
rect 301340 642370 301440 642470
rect 301564 642370 301664 642470
rect 301788 642370 301888 642470
rect 302012 642370 302112 642470
rect 302236 642370 302336 642470
rect 302460 642370 302560 642470
rect 302684 642370 302784 642470
rect 302908 642370 303008 642470
rect 303132 642370 303232 642470
rect 303356 642370 303456 642470
rect 303580 642370 303680 642470
rect 303804 642370 303904 642470
rect 304028 642370 304128 642470
rect 304252 642370 304352 642470
rect 304476 642370 304576 642470
rect 304700 642370 304800 642470
rect 304924 642370 305024 642470
rect 305148 642370 305248 642470
rect 305372 642370 305472 642470
rect 309346 642370 309446 642470
rect 309570 642370 309670 642470
rect 309794 642370 309894 642470
rect 310018 642370 310118 642470
rect 310242 642370 310342 642470
rect 310466 642370 310566 642470
rect 310690 642370 310790 642470
rect 310914 642370 311014 642470
rect 311138 642370 311238 642470
rect 311362 642370 311462 642470
rect 311586 642370 311686 642470
rect 311810 642370 311910 642470
rect 312034 642370 312134 642470
rect 312258 642370 312358 642470
rect 312482 642370 312582 642470
rect 312706 642370 312806 642470
rect 312930 642370 313030 642470
rect 313154 642370 313254 642470
rect 313378 642370 313478 642470
rect 313602 642370 313702 642470
rect 313826 642370 313926 642470
rect 314050 642370 314150 642470
rect 314274 642370 314374 642470
rect 314498 642370 314598 642470
rect 314722 642370 314822 642470
rect 314946 642370 315046 642470
rect 315170 642370 315270 642470
rect 315394 642370 315494 642470
rect 315618 642370 315718 642470
rect 315842 642370 315942 642470
rect 335616 642390 335716 642490
rect 335840 642390 335940 642490
rect 336064 642390 336164 642490
rect 336288 642390 336388 642490
rect 336512 642390 336612 642490
rect 336736 642390 336836 642490
rect 336960 642390 337060 642490
rect 337184 642390 337284 642490
rect 337408 642390 337508 642490
rect 337632 642390 337732 642490
rect 337856 642390 337956 642490
rect 338080 642390 338180 642490
rect 338304 642390 338404 642490
rect 338528 642390 338628 642490
rect 338752 642390 338852 642490
rect 338976 642390 339076 642490
rect 339200 642390 339300 642490
rect 339424 642390 339524 642490
rect 339648 642390 339748 642490
rect 339872 642390 339972 642490
rect 340096 642390 340196 642490
rect 340320 642390 340420 642490
rect 340544 642390 340644 642490
rect 340768 642390 340868 642490
rect 340992 642390 341092 642490
rect 341216 642390 341316 642490
rect 341440 642390 341540 642490
rect 341664 642390 341764 642490
rect 341888 642390 341988 642490
rect 342112 642390 342212 642490
rect 298876 642146 298976 642246
rect 299100 642146 299200 642246
rect 299324 642146 299424 642246
rect 299548 642146 299648 642246
rect 299772 642146 299872 642246
rect 299996 642146 300096 642246
rect 300220 642146 300320 642246
rect 300444 642146 300544 642246
rect 300668 642146 300768 642246
rect 300892 642146 300992 642246
rect 301116 642146 301216 642246
rect 301340 642146 301440 642246
rect 301564 642146 301664 642246
rect 301788 642146 301888 642246
rect 302012 642146 302112 642246
rect 302236 642146 302336 642246
rect 302460 642146 302560 642246
rect 302684 642146 302784 642246
rect 302908 642146 303008 642246
rect 303132 642146 303232 642246
rect 303356 642146 303456 642246
rect 303580 642146 303680 642246
rect 303804 642146 303904 642246
rect 304028 642146 304128 642246
rect 304252 642146 304352 642246
rect 304476 642146 304576 642246
rect 304700 642146 304800 642246
rect 304924 642146 305024 642246
rect 305148 642146 305248 642246
rect 305372 642146 305472 642246
rect 309346 642146 309446 642246
rect 309570 642146 309670 642246
rect 309794 642146 309894 642246
rect 310018 642146 310118 642246
rect 310242 642146 310342 642246
rect 310466 642146 310566 642246
rect 310690 642146 310790 642246
rect 310914 642146 311014 642246
rect 311138 642146 311238 642246
rect 311362 642146 311462 642246
rect 311586 642146 311686 642246
rect 311810 642146 311910 642246
rect 312034 642146 312134 642246
rect 312258 642146 312358 642246
rect 312482 642146 312582 642246
rect 312706 642146 312806 642246
rect 312930 642146 313030 642246
rect 313154 642146 313254 642246
rect 313378 642146 313478 642246
rect 313602 642146 313702 642246
rect 313826 642146 313926 642246
rect 314050 642146 314150 642246
rect 314274 642146 314374 642246
rect 314498 642146 314598 642246
rect 314722 642146 314822 642246
rect 314946 642146 315046 642246
rect 315170 642146 315270 642246
rect 315394 642146 315494 642246
rect 315618 642146 315718 642246
rect 315842 642146 315942 642246
rect 335616 642166 335716 642266
rect 335840 642166 335940 642266
rect 336064 642166 336164 642266
rect 336288 642166 336388 642266
rect 336512 642166 336612 642266
rect 336736 642166 336836 642266
rect 336960 642166 337060 642266
rect 337184 642166 337284 642266
rect 337408 642166 337508 642266
rect 337632 642166 337732 642266
rect 337856 642166 337956 642266
rect 338080 642166 338180 642266
rect 338304 642166 338404 642266
rect 338528 642166 338628 642266
rect 338752 642166 338852 642266
rect 338976 642166 339076 642266
rect 339200 642166 339300 642266
rect 339424 642166 339524 642266
rect 339648 642166 339748 642266
rect 339872 642166 339972 642266
rect 340096 642166 340196 642266
rect 340320 642166 340420 642266
rect 340544 642166 340644 642266
rect 340768 642166 340868 642266
rect 340992 642166 341092 642266
rect 341216 642166 341316 642266
rect 341440 642166 341540 642266
rect 341664 642166 341764 642266
rect 341888 642166 341988 642266
rect 342112 642166 342212 642266
rect 298876 641922 298976 642022
rect 299100 641922 299200 642022
rect 299324 641922 299424 642022
rect 299548 641922 299648 642022
rect 299772 641922 299872 642022
rect 299996 641922 300096 642022
rect 300220 641922 300320 642022
rect 300444 641922 300544 642022
rect 300668 641922 300768 642022
rect 300892 641922 300992 642022
rect 301116 641922 301216 642022
rect 301340 641922 301440 642022
rect 301564 641922 301664 642022
rect 301788 641922 301888 642022
rect 302012 641922 302112 642022
rect 302236 641922 302336 642022
rect 302460 641922 302560 642022
rect 302684 641922 302784 642022
rect 302908 641922 303008 642022
rect 303132 641922 303232 642022
rect 303356 641922 303456 642022
rect 303580 641922 303680 642022
rect 303804 641922 303904 642022
rect 304028 641922 304128 642022
rect 304252 641922 304352 642022
rect 304476 641922 304576 642022
rect 304700 641922 304800 642022
rect 304924 641922 305024 642022
rect 305148 641922 305248 642022
rect 305372 641922 305472 642022
rect 309346 641922 309446 642022
rect 309570 641922 309670 642022
rect 309794 641922 309894 642022
rect 310018 641922 310118 642022
rect 310242 641922 310342 642022
rect 310466 641922 310566 642022
rect 310690 641922 310790 642022
rect 310914 641922 311014 642022
rect 311138 641922 311238 642022
rect 311362 641922 311462 642022
rect 311586 641922 311686 642022
rect 311810 641922 311910 642022
rect 312034 641922 312134 642022
rect 312258 641922 312358 642022
rect 312482 641922 312582 642022
rect 312706 641922 312806 642022
rect 312930 641922 313030 642022
rect 313154 641922 313254 642022
rect 313378 641922 313478 642022
rect 313602 641922 313702 642022
rect 313826 641922 313926 642022
rect 314050 641922 314150 642022
rect 314274 641922 314374 642022
rect 314498 641922 314598 642022
rect 314722 641922 314822 642022
rect 314946 641922 315046 642022
rect 315170 641922 315270 642022
rect 315394 641922 315494 642022
rect 315618 641922 315718 642022
rect 315842 641922 315942 642022
rect 335616 641942 335716 642042
rect 335840 641942 335940 642042
rect 336064 641942 336164 642042
rect 336288 641942 336388 642042
rect 336512 641942 336612 642042
rect 336736 641942 336836 642042
rect 336960 641942 337060 642042
rect 337184 641942 337284 642042
rect 337408 641942 337508 642042
rect 337632 641942 337732 642042
rect 337856 641942 337956 642042
rect 338080 641942 338180 642042
rect 338304 641942 338404 642042
rect 338528 641942 338628 642042
rect 338752 641942 338852 642042
rect 338976 641942 339076 642042
rect 339200 641942 339300 642042
rect 339424 641942 339524 642042
rect 339648 641942 339748 642042
rect 339872 641942 339972 642042
rect 340096 641942 340196 642042
rect 340320 641942 340420 642042
rect 340544 641942 340644 642042
rect 340768 641942 340868 642042
rect 340992 641942 341092 642042
rect 341216 641942 341316 642042
rect 341440 641942 341540 642042
rect 341664 641942 341764 642042
rect 341888 641942 341988 642042
rect 342112 641942 342212 642042
rect 298876 641698 298976 641798
rect 299100 641698 299200 641798
rect 299324 641698 299424 641798
rect 299548 641698 299648 641798
rect 299772 641698 299872 641798
rect 299996 641698 300096 641798
rect 300220 641698 300320 641798
rect 300444 641698 300544 641798
rect 300668 641698 300768 641798
rect 300892 641698 300992 641798
rect 301116 641698 301216 641798
rect 301340 641698 301440 641798
rect 301564 641698 301664 641798
rect 301788 641698 301888 641798
rect 302012 641698 302112 641798
rect 302236 641698 302336 641798
rect 302460 641698 302560 641798
rect 302684 641698 302784 641798
rect 302908 641698 303008 641798
rect 303132 641698 303232 641798
rect 303356 641698 303456 641798
rect 303580 641698 303680 641798
rect 303804 641698 303904 641798
rect 304028 641698 304128 641798
rect 304252 641698 304352 641798
rect 304476 641698 304576 641798
rect 304700 641698 304800 641798
rect 304924 641698 305024 641798
rect 305148 641698 305248 641798
rect 305372 641698 305472 641798
rect 309346 641698 309446 641798
rect 309570 641698 309670 641798
rect 309794 641698 309894 641798
rect 310018 641698 310118 641798
rect 310242 641698 310342 641798
rect 310466 641698 310566 641798
rect 310690 641698 310790 641798
rect 310914 641698 311014 641798
rect 311138 641698 311238 641798
rect 311362 641698 311462 641798
rect 311586 641698 311686 641798
rect 311810 641698 311910 641798
rect 312034 641698 312134 641798
rect 312258 641698 312358 641798
rect 312482 641698 312582 641798
rect 312706 641698 312806 641798
rect 312930 641698 313030 641798
rect 313154 641698 313254 641798
rect 313378 641698 313478 641798
rect 313602 641698 313702 641798
rect 313826 641698 313926 641798
rect 314050 641698 314150 641798
rect 314274 641698 314374 641798
rect 314498 641698 314598 641798
rect 314722 641698 314822 641798
rect 314946 641698 315046 641798
rect 315170 641698 315270 641798
rect 315394 641698 315494 641798
rect 315618 641698 315718 641798
rect 315842 641698 315942 641798
rect 335616 641718 335716 641818
rect 335840 641718 335940 641818
rect 336064 641718 336164 641818
rect 336288 641718 336388 641818
rect 336512 641718 336612 641818
rect 336736 641718 336836 641818
rect 336960 641718 337060 641818
rect 337184 641718 337284 641818
rect 337408 641718 337508 641818
rect 337632 641718 337732 641818
rect 337856 641718 337956 641818
rect 338080 641718 338180 641818
rect 338304 641718 338404 641818
rect 338528 641718 338628 641818
rect 338752 641718 338852 641818
rect 338976 641718 339076 641818
rect 339200 641718 339300 641818
rect 339424 641718 339524 641818
rect 339648 641718 339748 641818
rect 339872 641718 339972 641818
rect 340096 641718 340196 641818
rect 340320 641718 340420 641818
rect 340544 641718 340644 641818
rect 340768 641718 340868 641818
rect 340992 641718 341092 641818
rect 341216 641718 341316 641818
rect 341440 641718 341540 641818
rect 341664 641718 341764 641818
rect 341888 641718 341988 641818
rect 342112 641718 342212 641818
rect 297850 637896 297950 637996
rect 298074 637896 298174 637996
rect 298298 637896 298398 637996
rect 298522 637896 298622 637996
rect 298746 637896 298846 637996
rect 342130 637896 342230 637996
rect 342354 637896 342454 637996
rect 342578 637896 342678 637996
rect 342802 637896 342902 637996
rect 343026 637896 343126 637996
rect 297850 637672 297950 637772
rect 298074 637672 298174 637772
rect 298298 637672 298398 637772
rect 298522 637672 298622 637772
rect 298746 637672 298846 637772
rect 342130 637672 342230 637772
rect 342354 637672 342454 637772
rect 342578 637672 342678 637772
rect 342802 637672 342902 637772
rect 343026 637672 343126 637772
rect 297850 637448 297950 637548
rect 298074 637448 298174 637548
rect 298298 637448 298398 637548
rect 298522 637448 298622 637548
rect 298746 637448 298846 637548
rect 342130 637448 342230 637548
rect 342354 637448 342454 637548
rect 342578 637448 342678 637548
rect 342802 637448 342902 637548
rect 343026 637448 343126 637548
rect 297850 637224 297950 637324
rect 298074 637224 298174 637324
rect 298298 637224 298398 637324
rect 298522 637224 298622 637324
rect 298746 637224 298846 637324
rect 342130 637224 342230 637324
rect 342354 637224 342454 637324
rect 342578 637224 342678 637324
rect 342802 637224 342902 637324
rect 343026 637224 343126 637324
rect 297850 637000 297950 637100
rect 298074 637000 298174 637100
rect 298298 637000 298398 637100
rect 298522 637000 298622 637100
rect 298746 637000 298846 637100
rect 342130 637000 342230 637100
rect 342354 637000 342454 637100
rect 342578 637000 342678 637100
rect 342802 637000 342902 637100
rect 343026 637000 343126 637100
rect 297850 636776 297950 636876
rect 298074 636776 298174 636876
rect 298298 636776 298398 636876
rect 298522 636776 298622 636876
rect 298746 636776 298846 636876
rect 342130 636776 342230 636876
rect 342354 636776 342454 636876
rect 342578 636776 342678 636876
rect 342802 636776 342902 636876
rect 343026 636776 343126 636876
rect 297850 636552 297950 636652
rect 298074 636552 298174 636652
rect 298298 636552 298398 636652
rect 298522 636552 298622 636652
rect 298746 636552 298846 636652
rect 342130 636552 342230 636652
rect 342354 636552 342454 636652
rect 342578 636552 342678 636652
rect 342802 636552 342902 636652
rect 343026 636552 343126 636652
rect 297850 636328 297950 636428
rect 298074 636328 298174 636428
rect 298298 636328 298398 636428
rect 298522 636328 298622 636428
rect 298746 636328 298846 636428
rect 342130 636328 342230 636428
rect 342354 636328 342454 636428
rect 342578 636328 342678 636428
rect 342802 636328 342902 636428
rect 343026 636328 343126 636428
rect 297850 636104 297950 636204
rect 298074 636104 298174 636204
rect 298298 636104 298398 636204
rect 298522 636104 298622 636204
rect 298746 636104 298846 636204
rect 342130 636104 342230 636204
rect 342354 636104 342454 636204
rect 342578 636104 342678 636204
rect 342802 636104 342902 636204
rect 343026 636104 343126 636204
rect 297850 635880 297950 635980
rect 298074 635880 298174 635980
rect 298298 635880 298398 635980
rect 298522 635880 298622 635980
rect 298746 635880 298846 635980
rect 342130 635880 342230 635980
rect 342354 635880 342454 635980
rect 342578 635880 342678 635980
rect 342802 635880 342902 635980
rect 343026 635880 343126 635980
rect 297850 635656 297950 635756
rect 298074 635656 298174 635756
rect 298298 635656 298398 635756
rect 298522 635656 298622 635756
rect 298746 635656 298846 635756
rect 342130 635656 342230 635756
rect 342354 635656 342454 635756
rect 342578 635656 342678 635756
rect 342802 635656 342902 635756
rect 343026 635656 343126 635756
rect 297850 635432 297950 635532
rect 298074 635432 298174 635532
rect 298298 635432 298398 635532
rect 298522 635432 298622 635532
rect 298746 635432 298846 635532
rect 342130 635432 342230 635532
rect 342354 635432 342454 635532
rect 342578 635432 342678 635532
rect 342802 635432 342902 635532
rect 343026 635432 343126 635532
rect 297850 635208 297950 635308
rect 298074 635208 298174 635308
rect 298298 635208 298398 635308
rect 298522 635208 298622 635308
rect 298746 635208 298846 635308
rect 342130 635208 342230 635308
rect 342354 635208 342454 635308
rect 342578 635208 342678 635308
rect 342802 635208 342902 635308
rect 343026 635208 343126 635308
rect 297850 634984 297950 635084
rect 298074 634984 298174 635084
rect 298298 634984 298398 635084
rect 298522 634984 298622 635084
rect 298746 634984 298846 635084
rect 342130 634984 342230 635084
rect 342354 634984 342454 635084
rect 342578 634984 342678 635084
rect 342802 634984 342902 635084
rect 343026 634984 343126 635084
rect 297850 634760 297950 634860
rect 298074 634760 298174 634860
rect 298298 634760 298398 634860
rect 298522 634760 298622 634860
rect 298746 634760 298846 634860
rect 342130 634760 342230 634860
rect 342354 634760 342454 634860
rect 342578 634760 342678 634860
rect 342802 634760 342902 634860
rect 343026 634760 343126 634860
rect 297850 634536 297950 634636
rect 298074 634536 298174 634636
rect 298298 634536 298398 634636
rect 298522 634536 298622 634636
rect 298746 634536 298846 634636
rect 342130 634536 342230 634636
rect 342354 634536 342454 634636
rect 342578 634536 342678 634636
rect 342802 634536 342902 634636
rect 343026 634536 343126 634636
rect 297850 634312 297950 634412
rect 298074 634312 298174 634412
rect 298298 634312 298398 634412
rect 298522 634312 298622 634412
rect 298746 634312 298846 634412
rect 342130 634312 342230 634412
rect 342354 634312 342454 634412
rect 342578 634312 342678 634412
rect 342802 634312 342902 634412
rect 343026 634312 343126 634412
rect 297850 634088 297950 634188
rect 298074 634088 298174 634188
rect 298298 634088 298398 634188
rect 298522 634088 298622 634188
rect 298746 634088 298846 634188
rect 342130 634088 342230 634188
rect 342354 634088 342454 634188
rect 342578 634088 342678 634188
rect 342802 634088 342902 634188
rect 343026 634088 343126 634188
rect 297850 633864 297950 633964
rect 298074 633864 298174 633964
rect 298298 633864 298398 633964
rect 298522 633864 298622 633964
rect 298746 633864 298846 633964
rect 342130 633864 342230 633964
rect 342354 633864 342454 633964
rect 342578 633864 342678 633964
rect 342802 633864 342902 633964
rect 343026 633864 343126 633964
rect 297850 633640 297950 633740
rect 298074 633640 298174 633740
rect 298298 633640 298398 633740
rect 298522 633640 298622 633740
rect 298746 633640 298846 633740
rect 342130 633640 342230 633740
rect 342354 633640 342454 633740
rect 342578 633640 342678 633740
rect 342802 633640 342902 633740
rect 343026 633640 343126 633740
rect 297850 633416 297950 633516
rect 298074 633416 298174 633516
rect 298298 633416 298398 633516
rect 298522 633416 298622 633516
rect 298746 633416 298846 633516
rect 342130 633416 342230 633516
rect 342354 633416 342454 633516
rect 342578 633416 342678 633516
rect 342802 633416 342902 633516
rect 343026 633416 343126 633516
rect 297850 633192 297950 633292
rect 298074 633192 298174 633292
rect 298298 633192 298398 633292
rect 298522 633192 298622 633292
rect 298746 633192 298846 633292
rect 342130 633192 342230 633292
rect 342354 633192 342454 633292
rect 342578 633192 342678 633292
rect 342802 633192 342902 633292
rect 343026 633192 343126 633292
rect 297850 632968 297950 633068
rect 298074 632968 298174 633068
rect 298298 632968 298398 633068
rect 298522 632968 298622 633068
rect 298746 632968 298846 633068
rect 342130 632968 342230 633068
rect 342354 632968 342454 633068
rect 342578 632968 342678 633068
rect 342802 632968 342902 633068
rect 343026 632968 343126 633068
rect 297850 632744 297950 632844
rect 298074 632744 298174 632844
rect 298298 632744 298398 632844
rect 298522 632744 298622 632844
rect 298746 632744 298846 632844
rect 342130 632744 342230 632844
rect 342354 632744 342454 632844
rect 342578 632744 342678 632844
rect 342802 632744 342902 632844
rect 343026 632744 343126 632844
rect 297850 632520 297950 632620
rect 298074 632520 298174 632620
rect 298298 632520 298398 632620
rect 298522 632520 298622 632620
rect 298746 632520 298846 632620
rect 342130 632520 342230 632620
rect 342354 632520 342454 632620
rect 342578 632520 342678 632620
rect 342802 632520 342902 632620
rect 343026 632520 343126 632620
rect 297850 632296 297950 632396
rect 298074 632296 298174 632396
rect 298298 632296 298398 632396
rect 298522 632296 298622 632396
rect 298746 632296 298846 632396
rect 342130 632296 342230 632396
rect 342354 632296 342454 632396
rect 342578 632296 342678 632396
rect 342802 632296 342902 632396
rect 343026 632296 343126 632396
rect 297850 632072 297950 632172
rect 298074 632072 298174 632172
rect 298298 632072 298398 632172
rect 298522 632072 298622 632172
rect 298746 632072 298846 632172
rect 342130 632072 342230 632172
rect 342354 632072 342454 632172
rect 342578 632072 342678 632172
rect 342802 632072 342902 632172
rect 343026 632072 343126 632172
rect 297850 631848 297950 631948
rect 298074 631848 298174 631948
rect 298298 631848 298398 631948
rect 298522 631848 298622 631948
rect 298746 631848 298846 631948
rect 342130 631848 342230 631948
rect 342354 631848 342454 631948
rect 342578 631848 342678 631948
rect 342802 631848 342902 631948
rect 343026 631848 343126 631948
rect 297850 631624 297950 631724
rect 298074 631624 298174 631724
rect 298298 631624 298398 631724
rect 298522 631624 298622 631724
rect 298746 631624 298846 631724
rect 342130 631624 342230 631724
rect 342354 631624 342454 631724
rect 342578 631624 342678 631724
rect 342802 631624 342902 631724
rect 343026 631624 343126 631724
rect 297850 631400 297950 631500
rect 298074 631400 298174 631500
rect 298298 631400 298398 631500
rect 298522 631400 298622 631500
rect 298746 631400 298846 631500
rect 342130 631400 342230 631500
rect 342354 631400 342454 631500
rect 342578 631400 342678 631500
rect 342802 631400 342902 631500
rect 343026 631400 343126 631500
rect 297850 624496 297950 624596
rect 298074 624496 298174 624596
rect 298298 624496 298398 624596
rect 298522 624496 298622 624596
rect 298746 624496 298846 624596
rect 297850 624272 297950 624372
rect 298074 624272 298174 624372
rect 298298 624272 298398 624372
rect 298522 624272 298622 624372
rect 298746 624272 298846 624372
rect 297850 624048 297950 624148
rect 298074 624048 298174 624148
rect 298298 624048 298398 624148
rect 298522 624048 298622 624148
rect 298746 624048 298846 624148
rect 297850 623824 297950 623924
rect 298074 623824 298174 623924
rect 298298 623824 298398 623924
rect 298522 623824 298622 623924
rect 298746 623824 298846 623924
rect 297850 623600 297950 623700
rect 298074 623600 298174 623700
rect 298298 623600 298398 623700
rect 298522 623600 298622 623700
rect 298746 623600 298846 623700
rect 297850 623376 297950 623476
rect 298074 623376 298174 623476
rect 298298 623376 298398 623476
rect 298522 623376 298622 623476
rect 298746 623376 298846 623476
rect 297850 623152 297950 623252
rect 298074 623152 298174 623252
rect 298298 623152 298398 623252
rect 298522 623152 298622 623252
rect 298746 623152 298846 623252
rect 297850 622928 297950 623028
rect 298074 622928 298174 623028
rect 298298 622928 298398 623028
rect 298522 622928 298622 623028
rect 298746 622928 298846 623028
rect 297850 622704 297950 622804
rect 298074 622704 298174 622804
rect 298298 622704 298398 622804
rect 298522 622704 298622 622804
rect 298746 622704 298846 622804
rect 297850 622480 297950 622580
rect 298074 622480 298174 622580
rect 298298 622480 298398 622580
rect 298522 622480 298622 622580
rect 298746 622480 298846 622580
rect 297850 622256 297950 622356
rect 298074 622256 298174 622356
rect 298298 622256 298398 622356
rect 298522 622256 298622 622356
rect 298746 622256 298846 622356
rect 297850 622032 297950 622132
rect 298074 622032 298174 622132
rect 298298 622032 298398 622132
rect 298522 622032 298622 622132
rect 298746 622032 298846 622132
rect 297850 621808 297950 621908
rect 298074 621808 298174 621908
rect 298298 621808 298398 621908
rect 298522 621808 298622 621908
rect 298746 621808 298846 621908
rect 297850 621584 297950 621684
rect 298074 621584 298174 621684
rect 298298 621584 298398 621684
rect 298522 621584 298622 621684
rect 298746 621584 298846 621684
rect 297850 621360 297950 621460
rect 298074 621360 298174 621460
rect 298298 621360 298398 621460
rect 298522 621360 298622 621460
rect 298746 621360 298846 621460
rect 297850 621136 297950 621236
rect 298074 621136 298174 621236
rect 298298 621136 298398 621236
rect 298522 621136 298622 621236
rect 298746 621136 298846 621236
rect 297850 620912 297950 621012
rect 298074 620912 298174 621012
rect 298298 620912 298398 621012
rect 298522 620912 298622 621012
rect 298746 620912 298846 621012
rect 297850 620688 297950 620788
rect 298074 620688 298174 620788
rect 298298 620688 298398 620788
rect 298522 620688 298622 620788
rect 298746 620688 298846 620788
rect 297850 620464 297950 620564
rect 298074 620464 298174 620564
rect 298298 620464 298398 620564
rect 298522 620464 298622 620564
rect 298746 620464 298846 620564
rect 297850 620240 297950 620340
rect 298074 620240 298174 620340
rect 298298 620240 298398 620340
rect 298522 620240 298622 620340
rect 298746 620240 298846 620340
rect 297850 620016 297950 620116
rect 298074 620016 298174 620116
rect 298298 620016 298398 620116
rect 298522 620016 298622 620116
rect 298746 620016 298846 620116
rect 297850 619792 297950 619892
rect 298074 619792 298174 619892
rect 298298 619792 298398 619892
rect 298522 619792 298622 619892
rect 298746 619792 298846 619892
rect 297850 619568 297950 619668
rect 298074 619568 298174 619668
rect 298298 619568 298398 619668
rect 298522 619568 298622 619668
rect 298746 619568 298846 619668
rect 297850 619344 297950 619444
rect 298074 619344 298174 619444
rect 298298 619344 298398 619444
rect 298522 619344 298622 619444
rect 298746 619344 298846 619444
rect 297850 619120 297950 619220
rect 298074 619120 298174 619220
rect 298298 619120 298398 619220
rect 298522 619120 298622 619220
rect 298746 619120 298846 619220
rect 297850 618896 297950 618996
rect 298074 618896 298174 618996
rect 298298 618896 298398 618996
rect 298522 618896 298622 618996
rect 298746 618896 298846 618996
rect 297850 618672 297950 618772
rect 298074 618672 298174 618772
rect 298298 618672 298398 618772
rect 298522 618672 298622 618772
rect 298746 618672 298846 618772
rect 297850 618448 297950 618548
rect 298074 618448 298174 618548
rect 298298 618448 298398 618548
rect 298522 618448 298622 618548
rect 298746 618448 298846 618548
rect 297850 618224 297950 618324
rect 298074 618224 298174 618324
rect 298298 618224 298398 618324
rect 298522 618224 298622 618324
rect 298746 618224 298846 618324
rect 297850 618000 297950 618100
rect 298074 618000 298174 618100
rect 298298 618000 298398 618100
rect 298522 618000 298622 618100
rect 298746 618000 298846 618100
rect 342130 624496 342230 624596
rect 342354 624496 342454 624596
rect 342578 624496 342678 624596
rect 342802 624496 342902 624596
rect 343026 624496 343126 624596
rect 342130 624272 342230 624372
rect 342354 624272 342454 624372
rect 342578 624272 342678 624372
rect 342802 624272 342902 624372
rect 343026 624272 343126 624372
rect 342130 624048 342230 624148
rect 342354 624048 342454 624148
rect 342578 624048 342678 624148
rect 342802 624048 342902 624148
rect 343026 624048 343126 624148
rect 342130 623824 342230 623924
rect 342354 623824 342454 623924
rect 342578 623824 342678 623924
rect 342802 623824 342902 623924
rect 343026 623824 343126 623924
rect 342130 623600 342230 623700
rect 342354 623600 342454 623700
rect 342578 623600 342678 623700
rect 342802 623600 342902 623700
rect 343026 623600 343126 623700
rect 342130 623376 342230 623476
rect 342354 623376 342454 623476
rect 342578 623376 342678 623476
rect 342802 623376 342902 623476
rect 343026 623376 343126 623476
rect 342130 623152 342230 623252
rect 342354 623152 342454 623252
rect 342578 623152 342678 623252
rect 342802 623152 342902 623252
rect 343026 623152 343126 623252
rect 342130 622928 342230 623028
rect 342354 622928 342454 623028
rect 342578 622928 342678 623028
rect 342802 622928 342902 623028
rect 343026 622928 343126 623028
rect 342130 622704 342230 622804
rect 342354 622704 342454 622804
rect 342578 622704 342678 622804
rect 342802 622704 342902 622804
rect 343026 622704 343126 622804
rect 342130 622480 342230 622580
rect 342354 622480 342454 622580
rect 342578 622480 342678 622580
rect 342802 622480 342902 622580
rect 343026 622480 343126 622580
rect 342130 622256 342230 622356
rect 342354 622256 342454 622356
rect 342578 622256 342678 622356
rect 342802 622256 342902 622356
rect 343026 622256 343126 622356
rect 342130 622032 342230 622132
rect 342354 622032 342454 622132
rect 342578 622032 342678 622132
rect 342802 622032 342902 622132
rect 343026 622032 343126 622132
rect 342130 621808 342230 621908
rect 342354 621808 342454 621908
rect 342578 621808 342678 621908
rect 342802 621808 342902 621908
rect 343026 621808 343126 621908
rect 342130 621584 342230 621684
rect 342354 621584 342454 621684
rect 342578 621584 342678 621684
rect 342802 621584 342902 621684
rect 343026 621584 343126 621684
rect 342130 621360 342230 621460
rect 342354 621360 342454 621460
rect 342578 621360 342678 621460
rect 342802 621360 342902 621460
rect 343026 621360 343126 621460
rect 342130 621136 342230 621236
rect 342354 621136 342454 621236
rect 342578 621136 342678 621236
rect 342802 621136 342902 621236
rect 343026 621136 343126 621236
rect 342130 620912 342230 621012
rect 342354 620912 342454 621012
rect 342578 620912 342678 621012
rect 342802 620912 342902 621012
rect 343026 620912 343126 621012
rect 342130 620688 342230 620788
rect 342354 620688 342454 620788
rect 342578 620688 342678 620788
rect 342802 620688 342902 620788
rect 343026 620688 343126 620788
rect 342130 620464 342230 620564
rect 342354 620464 342454 620564
rect 342578 620464 342678 620564
rect 342802 620464 342902 620564
rect 343026 620464 343126 620564
rect 342130 620240 342230 620340
rect 342354 620240 342454 620340
rect 342578 620240 342678 620340
rect 342802 620240 342902 620340
rect 343026 620240 343126 620340
rect 342130 620016 342230 620116
rect 342354 620016 342454 620116
rect 342578 620016 342678 620116
rect 342802 620016 342902 620116
rect 343026 620016 343126 620116
rect 342130 619792 342230 619892
rect 342354 619792 342454 619892
rect 342578 619792 342678 619892
rect 342802 619792 342902 619892
rect 343026 619792 343126 619892
rect 342130 619568 342230 619668
rect 342354 619568 342454 619668
rect 342578 619568 342678 619668
rect 342802 619568 342902 619668
rect 343026 619568 343126 619668
rect 342130 619344 342230 619444
rect 342354 619344 342454 619444
rect 342578 619344 342678 619444
rect 342802 619344 342902 619444
rect 343026 619344 343126 619444
rect 342130 619120 342230 619220
rect 342354 619120 342454 619220
rect 342578 619120 342678 619220
rect 342802 619120 342902 619220
rect 343026 619120 343126 619220
rect 342130 618896 342230 618996
rect 342354 618896 342454 618996
rect 342578 618896 342678 618996
rect 342802 618896 342902 618996
rect 343026 618896 343126 618996
rect 342130 618672 342230 618772
rect 342354 618672 342454 618772
rect 342578 618672 342678 618772
rect 342802 618672 342902 618772
rect 343026 618672 343126 618772
rect 342130 618448 342230 618548
rect 342354 618448 342454 618548
rect 342578 618448 342678 618548
rect 342802 618448 342902 618548
rect 343026 618448 343126 618548
rect 342130 618224 342230 618324
rect 342354 618224 342454 618324
rect 342578 618224 342678 618324
rect 342802 618224 342902 618324
rect 343026 618224 343126 618324
rect 342130 618000 342230 618100
rect 342354 618000 342454 618100
rect 342578 618000 342678 618100
rect 342802 618000 342902 618100
rect 343026 618000 343126 618100
rect 298876 615374 298976 615474
rect 299100 615374 299200 615474
rect 299324 615374 299424 615474
rect 299548 615374 299648 615474
rect 299772 615374 299872 615474
rect 299996 615374 300096 615474
rect 300220 615374 300320 615474
rect 300444 615374 300544 615474
rect 300668 615374 300768 615474
rect 300892 615374 300992 615474
rect 301116 615374 301216 615474
rect 301340 615374 301440 615474
rect 301564 615374 301664 615474
rect 301788 615374 301888 615474
rect 302012 615374 302112 615474
rect 302236 615374 302336 615474
rect 302460 615374 302560 615474
rect 302684 615374 302784 615474
rect 302908 615374 303008 615474
rect 303132 615374 303232 615474
rect 303356 615374 303456 615474
rect 303580 615374 303680 615474
rect 303804 615374 303904 615474
rect 304028 615374 304128 615474
rect 304252 615374 304352 615474
rect 304476 615374 304576 615474
rect 304700 615374 304800 615474
rect 304924 615374 305024 615474
rect 305148 615374 305248 615474
rect 305372 615374 305472 615474
rect 309346 615374 309446 615474
rect 309570 615374 309670 615474
rect 309794 615374 309894 615474
rect 310018 615374 310118 615474
rect 310242 615374 310342 615474
rect 310466 615374 310566 615474
rect 310690 615374 310790 615474
rect 310914 615374 311014 615474
rect 311138 615374 311238 615474
rect 311362 615374 311462 615474
rect 311586 615374 311686 615474
rect 311810 615374 311910 615474
rect 312034 615374 312134 615474
rect 312258 615374 312358 615474
rect 312482 615374 312582 615474
rect 312706 615374 312806 615474
rect 312930 615374 313030 615474
rect 313154 615374 313254 615474
rect 313378 615374 313478 615474
rect 313602 615374 313702 615474
rect 313826 615374 313926 615474
rect 314050 615374 314150 615474
rect 314274 615374 314374 615474
rect 314498 615374 314598 615474
rect 314722 615374 314822 615474
rect 314946 615374 315046 615474
rect 315170 615374 315270 615474
rect 315394 615374 315494 615474
rect 315618 615374 315718 615474
rect 315842 615374 315942 615474
rect 335616 615394 335716 615494
rect 335840 615394 335940 615494
rect 336064 615394 336164 615494
rect 336288 615394 336388 615494
rect 336512 615394 336612 615494
rect 336736 615394 336836 615494
rect 336960 615394 337060 615494
rect 337184 615394 337284 615494
rect 337408 615394 337508 615494
rect 337632 615394 337732 615494
rect 337856 615394 337956 615494
rect 338080 615394 338180 615494
rect 338304 615394 338404 615494
rect 338528 615394 338628 615494
rect 338752 615394 338852 615494
rect 338976 615394 339076 615494
rect 339200 615394 339300 615494
rect 339424 615394 339524 615494
rect 339648 615394 339748 615494
rect 339872 615394 339972 615494
rect 340096 615394 340196 615494
rect 340320 615394 340420 615494
rect 340544 615394 340644 615494
rect 340768 615394 340868 615494
rect 340992 615394 341092 615494
rect 341216 615394 341316 615494
rect 341440 615394 341540 615494
rect 341664 615394 341764 615494
rect 341888 615394 341988 615494
rect 342112 615394 342212 615494
rect 298876 615150 298976 615250
rect 299100 615150 299200 615250
rect 299324 615150 299424 615250
rect 299548 615150 299648 615250
rect 299772 615150 299872 615250
rect 299996 615150 300096 615250
rect 300220 615150 300320 615250
rect 300444 615150 300544 615250
rect 300668 615150 300768 615250
rect 300892 615150 300992 615250
rect 301116 615150 301216 615250
rect 301340 615150 301440 615250
rect 301564 615150 301664 615250
rect 301788 615150 301888 615250
rect 302012 615150 302112 615250
rect 302236 615150 302336 615250
rect 302460 615150 302560 615250
rect 302684 615150 302784 615250
rect 302908 615150 303008 615250
rect 303132 615150 303232 615250
rect 303356 615150 303456 615250
rect 303580 615150 303680 615250
rect 303804 615150 303904 615250
rect 304028 615150 304128 615250
rect 304252 615150 304352 615250
rect 304476 615150 304576 615250
rect 304700 615150 304800 615250
rect 304924 615150 305024 615250
rect 305148 615150 305248 615250
rect 305372 615150 305472 615250
rect 309346 615150 309446 615250
rect 309570 615150 309670 615250
rect 309794 615150 309894 615250
rect 310018 615150 310118 615250
rect 310242 615150 310342 615250
rect 310466 615150 310566 615250
rect 310690 615150 310790 615250
rect 310914 615150 311014 615250
rect 311138 615150 311238 615250
rect 311362 615150 311462 615250
rect 311586 615150 311686 615250
rect 311810 615150 311910 615250
rect 312034 615150 312134 615250
rect 312258 615150 312358 615250
rect 312482 615150 312582 615250
rect 312706 615150 312806 615250
rect 312930 615150 313030 615250
rect 313154 615150 313254 615250
rect 313378 615150 313478 615250
rect 313602 615150 313702 615250
rect 313826 615150 313926 615250
rect 314050 615150 314150 615250
rect 314274 615150 314374 615250
rect 314498 615150 314598 615250
rect 314722 615150 314822 615250
rect 314946 615150 315046 615250
rect 315170 615150 315270 615250
rect 315394 615150 315494 615250
rect 315618 615150 315718 615250
rect 315842 615150 315942 615250
rect 335616 615170 335716 615270
rect 335840 615170 335940 615270
rect 336064 615170 336164 615270
rect 336288 615170 336388 615270
rect 336512 615170 336612 615270
rect 336736 615170 336836 615270
rect 336960 615170 337060 615270
rect 337184 615170 337284 615270
rect 337408 615170 337508 615270
rect 337632 615170 337732 615270
rect 337856 615170 337956 615270
rect 338080 615170 338180 615270
rect 338304 615170 338404 615270
rect 338528 615170 338628 615270
rect 338752 615170 338852 615270
rect 338976 615170 339076 615270
rect 339200 615170 339300 615270
rect 339424 615170 339524 615270
rect 339648 615170 339748 615270
rect 339872 615170 339972 615270
rect 340096 615170 340196 615270
rect 340320 615170 340420 615270
rect 340544 615170 340644 615270
rect 340768 615170 340868 615270
rect 340992 615170 341092 615270
rect 341216 615170 341316 615270
rect 341440 615170 341540 615270
rect 341664 615170 341764 615270
rect 341888 615170 341988 615270
rect 342112 615170 342212 615270
rect 298876 614926 298976 615026
rect 299100 614926 299200 615026
rect 299324 614926 299424 615026
rect 299548 614926 299648 615026
rect 299772 614926 299872 615026
rect 299996 614926 300096 615026
rect 300220 614926 300320 615026
rect 300444 614926 300544 615026
rect 300668 614926 300768 615026
rect 300892 614926 300992 615026
rect 301116 614926 301216 615026
rect 301340 614926 301440 615026
rect 301564 614926 301664 615026
rect 301788 614926 301888 615026
rect 302012 614926 302112 615026
rect 302236 614926 302336 615026
rect 302460 614926 302560 615026
rect 302684 614926 302784 615026
rect 302908 614926 303008 615026
rect 303132 614926 303232 615026
rect 303356 614926 303456 615026
rect 303580 614926 303680 615026
rect 303804 614926 303904 615026
rect 304028 614926 304128 615026
rect 304252 614926 304352 615026
rect 304476 614926 304576 615026
rect 304700 614926 304800 615026
rect 304924 614926 305024 615026
rect 305148 614926 305248 615026
rect 305372 614926 305472 615026
rect 309346 614926 309446 615026
rect 309570 614926 309670 615026
rect 309794 614926 309894 615026
rect 310018 614926 310118 615026
rect 310242 614926 310342 615026
rect 310466 614926 310566 615026
rect 310690 614926 310790 615026
rect 310914 614926 311014 615026
rect 311138 614926 311238 615026
rect 311362 614926 311462 615026
rect 311586 614926 311686 615026
rect 311810 614926 311910 615026
rect 312034 614926 312134 615026
rect 312258 614926 312358 615026
rect 312482 614926 312582 615026
rect 312706 614926 312806 615026
rect 312930 614926 313030 615026
rect 313154 614926 313254 615026
rect 313378 614926 313478 615026
rect 313602 614926 313702 615026
rect 313826 614926 313926 615026
rect 314050 614926 314150 615026
rect 314274 614926 314374 615026
rect 314498 614926 314598 615026
rect 314722 614926 314822 615026
rect 314946 614926 315046 615026
rect 315170 614926 315270 615026
rect 315394 614926 315494 615026
rect 315618 614926 315718 615026
rect 315842 614926 315942 615026
rect 335616 614946 335716 615046
rect 335840 614946 335940 615046
rect 336064 614946 336164 615046
rect 336288 614946 336388 615046
rect 336512 614946 336612 615046
rect 336736 614946 336836 615046
rect 336960 614946 337060 615046
rect 337184 614946 337284 615046
rect 337408 614946 337508 615046
rect 337632 614946 337732 615046
rect 337856 614946 337956 615046
rect 338080 614946 338180 615046
rect 338304 614946 338404 615046
rect 338528 614946 338628 615046
rect 338752 614946 338852 615046
rect 338976 614946 339076 615046
rect 339200 614946 339300 615046
rect 339424 614946 339524 615046
rect 339648 614946 339748 615046
rect 339872 614946 339972 615046
rect 340096 614946 340196 615046
rect 340320 614946 340420 615046
rect 340544 614946 340644 615046
rect 340768 614946 340868 615046
rect 340992 614946 341092 615046
rect 341216 614946 341316 615046
rect 341440 614946 341540 615046
rect 341664 614946 341764 615046
rect 341888 614946 341988 615046
rect 342112 614946 342212 615046
rect 298876 614702 298976 614802
rect 299100 614702 299200 614802
rect 299324 614702 299424 614802
rect 299548 614702 299648 614802
rect 299772 614702 299872 614802
rect 299996 614702 300096 614802
rect 300220 614702 300320 614802
rect 300444 614702 300544 614802
rect 300668 614702 300768 614802
rect 300892 614702 300992 614802
rect 301116 614702 301216 614802
rect 301340 614702 301440 614802
rect 301564 614702 301664 614802
rect 301788 614702 301888 614802
rect 302012 614702 302112 614802
rect 302236 614702 302336 614802
rect 302460 614702 302560 614802
rect 302684 614702 302784 614802
rect 302908 614702 303008 614802
rect 303132 614702 303232 614802
rect 303356 614702 303456 614802
rect 303580 614702 303680 614802
rect 303804 614702 303904 614802
rect 304028 614702 304128 614802
rect 304252 614702 304352 614802
rect 304476 614702 304576 614802
rect 304700 614702 304800 614802
rect 304924 614702 305024 614802
rect 305148 614702 305248 614802
rect 305372 614702 305472 614802
rect 309346 614702 309446 614802
rect 309570 614702 309670 614802
rect 309794 614702 309894 614802
rect 310018 614702 310118 614802
rect 310242 614702 310342 614802
rect 310466 614702 310566 614802
rect 310690 614702 310790 614802
rect 310914 614702 311014 614802
rect 311138 614702 311238 614802
rect 311362 614702 311462 614802
rect 311586 614702 311686 614802
rect 311810 614702 311910 614802
rect 312034 614702 312134 614802
rect 312258 614702 312358 614802
rect 312482 614702 312582 614802
rect 312706 614702 312806 614802
rect 312930 614702 313030 614802
rect 313154 614702 313254 614802
rect 313378 614702 313478 614802
rect 313602 614702 313702 614802
rect 313826 614702 313926 614802
rect 314050 614702 314150 614802
rect 314274 614702 314374 614802
rect 314498 614702 314598 614802
rect 314722 614702 314822 614802
rect 314946 614702 315046 614802
rect 315170 614702 315270 614802
rect 315394 614702 315494 614802
rect 315618 614702 315718 614802
rect 315842 614702 315942 614802
rect 335616 614722 335716 614822
rect 335840 614722 335940 614822
rect 336064 614722 336164 614822
rect 336288 614722 336388 614822
rect 336512 614722 336612 614822
rect 336736 614722 336836 614822
rect 336960 614722 337060 614822
rect 337184 614722 337284 614822
rect 337408 614722 337508 614822
rect 337632 614722 337732 614822
rect 337856 614722 337956 614822
rect 338080 614722 338180 614822
rect 338304 614722 338404 614822
rect 338528 614722 338628 614822
rect 338752 614722 338852 614822
rect 338976 614722 339076 614822
rect 339200 614722 339300 614822
rect 339424 614722 339524 614822
rect 339648 614722 339748 614822
rect 339872 614722 339972 614822
rect 340096 614722 340196 614822
rect 340320 614722 340420 614822
rect 340544 614722 340644 614822
rect 340768 614722 340868 614822
rect 340992 614722 341092 614822
rect 341216 614722 341316 614822
rect 341440 614722 341540 614822
rect 341664 614722 341764 614822
rect 341888 614722 341988 614822
rect 342112 614722 342212 614822
rect 298876 614478 298976 614578
rect 299100 614478 299200 614578
rect 299324 614478 299424 614578
rect 299548 614478 299648 614578
rect 299772 614478 299872 614578
rect 299996 614478 300096 614578
rect 300220 614478 300320 614578
rect 300444 614478 300544 614578
rect 300668 614478 300768 614578
rect 300892 614478 300992 614578
rect 301116 614478 301216 614578
rect 301340 614478 301440 614578
rect 301564 614478 301664 614578
rect 301788 614478 301888 614578
rect 302012 614478 302112 614578
rect 302236 614478 302336 614578
rect 302460 614478 302560 614578
rect 302684 614478 302784 614578
rect 302908 614478 303008 614578
rect 303132 614478 303232 614578
rect 303356 614478 303456 614578
rect 303580 614478 303680 614578
rect 303804 614478 303904 614578
rect 304028 614478 304128 614578
rect 304252 614478 304352 614578
rect 304476 614478 304576 614578
rect 304700 614478 304800 614578
rect 304924 614478 305024 614578
rect 305148 614478 305248 614578
rect 305372 614478 305472 614578
rect 309346 614478 309446 614578
rect 309570 614478 309670 614578
rect 309794 614478 309894 614578
rect 310018 614478 310118 614578
rect 310242 614478 310342 614578
rect 310466 614478 310566 614578
rect 310690 614478 310790 614578
rect 310914 614478 311014 614578
rect 311138 614478 311238 614578
rect 311362 614478 311462 614578
rect 311586 614478 311686 614578
rect 311810 614478 311910 614578
rect 312034 614478 312134 614578
rect 312258 614478 312358 614578
rect 312482 614478 312582 614578
rect 312706 614478 312806 614578
rect 312930 614478 313030 614578
rect 313154 614478 313254 614578
rect 313378 614478 313478 614578
rect 313602 614478 313702 614578
rect 313826 614478 313926 614578
rect 314050 614478 314150 614578
rect 314274 614478 314374 614578
rect 314498 614478 314598 614578
rect 314722 614478 314822 614578
rect 314946 614478 315046 614578
rect 315170 614478 315270 614578
rect 315394 614478 315494 614578
rect 315618 614478 315718 614578
rect 315842 614478 315942 614578
rect 335616 614498 335716 614598
rect 335840 614498 335940 614598
rect 336064 614498 336164 614598
rect 336288 614498 336388 614598
rect 336512 614498 336612 614598
rect 336736 614498 336836 614598
rect 336960 614498 337060 614598
rect 337184 614498 337284 614598
rect 337408 614498 337508 614598
rect 337632 614498 337732 614598
rect 337856 614498 337956 614598
rect 338080 614498 338180 614598
rect 338304 614498 338404 614598
rect 338528 614498 338628 614598
rect 338752 614498 338852 614598
rect 338976 614498 339076 614598
rect 339200 614498 339300 614598
rect 339424 614498 339524 614598
rect 339648 614498 339748 614598
rect 339872 614498 339972 614598
rect 340096 614498 340196 614598
rect 340320 614498 340420 614598
rect 340544 614498 340644 614598
rect 340768 614498 340868 614598
rect 340992 614498 341092 614598
rect 341216 614498 341316 614598
rect 341440 614498 341540 614598
rect 341664 614498 341764 614598
rect 341888 614498 341988 614598
rect 342112 614498 342212 614598
<< metal1 >>
rect 298836 642694 305496 642724
rect 298836 642594 298876 642694
rect 298976 642594 299100 642694
rect 299200 642594 299324 642694
rect 299424 642594 299548 642694
rect 299648 642594 299772 642694
rect 299872 642594 299996 642694
rect 300096 642594 300220 642694
rect 300320 642594 300444 642694
rect 300544 642594 300668 642694
rect 300768 642594 300892 642694
rect 300992 642594 301116 642694
rect 301216 642594 301340 642694
rect 301440 642594 301564 642694
rect 301664 642594 301788 642694
rect 301888 642594 302012 642694
rect 302112 642594 302236 642694
rect 302336 642594 302460 642694
rect 302560 642594 302684 642694
rect 302784 642594 302908 642694
rect 303008 642594 303132 642694
rect 303232 642594 303356 642694
rect 303456 642594 303580 642694
rect 303680 642594 303804 642694
rect 303904 642594 304028 642694
rect 304128 642594 304252 642694
rect 304352 642594 304476 642694
rect 304576 642594 304700 642694
rect 304800 642594 304924 642694
rect 305024 642594 305148 642694
rect 305248 642594 305372 642694
rect 305472 642594 305496 642694
rect 298836 642470 305496 642594
rect 298836 642370 298876 642470
rect 298976 642370 299100 642470
rect 299200 642370 299324 642470
rect 299424 642370 299548 642470
rect 299648 642370 299772 642470
rect 299872 642370 299996 642470
rect 300096 642370 300220 642470
rect 300320 642370 300444 642470
rect 300544 642370 300668 642470
rect 300768 642370 300892 642470
rect 300992 642370 301116 642470
rect 301216 642370 301340 642470
rect 301440 642370 301564 642470
rect 301664 642370 301788 642470
rect 301888 642370 302012 642470
rect 302112 642370 302236 642470
rect 302336 642370 302460 642470
rect 302560 642370 302684 642470
rect 302784 642370 302908 642470
rect 303008 642370 303132 642470
rect 303232 642370 303356 642470
rect 303456 642370 303580 642470
rect 303680 642370 303804 642470
rect 303904 642370 304028 642470
rect 304128 642370 304252 642470
rect 304352 642370 304476 642470
rect 304576 642370 304700 642470
rect 304800 642370 304924 642470
rect 305024 642370 305148 642470
rect 305248 642370 305372 642470
rect 305472 642370 305496 642470
rect 298836 642246 305496 642370
rect 298836 642146 298876 642246
rect 298976 642146 299100 642246
rect 299200 642146 299324 642246
rect 299424 642146 299548 642246
rect 299648 642146 299772 642246
rect 299872 642146 299996 642246
rect 300096 642146 300220 642246
rect 300320 642146 300444 642246
rect 300544 642146 300668 642246
rect 300768 642146 300892 642246
rect 300992 642146 301116 642246
rect 301216 642146 301340 642246
rect 301440 642146 301564 642246
rect 301664 642146 301788 642246
rect 301888 642146 302012 642246
rect 302112 642146 302236 642246
rect 302336 642146 302460 642246
rect 302560 642146 302684 642246
rect 302784 642146 302908 642246
rect 303008 642146 303132 642246
rect 303232 642146 303356 642246
rect 303456 642146 303580 642246
rect 303680 642146 303804 642246
rect 303904 642146 304028 642246
rect 304128 642146 304252 642246
rect 304352 642146 304476 642246
rect 304576 642146 304700 642246
rect 304800 642146 304924 642246
rect 305024 642146 305148 642246
rect 305248 642146 305372 642246
rect 305472 642146 305496 642246
rect 298836 642022 305496 642146
rect 298836 641922 298876 642022
rect 298976 641922 299100 642022
rect 299200 641922 299324 642022
rect 299424 641922 299548 642022
rect 299648 641922 299772 642022
rect 299872 641922 299996 642022
rect 300096 641922 300220 642022
rect 300320 641922 300444 642022
rect 300544 641922 300668 642022
rect 300768 641922 300892 642022
rect 300992 641922 301116 642022
rect 301216 641922 301340 642022
rect 301440 641922 301564 642022
rect 301664 641922 301788 642022
rect 301888 641922 302012 642022
rect 302112 641922 302236 642022
rect 302336 641922 302460 642022
rect 302560 641922 302684 642022
rect 302784 641922 302908 642022
rect 303008 641922 303132 642022
rect 303232 641922 303356 642022
rect 303456 641922 303580 642022
rect 303680 641922 303804 642022
rect 303904 641922 304028 642022
rect 304128 641922 304252 642022
rect 304352 641922 304476 642022
rect 304576 641922 304700 642022
rect 304800 641922 304924 642022
rect 305024 641922 305148 642022
rect 305248 641922 305372 642022
rect 305472 641922 305496 642022
rect 298836 641798 305496 641922
rect 298836 641698 298876 641798
rect 298976 641698 299100 641798
rect 299200 641698 299324 641798
rect 299424 641698 299548 641798
rect 299648 641698 299772 641798
rect 299872 641698 299996 641798
rect 300096 641698 300220 641798
rect 300320 641698 300444 641798
rect 300544 641698 300668 641798
rect 300768 641698 300892 641798
rect 300992 641698 301116 641798
rect 301216 641698 301340 641798
rect 301440 641698 301564 641798
rect 301664 641698 301788 641798
rect 301888 641698 302012 641798
rect 302112 641698 302236 641798
rect 302336 641698 302460 641798
rect 302560 641698 302684 641798
rect 302784 641698 302908 641798
rect 303008 641698 303132 641798
rect 303232 641698 303356 641798
rect 303456 641698 303580 641798
rect 303680 641698 303804 641798
rect 303904 641698 304028 641798
rect 304128 641698 304252 641798
rect 304352 641698 304476 641798
rect 304576 641698 304700 641798
rect 304800 641698 304924 641798
rect 305024 641698 305148 641798
rect 305248 641698 305372 641798
rect 305472 641698 305496 641798
rect 298836 641664 305496 641698
rect 309306 642694 315966 642724
rect 309306 642594 309346 642694
rect 309446 642594 309570 642694
rect 309670 642594 309794 642694
rect 309894 642594 310018 642694
rect 310118 642594 310242 642694
rect 310342 642594 310466 642694
rect 310566 642594 310690 642694
rect 310790 642594 310914 642694
rect 311014 642594 311138 642694
rect 311238 642594 311362 642694
rect 311462 642594 311586 642694
rect 311686 642594 311810 642694
rect 311910 642594 312034 642694
rect 312134 642594 312258 642694
rect 312358 642594 312482 642694
rect 312582 642594 312706 642694
rect 312806 642594 312930 642694
rect 313030 642594 313154 642694
rect 313254 642594 313378 642694
rect 313478 642594 313602 642694
rect 313702 642594 313826 642694
rect 313926 642594 314050 642694
rect 314150 642594 314274 642694
rect 314374 642594 314498 642694
rect 314598 642594 314722 642694
rect 314822 642594 314946 642694
rect 315046 642594 315170 642694
rect 315270 642594 315394 642694
rect 315494 642594 315618 642694
rect 315718 642594 315842 642694
rect 315942 642594 315966 642694
rect 309306 642470 315966 642594
rect 309306 642370 309346 642470
rect 309446 642370 309570 642470
rect 309670 642370 309794 642470
rect 309894 642370 310018 642470
rect 310118 642370 310242 642470
rect 310342 642370 310466 642470
rect 310566 642370 310690 642470
rect 310790 642370 310914 642470
rect 311014 642370 311138 642470
rect 311238 642370 311362 642470
rect 311462 642370 311586 642470
rect 311686 642370 311810 642470
rect 311910 642370 312034 642470
rect 312134 642370 312258 642470
rect 312358 642370 312482 642470
rect 312582 642370 312706 642470
rect 312806 642370 312930 642470
rect 313030 642370 313154 642470
rect 313254 642370 313378 642470
rect 313478 642370 313602 642470
rect 313702 642370 313826 642470
rect 313926 642370 314050 642470
rect 314150 642370 314274 642470
rect 314374 642370 314498 642470
rect 314598 642370 314722 642470
rect 314822 642370 314946 642470
rect 315046 642370 315170 642470
rect 315270 642370 315394 642470
rect 315494 642370 315618 642470
rect 315718 642370 315842 642470
rect 315942 642370 315966 642470
rect 309306 642246 315966 642370
rect 309306 642146 309346 642246
rect 309446 642146 309570 642246
rect 309670 642146 309794 642246
rect 309894 642146 310018 642246
rect 310118 642146 310242 642246
rect 310342 642146 310466 642246
rect 310566 642146 310690 642246
rect 310790 642146 310914 642246
rect 311014 642146 311138 642246
rect 311238 642146 311362 642246
rect 311462 642146 311586 642246
rect 311686 642146 311810 642246
rect 311910 642146 312034 642246
rect 312134 642146 312258 642246
rect 312358 642146 312482 642246
rect 312582 642146 312706 642246
rect 312806 642146 312930 642246
rect 313030 642146 313154 642246
rect 313254 642146 313378 642246
rect 313478 642146 313602 642246
rect 313702 642146 313826 642246
rect 313926 642146 314050 642246
rect 314150 642146 314274 642246
rect 314374 642146 314498 642246
rect 314598 642146 314722 642246
rect 314822 642146 314946 642246
rect 315046 642146 315170 642246
rect 315270 642146 315394 642246
rect 315494 642146 315618 642246
rect 315718 642146 315842 642246
rect 315942 642146 315966 642246
rect 309306 642022 315966 642146
rect 309306 641922 309346 642022
rect 309446 641922 309570 642022
rect 309670 641922 309794 642022
rect 309894 641922 310018 642022
rect 310118 641922 310242 642022
rect 310342 641922 310466 642022
rect 310566 641922 310690 642022
rect 310790 641922 310914 642022
rect 311014 641922 311138 642022
rect 311238 641922 311362 642022
rect 311462 641922 311586 642022
rect 311686 641922 311810 642022
rect 311910 641922 312034 642022
rect 312134 641922 312258 642022
rect 312358 641922 312482 642022
rect 312582 641922 312706 642022
rect 312806 641922 312930 642022
rect 313030 641922 313154 642022
rect 313254 641922 313378 642022
rect 313478 641922 313602 642022
rect 313702 641922 313826 642022
rect 313926 641922 314050 642022
rect 314150 641922 314274 642022
rect 314374 641922 314498 642022
rect 314598 641922 314722 642022
rect 314822 641922 314946 642022
rect 315046 641922 315170 642022
rect 315270 641922 315394 642022
rect 315494 641922 315618 642022
rect 315718 641922 315842 642022
rect 315942 641922 315966 642022
rect 309306 641798 315966 641922
rect 309306 641698 309346 641798
rect 309446 641698 309570 641798
rect 309670 641698 309794 641798
rect 309894 641698 310018 641798
rect 310118 641698 310242 641798
rect 310342 641698 310466 641798
rect 310566 641698 310690 641798
rect 310790 641698 310914 641798
rect 311014 641698 311138 641798
rect 311238 641698 311362 641798
rect 311462 641698 311586 641798
rect 311686 641698 311810 641798
rect 311910 641698 312034 641798
rect 312134 641698 312258 641798
rect 312358 641698 312482 641798
rect 312582 641698 312706 641798
rect 312806 641698 312930 641798
rect 313030 641698 313154 641798
rect 313254 641698 313378 641798
rect 313478 641698 313602 641798
rect 313702 641698 313826 641798
rect 313926 641698 314050 641798
rect 314150 641698 314274 641798
rect 314374 641698 314498 641798
rect 314598 641698 314722 641798
rect 314822 641698 314946 641798
rect 315046 641698 315170 641798
rect 315270 641698 315394 641798
rect 315494 641698 315618 641798
rect 315718 641698 315842 641798
rect 315942 641698 315966 641798
rect 309306 641664 315966 641698
rect 335576 642714 342236 642744
rect 335576 642614 335616 642714
rect 335716 642614 335840 642714
rect 335940 642614 336064 642714
rect 336164 642614 336288 642714
rect 336388 642614 336512 642714
rect 336612 642614 336736 642714
rect 336836 642614 336960 642714
rect 337060 642614 337184 642714
rect 337284 642614 337408 642714
rect 337508 642614 337632 642714
rect 337732 642614 337856 642714
rect 337956 642614 338080 642714
rect 338180 642614 338304 642714
rect 338404 642614 338528 642714
rect 338628 642614 338752 642714
rect 338852 642614 338976 642714
rect 339076 642614 339200 642714
rect 339300 642614 339424 642714
rect 339524 642614 339648 642714
rect 339748 642614 339872 642714
rect 339972 642614 340096 642714
rect 340196 642614 340320 642714
rect 340420 642614 340544 642714
rect 340644 642614 340768 642714
rect 340868 642614 340992 642714
rect 341092 642614 341216 642714
rect 341316 642614 341440 642714
rect 341540 642614 341664 642714
rect 341764 642614 341888 642714
rect 341988 642614 342112 642714
rect 342212 642614 342236 642714
rect 335576 642490 342236 642614
rect 335576 642390 335616 642490
rect 335716 642390 335840 642490
rect 335940 642390 336064 642490
rect 336164 642390 336288 642490
rect 336388 642390 336512 642490
rect 336612 642390 336736 642490
rect 336836 642390 336960 642490
rect 337060 642390 337184 642490
rect 337284 642390 337408 642490
rect 337508 642390 337632 642490
rect 337732 642390 337856 642490
rect 337956 642390 338080 642490
rect 338180 642390 338304 642490
rect 338404 642390 338528 642490
rect 338628 642390 338752 642490
rect 338852 642390 338976 642490
rect 339076 642390 339200 642490
rect 339300 642390 339424 642490
rect 339524 642390 339648 642490
rect 339748 642390 339872 642490
rect 339972 642390 340096 642490
rect 340196 642390 340320 642490
rect 340420 642390 340544 642490
rect 340644 642390 340768 642490
rect 340868 642390 340992 642490
rect 341092 642390 341216 642490
rect 341316 642390 341440 642490
rect 341540 642390 341664 642490
rect 341764 642390 341888 642490
rect 341988 642390 342112 642490
rect 342212 642390 342236 642490
rect 335576 642266 342236 642390
rect 335576 642166 335616 642266
rect 335716 642166 335840 642266
rect 335940 642166 336064 642266
rect 336164 642166 336288 642266
rect 336388 642166 336512 642266
rect 336612 642166 336736 642266
rect 336836 642166 336960 642266
rect 337060 642166 337184 642266
rect 337284 642166 337408 642266
rect 337508 642166 337632 642266
rect 337732 642166 337856 642266
rect 337956 642166 338080 642266
rect 338180 642166 338304 642266
rect 338404 642166 338528 642266
rect 338628 642166 338752 642266
rect 338852 642166 338976 642266
rect 339076 642166 339200 642266
rect 339300 642166 339424 642266
rect 339524 642166 339648 642266
rect 339748 642166 339872 642266
rect 339972 642166 340096 642266
rect 340196 642166 340320 642266
rect 340420 642166 340544 642266
rect 340644 642166 340768 642266
rect 340868 642166 340992 642266
rect 341092 642166 341216 642266
rect 341316 642166 341440 642266
rect 341540 642166 341664 642266
rect 341764 642166 341888 642266
rect 341988 642166 342112 642266
rect 342212 642166 342236 642266
rect 335576 642042 342236 642166
rect 335576 641942 335616 642042
rect 335716 641942 335840 642042
rect 335940 641942 336064 642042
rect 336164 641942 336288 642042
rect 336388 641942 336512 642042
rect 336612 641942 336736 642042
rect 336836 641942 336960 642042
rect 337060 641942 337184 642042
rect 337284 641942 337408 642042
rect 337508 641942 337632 642042
rect 337732 641942 337856 642042
rect 337956 641942 338080 642042
rect 338180 641942 338304 642042
rect 338404 641942 338528 642042
rect 338628 641942 338752 642042
rect 338852 641942 338976 642042
rect 339076 641942 339200 642042
rect 339300 641942 339424 642042
rect 339524 641942 339648 642042
rect 339748 641942 339872 642042
rect 339972 641942 340096 642042
rect 340196 641942 340320 642042
rect 340420 641942 340544 642042
rect 340644 641942 340768 642042
rect 340868 641942 340992 642042
rect 341092 641942 341216 642042
rect 341316 641942 341440 642042
rect 341540 641942 341664 642042
rect 341764 641942 341888 642042
rect 341988 641942 342112 642042
rect 342212 641942 342236 642042
rect 335576 641818 342236 641942
rect 335576 641718 335616 641818
rect 335716 641718 335840 641818
rect 335940 641718 336064 641818
rect 336164 641718 336288 641818
rect 336388 641718 336512 641818
rect 336612 641718 336736 641818
rect 336836 641718 336960 641818
rect 337060 641718 337184 641818
rect 337284 641718 337408 641818
rect 337508 641718 337632 641818
rect 337732 641718 337856 641818
rect 337956 641718 338080 641818
rect 338180 641718 338304 641818
rect 338404 641718 338528 641818
rect 338628 641718 338752 641818
rect 338852 641718 338976 641818
rect 339076 641718 339200 641818
rect 339300 641718 339424 641818
rect 339524 641718 339648 641818
rect 339748 641718 339872 641818
rect 339972 641718 340096 641818
rect 340196 641718 340320 641818
rect 340420 641718 340544 641818
rect 340644 641718 340768 641818
rect 340868 641718 340992 641818
rect 341092 641718 341216 641818
rect 341316 641718 341440 641818
rect 341540 641718 341664 641818
rect 341764 641718 341888 641818
rect 341988 641718 342112 641818
rect 342212 641718 342236 641818
rect 335576 641684 342236 641718
rect 297820 637996 298880 638020
rect 297820 637896 297850 637996
rect 297950 637896 298074 637996
rect 298174 637896 298298 637996
rect 298398 637896 298522 637996
rect 298622 637896 298746 637996
rect 298846 637896 298880 637996
rect 297820 637772 298880 637896
rect 297820 637672 297850 637772
rect 297950 637672 298074 637772
rect 298174 637672 298298 637772
rect 298398 637672 298522 637772
rect 298622 637672 298746 637772
rect 298846 637672 298880 637772
rect 297820 637548 298880 637672
rect 297820 637448 297850 637548
rect 297950 637448 298074 637548
rect 298174 637448 298298 637548
rect 298398 637448 298522 637548
rect 298622 637448 298746 637548
rect 298846 637448 298880 637548
rect 297820 637324 298880 637448
rect 297820 637224 297850 637324
rect 297950 637224 298074 637324
rect 298174 637224 298298 637324
rect 298398 637224 298522 637324
rect 298622 637224 298746 637324
rect 298846 637224 298880 637324
rect 297820 637100 298880 637224
rect 297820 637000 297850 637100
rect 297950 637000 298074 637100
rect 298174 637000 298298 637100
rect 298398 637000 298522 637100
rect 298622 637000 298746 637100
rect 298846 637000 298880 637100
rect 297820 636876 298880 637000
rect 297820 636776 297850 636876
rect 297950 636776 298074 636876
rect 298174 636776 298298 636876
rect 298398 636776 298522 636876
rect 298622 636776 298746 636876
rect 298846 636776 298880 636876
rect 297820 636652 298880 636776
rect 297820 636552 297850 636652
rect 297950 636552 298074 636652
rect 298174 636552 298298 636652
rect 298398 636552 298522 636652
rect 298622 636552 298746 636652
rect 298846 636552 298880 636652
rect 297820 636428 298880 636552
rect 297820 636328 297850 636428
rect 297950 636328 298074 636428
rect 298174 636328 298298 636428
rect 298398 636328 298522 636428
rect 298622 636328 298746 636428
rect 298846 636328 298880 636428
rect 297820 636204 298880 636328
rect 297820 636104 297850 636204
rect 297950 636104 298074 636204
rect 298174 636104 298298 636204
rect 298398 636104 298522 636204
rect 298622 636104 298746 636204
rect 298846 636104 298880 636204
rect 297820 635980 298880 636104
rect 297820 635880 297850 635980
rect 297950 635880 298074 635980
rect 298174 635880 298298 635980
rect 298398 635880 298522 635980
rect 298622 635880 298746 635980
rect 298846 635880 298880 635980
rect 297820 635756 298880 635880
rect 297820 635656 297850 635756
rect 297950 635656 298074 635756
rect 298174 635656 298298 635756
rect 298398 635656 298522 635756
rect 298622 635656 298746 635756
rect 298846 635656 298880 635756
rect 297820 635532 298880 635656
rect 297820 635432 297850 635532
rect 297950 635432 298074 635532
rect 298174 635432 298298 635532
rect 298398 635432 298522 635532
rect 298622 635432 298746 635532
rect 298846 635432 298880 635532
rect 297820 635308 298880 635432
rect 297820 635208 297850 635308
rect 297950 635208 298074 635308
rect 298174 635208 298298 635308
rect 298398 635208 298522 635308
rect 298622 635208 298746 635308
rect 298846 635208 298880 635308
rect 297820 635084 298880 635208
rect 297820 634984 297850 635084
rect 297950 634984 298074 635084
rect 298174 634984 298298 635084
rect 298398 634984 298522 635084
rect 298622 634984 298746 635084
rect 298846 634984 298880 635084
rect 297820 634860 298880 634984
rect 297820 634760 297850 634860
rect 297950 634760 298074 634860
rect 298174 634760 298298 634860
rect 298398 634760 298522 634860
rect 298622 634760 298746 634860
rect 298846 634760 298880 634860
rect 297820 634636 298880 634760
rect 297820 634536 297850 634636
rect 297950 634536 298074 634636
rect 298174 634536 298298 634636
rect 298398 634536 298522 634636
rect 298622 634536 298746 634636
rect 298846 634536 298880 634636
rect 297820 634412 298880 634536
rect 297820 634312 297850 634412
rect 297950 634312 298074 634412
rect 298174 634312 298298 634412
rect 298398 634312 298522 634412
rect 298622 634312 298746 634412
rect 298846 634312 298880 634412
rect 297820 634188 298880 634312
rect 297820 634088 297850 634188
rect 297950 634088 298074 634188
rect 298174 634088 298298 634188
rect 298398 634088 298522 634188
rect 298622 634088 298746 634188
rect 298846 634088 298880 634188
rect 297820 633964 298880 634088
rect 297820 633864 297850 633964
rect 297950 633864 298074 633964
rect 298174 633864 298298 633964
rect 298398 633864 298522 633964
rect 298622 633864 298746 633964
rect 298846 633864 298880 633964
rect 297820 633740 298880 633864
rect 297820 633640 297850 633740
rect 297950 633640 298074 633740
rect 298174 633640 298298 633740
rect 298398 633640 298522 633740
rect 298622 633640 298746 633740
rect 298846 633640 298880 633740
rect 297820 633516 298880 633640
rect 297820 633416 297850 633516
rect 297950 633416 298074 633516
rect 298174 633416 298298 633516
rect 298398 633416 298522 633516
rect 298622 633416 298746 633516
rect 298846 633416 298880 633516
rect 297820 633292 298880 633416
rect 297820 633192 297850 633292
rect 297950 633192 298074 633292
rect 298174 633192 298298 633292
rect 298398 633192 298522 633292
rect 298622 633192 298746 633292
rect 298846 633192 298880 633292
rect 297820 633068 298880 633192
rect 297820 632968 297850 633068
rect 297950 632968 298074 633068
rect 298174 632968 298298 633068
rect 298398 632968 298522 633068
rect 298622 632968 298746 633068
rect 298846 632968 298880 633068
rect 297820 632844 298880 632968
rect 297820 632744 297850 632844
rect 297950 632744 298074 632844
rect 298174 632744 298298 632844
rect 298398 632744 298522 632844
rect 298622 632744 298746 632844
rect 298846 632744 298880 632844
rect 297820 632620 298880 632744
rect 297820 632520 297850 632620
rect 297950 632520 298074 632620
rect 298174 632520 298298 632620
rect 298398 632520 298522 632620
rect 298622 632520 298746 632620
rect 298846 632520 298880 632620
rect 297820 632396 298880 632520
rect 297820 632296 297850 632396
rect 297950 632296 298074 632396
rect 298174 632296 298298 632396
rect 298398 632296 298522 632396
rect 298622 632296 298746 632396
rect 298846 632296 298880 632396
rect 297820 632172 298880 632296
rect 297820 632072 297850 632172
rect 297950 632072 298074 632172
rect 298174 632072 298298 632172
rect 298398 632072 298522 632172
rect 298622 632072 298746 632172
rect 298846 632072 298880 632172
rect 297820 631948 298880 632072
rect 297820 631848 297850 631948
rect 297950 631848 298074 631948
rect 298174 631848 298298 631948
rect 298398 631848 298522 631948
rect 298622 631848 298746 631948
rect 298846 631848 298880 631948
rect 297820 631724 298880 631848
rect 297820 631624 297850 631724
rect 297950 631624 298074 631724
rect 298174 631624 298298 631724
rect 298398 631624 298522 631724
rect 298622 631624 298746 631724
rect 298846 631624 298880 631724
rect 297820 631500 298880 631624
rect 297820 631400 297850 631500
rect 297950 631400 298074 631500
rect 298174 631400 298298 631500
rect 298398 631400 298522 631500
rect 298622 631400 298746 631500
rect 298846 631400 298880 631500
rect 297820 631360 298880 631400
rect 342100 637996 343160 638020
rect 342100 637896 342130 637996
rect 342230 637896 342354 637996
rect 342454 637896 342578 637996
rect 342678 637896 342802 637996
rect 342902 637896 343026 637996
rect 343126 637896 343160 637996
rect 342100 637772 343160 637896
rect 342100 637672 342130 637772
rect 342230 637672 342354 637772
rect 342454 637672 342578 637772
rect 342678 637672 342802 637772
rect 342902 637672 343026 637772
rect 343126 637672 343160 637772
rect 342100 637548 343160 637672
rect 342100 637448 342130 637548
rect 342230 637448 342354 637548
rect 342454 637448 342578 637548
rect 342678 637448 342802 637548
rect 342902 637448 343026 637548
rect 343126 637448 343160 637548
rect 342100 637324 343160 637448
rect 342100 637224 342130 637324
rect 342230 637224 342354 637324
rect 342454 637224 342578 637324
rect 342678 637224 342802 637324
rect 342902 637224 343026 637324
rect 343126 637224 343160 637324
rect 342100 637100 343160 637224
rect 342100 637000 342130 637100
rect 342230 637000 342354 637100
rect 342454 637000 342578 637100
rect 342678 637000 342802 637100
rect 342902 637000 343026 637100
rect 343126 637000 343160 637100
rect 342100 636876 343160 637000
rect 342100 636776 342130 636876
rect 342230 636776 342354 636876
rect 342454 636776 342578 636876
rect 342678 636776 342802 636876
rect 342902 636776 343026 636876
rect 343126 636776 343160 636876
rect 342100 636652 343160 636776
rect 342100 636552 342130 636652
rect 342230 636552 342354 636652
rect 342454 636552 342578 636652
rect 342678 636552 342802 636652
rect 342902 636552 343026 636652
rect 343126 636552 343160 636652
rect 342100 636428 343160 636552
rect 342100 636328 342130 636428
rect 342230 636328 342354 636428
rect 342454 636328 342578 636428
rect 342678 636328 342802 636428
rect 342902 636328 343026 636428
rect 343126 636328 343160 636428
rect 342100 636204 343160 636328
rect 342100 636104 342130 636204
rect 342230 636104 342354 636204
rect 342454 636104 342578 636204
rect 342678 636104 342802 636204
rect 342902 636104 343026 636204
rect 343126 636104 343160 636204
rect 342100 635980 343160 636104
rect 342100 635880 342130 635980
rect 342230 635880 342354 635980
rect 342454 635880 342578 635980
rect 342678 635880 342802 635980
rect 342902 635880 343026 635980
rect 343126 635880 343160 635980
rect 342100 635756 343160 635880
rect 342100 635656 342130 635756
rect 342230 635656 342354 635756
rect 342454 635656 342578 635756
rect 342678 635656 342802 635756
rect 342902 635656 343026 635756
rect 343126 635656 343160 635756
rect 342100 635532 343160 635656
rect 342100 635432 342130 635532
rect 342230 635432 342354 635532
rect 342454 635432 342578 635532
rect 342678 635432 342802 635532
rect 342902 635432 343026 635532
rect 343126 635432 343160 635532
rect 342100 635308 343160 635432
rect 342100 635208 342130 635308
rect 342230 635208 342354 635308
rect 342454 635208 342578 635308
rect 342678 635208 342802 635308
rect 342902 635208 343026 635308
rect 343126 635208 343160 635308
rect 342100 635084 343160 635208
rect 342100 634984 342130 635084
rect 342230 634984 342354 635084
rect 342454 634984 342578 635084
rect 342678 634984 342802 635084
rect 342902 634984 343026 635084
rect 343126 634984 343160 635084
rect 342100 634860 343160 634984
rect 342100 634760 342130 634860
rect 342230 634760 342354 634860
rect 342454 634760 342578 634860
rect 342678 634760 342802 634860
rect 342902 634760 343026 634860
rect 343126 634760 343160 634860
rect 342100 634636 343160 634760
rect 342100 634536 342130 634636
rect 342230 634536 342354 634636
rect 342454 634536 342578 634636
rect 342678 634536 342802 634636
rect 342902 634536 343026 634636
rect 343126 634536 343160 634636
rect 342100 634412 343160 634536
rect 342100 634312 342130 634412
rect 342230 634312 342354 634412
rect 342454 634312 342578 634412
rect 342678 634312 342802 634412
rect 342902 634312 343026 634412
rect 343126 634312 343160 634412
rect 342100 634188 343160 634312
rect 342100 634088 342130 634188
rect 342230 634088 342354 634188
rect 342454 634088 342578 634188
rect 342678 634088 342802 634188
rect 342902 634088 343026 634188
rect 343126 634088 343160 634188
rect 342100 633964 343160 634088
rect 342100 633864 342130 633964
rect 342230 633864 342354 633964
rect 342454 633864 342578 633964
rect 342678 633864 342802 633964
rect 342902 633864 343026 633964
rect 343126 633864 343160 633964
rect 342100 633740 343160 633864
rect 342100 633640 342130 633740
rect 342230 633640 342354 633740
rect 342454 633640 342578 633740
rect 342678 633640 342802 633740
rect 342902 633640 343026 633740
rect 343126 633640 343160 633740
rect 342100 633516 343160 633640
rect 342100 633416 342130 633516
rect 342230 633416 342354 633516
rect 342454 633416 342578 633516
rect 342678 633416 342802 633516
rect 342902 633416 343026 633516
rect 343126 633416 343160 633516
rect 342100 633292 343160 633416
rect 342100 633192 342130 633292
rect 342230 633192 342354 633292
rect 342454 633192 342578 633292
rect 342678 633192 342802 633292
rect 342902 633192 343026 633292
rect 343126 633192 343160 633292
rect 342100 633068 343160 633192
rect 342100 632968 342130 633068
rect 342230 632968 342354 633068
rect 342454 632968 342578 633068
rect 342678 632968 342802 633068
rect 342902 632968 343026 633068
rect 343126 632968 343160 633068
rect 342100 632844 343160 632968
rect 342100 632744 342130 632844
rect 342230 632744 342354 632844
rect 342454 632744 342578 632844
rect 342678 632744 342802 632844
rect 342902 632744 343026 632844
rect 343126 632744 343160 632844
rect 342100 632620 343160 632744
rect 342100 632520 342130 632620
rect 342230 632520 342354 632620
rect 342454 632520 342578 632620
rect 342678 632520 342802 632620
rect 342902 632520 343026 632620
rect 343126 632520 343160 632620
rect 342100 632396 343160 632520
rect 342100 632296 342130 632396
rect 342230 632296 342354 632396
rect 342454 632296 342578 632396
rect 342678 632296 342802 632396
rect 342902 632296 343026 632396
rect 343126 632296 343160 632396
rect 342100 632172 343160 632296
rect 342100 632072 342130 632172
rect 342230 632072 342354 632172
rect 342454 632072 342578 632172
rect 342678 632072 342802 632172
rect 342902 632072 343026 632172
rect 343126 632072 343160 632172
rect 342100 631948 343160 632072
rect 342100 631848 342130 631948
rect 342230 631848 342354 631948
rect 342454 631848 342578 631948
rect 342678 631848 342802 631948
rect 342902 631848 343026 631948
rect 343126 631848 343160 631948
rect 342100 631724 343160 631848
rect 342100 631624 342130 631724
rect 342230 631624 342354 631724
rect 342454 631624 342578 631724
rect 342678 631624 342802 631724
rect 342902 631624 343026 631724
rect 343126 631624 343160 631724
rect 342100 631500 343160 631624
rect 342100 631400 342130 631500
rect 342230 631400 342354 631500
rect 342454 631400 342578 631500
rect 342678 631400 342802 631500
rect 342902 631400 343026 631500
rect 343126 631400 343160 631500
rect 342100 631360 343160 631400
rect 297820 624596 298878 624606
rect 297820 624496 297850 624596
rect 297950 624496 298074 624596
rect 298174 624496 298298 624596
rect 298398 624496 298522 624596
rect 298622 624496 298746 624596
rect 298846 624496 298878 624596
rect 297820 624372 298878 624496
rect 297820 624272 297850 624372
rect 297950 624272 298074 624372
rect 298174 624272 298298 624372
rect 298398 624272 298522 624372
rect 298622 624272 298746 624372
rect 298846 624272 298878 624372
rect 297820 624148 298878 624272
rect 342100 624596 343158 624606
rect 342100 624496 342130 624596
rect 342230 624496 342354 624596
rect 342454 624496 342578 624596
rect 342678 624496 342802 624596
rect 342902 624496 343026 624596
rect 343126 624496 343158 624596
rect 342100 624372 343158 624496
rect 342100 624272 342130 624372
rect 342230 624272 342354 624372
rect 342454 624272 342578 624372
rect 342678 624272 342802 624372
rect 342902 624272 343026 624372
rect 343126 624272 343158 624372
rect 297820 624048 297850 624148
rect 297950 624048 298074 624148
rect 298174 624048 298298 624148
rect 298398 624048 298522 624148
rect 298622 624048 298746 624148
rect 298846 624048 298878 624148
rect 342100 624148 343158 624272
rect 297820 623924 298878 624048
rect 342100 624048 342130 624148
rect 342230 624048 342354 624148
rect 342454 624048 342578 624148
rect 342678 624048 342802 624148
rect 342902 624048 343026 624148
rect 343126 624048 343158 624148
rect 297820 623824 297850 623924
rect 297950 623824 298074 623924
rect 298174 623824 298298 623924
rect 298398 623824 298522 623924
rect 298622 623824 298746 623924
rect 298846 623824 298878 623924
rect 297820 623700 298878 623824
rect 297820 623600 297850 623700
rect 297950 623600 298074 623700
rect 298174 623600 298298 623700
rect 298398 623600 298522 623700
rect 298622 623600 298746 623700
rect 298846 623600 298878 623700
rect 297820 623476 298878 623600
rect 297820 623376 297850 623476
rect 297950 623376 298074 623476
rect 298174 623376 298298 623476
rect 298398 623376 298522 623476
rect 298622 623376 298746 623476
rect 298846 623376 298878 623476
rect 297820 623252 298878 623376
rect 297820 623152 297850 623252
rect 297950 623152 298074 623252
rect 298174 623152 298298 623252
rect 298398 623152 298522 623252
rect 298622 623152 298746 623252
rect 298846 623152 298878 623252
rect 297820 623028 298878 623152
rect 297820 622928 297850 623028
rect 297950 622928 298074 623028
rect 298174 622928 298298 623028
rect 298398 622928 298522 623028
rect 298622 622928 298746 623028
rect 298846 622928 298878 623028
rect 297820 622804 298878 622928
rect 297820 622704 297850 622804
rect 297950 622704 298074 622804
rect 298174 622704 298298 622804
rect 298398 622704 298522 622804
rect 298622 622704 298746 622804
rect 298846 622704 298878 622804
rect 297820 622580 298878 622704
rect 297820 622480 297850 622580
rect 297950 622480 298074 622580
rect 298174 622480 298298 622580
rect 298398 622480 298522 622580
rect 298622 622480 298746 622580
rect 298846 622480 298878 622580
rect 297820 622356 298878 622480
rect 297820 622256 297850 622356
rect 297950 622256 298074 622356
rect 298174 622256 298298 622356
rect 298398 622256 298522 622356
rect 298622 622256 298746 622356
rect 298846 622256 298878 622356
rect 297820 622132 298878 622256
rect 297820 622032 297850 622132
rect 297950 622032 298074 622132
rect 298174 622032 298298 622132
rect 298398 622032 298522 622132
rect 298622 622032 298746 622132
rect 298846 622032 298878 622132
rect 297820 621908 298878 622032
rect 297820 621808 297850 621908
rect 297950 621808 298074 621908
rect 298174 621808 298298 621908
rect 298398 621808 298522 621908
rect 298622 621808 298746 621908
rect 298846 621808 298878 621908
rect 297820 621684 298878 621808
rect 297820 621584 297850 621684
rect 297950 621584 298074 621684
rect 298174 621584 298298 621684
rect 298398 621584 298522 621684
rect 298622 621584 298746 621684
rect 298846 621584 298878 621684
rect 297820 621460 298878 621584
rect 297820 621360 297850 621460
rect 297950 621360 298074 621460
rect 298174 621360 298298 621460
rect 298398 621360 298522 621460
rect 298622 621360 298746 621460
rect 298846 621360 298878 621460
rect 297820 621236 298878 621360
rect 297820 621136 297850 621236
rect 297950 621136 298074 621236
rect 298174 621136 298298 621236
rect 298398 621136 298522 621236
rect 298622 621136 298746 621236
rect 298846 621136 298878 621236
rect 297820 621012 298878 621136
rect 297820 620912 297850 621012
rect 297950 620912 298074 621012
rect 298174 620912 298298 621012
rect 298398 620912 298522 621012
rect 298622 620912 298746 621012
rect 298846 620912 298878 621012
rect 297820 620788 298878 620912
rect 297820 620688 297850 620788
rect 297950 620688 298074 620788
rect 298174 620688 298298 620788
rect 298398 620688 298522 620788
rect 298622 620688 298746 620788
rect 298846 620688 298878 620788
rect 297820 620564 298878 620688
rect 297820 620464 297850 620564
rect 297950 620464 298074 620564
rect 298174 620464 298298 620564
rect 298398 620464 298522 620564
rect 298622 620464 298746 620564
rect 298846 620464 298878 620564
rect 297820 620340 298878 620464
rect 297820 620240 297850 620340
rect 297950 620240 298074 620340
rect 298174 620240 298298 620340
rect 298398 620240 298522 620340
rect 298622 620240 298746 620340
rect 298846 620240 298878 620340
rect 297820 620116 298878 620240
rect 297820 620016 297850 620116
rect 297950 620016 298074 620116
rect 298174 620016 298298 620116
rect 298398 620016 298522 620116
rect 298622 620016 298746 620116
rect 298846 620016 298878 620116
rect 297820 619892 298878 620016
rect 297820 619792 297850 619892
rect 297950 619792 298074 619892
rect 298174 619792 298298 619892
rect 298398 619792 298522 619892
rect 298622 619792 298746 619892
rect 298846 619792 298878 619892
rect 297820 619668 298878 619792
rect 297820 619568 297850 619668
rect 297950 619568 298074 619668
rect 298174 619568 298298 619668
rect 298398 619568 298522 619668
rect 298622 619568 298746 619668
rect 298846 619568 298878 619668
rect 297820 619444 298878 619568
rect 297820 619344 297850 619444
rect 297950 619344 298074 619444
rect 298174 619344 298298 619444
rect 298398 619344 298522 619444
rect 298622 619344 298746 619444
rect 298846 619344 298878 619444
rect 297820 619220 298878 619344
rect 297820 619120 297850 619220
rect 297950 619120 298074 619220
rect 298174 619120 298298 619220
rect 298398 619120 298522 619220
rect 298622 619120 298746 619220
rect 298846 619120 298878 619220
rect 297820 618996 298878 619120
rect 297820 618896 297850 618996
rect 297950 618896 298074 618996
rect 298174 618896 298298 618996
rect 298398 618896 298522 618996
rect 298622 618896 298746 618996
rect 298846 618896 298878 618996
rect 297820 618772 298878 618896
rect 297820 618672 297850 618772
rect 297950 618672 298074 618772
rect 298174 618672 298298 618772
rect 298398 618672 298522 618772
rect 298622 618672 298746 618772
rect 298846 618672 298878 618772
rect 297820 618548 298878 618672
rect 297820 618448 297850 618548
rect 297950 618448 298074 618548
rect 298174 618448 298298 618548
rect 298398 618448 298522 618548
rect 298622 618448 298746 618548
rect 298846 618448 298878 618548
rect 297820 618324 298878 618448
rect 297820 618224 297850 618324
rect 297950 618224 298074 618324
rect 298174 618224 298298 618324
rect 298398 618224 298522 618324
rect 298622 618224 298746 618324
rect 298846 618224 298878 618324
rect 297820 618100 298878 618224
rect 297820 618000 297850 618100
rect 297950 618000 298074 618100
rect 298174 618000 298298 618100
rect 298398 618000 298522 618100
rect 298622 618000 298746 618100
rect 298846 618000 298878 618100
rect 297820 617980 298878 618000
rect 342100 623924 343158 624048
rect 342100 623824 342130 623924
rect 342230 623824 342354 623924
rect 342454 623824 342578 623924
rect 342678 623824 342802 623924
rect 342902 623824 343026 623924
rect 343126 623824 343158 623924
rect 342100 623700 343158 623824
rect 342100 623600 342130 623700
rect 342230 623600 342354 623700
rect 342454 623600 342578 623700
rect 342678 623600 342802 623700
rect 342902 623600 343026 623700
rect 343126 623600 343158 623700
rect 342100 623476 343158 623600
rect 342100 623376 342130 623476
rect 342230 623376 342354 623476
rect 342454 623376 342578 623476
rect 342678 623376 342802 623476
rect 342902 623376 343026 623476
rect 343126 623376 343158 623476
rect 342100 623252 343158 623376
rect 342100 623152 342130 623252
rect 342230 623152 342354 623252
rect 342454 623152 342578 623252
rect 342678 623152 342802 623252
rect 342902 623152 343026 623252
rect 343126 623152 343158 623252
rect 342100 623028 343158 623152
rect 342100 622928 342130 623028
rect 342230 622928 342354 623028
rect 342454 622928 342578 623028
rect 342678 622928 342802 623028
rect 342902 622928 343026 623028
rect 343126 622928 343158 623028
rect 342100 622804 343158 622928
rect 342100 622704 342130 622804
rect 342230 622704 342354 622804
rect 342454 622704 342578 622804
rect 342678 622704 342802 622804
rect 342902 622704 343026 622804
rect 343126 622704 343158 622804
rect 342100 622580 343158 622704
rect 342100 622480 342130 622580
rect 342230 622480 342354 622580
rect 342454 622480 342578 622580
rect 342678 622480 342802 622580
rect 342902 622480 343026 622580
rect 343126 622480 343158 622580
rect 342100 622356 343158 622480
rect 342100 622256 342130 622356
rect 342230 622256 342354 622356
rect 342454 622256 342578 622356
rect 342678 622256 342802 622356
rect 342902 622256 343026 622356
rect 343126 622256 343158 622356
rect 342100 622132 343158 622256
rect 342100 622032 342130 622132
rect 342230 622032 342354 622132
rect 342454 622032 342578 622132
rect 342678 622032 342802 622132
rect 342902 622032 343026 622132
rect 343126 622032 343158 622132
rect 342100 621908 343158 622032
rect 342100 621808 342130 621908
rect 342230 621808 342354 621908
rect 342454 621808 342578 621908
rect 342678 621808 342802 621908
rect 342902 621808 343026 621908
rect 343126 621808 343158 621908
rect 342100 621684 343158 621808
rect 342100 621584 342130 621684
rect 342230 621584 342354 621684
rect 342454 621584 342578 621684
rect 342678 621584 342802 621684
rect 342902 621584 343026 621684
rect 343126 621584 343158 621684
rect 342100 621460 343158 621584
rect 342100 621360 342130 621460
rect 342230 621360 342354 621460
rect 342454 621360 342578 621460
rect 342678 621360 342802 621460
rect 342902 621360 343026 621460
rect 343126 621360 343158 621460
rect 342100 621236 343158 621360
rect 342100 621136 342130 621236
rect 342230 621136 342354 621236
rect 342454 621136 342578 621236
rect 342678 621136 342802 621236
rect 342902 621136 343026 621236
rect 343126 621136 343158 621236
rect 342100 621012 343158 621136
rect 342100 620912 342130 621012
rect 342230 620912 342354 621012
rect 342454 620912 342578 621012
rect 342678 620912 342802 621012
rect 342902 620912 343026 621012
rect 343126 620912 343158 621012
rect 342100 620788 343158 620912
rect 342100 620688 342130 620788
rect 342230 620688 342354 620788
rect 342454 620688 342578 620788
rect 342678 620688 342802 620788
rect 342902 620688 343026 620788
rect 343126 620688 343158 620788
rect 342100 620564 343158 620688
rect 342100 620464 342130 620564
rect 342230 620464 342354 620564
rect 342454 620464 342578 620564
rect 342678 620464 342802 620564
rect 342902 620464 343026 620564
rect 343126 620464 343158 620564
rect 342100 620340 343158 620464
rect 342100 620240 342130 620340
rect 342230 620240 342354 620340
rect 342454 620240 342578 620340
rect 342678 620240 342802 620340
rect 342902 620240 343026 620340
rect 343126 620240 343158 620340
rect 342100 620116 343158 620240
rect 342100 620016 342130 620116
rect 342230 620016 342354 620116
rect 342454 620016 342578 620116
rect 342678 620016 342802 620116
rect 342902 620016 343026 620116
rect 343126 620016 343158 620116
rect 342100 619892 343158 620016
rect 342100 619792 342130 619892
rect 342230 619792 342354 619892
rect 342454 619792 342578 619892
rect 342678 619792 342802 619892
rect 342902 619792 343026 619892
rect 343126 619792 343158 619892
rect 342100 619668 343158 619792
rect 342100 619568 342130 619668
rect 342230 619568 342354 619668
rect 342454 619568 342578 619668
rect 342678 619568 342802 619668
rect 342902 619568 343026 619668
rect 343126 619568 343158 619668
rect 342100 619444 343158 619568
rect 342100 619344 342130 619444
rect 342230 619344 342354 619444
rect 342454 619344 342578 619444
rect 342678 619344 342802 619444
rect 342902 619344 343026 619444
rect 343126 619344 343158 619444
rect 342100 619220 343158 619344
rect 342100 619120 342130 619220
rect 342230 619120 342354 619220
rect 342454 619120 342578 619220
rect 342678 619120 342802 619220
rect 342902 619120 343026 619220
rect 343126 619120 343158 619220
rect 342100 618996 343158 619120
rect 342100 618896 342130 618996
rect 342230 618896 342354 618996
rect 342454 618896 342578 618996
rect 342678 618896 342802 618996
rect 342902 618896 343026 618996
rect 343126 618896 343158 618996
rect 342100 618772 343158 618896
rect 342100 618672 342130 618772
rect 342230 618672 342354 618772
rect 342454 618672 342578 618772
rect 342678 618672 342802 618772
rect 342902 618672 343026 618772
rect 343126 618672 343158 618772
rect 342100 618548 343158 618672
rect 342100 618448 342130 618548
rect 342230 618448 342354 618548
rect 342454 618448 342578 618548
rect 342678 618448 342802 618548
rect 342902 618448 343026 618548
rect 343126 618448 343158 618548
rect 342100 618324 343158 618448
rect 342100 618224 342130 618324
rect 342230 618224 342354 618324
rect 342454 618224 342578 618324
rect 342678 618224 342802 618324
rect 342902 618224 343026 618324
rect 343126 618224 343158 618324
rect 342100 618100 343158 618224
rect 342100 618000 342130 618100
rect 342230 618000 342354 618100
rect 342454 618000 342578 618100
rect 342678 618000 342802 618100
rect 342902 618000 343026 618100
rect 343126 618000 343158 618100
rect 342100 617980 343158 618000
rect 298836 615474 305496 615504
rect 298836 615374 298876 615474
rect 298976 615374 299100 615474
rect 299200 615374 299324 615474
rect 299424 615374 299548 615474
rect 299648 615374 299772 615474
rect 299872 615374 299996 615474
rect 300096 615374 300220 615474
rect 300320 615374 300444 615474
rect 300544 615374 300668 615474
rect 300768 615374 300892 615474
rect 300992 615374 301116 615474
rect 301216 615374 301340 615474
rect 301440 615374 301564 615474
rect 301664 615374 301788 615474
rect 301888 615374 302012 615474
rect 302112 615374 302236 615474
rect 302336 615374 302460 615474
rect 302560 615374 302684 615474
rect 302784 615374 302908 615474
rect 303008 615374 303132 615474
rect 303232 615374 303356 615474
rect 303456 615374 303580 615474
rect 303680 615374 303804 615474
rect 303904 615374 304028 615474
rect 304128 615374 304252 615474
rect 304352 615374 304476 615474
rect 304576 615374 304700 615474
rect 304800 615374 304924 615474
rect 305024 615374 305148 615474
rect 305248 615374 305372 615474
rect 305472 615374 305496 615474
rect 298836 615250 305496 615374
rect 298836 615150 298876 615250
rect 298976 615150 299100 615250
rect 299200 615150 299324 615250
rect 299424 615150 299548 615250
rect 299648 615150 299772 615250
rect 299872 615150 299996 615250
rect 300096 615150 300220 615250
rect 300320 615150 300444 615250
rect 300544 615150 300668 615250
rect 300768 615150 300892 615250
rect 300992 615150 301116 615250
rect 301216 615150 301340 615250
rect 301440 615150 301564 615250
rect 301664 615150 301788 615250
rect 301888 615150 302012 615250
rect 302112 615150 302236 615250
rect 302336 615150 302460 615250
rect 302560 615150 302684 615250
rect 302784 615150 302908 615250
rect 303008 615150 303132 615250
rect 303232 615150 303356 615250
rect 303456 615150 303580 615250
rect 303680 615150 303804 615250
rect 303904 615150 304028 615250
rect 304128 615150 304252 615250
rect 304352 615150 304476 615250
rect 304576 615150 304700 615250
rect 304800 615150 304924 615250
rect 305024 615150 305148 615250
rect 305248 615150 305372 615250
rect 305472 615150 305496 615250
rect 298836 615026 305496 615150
rect 298836 614926 298876 615026
rect 298976 614926 299100 615026
rect 299200 614926 299324 615026
rect 299424 614926 299548 615026
rect 299648 614926 299772 615026
rect 299872 614926 299996 615026
rect 300096 614926 300220 615026
rect 300320 614926 300444 615026
rect 300544 614926 300668 615026
rect 300768 614926 300892 615026
rect 300992 614926 301116 615026
rect 301216 614926 301340 615026
rect 301440 614926 301564 615026
rect 301664 614926 301788 615026
rect 301888 614926 302012 615026
rect 302112 614926 302236 615026
rect 302336 614926 302460 615026
rect 302560 614926 302684 615026
rect 302784 614926 302908 615026
rect 303008 614926 303132 615026
rect 303232 614926 303356 615026
rect 303456 614926 303580 615026
rect 303680 614926 303804 615026
rect 303904 614926 304028 615026
rect 304128 614926 304252 615026
rect 304352 614926 304476 615026
rect 304576 614926 304700 615026
rect 304800 614926 304924 615026
rect 305024 614926 305148 615026
rect 305248 614926 305372 615026
rect 305472 614926 305496 615026
rect 298836 614802 305496 614926
rect 298836 614702 298876 614802
rect 298976 614702 299100 614802
rect 299200 614702 299324 614802
rect 299424 614702 299548 614802
rect 299648 614702 299772 614802
rect 299872 614702 299996 614802
rect 300096 614702 300220 614802
rect 300320 614702 300444 614802
rect 300544 614702 300668 614802
rect 300768 614702 300892 614802
rect 300992 614702 301116 614802
rect 301216 614702 301340 614802
rect 301440 614702 301564 614802
rect 301664 614702 301788 614802
rect 301888 614702 302012 614802
rect 302112 614702 302236 614802
rect 302336 614702 302460 614802
rect 302560 614702 302684 614802
rect 302784 614702 302908 614802
rect 303008 614702 303132 614802
rect 303232 614702 303356 614802
rect 303456 614702 303580 614802
rect 303680 614702 303804 614802
rect 303904 614702 304028 614802
rect 304128 614702 304252 614802
rect 304352 614702 304476 614802
rect 304576 614702 304700 614802
rect 304800 614702 304924 614802
rect 305024 614702 305148 614802
rect 305248 614702 305372 614802
rect 305472 614702 305496 614802
rect 298836 614578 305496 614702
rect 298836 614478 298876 614578
rect 298976 614478 299100 614578
rect 299200 614478 299324 614578
rect 299424 614478 299548 614578
rect 299648 614478 299772 614578
rect 299872 614478 299996 614578
rect 300096 614478 300220 614578
rect 300320 614478 300444 614578
rect 300544 614478 300668 614578
rect 300768 614478 300892 614578
rect 300992 614478 301116 614578
rect 301216 614478 301340 614578
rect 301440 614478 301564 614578
rect 301664 614478 301788 614578
rect 301888 614478 302012 614578
rect 302112 614478 302236 614578
rect 302336 614478 302460 614578
rect 302560 614478 302684 614578
rect 302784 614478 302908 614578
rect 303008 614478 303132 614578
rect 303232 614478 303356 614578
rect 303456 614478 303580 614578
rect 303680 614478 303804 614578
rect 303904 614478 304028 614578
rect 304128 614478 304252 614578
rect 304352 614478 304476 614578
rect 304576 614478 304700 614578
rect 304800 614478 304924 614578
rect 305024 614478 305148 614578
rect 305248 614478 305372 614578
rect 305472 614478 305496 614578
rect 298836 614444 305496 614478
rect 309306 615474 315966 615504
rect 309306 615374 309346 615474
rect 309446 615374 309570 615474
rect 309670 615374 309794 615474
rect 309894 615374 310018 615474
rect 310118 615374 310242 615474
rect 310342 615374 310466 615474
rect 310566 615374 310690 615474
rect 310790 615374 310914 615474
rect 311014 615374 311138 615474
rect 311238 615374 311362 615474
rect 311462 615374 311586 615474
rect 311686 615374 311810 615474
rect 311910 615374 312034 615474
rect 312134 615374 312258 615474
rect 312358 615374 312482 615474
rect 312582 615374 312706 615474
rect 312806 615374 312930 615474
rect 313030 615374 313154 615474
rect 313254 615374 313378 615474
rect 313478 615374 313602 615474
rect 313702 615374 313826 615474
rect 313926 615374 314050 615474
rect 314150 615374 314274 615474
rect 314374 615374 314498 615474
rect 314598 615374 314722 615474
rect 314822 615374 314946 615474
rect 315046 615374 315170 615474
rect 315270 615374 315394 615474
rect 315494 615374 315618 615474
rect 315718 615374 315842 615474
rect 315942 615374 315966 615474
rect 309306 615250 315966 615374
rect 309306 615150 309346 615250
rect 309446 615150 309570 615250
rect 309670 615150 309794 615250
rect 309894 615150 310018 615250
rect 310118 615150 310242 615250
rect 310342 615150 310466 615250
rect 310566 615150 310690 615250
rect 310790 615150 310914 615250
rect 311014 615150 311138 615250
rect 311238 615150 311362 615250
rect 311462 615150 311586 615250
rect 311686 615150 311810 615250
rect 311910 615150 312034 615250
rect 312134 615150 312258 615250
rect 312358 615150 312482 615250
rect 312582 615150 312706 615250
rect 312806 615150 312930 615250
rect 313030 615150 313154 615250
rect 313254 615150 313378 615250
rect 313478 615150 313602 615250
rect 313702 615150 313826 615250
rect 313926 615150 314050 615250
rect 314150 615150 314274 615250
rect 314374 615150 314498 615250
rect 314598 615150 314722 615250
rect 314822 615150 314946 615250
rect 315046 615150 315170 615250
rect 315270 615150 315394 615250
rect 315494 615150 315618 615250
rect 315718 615150 315842 615250
rect 315942 615150 315966 615250
rect 309306 615026 315966 615150
rect 309306 614926 309346 615026
rect 309446 614926 309570 615026
rect 309670 614926 309794 615026
rect 309894 614926 310018 615026
rect 310118 614926 310242 615026
rect 310342 614926 310466 615026
rect 310566 614926 310690 615026
rect 310790 614926 310914 615026
rect 311014 614926 311138 615026
rect 311238 614926 311362 615026
rect 311462 614926 311586 615026
rect 311686 614926 311810 615026
rect 311910 614926 312034 615026
rect 312134 614926 312258 615026
rect 312358 614926 312482 615026
rect 312582 614926 312706 615026
rect 312806 614926 312930 615026
rect 313030 614926 313154 615026
rect 313254 614926 313378 615026
rect 313478 614926 313602 615026
rect 313702 614926 313826 615026
rect 313926 614926 314050 615026
rect 314150 614926 314274 615026
rect 314374 614926 314498 615026
rect 314598 614926 314722 615026
rect 314822 614926 314946 615026
rect 315046 614926 315170 615026
rect 315270 614926 315394 615026
rect 315494 614926 315618 615026
rect 315718 614926 315842 615026
rect 315942 614926 315966 615026
rect 309306 614802 315966 614926
rect 309306 614702 309346 614802
rect 309446 614702 309570 614802
rect 309670 614702 309794 614802
rect 309894 614702 310018 614802
rect 310118 614702 310242 614802
rect 310342 614702 310466 614802
rect 310566 614702 310690 614802
rect 310790 614702 310914 614802
rect 311014 614702 311138 614802
rect 311238 614702 311362 614802
rect 311462 614702 311586 614802
rect 311686 614702 311810 614802
rect 311910 614702 312034 614802
rect 312134 614702 312258 614802
rect 312358 614702 312482 614802
rect 312582 614702 312706 614802
rect 312806 614702 312930 614802
rect 313030 614702 313154 614802
rect 313254 614702 313378 614802
rect 313478 614702 313602 614802
rect 313702 614702 313826 614802
rect 313926 614702 314050 614802
rect 314150 614702 314274 614802
rect 314374 614702 314498 614802
rect 314598 614702 314722 614802
rect 314822 614702 314946 614802
rect 315046 614702 315170 614802
rect 315270 614702 315394 614802
rect 315494 614702 315618 614802
rect 315718 614702 315842 614802
rect 315942 614702 315966 614802
rect 309306 614578 315966 614702
rect 309306 614478 309346 614578
rect 309446 614478 309570 614578
rect 309670 614478 309794 614578
rect 309894 614478 310018 614578
rect 310118 614478 310242 614578
rect 310342 614478 310466 614578
rect 310566 614478 310690 614578
rect 310790 614478 310914 614578
rect 311014 614478 311138 614578
rect 311238 614478 311362 614578
rect 311462 614478 311586 614578
rect 311686 614478 311810 614578
rect 311910 614478 312034 614578
rect 312134 614478 312258 614578
rect 312358 614478 312482 614578
rect 312582 614478 312706 614578
rect 312806 614478 312930 614578
rect 313030 614478 313154 614578
rect 313254 614478 313378 614578
rect 313478 614478 313602 614578
rect 313702 614478 313826 614578
rect 313926 614478 314050 614578
rect 314150 614478 314274 614578
rect 314374 614478 314498 614578
rect 314598 614478 314722 614578
rect 314822 614478 314946 614578
rect 315046 614478 315170 614578
rect 315270 614478 315394 614578
rect 315494 614478 315618 614578
rect 315718 614478 315842 614578
rect 315942 614478 315966 614578
rect 309306 614444 315966 614478
rect 335576 615494 342236 615524
rect 335576 615394 335616 615494
rect 335716 615394 335840 615494
rect 335940 615394 336064 615494
rect 336164 615394 336288 615494
rect 336388 615394 336512 615494
rect 336612 615394 336736 615494
rect 336836 615394 336960 615494
rect 337060 615394 337184 615494
rect 337284 615394 337408 615494
rect 337508 615394 337632 615494
rect 337732 615394 337856 615494
rect 337956 615394 338080 615494
rect 338180 615394 338304 615494
rect 338404 615394 338528 615494
rect 338628 615394 338752 615494
rect 338852 615394 338976 615494
rect 339076 615394 339200 615494
rect 339300 615394 339424 615494
rect 339524 615394 339648 615494
rect 339748 615394 339872 615494
rect 339972 615394 340096 615494
rect 340196 615394 340320 615494
rect 340420 615394 340544 615494
rect 340644 615394 340768 615494
rect 340868 615394 340992 615494
rect 341092 615394 341216 615494
rect 341316 615394 341440 615494
rect 341540 615394 341664 615494
rect 341764 615394 341888 615494
rect 341988 615394 342112 615494
rect 342212 615394 342236 615494
rect 335576 615270 342236 615394
rect 335576 615170 335616 615270
rect 335716 615170 335840 615270
rect 335940 615170 336064 615270
rect 336164 615170 336288 615270
rect 336388 615170 336512 615270
rect 336612 615170 336736 615270
rect 336836 615170 336960 615270
rect 337060 615170 337184 615270
rect 337284 615170 337408 615270
rect 337508 615170 337632 615270
rect 337732 615170 337856 615270
rect 337956 615170 338080 615270
rect 338180 615170 338304 615270
rect 338404 615170 338528 615270
rect 338628 615170 338752 615270
rect 338852 615170 338976 615270
rect 339076 615170 339200 615270
rect 339300 615170 339424 615270
rect 339524 615170 339648 615270
rect 339748 615170 339872 615270
rect 339972 615170 340096 615270
rect 340196 615170 340320 615270
rect 340420 615170 340544 615270
rect 340644 615170 340768 615270
rect 340868 615170 340992 615270
rect 341092 615170 341216 615270
rect 341316 615170 341440 615270
rect 341540 615170 341664 615270
rect 341764 615170 341888 615270
rect 341988 615170 342112 615270
rect 342212 615170 342236 615270
rect 335576 615046 342236 615170
rect 335576 614946 335616 615046
rect 335716 614946 335840 615046
rect 335940 614946 336064 615046
rect 336164 614946 336288 615046
rect 336388 614946 336512 615046
rect 336612 614946 336736 615046
rect 336836 614946 336960 615046
rect 337060 614946 337184 615046
rect 337284 614946 337408 615046
rect 337508 614946 337632 615046
rect 337732 614946 337856 615046
rect 337956 614946 338080 615046
rect 338180 614946 338304 615046
rect 338404 614946 338528 615046
rect 338628 614946 338752 615046
rect 338852 614946 338976 615046
rect 339076 614946 339200 615046
rect 339300 614946 339424 615046
rect 339524 614946 339648 615046
rect 339748 614946 339872 615046
rect 339972 614946 340096 615046
rect 340196 614946 340320 615046
rect 340420 614946 340544 615046
rect 340644 614946 340768 615046
rect 340868 614946 340992 615046
rect 341092 614946 341216 615046
rect 341316 614946 341440 615046
rect 341540 614946 341664 615046
rect 341764 614946 341888 615046
rect 341988 614946 342112 615046
rect 342212 614946 342236 615046
rect 335576 614822 342236 614946
rect 335576 614722 335616 614822
rect 335716 614722 335840 614822
rect 335940 614722 336064 614822
rect 336164 614722 336288 614822
rect 336388 614722 336512 614822
rect 336612 614722 336736 614822
rect 336836 614722 336960 614822
rect 337060 614722 337184 614822
rect 337284 614722 337408 614822
rect 337508 614722 337632 614822
rect 337732 614722 337856 614822
rect 337956 614722 338080 614822
rect 338180 614722 338304 614822
rect 338404 614722 338528 614822
rect 338628 614722 338752 614822
rect 338852 614722 338976 614822
rect 339076 614722 339200 614822
rect 339300 614722 339424 614822
rect 339524 614722 339648 614822
rect 339748 614722 339872 614822
rect 339972 614722 340096 614822
rect 340196 614722 340320 614822
rect 340420 614722 340544 614822
rect 340644 614722 340768 614822
rect 340868 614722 340992 614822
rect 341092 614722 341216 614822
rect 341316 614722 341440 614822
rect 341540 614722 341664 614822
rect 341764 614722 341888 614822
rect 341988 614722 342112 614822
rect 342212 614722 342236 614822
rect 335576 614598 342236 614722
rect 335576 614498 335616 614598
rect 335716 614498 335840 614598
rect 335940 614498 336064 614598
rect 336164 614498 336288 614598
rect 336388 614498 336512 614598
rect 336612 614498 336736 614598
rect 336836 614498 336960 614598
rect 337060 614498 337184 614598
rect 337284 614498 337408 614598
rect 337508 614498 337632 614598
rect 337732 614498 337856 614598
rect 337956 614498 338080 614598
rect 338180 614498 338304 614598
rect 338404 614498 338528 614598
rect 338628 614498 338752 614598
rect 338852 614498 338976 614598
rect 339076 614498 339200 614598
rect 339300 614498 339424 614598
rect 339524 614498 339648 614598
rect 339748 614498 339872 614598
rect 339972 614498 340096 614598
rect 340196 614498 340320 614598
rect 340420 614498 340544 614598
rect 340644 614498 340768 614598
rect 340868 614498 340992 614598
rect 341092 614498 341216 614598
rect 341316 614498 341440 614598
rect 341540 614498 341664 614598
rect 341764 614498 341888 614598
rect 341988 614498 342112 614598
rect 342212 614498 342236 614598
rect 335576 614464 342236 614498
<< via1 >>
rect 298876 642594 298976 642694
rect 299100 642594 299200 642694
rect 299324 642594 299424 642694
rect 299548 642594 299648 642694
rect 299772 642594 299872 642694
rect 299996 642594 300096 642694
rect 300220 642594 300320 642694
rect 300444 642594 300544 642694
rect 300668 642594 300768 642694
rect 300892 642594 300992 642694
rect 301116 642594 301216 642694
rect 301340 642594 301440 642694
rect 301564 642594 301664 642694
rect 301788 642594 301888 642694
rect 302012 642594 302112 642694
rect 302236 642594 302336 642694
rect 302460 642594 302560 642694
rect 302684 642594 302784 642694
rect 302908 642594 303008 642694
rect 303132 642594 303232 642694
rect 303356 642594 303456 642694
rect 303580 642594 303680 642694
rect 303804 642594 303904 642694
rect 304028 642594 304128 642694
rect 304252 642594 304352 642694
rect 304476 642594 304576 642694
rect 304700 642594 304800 642694
rect 304924 642594 305024 642694
rect 305148 642594 305248 642694
rect 305372 642594 305472 642694
rect 298876 642370 298976 642470
rect 299100 642370 299200 642470
rect 299324 642370 299424 642470
rect 299548 642370 299648 642470
rect 299772 642370 299872 642470
rect 299996 642370 300096 642470
rect 300220 642370 300320 642470
rect 300444 642370 300544 642470
rect 300668 642370 300768 642470
rect 300892 642370 300992 642470
rect 301116 642370 301216 642470
rect 301340 642370 301440 642470
rect 301564 642370 301664 642470
rect 301788 642370 301888 642470
rect 302012 642370 302112 642470
rect 302236 642370 302336 642470
rect 302460 642370 302560 642470
rect 302684 642370 302784 642470
rect 302908 642370 303008 642470
rect 303132 642370 303232 642470
rect 303356 642370 303456 642470
rect 303580 642370 303680 642470
rect 303804 642370 303904 642470
rect 304028 642370 304128 642470
rect 304252 642370 304352 642470
rect 304476 642370 304576 642470
rect 304700 642370 304800 642470
rect 304924 642370 305024 642470
rect 305148 642370 305248 642470
rect 305372 642370 305472 642470
rect 298876 642146 298976 642246
rect 299100 642146 299200 642246
rect 299324 642146 299424 642246
rect 299548 642146 299648 642246
rect 299772 642146 299872 642246
rect 299996 642146 300096 642246
rect 300220 642146 300320 642246
rect 300444 642146 300544 642246
rect 300668 642146 300768 642246
rect 300892 642146 300992 642246
rect 301116 642146 301216 642246
rect 301340 642146 301440 642246
rect 301564 642146 301664 642246
rect 301788 642146 301888 642246
rect 302012 642146 302112 642246
rect 302236 642146 302336 642246
rect 302460 642146 302560 642246
rect 302684 642146 302784 642246
rect 302908 642146 303008 642246
rect 303132 642146 303232 642246
rect 303356 642146 303456 642246
rect 303580 642146 303680 642246
rect 303804 642146 303904 642246
rect 304028 642146 304128 642246
rect 304252 642146 304352 642246
rect 304476 642146 304576 642246
rect 304700 642146 304800 642246
rect 304924 642146 305024 642246
rect 305148 642146 305248 642246
rect 305372 642146 305472 642246
rect 298876 641922 298976 642022
rect 299100 641922 299200 642022
rect 299324 641922 299424 642022
rect 299548 641922 299648 642022
rect 299772 641922 299872 642022
rect 299996 641922 300096 642022
rect 300220 641922 300320 642022
rect 300444 641922 300544 642022
rect 300668 641922 300768 642022
rect 300892 641922 300992 642022
rect 301116 641922 301216 642022
rect 301340 641922 301440 642022
rect 301564 641922 301664 642022
rect 301788 641922 301888 642022
rect 302012 641922 302112 642022
rect 302236 641922 302336 642022
rect 302460 641922 302560 642022
rect 302684 641922 302784 642022
rect 302908 641922 303008 642022
rect 303132 641922 303232 642022
rect 303356 641922 303456 642022
rect 303580 641922 303680 642022
rect 303804 641922 303904 642022
rect 304028 641922 304128 642022
rect 304252 641922 304352 642022
rect 304476 641922 304576 642022
rect 304700 641922 304800 642022
rect 304924 641922 305024 642022
rect 305148 641922 305248 642022
rect 305372 641922 305472 642022
rect 298876 641698 298976 641798
rect 299100 641698 299200 641798
rect 299324 641698 299424 641798
rect 299548 641698 299648 641798
rect 299772 641698 299872 641798
rect 299996 641698 300096 641798
rect 300220 641698 300320 641798
rect 300444 641698 300544 641798
rect 300668 641698 300768 641798
rect 300892 641698 300992 641798
rect 301116 641698 301216 641798
rect 301340 641698 301440 641798
rect 301564 641698 301664 641798
rect 301788 641698 301888 641798
rect 302012 641698 302112 641798
rect 302236 641698 302336 641798
rect 302460 641698 302560 641798
rect 302684 641698 302784 641798
rect 302908 641698 303008 641798
rect 303132 641698 303232 641798
rect 303356 641698 303456 641798
rect 303580 641698 303680 641798
rect 303804 641698 303904 641798
rect 304028 641698 304128 641798
rect 304252 641698 304352 641798
rect 304476 641698 304576 641798
rect 304700 641698 304800 641798
rect 304924 641698 305024 641798
rect 305148 641698 305248 641798
rect 305372 641698 305472 641798
rect 309346 642594 309446 642694
rect 309570 642594 309670 642694
rect 309794 642594 309894 642694
rect 310018 642594 310118 642694
rect 310242 642594 310342 642694
rect 310466 642594 310566 642694
rect 310690 642594 310790 642694
rect 310914 642594 311014 642694
rect 311138 642594 311238 642694
rect 311362 642594 311462 642694
rect 311586 642594 311686 642694
rect 311810 642594 311910 642694
rect 312034 642594 312134 642694
rect 312258 642594 312358 642694
rect 312482 642594 312582 642694
rect 312706 642594 312806 642694
rect 312930 642594 313030 642694
rect 313154 642594 313254 642694
rect 313378 642594 313478 642694
rect 313602 642594 313702 642694
rect 313826 642594 313926 642694
rect 314050 642594 314150 642694
rect 314274 642594 314374 642694
rect 314498 642594 314598 642694
rect 314722 642594 314822 642694
rect 314946 642594 315046 642694
rect 315170 642594 315270 642694
rect 315394 642594 315494 642694
rect 315618 642594 315718 642694
rect 315842 642594 315942 642694
rect 309346 642370 309446 642470
rect 309570 642370 309670 642470
rect 309794 642370 309894 642470
rect 310018 642370 310118 642470
rect 310242 642370 310342 642470
rect 310466 642370 310566 642470
rect 310690 642370 310790 642470
rect 310914 642370 311014 642470
rect 311138 642370 311238 642470
rect 311362 642370 311462 642470
rect 311586 642370 311686 642470
rect 311810 642370 311910 642470
rect 312034 642370 312134 642470
rect 312258 642370 312358 642470
rect 312482 642370 312582 642470
rect 312706 642370 312806 642470
rect 312930 642370 313030 642470
rect 313154 642370 313254 642470
rect 313378 642370 313478 642470
rect 313602 642370 313702 642470
rect 313826 642370 313926 642470
rect 314050 642370 314150 642470
rect 314274 642370 314374 642470
rect 314498 642370 314598 642470
rect 314722 642370 314822 642470
rect 314946 642370 315046 642470
rect 315170 642370 315270 642470
rect 315394 642370 315494 642470
rect 315618 642370 315718 642470
rect 315842 642370 315942 642470
rect 309346 642146 309446 642246
rect 309570 642146 309670 642246
rect 309794 642146 309894 642246
rect 310018 642146 310118 642246
rect 310242 642146 310342 642246
rect 310466 642146 310566 642246
rect 310690 642146 310790 642246
rect 310914 642146 311014 642246
rect 311138 642146 311238 642246
rect 311362 642146 311462 642246
rect 311586 642146 311686 642246
rect 311810 642146 311910 642246
rect 312034 642146 312134 642246
rect 312258 642146 312358 642246
rect 312482 642146 312582 642246
rect 312706 642146 312806 642246
rect 312930 642146 313030 642246
rect 313154 642146 313254 642246
rect 313378 642146 313478 642246
rect 313602 642146 313702 642246
rect 313826 642146 313926 642246
rect 314050 642146 314150 642246
rect 314274 642146 314374 642246
rect 314498 642146 314598 642246
rect 314722 642146 314822 642246
rect 314946 642146 315046 642246
rect 315170 642146 315270 642246
rect 315394 642146 315494 642246
rect 315618 642146 315718 642246
rect 315842 642146 315942 642246
rect 309346 641922 309446 642022
rect 309570 641922 309670 642022
rect 309794 641922 309894 642022
rect 310018 641922 310118 642022
rect 310242 641922 310342 642022
rect 310466 641922 310566 642022
rect 310690 641922 310790 642022
rect 310914 641922 311014 642022
rect 311138 641922 311238 642022
rect 311362 641922 311462 642022
rect 311586 641922 311686 642022
rect 311810 641922 311910 642022
rect 312034 641922 312134 642022
rect 312258 641922 312358 642022
rect 312482 641922 312582 642022
rect 312706 641922 312806 642022
rect 312930 641922 313030 642022
rect 313154 641922 313254 642022
rect 313378 641922 313478 642022
rect 313602 641922 313702 642022
rect 313826 641922 313926 642022
rect 314050 641922 314150 642022
rect 314274 641922 314374 642022
rect 314498 641922 314598 642022
rect 314722 641922 314822 642022
rect 314946 641922 315046 642022
rect 315170 641922 315270 642022
rect 315394 641922 315494 642022
rect 315618 641922 315718 642022
rect 315842 641922 315942 642022
rect 309346 641698 309446 641798
rect 309570 641698 309670 641798
rect 309794 641698 309894 641798
rect 310018 641698 310118 641798
rect 310242 641698 310342 641798
rect 310466 641698 310566 641798
rect 310690 641698 310790 641798
rect 310914 641698 311014 641798
rect 311138 641698 311238 641798
rect 311362 641698 311462 641798
rect 311586 641698 311686 641798
rect 311810 641698 311910 641798
rect 312034 641698 312134 641798
rect 312258 641698 312358 641798
rect 312482 641698 312582 641798
rect 312706 641698 312806 641798
rect 312930 641698 313030 641798
rect 313154 641698 313254 641798
rect 313378 641698 313478 641798
rect 313602 641698 313702 641798
rect 313826 641698 313926 641798
rect 314050 641698 314150 641798
rect 314274 641698 314374 641798
rect 314498 641698 314598 641798
rect 314722 641698 314822 641798
rect 314946 641698 315046 641798
rect 315170 641698 315270 641798
rect 315394 641698 315494 641798
rect 315618 641698 315718 641798
rect 315842 641698 315942 641798
rect 335616 642614 335716 642714
rect 335840 642614 335940 642714
rect 336064 642614 336164 642714
rect 336288 642614 336388 642714
rect 336512 642614 336612 642714
rect 336736 642614 336836 642714
rect 336960 642614 337060 642714
rect 337184 642614 337284 642714
rect 337408 642614 337508 642714
rect 337632 642614 337732 642714
rect 337856 642614 337956 642714
rect 338080 642614 338180 642714
rect 338304 642614 338404 642714
rect 338528 642614 338628 642714
rect 338752 642614 338852 642714
rect 338976 642614 339076 642714
rect 339200 642614 339300 642714
rect 339424 642614 339524 642714
rect 339648 642614 339748 642714
rect 339872 642614 339972 642714
rect 340096 642614 340196 642714
rect 340320 642614 340420 642714
rect 340544 642614 340644 642714
rect 340768 642614 340868 642714
rect 340992 642614 341092 642714
rect 341216 642614 341316 642714
rect 341440 642614 341540 642714
rect 341664 642614 341764 642714
rect 341888 642614 341988 642714
rect 342112 642614 342212 642714
rect 335616 642390 335716 642490
rect 335840 642390 335940 642490
rect 336064 642390 336164 642490
rect 336288 642390 336388 642490
rect 336512 642390 336612 642490
rect 336736 642390 336836 642490
rect 336960 642390 337060 642490
rect 337184 642390 337284 642490
rect 337408 642390 337508 642490
rect 337632 642390 337732 642490
rect 337856 642390 337956 642490
rect 338080 642390 338180 642490
rect 338304 642390 338404 642490
rect 338528 642390 338628 642490
rect 338752 642390 338852 642490
rect 338976 642390 339076 642490
rect 339200 642390 339300 642490
rect 339424 642390 339524 642490
rect 339648 642390 339748 642490
rect 339872 642390 339972 642490
rect 340096 642390 340196 642490
rect 340320 642390 340420 642490
rect 340544 642390 340644 642490
rect 340768 642390 340868 642490
rect 340992 642390 341092 642490
rect 341216 642390 341316 642490
rect 341440 642390 341540 642490
rect 341664 642390 341764 642490
rect 341888 642390 341988 642490
rect 342112 642390 342212 642490
rect 335616 642166 335716 642266
rect 335840 642166 335940 642266
rect 336064 642166 336164 642266
rect 336288 642166 336388 642266
rect 336512 642166 336612 642266
rect 336736 642166 336836 642266
rect 336960 642166 337060 642266
rect 337184 642166 337284 642266
rect 337408 642166 337508 642266
rect 337632 642166 337732 642266
rect 337856 642166 337956 642266
rect 338080 642166 338180 642266
rect 338304 642166 338404 642266
rect 338528 642166 338628 642266
rect 338752 642166 338852 642266
rect 338976 642166 339076 642266
rect 339200 642166 339300 642266
rect 339424 642166 339524 642266
rect 339648 642166 339748 642266
rect 339872 642166 339972 642266
rect 340096 642166 340196 642266
rect 340320 642166 340420 642266
rect 340544 642166 340644 642266
rect 340768 642166 340868 642266
rect 340992 642166 341092 642266
rect 341216 642166 341316 642266
rect 341440 642166 341540 642266
rect 341664 642166 341764 642266
rect 341888 642166 341988 642266
rect 342112 642166 342212 642266
rect 335616 641942 335716 642042
rect 335840 641942 335940 642042
rect 336064 641942 336164 642042
rect 336288 641942 336388 642042
rect 336512 641942 336612 642042
rect 336736 641942 336836 642042
rect 336960 641942 337060 642042
rect 337184 641942 337284 642042
rect 337408 641942 337508 642042
rect 337632 641942 337732 642042
rect 337856 641942 337956 642042
rect 338080 641942 338180 642042
rect 338304 641942 338404 642042
rect 338528 641942 338628 642042
rect 338752 641942 338852 642042
rect 338976 641942 339076 642042
rect 339200 641942 339300 642042
rect 339424 641942 339524 642042
rect 339648 641942 339748 642042
rect 339872 641942 339972 642042
rect 340096 641942 340196 642042
rect 340320 641942 340420 642042
rect 340544 641942 340644 642042
rect 340768 641942 340868 642042
rect 340992 641942 341092 642042
rect 341216 641942 341316 642042
rect 341440 641942 341540 642042
rect 341664 641942 341764 642042
rect 341888 641942 341988 642042
rect 342112 641942 342212 642042
rect 335616 641718 335716 641818
rect 335840 641718 335940 641818
rect 336064 641718 336164 641818
rect 336288 641718 336388 641818
rect 336512 641718 336612 641818
rect 336736 641718 336836 641818
rect 336960 641718 337060 641818
rect 337184 641718 337284 641818
rect 337408 641718 337508 641818
rect 337632 641718 337732 641818
rect 337856 641718 337956 641818
rect 338080 641718 338180 641818
rect 338304 641718 338404 641818
rect 338528 641718 338628 641818
rect 338752 641718 338852 641818
rect 338976 641718 339076 641818
rect 339200 641718 339300 641818
rect 339424 641718 339524 641818
rect 339648 641718 339748 641818
rect 339872 641718 339972 641818
rect 340096 641718 340196 641818
rect 340320 641718 340420 641818
rect 340544 641718 340644 641818
rect 340768 641718 340868 641818
rect 340992 641718 341092 641818
rect 341216 641718 341316 641818
rect 341440 641718 341540 641818
rect 341664 641718 341764 641818
rect 341888 641718 341988 641818
rect 342112 641718 342212 641818
rect 297850 637896 297950 637996
rect 298074 637896 298174 637996
rect 298298 637896 298398 637996
rect 298522 637896 298622 637996
rect 298746 637896 298846 637996
rect 297850 637672 297950 637772
rect 298074 637672 298174 637772
rect 298298 637672 298398 637772
rect 298522 637672 298622 637772
rect 298746 637672 298846 637772
rect 297850 637448 297950 637548
rect 298074 637448 298174 637548
rect 298298 637448 298398 637548
rect 298522 637448 298622 637548
rect 298746 637448 298846 637548
rect 297850 637224 297950 637324
rect 298074 637224 298174 637324
rect 298298 637224 298398 637324
rect 298522 637224 298622 637324
rect 298746 637224 298846 637324
rect 297850 637000 297950 637100
rect 298074 637000 298174 637100
rect 298298 637000 298398 637100
rect 298522 637000 298622 637100
rect 298746 637000 298846 637100
rect 297850 636776 297950 636876
rect 298074 636776 298174 636876
rect 298298 636776 298398 636876
rect 298522 636776 298622 636876
rect 298746 636776 298846 636876
rect 297850 636552 297950 636652
rect 298074 636552 298174 636652
rect 298298 636552 298398 636652
rect 298522 636552 298622 636652
rect 298746 636552 298846 636652
rect 297850 636328 297950 636428
rect 298074 636328 298174 636428
rect 298298 636328 298398 636428
rect 298522 636328 298622 636428
rect 298746 636328 298846 636428
rect 297850 636104 297950 636204
rect 298074 636104 298174 636204
rect 298298 636104 298398 636204
rect 298522 636104 298622 636204
rect 298746 636104 298846 636204
rect 297850 635880 297950 635980
rect 298074 635880 298174 635980
rect 298298 635880 298398 635980
rect 298522 635880 298622 635980
rect 298746 635880 298846 635980
rect 297850 635656 297950 635756
rect 298074 635656 298174 635756
rect 298298 635656 298398 635756
rect 298522 635656 298622 635756
rect 298746 635656 298846 635756
rect 297850 635432 297950 635532
rect 298074 635432 298174 635532
rect 298298 635432 298398 635532
rect 298522 635432 298622 635532
rect 298746 635432 298846 635532
rect 297850 635208 297950 635308
rect 298074 635208 298174 635308
rect 298298 635208 298398 635308
rect 298522 635208 298622 635308
rect 298746 635208 298846 635308
rect 297850 634984 297950 635084
rect 298074 634984 298174 635084
rect 298298 634984 298398 635084
rect 298522 634984 298622 635084
rect 298746 634984 298846 635084
rect 297850 634760 297950 634860
rect 298074 634760 298174 634860
rect 298298 634760 298398 634860
rect 298522 634760 298622 634860
rect 298746 634760 298846 634860
rect 297850 634536 297950 634636
rect 298074 634536 298174 634636
rect 298298 634536 298398 634636
rect 298522 634536 298622 634636
rect 298746 634536 298846 634636
rect 297850 634312 297950 634412
rect 298074 634312 298174 634412
rect 298298 634312 298398 634412
rect 298522 634312 298622 634412
rect 298746 634312 298846 634412
rect 297850 634088 297950 634188
rect 298074 634088 298174 634188
rect 298298 634088 298398 634188
rect 298522 634088 298622 634188
rect 298746 634088 298846 634188
rect 297850 633864 297950 633964
rect 298074 633864 298174 633964
rect 298298 633864 298398 633964
rect 298522 633864 298622 633964
rect 298746 633864 298846 633964
rect 297850 633640 297950 633740
rect 298074 633640 298174 633740
rect 298298 633640 298398 633740
rect 298522 633640 298622 633740
rect 298746 633640 298846 633740
rect 297850 633416 297950 633516
rect 298074 633416 298174 633516
rect 298298 633416 298398 633516
rect 298522 633416 298622 633516
rect 298746 633416 298846 633516
rect 297850 633192 297950 633292
rect 298074 633192 298174 633292
rect 298298 633192 298398 633292
rect 298522 633192 298622 633292
rect 298746 633192 298846 633292
rect 297850 632968 297950 633068
rect 298074 632968 298174 633068
rect 298298 632968 298398 633068
rect 298522 632968 298622 633068
rect 298746 632968 298846 633068
rect 297850 632744 297950 632844
rect 298074 632744 298174 632844
rect 298298 632744 298398 632844
rect 298522 632744 298622 632844
rect 298746 632744 298846 632844
rect 297850 632520 297950 632620
rect 298074 632520 298174 632620
rect 298298 632520 298398 632620
rect 298522 632520 298622 632620
rect 298746 632520 298846 632620
rect 297850 632296 297950 632396
rect 298074 632296 298174 632396
rect 298298 632296 298398 632396
rect 298522 632296 298622 632396
rect 298746 632296 298846 632396
rect 297850 632072 297950 632172
rect 298074 632072 298174 632172
rect 298298 632072 298398 632172
rect 298522 632072 298622 632172
rect 298746 632072 298846 632172
rect 297850 631848 297950 631948
rect 298074 631848 298174 631948
rect 298298 631848 298398 631948
rect 298522 631848 298622 631948
rect 298746 631848 298846 631948
rect 297850 631624 297950 631724
rect 298074 631624 298174 631724
rect 298298 631624 298398 631724
rect 298522 631624 298622 631724
rect 298746 631624 298846 631724
rect 297850 631400 297950 631500
rect 298074 631400 298174 631500
rect 298298 631400 298398 631500
rect 298522 631400 298622 631500
rect 298746 631400 298846 631500
rect 342130 637896 342230 637996
rect 342354 637896 342454 637996
rect 342578 637896 342678 637996
rect 342802 637896 342902 637996
rect 343026 637896 343126 637996
rect 342130 637672 342230 637772
rect 342354 637672 342454 637772
rect 342578 637672 342678 637772
rect 342802 637672 342902 637772
rect 343026 637672 343126 637772
rect 342130 637448 342230 637548
rect 342354 637448 342454 637548
rect 342578 637448 342678 637548
rect 342802 637448 342902 637548
rect 343026 637448 343126 637548
rect 342130 637224 342230 637324
rect 342354 637224 342454 637324
rect 342578 637224 342678 637324
rect 342802 637224 342902 637324
rect 343026 637224 343126 637324
rect 342130 637000 342230 637100
rect 342354 637000 342454 637100
rect 342578 637000 342678 637100
rect 342802 637000 342902 637100
rect 343026 637000 343126 637100
rect 342130 636776 342230 636876
rect 342354 636776 342454 636876
rect 342578 636776 342678 636876
rect 342802 636776 342902 636876
rect 343026 636776 343126 636876
rect 342130 636552 342230 636652
rect 342354 636552 342454 636652
rect 342578 636552 342678 636652
rect 342802 636552 342902 636652
rect 343026 636552 343126 636652
rect 342130 636328 342230 636428
rect 342354 636328 342454 636428
rect 342578 636328 342678 636428
rect 342802 636328 342902 636428
rect 343026 636328 343126 636428
rect 342130 636104 342230 636204
rect 342354 636104 342454 636204
rect 342578 636104 342678 636204
rect 342802 636104 342902 636204
rect 343026 636104 343126 636204
rect 342130 635880 342230 635980
rect 342354 635880 342454 635980
rect 342578 635880 342678 635980
rect 342802 635880 342902 635980
rect 343026 635880 343126 635980
rect 342130 635656 342230 635756
rect 342354 635656 342454 635756
rect 342578 635656 342678 635756
rect 342802 635656 342902 635756
rect 343026 635656 343126 635756
rect 342130 635432 342230 635532
rect 342354 635432 342454 635532
rect 342578 635432 342678 635532
rect 342802 635432 342902 635532
rect 343026 635432 343126 635532
rect 342130 635208 342230 635308
rect 342354 635208 342454 635308
rect 342578 635208 342678 635308
rect 342802 635208 342902 635308
rect 343026 635208 343126 635308
rect 342130 634984 342230 635084
rect 342354 634984 342454 635084
rect 342578 634984 342678 635084
rect 342802 634984 342902 635084
rect 343026 634984 343126 635084
rect 342130 634760 342230 634860
rect 342354 634760 342454 634860
rect 342578 634760 342678 634860
rect 342802 634760 342902 634860
rect 343026 634760 343126 634860
rect 342130 634536 342230 634636
rect 342354 634536 342454 634636
rect 342578 634536 342678 634636
rect 342802 634536 342902 634636
rect 343026 634536 343126 634636
rect 342130 634312 342230 634412
rect 342354 634312 342454 634412
rect 342578 634312 342678 634412
rect 342802 634312 342902 634412
rect 343026 634312 343126 634412
rect 342130 634088 342230 634188
rect 342354 634088 342454 634188
rect 342578 634088 342678 634188
rect 342802 634088 342902 634188
rect 343026 634088 343126 634188
rect 342130 633864 342230 633964
rect 342354 633864 342454 633964
rect 342578 633864 342678 633964
rect 342802 633864 342902 633964
rect 343026 633864 343126 633964
rect 342130 633640 342230 633740
rect 342354 633640 342454 633740
rect 342578 633640 342678 633740
rect 342802 633640 342902 633740
rect 343026 633640 343126 633740
rect 342130 633416 342230 633516
rect 342354 633416 342454 633516
rect 342578 633416 342678 633516
rect 342802 633416 342902 633516
rect 343026 633416 343126 633516
rect 342130 633192 342230 633292
rect 342354 633192 342454 633292
rect 342578 633192 342678 633292
rect 342802 633192 342902 633292
rect 343026 633192 343126 633292
rect 342130 632968 342230 633068
rect 342354 632968 342454 633068
rect 342578 632968 342678 633068
rect 342802 632968 342902 633068
rect 343026 632968 343126 633068
rect 342130 632744 342230 632844
rect 342354 632744 342454 632844
rect 342578 632744 342678 632844
rect 342802 632744 342902 632844
rect 343026 632744 343126 632844
rect 342130 632520 342230 632620
rect 342354 632520 342454 632620
rect 342578 632520 342678 632620
rect 342802 632520 342902 632620
rect 343026 632520 343126 632620
rect 342130 632296 342230 632396
rect 342354 632296 342454 632396
rect 342578 632296 342678 632396
rect 342802 632296 342902 632396
rect 343026 632296 343126 632396
rect 342130 632072 342230 632172
rect 342354 632072 342454 632172
rect 342578 632072 342678 632172
rect 342802 632072 342902 632172
rect 343026 632072 343126 632172
rect 342130 631848 342230 631948
rect 342354 631848 342454 631948
rect 342578 631848 342678 631948
rect 342802 631848 342902 631948
rect 343026 631848 343126 631948
rect 342130 631624 342230 631724
rect 342354 631624 342454 631724
rect 342578 631624 342678 631724
rect 342802 631624 342902 631724
rect 343026 631624 343126 631724
rect 342130 631400 342230 631500
rect 342354 631400 342454 631500
rect 342578 631400 342678 631500
rect 342802 631400 342902 631500
rect 343026 631400 343126 631500
rect 319400 628668 319600 628868
rect 319834 628668 320034 628868
rect 320268 628668 320468 628868
rect 320702 628668 320902 628868
rect 321136 628668 321336 628868
rect 321570 628668 321770 628868
rect 322004 628668 322204 628868
rect 322438 628668 322638 628868
rect 322872 628668 323072 628868
rect 323306 628668 323506 628868
rect 323740 628668 323940 628868
rect 324140 628668 324340 628868
rect 324540 628668 324740 628868
rect 324940 628668 325140 628868
rect 325340 628668 325540 628868
rect 325740 628668 325940 628868
rect 326140 628668 326340 628868
rect 326540 628668 326740 628868
rect 326940 628668 327140 628868
rect 327340 628668 327540 628868
rect 328940 628668 329140 628868
rect 329340 628668 329540 628868
rect 329740 628668 329940 628868
rect 330140 628668 330340 628868
rect 330540 628668 330740 628868
rect 330940 628668 331140 628868
rect 331340 628668 331540 628868
rect 331740 628668 331940 628868
rect 332140 628668 332340 628868
rect 319400 628234 319600 628434
rect 319834 628234 320034 628434
rect 320268 628234 320468 628434
rect 320702 628234 320902 628434
rect 321136 628234 321336 628434
rect 321570 628234 321770 628434
rect 322004 628234 322204 628434
rect 322438 628234 322638 628434
rect 322872 628234 323072 628434
rect 323306 628234 323506 628434
rect 323740 628234 323940 628434
rect 319400 627800 319600 628000
rect 319834 627800 320034 628000
rect 320268 627800 320468 628000
rect 320702 627800 320902 628000
rect 321136 627800 321336 628000
rect 321570 627800 321770 628000
rect 322004 627800 322204 628000
rect 322438 627800 322638 628000
rect 322872 627800 323072 628000
rect 323306 627800 323506 628000
rect 323740 627800 323940 628000
rect 297850 624496 297950 624596
rect 298074 624496 298174 624596
rect 298298 624496 298398 624596
rect 298522 624496 298622 624596
rect 298746 624496 298846 624596
rect 297850 624272 297950 624372
rect 298074 624272 298174 624372
rect 298298 624272 298398 624372
rect 298522 624272 298622 624372
rect 298746 624272 298846 624372
rect 342130 624496 342230 624596
rect 342354 624496 342454 624596
rect 342578 624496 342678 624596
rect 342802 624496 342902 624596
rect 343026 624496 343126 624596
rect 342130 624272 342230 624372
rect 342354 624272 342454 624372
rect 342578 624272 342678 624372
rect 342802 624272 342902 624372
rect 343026 624272 343126 624372
rect 297850 624048 297950 624148
rect 298074 624048 298174 624148
rect 298298 624048 298398 624148
rect 298522 624048 298622 624148
rect 298746 624048 298846 624148
rect 302972 624114 303032 624184
rect 303044 624114 303104 624184
rect 303116 624114 303176 624184
rect 303188 624114 303248 624184
rect 303260 624114 303320 624184
rect 303332 624114 303392 624184
rect 303404 624114 303464 624184
rect 303476 624114 303536 624184
rect 302972 624020 303032 624090
rect 303044 624020 303104 624090
rect 303116 624020 303176 624090
rect 303188 624020 303248 624090
rect 303260 624020 303320 624090
rect 303332 624020 303392 624090
rect 303404 624020 303464 624090
rect 303476 624020 303536 624090
rect 342130 624048 342230 624148
rect 342354 624048 342454 624148
rect 342578 624048 342678 624148
rect 342802 624048 342902 624148
rect 343026 624048 343126 624148
rect 297850 623824 297950 623924
rect 298074 623824 298174 623924
rect 298298 623824 298398 623924
rect 298522 623824 298622 623924
rect 298746 623824 298846 623924
rect 297850 623600 297950 623700
rect 298074 623600 298174 623700
rect 298298 623600 298398 623700
rect 298522 623600 298622 623700
rect 298746 623600 298846 623700
rect 297850 623376 297950 623476
rect 298074 623376 298174 623476
rect 298298 623376 298398 623476
rect 298522 623376 298622 623476
rect 298746 623376 298846 623476
rect 297850 623152 297950 623252
rect 298074 623152 298174 623252
rect 298298 623152 298398 623252
rect 298522 623152 298622 623252
rect 298746 623152 298846 623252
rect 297850 622928 297950 623028
rect 298074 622928 298174 623028
rect 298298 622928 298398 623028
rect 298522 622928 298622 623028
rect 298746 622928 298846 623028
rect 297850 622704 297950 622804
rect 298074 622704 298174 622804
rect 298298 622704 298398 622804
rect 298522 622704 298622 622804
rect 298746 622704 298846 622804
rect 297850 622480 297950 622580
rect 298074 622480 298174 622580
rect 298298 622480 298398 622580
rect 298522 622480 298622 622580
rect 298746 622480 298846 622580
rect 297850 622256 297950 622356
rect 298074 622256 298174 622356
rect 298298 622256 298398 622356
rect 298522 622256 298622 622356
rect 298746 622256 298846 622356
rect 297850 622032 297950 622132
rect 298074 622032 298174 622132
rect 298298 622032 298398 622132
rect 298522 622032 298622 622132
rect 298746 622032 298846 622132
rect 297850 621808 297950 621908
rect 298074 621808 298174 621908
rect 298298 621808 298398 621908
rect 298522 621808 298622 621908
rect 298746 621808 298846 621908
rect 297850 621584 297950 621684
rect 298074 621584 298174 621684
rect 298298 621584 298398 621684
rect 298522 621584 298622 621684
rect 298746 621584 298846 621684
rect 297850 621360 297950 621460
rect 298074 621360 298174 621460
rect 298298 621360 298398 621460
rect 298522 621360 298622 621460
rect 298746 621360 298846 621460
rect 297850 621136 297950 621236
rect 298074 621136 298174 621236
rect 298298 621136 298398 621236
rect 298522 621136 298622 621236
rect 298746 621136 298846 621236
rect 297850 620912 297950 621012
rect 298074 620912 298174 621012
rect 298298 620912 298398 621012
rect 298522 620912 298622 621012
rect 298746 620912 298846 621012
rect 297850 620688 297950 620788
rect 298074 620688 298174 620788
rect 298298 620688 298398 620788
rect 298522 620688 298622 620788
rect 298746 620688 298846 620788
rect 297850 620464 297950 620564
rect 298074 620464 298174 620564
rect 298298 620464 298398 620564
rect 298522 620464 298622 620564
rect 298746 620464 298846 620564
rect 297850 620240 297950 620340
rect 298074 620240 298174 620340
rect 298298 620240 298398 620340
rect 298522 620240 298622 620340
rect 298746 620240 298846 620340
rect 297850 620016 297950 620116
rect 298074 620016 298174 620116
rect 298298 620016 298398 620116
rect 298522 620016 298622 620116
rect 298746 620016 298846 620116
rect 297850 619792 297950 619892
rect 298074 619792 298174 619892
rect 298298 619792 298398 619892
rect 298522 619792 298622 619892
rect 298746 619792 298846 619892
rect 297850 619568 297950 619668
rect 298074 619568 298174 619668
rect 298298 619568 298398 619668
rect 298522 619568 298622 619668
rect 298746 619568 298846 619668
rect 297850 619344 297950 619444
rect 298074 619344 298174 619444
rect 298298 619344 298398 619444
rect 298522 619344 298622 619444
rect 298746 619344 298846 619444
rect 297850 619120 297950 619220
rect 298074 619120 298174 619220
rect 298298 619120 298398 619220
rect 298522 619120 298622 619220
rect 298746 619120 298846 619220
rect 297850 618896 297950 618996
rect 298074 618896 298174 618996
rect 298298 618896 298398 618996
rect 298522 618896 298622 618996
rect 298746 618896 298846 618996
rect 297850 618672 297950 618772
rect 298074 618672 298174 618772
rect 298298 618672 298398 618772
rect 298522 618672 298622 618772
rect 298746 618672 298846 618772
rect 297850 618448 297950 618548
rect 298074 618448 298174 618548
rect 298298 618448 298398 618548
rect 298522 618448 298622 618548
rect 298746 618448 298846 618548
rect 297850 618224 297950 618324
rect 298074 618224 298174 618324
rect 298298 618224 298398 618324
rect 298522 618224 298622 618324
rect 298746 618224 298846 618324
rect 297850 618000 297950 618100
rect 298074 618000 298174 618100
rect 298298 618000 298398 618100
rect 298522 618000 298622 618100
rect 298746 618000 298846 618100
rect 342130 623824 342230 623924
rect 342354 623824 342454 623924
rect 342578 623824 342678 623924
rect 342802 623824 342902 623924
rect 343026 623824 343126 623924
rect 342130 623600 342230 623700
rect 342354 623600 342454 623700
rect 342578 623600 342678 623700
rect 342802 623600 342902 623700
rect 343026 623600 343126 623700
rect 342130 623376 342230 623476
rect 342354 623376 342454 623476
rect 342578 623376 342678 623476
rect 342802 623376 342902 623476
rect 343026 623376 343126 623476
rect 342130 623152 342230 623252
rect 342354 623152 342454 623252
rect 342578 623152 342678 623252
rect 342802 623152 342902 623252
rect 343026 623152 343126 623252
rect 342130 622928 342230 623028
rect 342354 622928 342454 623028
rect 342578 622928 342678 623028
rect 342802 622928 342902 623028
rect 343026 622928 343126 623028
rect 342130 622704 342230 622804
rect 342354 622704 342454 622804
rect 342578 622704 342678 622804
rect 342802 622704 342902 622804
rect 343026 622704 343126 622804
rect 342130 622480 342230 622580
rect 342354 622480 342454 622580
rect 342578 622480 342678 622580
rect 342802 622480 342902 622580
rect 343026 622480 343126 622580
rect 342130 622256 342230 622356
rect 342354 622256 342454 622356
rect 342578 622256 342678 622356
rect 342802 622256 342902 622356
rect 343026 622256 343126 622356
rect 342130 622032 342230 622132
rect 342354 622032 342454 622132
rect 342578 622032 342678 622132
rect 342802 622032 342902 622132
rect 343026 622032 343126 622132
rect 342130 621808 342230 621908
rect 342354 621808 342454 621908
rect 342578 621808 342678 621908
rect 342802 621808 342902 621908
rect 343026 621808 343126 621908
rect 342130 621584 342230 621684
rect 342354 621584 342454 621684
rect 342578 621584 342678 621684
rect 342802 621584 342902 621684
rect 343026 621584 343126 621684
rect 342130 621360 342230 621460
rect 342354 621360 342454 621460
rect 342578 621360 342678 621460
rect 342802 621360 342902 621460
rect 343026 621360 343126 621460
rect 342130 621136 342230 621236
rect 342354 621136 342454 621236
rect 342578 621136 342678 621236
rect 342802 621136 342902 621236
rect 343026 621136 343126 621236
rect 342130 620912 342230 621012
rect 342354 620912 342454 621012
rect 342578 620912 342678 621012
rect 342802 620912 342902 621012
rect 343026 620912 343126 621012
rect 342130 620688 342230 620788
rect 342354 620688 342454 620788
rect 342578 620688 342678 620788
rect 342802 620688 342902 620788
rect 343026 620688 343126 620788
rect 342130 620464 342230 620564
rect 342354 620464 342454 620564
rect 342578 620464 342678 620564
rect 342802 620464 342902 620564
rect 343026 620464 343126 620564
rect 342130 620240 342230 620340
rect 342354 620240 342454 620340
rect 342578 620240 342678 620340
rect 342802 620240 342902 620340
rect 343026 620240 343126 620340
rect 342130 620016 342230 620116
rect 342354 620016 342454 620116
rect 342578 620016 342678 620116
rect 342802 620016 342902 620116
rect 343026 620016 343126 620116
rect 342130 619792 342230 619892
rect 342354 619792 342454 619892
rect 342578 619792 342678 619892
rect 342802 619792 342902 619892
rect 343026 619792 343126 619892
rect 342130 619568 342230 619668
rect 342354 619568 342454 619668
rect 342578 619568 342678 619668
rect 342802 619568 342902 619668
rect 343026 619568 343126 619668
rect 342130 619344 342230 619444
rect 342354 619344 342454 619444
rect 342578 619344 342678 619444
rect 342802 619344 342902 619444
rect 343026 619344 343126 619444
rect 342130 619120 342230 619220
rect 342354 619120 342454 619220
rect 342578 619120 342678 619220
rect 342802 619120 342902 619220
rect 343026 619120 343126 619220
rect 342130 618896 342230 618996
rect 342354 618896 342454 618996
rect 342578 618896 342678 618996
rect 342802 618896 342902 618996
rect 343026 618896 343126 618996
rect 342130 618672 342230 618772
rect 342354 618672 342454 618772
rect 342578 618672 342678 618772
rect 342802 618672 342902 618772
rect 343026 618672 343126 618772
rect 342130 618448 342230 618548
rect 342354 618448 342454 618548
rect 342578 618448 342678 618548
rect 342802 618448 342902 618548
rect 343026 618448 343126 618548
rect 342130 618224 342230 618324
rect 342354 618224 342454 618324
rect 342578 618224 342678 618324
rect 342802 618224 342902 618324
rect 343026 618224 343126 618324
rect 342130 618000 342230 618100
rect 342354 618000 342454 618100
rect 342578 618000 342678 618100
rect 342802 618000 342902 618100
rect 343026 618000 343126 618100
rect 298876 615374 298976 615474
rect 299100 615374 299200 615474
rect 299324 615374 299424 615474
rect 299548 615374 299648 615474
rect 299772 615374 299872 615474
rect 299996 615374 300096 615474
rect 300220 615374 300320 615474
rect 300444 615374 300544 615474
rect 300668 615374 300768 615474
rect 300892 615374 300992 615474
rect 301116 615374 301216 615474
rect 301340 615374 301440 615474
rect 301564 615374 301664 615474
rect 301788 615374 301888 615474
rect 302012 615374 302112 615474
rect 302236 615374 302336 615474
rect 302460 615374 302560 615474
rect 302684 615374 302784 615474
rect 302908 615374 303008 615474
rect 303132 615374 303232 615474
rect 303356 615374 303456 615474
rect 303580 615374 303680 615474
rect 303804 615374 303904 615474
rect 304028 615374 304128 615474
rect 304252 615374 304352 615474
rect 304476 615374 304576 615474
rect 304700 615374 304800 615474
rect 304924 615374 305024 615474
rect 305148 615374 305248 615474
rect 305372 615374 305472 615474
rect 298876 615150 298976 615250
rect 299100 615150 299200 615250
rect 299324 615150 299424 615250
rect 299548 615150 299648 615250
rect 299772 615150 299872 615250
rect 299996 615150 300096 615250
rect 300220 615150 300320 615250
rect 300444 615150 300544 615250
rect 300668 615150 300768 615250
rect 300892 615150 300992 615250
rect 301116 615150 301216 615250
rect 301340 615150 301440 615250
rect 301564 615150 301664 615250
rect 301788 615150 301888 615250
rect 302012 615150 302112 615250
rect 302236 615150 302336 615250
rect 302460 615150 302560 615250
rect 302684 615150 302784 615250
rect 302908 615150 303008 615250
rect 303132 615150 303232 615250
rect 303356 615150 303456 615250
rect 303580 615150 303680 615250
rect 303804 615150 303904 615250
rect 304028 615150 304128 615250
rect 304252 615150 304352 615250
rect 304476 615150 304576 615250
rect 304700 615150 304800 615250
rect 304924 615150 305024 615250
rect 305148 615150 305248 615250
rect 305372 615150 305472 615250
rect 298876 614926 298976 615026
rect 299100 614926 299200 615026
rect 299324 614926 299424 615026
rect 299548 614926 299648 615026
rect 299772 614926 299872 615026
rect 299996 614926 300096 615026
rect 300220 614926 300320 615026
rect 300444 614926 300544 615026
rect 300668 614926 300768 615026
rect 300892 614926 300992 615026
rect 301116 614926 301216 615026
rect 301340 614926 301440 615026
rect 301564 614926 301664 615026
rect 301788 614926 301888 615026
rect 302012 614926 302112 615026
rect 302236 614926 302336 615026
rect 302460 614926 302560 615026
rect 302684 614926 302784 615026
rect 302908 614926 303008 615026
rect 303132 614926 303232 615026
rect 303356 614926 303456 615026
rect 303580 614926 303680 615026
rect 303804 614926 303904 615026
rect 304028 614926 304128 615026
rect 304252 614926 304352 615026
rect 304476 614926 304576 615026
rect 304700 614926 304800 615026
rect 304924 614926 305024 615026
rect 305148 614926 305248 615026
rect 305372 614926 305472 615026
rect 298876 614702 298976 614802
rect 299100 614702 299200 614802
rect 299324 614702 299424 614802
rect 299548 614702 299648 614802
rect 299772 614702 299872 614802
rect 299996 614702 300096 614802
rect 300220 614702 300320 614802
rect 300444 614702 300544 614802
rect 300668 614702 300768 614802
rect 300892 614702 300992 614802
rect 301116 614702 301216 614802
rect 301340 614702 301440 614802
rect 301564 614702 301664 614802
rect 301788 614702 301888 614802
rect 302012 614702 302112 614802
rect 302236 614702 302336 614802
rect 302460 614702 302560 614802
rect 302684 614702 302784 614802
rect 302908 614702 303008 614802
rect 303132 614702 303232 614802
rect 303356 614702 303456 614802
rect 303580 614702 303680 614802
rect 303804 614702 303904 614802
rect 304028 614702 304128 614802
rect 304252 614702 304352 614802
rect 304476 614702 304576 614802
rect 304700 614702 304800 614802
rect 304924 614702 305024 614802
rect 305148 614702 305248 614802
rect 305372 614702 305472 614802
rect 298876 614478 298976 614578
rect 299100 614478 299200 614578
rect 299324 614478 299424 614578
rect 299548 614478 299648 614578
rect 299772 614478 299872 614578
rect 299996 614478 300096 614578
rect 300220 614478 300320 614578
rect 300444 614478 300544 614578
rect 300668 614478 300768 614578
rect 300892 614478 300992 614578
rect 301116 614478 301216 614578
rect 301340 614478 301440 614578
rect 301564 614478 301664 614578
rect 301788 614478 301888 614578
rect 302012 614478 302112 614578
rect 302236 614478 302336 614578
rect 302460 614478 302560 614578
rect 302684 614478 302784 614578
rect 302908 614478 303008 614578
rect 303132 614478 303232 614578
rect 303356 614478 303456 614578
rect 303580 614478 303680 614578
rect 303804 614478 303904 614578
rect 304028 614478 304128 614578
rect 304252 614478 304352 614578
rect 304476 614478 304576 614578
rect 304700 614478 304800 614578
rect 304924 614478 305024 614578
rect 305148 614478 305248 614578
rect 305372 614478 305472 614578
rect 309346 615374 309446 615474
rect 309570 615374 309670 615474
rect 309794 615374 309894 615474
rect 310018 615374 310118 615474
rect 310242 615374 310342 615474
rect 310466 615374 310566 615474
rect 310690 615374 310790 615474
rect 310914 615374 311014 615474
rect 311138 615374 311238 615474
rect 311362 615374 311462 615474
rect 311586 615374 311686 615474
rect 311810 615374 311910 615474
rect 312034 615374 312134 615474
rect 312258 615374 312358 615474
rect 312482 615374 312582 615474
rect 312706 615374 312806 615474
rect 312930 615374 313030 615474
rect 313154 615374 313254 615474
rect 313378 615374 313478 615474
rect 313602 615374 313702 615474
rect 313826 615374 313926 615474
rect 314050 615374 314150 615474
rect 314274 615374 314374 615474
rect 314498 615374 314598 615474
rect 314722 615374 314822 615474
rect 314946 615374 315046 615474
rect 315170 615374 315270 615474
rect 315394 615374 315494 615474
rect 315618 615374 315718 615474
rect 315842 615374 315942 615474
rect 309346 615150 309446 615250
rect 309570 615150 309670 615250
rect 309794 615150 309894 615250
rect 310018 615150 310118 615250
rect 310242 615150 310342 615250
rect 310466 615150 310566 615250
rect 310690 615150 310790 615250
rect 310914 615150 311014 615250
rect 311138 615150 311238 615250
rect 311362 615150 311462 615250
rect 311586 615150 311686 615250
rect 311810 615150 311910 615250
rect 312034 615150 312134 615250
rect 312258 615150 312358 615250
rect 312482 615150 312582 615250
rect 312706 615150 312806 615250
rect 312930 615150 313030 615250
rect 313154 615150 313254 615250
rect 313378 615150 313478 615250
rect 313602 615150 313702 615250
rect 313826 615150 313926 615250
rect 314050 615150 314150 615250
rect 314274 615150 314374 615250
rect 314498 615150 314598 615250
rect 314722 615150 314822 615250
rect 314946 615150 315046 615250
rect 315170 615150 315270 615250
rect 315394 615150 315494 615250
rect 315618 615150 315718 615250
rect 315842 615150 315942 615250
rect 309346 614926 309446 615026
rect 309570 614926 309670 615026
rect 309794 614926 309894 615026
rect 310018 614926 310118 615026
rect 310242 614926 310342 615026
rect 310466 614926 310566 615026
rect 310690 614926 310790 615026
rect 310914 614926 311014 615026
rect 311138 614926 311238 615026
rect 311362 614926 311462 615026
rect 311586 614926 311686 615026
rect 311810 614926 311910 615026
rect 312034 614926 312134 615026
rect 312258 614926 312358 615026
rect 312482 614926 312582 615026
rect 312706 614926 312806 615026
rect 312930 614926 313030 615026
rect 313154 614926 313254 615026
rect 313378 614926 313478 615026
rect 313602 614926 313702 615026
rect 313826 614926 313926 615026
rect 314050 614926 314150 615026
rect 314274 614926 314374 615026
rect 314498 614926 314598 615026
rect 314722 614926 314822 615026
rect 314946 614926 315046 615026
rect 315170 614926 315270 615026
rect 315394 614926 315494 615026
rect 315618 614926 315718 615026
rect 315842 614926 315942 615026
rect 309346 614702 309446 614802
rect 309570 614702 309670 614802
rect 309794 614702 309894 614802
rect 310018 614702 310118 614802
rect 310242 614702 310342 614802
rect 310466 614702 310566 614802
rect 310690 614702 310790 614802
rect 310914 614702 311014 614802
rect 311138 614702 311238 614802
rect 311362 614702 311462 614802
rect 311586 614702 311686 614802
rect 311810 614702 311910 614802
rect 312034 614702 312134 614802
rect 312258 614702 312358 614802
rect 312482 614702 312582 614802
rect 312706 614702 312806 614802
rect 312930 614702 313030 614802
rect 313154 614702 313254 614802
rect 313378 614702 313478 614802
rect 313602 614702 313702 614802
rect 313826 614702 313926 614802
rect 314050 614702 314150 614802
rect 314274 614702 314374 614802
rect 314498 614702 314598 614802
rect 314722 614702 314822 614802
rect 314946 614702 315046 614802
rect 315170 614702 315270 614802
rect 315394 614702 315494 614802
rect 315618 614702 315718 614802
rect 315842 614702 315942 614802
rect 309346 614478 309446 614578
rect 309570 614478 309670 614578
rect 309794 614478 309894 614578
rect 310018 614478 310118 614578
rect 310242 614478 310342 614578
rect 310466 614478 310566 614578
rect 310690 614478 310790 614578
rect 310914 614478 311014 614578
rect 311138 614478 311238 614578
rect 311362 614478 311462 614578
rect 311586 614478 311686 614578
rect 311810 614478 311910 614578
rect 312034 614478 312134 614578
rect 312258 614478 312358 614578
rect 312482 614478 312582 614578
rect 312706 614478 312806 614578
rect 312930 614478 313030 614578
rect 313154 614478 313254 614578
rect 313378 614478 313478 614578
rect 313602 614478 313702 614578
rect 313826 614478 313926 614578
rect 314050 614478 314150 614578
rect 314274 614478 314374 614578
rect 314498 614478 314598 614578
rect 314722 614478 314822 614578
rect 314946 614478 315046 614578
rect 315170 614478 315270 614578
rect 315394 614478 315494 614578
rect 315618 614478 315718 614578
rect 315842 614478 315942 614578
rect 335616 615394 335716 615494
rect 335840 615394 335940 615494
rect 336064 615394 336164 615494
rect 336288 615394 336388 615494
rect 336512 615394 336612 615494
rect 336736 615394 336836 615494
rect 336960 615394 337060 615494
rect 337184 615394 337284 615494
rect 337408 615394 337508 615494
rect 337632 615394 337732 615494
rect 337856 615394 337956 615494
rect 338080 615394 338180 615494
rect 338304 615394 338404 615494
rect 338528 615394 338628 615494
rect 338752 615394 338852 615494
rect 338976 615394 339076 615494
rect 339200 615394 339300 615494
rect 339424 615394 339524 615494
rect 339648 615394 339748 615494
rect 339872 615394 339972 615494
rect 340096 615394 340196 615494
rect 340320 615394 340420 615494
rect 340544 615394 340644 615494
rect 340768 615394 340868 615494
rect 340992 615394 341092 615494
rect 341216 615394 341316 615494
rect 341440 615394 341540 615494
rect 341664 615394 341764 615494
rect 341888 615394 341988 615494
rect 342112 615394 342212 615494
rect 335616 615170 335716 615270
rect 335840 615170 335940 615270
rect 336064 615170 336164 615270
rect 336288 615170 336388 615270
rect 336512 615170 336612 615270
rect 336736 615170 336836 615270
rect 336960 615170 337060 615270
rect 337184 615170 337284 615270
rect 337408 615170 337508 615270
rect 337632 615170 337732 615270
rect 337856 615170 337956 615270
rect 338080 615170 338180 615270
rect 338304 615170 338404 615270
rect 338528 615170 338628 615270
rect 338752 615170 338852 615270
rect 338976 615170 339076 615270
rect 339200 615170 339300 615270
rect 339424 615170 339524 615270
rect 339648 615170 339748 615270
rect 339872 615170 339972 615270
rect 340096 615170 340196 615270
rect 340320 615170 340420 615270
rect 340544 615170 340644 615270
rect 340768 615170 340868 615270
rect 340992 615170 341092 615270
rect 341216 615170 341316 615270
rect 341440 615170 341540 615270
rect 341664 615170 341764 615270
rect 341888 615170 341988 615270
rect 342112 615170 342212 615270
rect 335616 614946 335716 615046
rect 335840 614946 335940 615046
rect 336064 614946 336164 615046
rect 336288 614946 336388 615046
rect 336512 614946 336612 615046
rect 336736 614946 336836 615046
rect 336960 614946 337060 615046
rect 337184 614946 337284 615046
rect 337408 614946 337508 615046
rect 337632 614946 337732 615046
rect 337856 614946 337956 615046
rect 338080 614946 338180 615046
rect 338304 614946 338404 615046
rect 338528 614946 338628 615046
rect 338752 614946 338852 615046
rect 338976 614946 339076 615046
rect 339200 614946 339300 615046
rect 339424 614946 339524 615046
rect 339648 614946 339748 615046
rect 339872 614946 339972 615046
rect 340096 614946 340196 615046
rect 340320 614946 340420 615046
rect 340544 614946 340644 615046
rect 340768 614946 340868 615046
rect 340992 614946 341092 615046
rect 341216 614946 341316 615046
rect 341440 614946 341540 615046
rect 341664 614946 341764 615046
rect 341888 614946 341988 615046
rect 342112 614946 342212 615046
rect 335616 614722 335716 614822
rect 335840 614722 335940 614822
rect 336064 614722 336164 614822
rect 336288 614722 336388 614822
rect 336512 614722 336612 614822
rect 336736 614722 336836 614822
rect 336960 614722 337060 614822
rect 337184 614722 337284 614822
rect 337408 614722 337508 614822
rect 337632 614722 337732 614822
rect 337856 614722 337956 614822
rect 338080 614722 338180 614822
rect 338304 614722 338404 614822
rect 338528 614722 338628 614822
rect 338752 614722 338852 614822
rect 338976 614722 339076 614822
rect 339200 614722 339300 614822
rect 339424 614722 339524 614822
rect 339648 614722 339748 614822
rect 339872 614722 339972 614822
rect 340096 614722 340196 614822
rect 340320 614722 340420 614822
rect 340544 614722 340644 614822
rect 340768 614722 340868 614822
rect 340992 614722 341092 614822
rect 341216 614722 341316 614822
rect 341440 614722 341540 614822
rect 341664 614722 341764 614822
rect 341888 614722 341988 614822
rect 342112 614722 342212 614822
rect 335616 614498 335716 614598
rect 335840 614498 335940 614598
rect 336064 614498 336164 614598
rect 336288 614498 336388 614598
rect 336512 614498 336612 614598
rect 336736 614498 336836 614598
rect 336960 614498 337060 614598
rect 337184 614498 337284 614598
rect 337408 614498 337508 614598
rect 337632 614498 337732 614598
rect 337856 614498 337956 614598
rect 338080 614498 338180 614598
rect 338304 614498 338404 614598
rect 338528 614498 338628 614598
rect 338752 614498 338852 614598
rect 338976 614498 339076 614598
rect 339200 614498 339300 614598
rect 339424 614498 339524 614598
rect 339648 614498 339748 614598
rect 339872 614498 339972 614598
rect 340096 614498 340196 614598
rect 340320 614498 340420 614598
rect 340544 614498 340644 614598
rect 340768 614498 340868 614598
rect 340992 614498 341092 614598
rect 341216 614498 341316 614598
rect 341440 614498 341540 614598
rect 341664 614498 341764 614598
rect 341888 614498 341988 614598
rect 342112 614498 342212 614598
<< metal2 >>
rect 298836 642694 305496 642724
rect 298836 642594 298876 642694
rect 298976 642594 299100 642694
rect 299200 642594 299324 642694
rect 299424 642594 299548 642694
rect 299648 642594 299772 642694
rect 299872 642594 299996 642694
rect 300096 642594 300220 642694
rect 300320 642594 300444 642694
rect 300544 642594 300668 642694
rect 300768 642594 300892 642694
rect 300992 642594 301116 642694
rect 301216 642594 301340 642694
rect 301440 642594 301564 642694
rect 301664 642594 301788 642694
rect 301888 642594 302012 642694
rect 302112 642594 302236 642694
rect 302336 642594 302460 642694
rect 302560 642594 302684 642694
rect 302784 642594 302908 642694
rect 303008 642594 303132 642694
rect 303232 642594 303356 642694
rect 303456 642594 303580 642694
rect 303680 642594 303804 642694
rect 303904 642594 304028 642694
rect 304128 642594 304252 642694
rect 304352 642594 304476 642694
rect 304576 642594 304700 642694
rect 304800 642594 304924 642694
rect 305024 642594 305148 642694
rect 305248 642594 305372 642694
rect 305472 642594 305496 642694
rect 298836 642470 305496 642594
rect 298836 642370 298876 642470
rect 298976 642370 299100 642470
rect 299200 642370 299324 642470
rect 299424 642370 299548 642470
rect 299648 642370 299772 642470
rect 299872 642370 299996 642470
rect 300096 642370 300220 642470
rect 300320 642370 300444 642470
rect 300544 642370 300668 642470
rect 300768 642370 300892 642470
rect 300992 642370 301116 642470
rect 301216 642370 301340 642470
rect 301440 642370 301564 642470
rect 301664 642370 301788 642470
rect 301888 642370 302012 642470
rect 302112 642370 302236 642470
rect 302336 642370 302460 642470
rect 302560 642370 302684 642470
rect 302784 642370 302908 642470
rect 303008 642370 303132 642470
rect 303232 642370 303356 642470
rect 303456 642370 303580 642470
rect 303680 642370 303804 642470
rect 303904 642370 304028 642470
rect 304128 642370 304252 642470
rect 304352 642370 304476 642470
rect 304576 642370 304700 642470
rect 304800 642370 304924 642470
rect 305024 642370 305148 642470
rect 305248 642370 305372 642470
rect 305472 642370 305496 642470
rect 298836 642246 305496 642370
rect 298836 642146 298876 642246
rect 298976 642146 299100 642246
rect 299200 642146 299324 642246
rect 299424 642146 299548 642246
rect 299648 642146 299772 642246
rect 299872 642146 299996 642246
rect 300096 642146 300220 642246
rect 300320 642146 300444 642246
rect 300544 642146 300668 642246
rect 300768 642146 300892 642246
rect 300992 642146 301116 642246
rect 301216 642146 301340 642246
rect 301440 642146 301564 642246
rect 301664 642146 301788 642246
rect 301888 642146 302012 642246
rect 302112 642146 302236 642246
rect 302336 642146 302460 642246
rect 302560 642146 302684 642246
rect 302784 642146 302908 642246
rect 303008 642146 303132 642246
rect 303232 642146 303356 642246
rect 303456 642146 303580 642246
rect 303680 642146 303804 642246
rect 303904 642146 304028 642246
rect 304128 642146 304252 642246
rect 304352 642146 304476 642246
rect 304576 642146 304700 642246
rect 304800 642146 304924 642246
rect 305024 642146 305148 642246
rect 305248 642146 305372 642246
rect 305472 642146 305496 642246
rect 298836 642022 305496 642146
rect 298836 641922 298876 642022
rect 298976 641922 299100 642022
rect 299200 641922 299324 642022
rect 299424 641922 299548 642022
rect 299648 641922 299772 642022
rect 299872 641922 299996 642022
rect 300096 641922 300220 642022
rect 300320 641922 300444 642022
rect 300544 641922 300668 642022
rect 300768 641922 300892 642022
rect 300992 641922 301116 642022
rect 301216 641922 301340 642022
rect 301440 641922 301564 642022
rect 301664 641922 301788 642022
rect 301888 641922 302012 642022
rect 302112 641922 302236 642022
rect 302336 641922 302460 642022
rect 302560 641922 302684 642022
rect 302784 641922 302908 642022
rect 303008 641922 303132 642022
rect 303232 641922 303356 642022
rect 303456 641922 303580 642022
rect 303680 641922 303804 642022
rect 303904 641922 304028 642022
rect 304128 641922 304252 642022
rect 304352 641922 304476 642022
rect 304576 641922 304700 642022
rect 304800 641922 304924 642022
rect 305024 641922 305148 642022
rect 305248 641922 305372 642022
rect 305472 641922 305496 642022
rect 298836 641798 305496 641922
rect 298836 641698 298876 641798
rect 298976 641698 299100 641798
rect 299200 641698 299324 641798
rect 299424 641698 299548 641798
rect 299648 641698 299772 641798
rect 299872 641698 299996 641798
rect 300096 641698 300220 641798
rect 300320 641698 300444 641798
rect 300544 641698 300668 641798
rect 300768 641698 300892 641798
rect 300992 641698 301116 641798
rect 301216 641698 301340 641798
rect 301440 641698 301564 641798
rect 301664 641698 301788 641798
rect 301888 641698 302012 641798
rect 302112 641698 302236 641798
rect 302336 641698 302460 641798
rect 302560 641698 302684 641798
rect 302784 641698 302908 641798
rect 303008 641698 303132 641798
rect 303232 641698 303356 641798
rect 303456 641698 303580 641798
rect 303680 641698 303804 641798
rect 303904 641698 304028 641798
rect 304128 641698 304252 641798
rect 304352 641698 304476 641798
rect 304576 641698 304700 641798
rect 304800 641698 304924 641798
rect 305024 641698 305148 641798
rect 305248 641698 305372 641798
rect 305472 641698 305496 641798
rect 298836 641664 305496 641698
rect 309306 642694 315966 642724
rect 309306 642594 309346 642694
rect 309446 642594 309570 642694
rect 309670 642594 309794 642694
rect 309894 642594 310018 642694
rect 310118 642594 310242 642694
rect 310342 642594 310466 642694
rect 310566 642594 310690 642694
rect 310790 642594 310914 642694
rect 311014 642594 311138 642694
rect 311238 642594 311362 642694
rect 311462 642594 311586 642694
rect 311686 642594 311810 642694
rect 311910 642594 312034 642694
rect 312134 642594 312258 642694
rect 312358 642594 312482 642694
rect 312582 642594 312706 642694
rect 312806 642594 312930 642694
rect 313030 642594 313154 642694
rect 313254 642594 313378 642694
rect 313478 642594 313602 642694
rect 313702 642594 313826 642694
rect 313926 642594 314050 642694
rect 314150 642594 314274 642694
rect 314374 642594 314498 642694
rect 314598 642594 314722 642694
rect 314822 642594 314946 642694
rect 315046 642594 315170 642694
rect 315270 642594 315394 642694
rect 315494 642594 315618 642694
rect 315718 642594 315842 642694
rect 315942 642594 315966 642694
rect 309306 642470 315966 642594
rect 309306 642370 309346 642470
rect 309446 642370 309570 642470
rect 309670 642370 309794 642470
rect 309894 642370 310018 642470
rect 310118 642370 310242 642470
rect 310342 642370 310466 642470
rect 310566 642370 310690 642470
rect 310790 642370 310914 642470
rect 311014 642370 311138 642470
rect 311238 642370 311362 642470
rect 311462 642370 311586 642470
rect 311686 642370 311810 642470
rect 311910 642370 312034 642470
rect 312134 642370 312258 642470
rect 312358 642370 312482 642470
rect 312582 642370 312706 642470
rect 312806 642370 312930 642470
rect 313030 642370 313154 642470
rect 313254 642370 313378 642470
rect 313478 642370 313602 642470
rect 313702 642370 313826 642470
rect 313926 642370 314050 642470
rect 314150 642370 314274 642470
rect 314374 642370 314498 642470
rect 314598 642370 314722 642470
rect 314822 642370 314946 642470
rect 315046 642370 315170 642470
rect 315270 642370 315394 642470
rect 315494 642370 315618 642470
rect 315718 642370 315842 642470
rect 315942 642370 315966 642470
rect 309306 642246 315966 642370
rect 309306 642146 309346 642246
rect 309446 642146 309570 642246
rect 309670 642146 309794 642246
rect 309894 642146 310018 642246
rect 310118 642146 310242 642246
rect 310342 642146 310466 642246
rect 310566 642146 310690 642246
rect 310790 642146 310914 642246
rect 311014 642146 311138 642246
rect 311238 642146 311362 642246
rect 311462 642146 311586 642246
rect 311686 642146 311810 642246
rect 311910 642146 312034 642246
rect 312134 642146 312258 642246
rect 312358 642146 312482 642246
rect 312582 642146 312706 642246
rect 312806 642146 312930 642246
rect 313030 642146 313154 642246
rect 313254 642146 313378 642246
rect 313478 642146 313602 642246
rect 313702 642146 313826 642246
rect 313926 642146 314050 642246
rect 314150 642146 314274 642246
rect 314374 642146 314498 642246
rect 314598 642146 314722 642246
rect 314822 642146 314946 642246
rect 315046 642146 315170 642246
rect 315270 642146 315394 642246
rect 315494 642146 315618 642246
rect 315718 642146 315842 642246
rect 315942 642146 315966 642246
rect 309306 642022 315966 642146
rect 309306 641922 309346 642022
rect 309446 641922 309570 642022
rect 309670 641922 309794 642022
rect 309894 641922 310018 642022
rect 310118 641922 310242 642022
rect 310342 641922 310466 642022
rect 310566 641922 310690 642022
rect 310790 641922 310914 642022
rect 311014 641922 311138 642022
rect 311238 641922 311362 642022
rect 311462 641922 311586 642022
rect 311686 641922 311810 642022
rect 311910 641922 312034 642022
rect 312134 641922 312258 642022
rect 312358 641922 312482 642022
rect 312582 641922 312706 642022
rect 312806 641922 312930 642022
rect 313030 641922 313154 642022
rect 313254 641922 313378 642022
rect 313478 641922 313602 642022
rect 313702 641922 313826 642022
rect 313926 641922 314050 642022
rect 314150 641922 314274 642022
rect 314374 641922 314498 642022
rect 314598 641922 314722 642022
rect 314822 641922 314946 642022
rect 315046 641922 315170 642022
rect 315270 641922 315394 642022
rect 315494 641922 315618 642022
rect 315718 641922 315842 642022
rect 315942 641922 315966 642022
rect 309306 641798 315966 641922
rect 309306 641698 309346 641798
rect 309446 641698 309570 641798
rect 309670 641698 309794 641798
rect 309894 641698 310018 641798
rect 310118 641698 310242 641798
rect 310342 641698 310466 641798
rect 310566 641698 310690 641798
rect 310790 641698 310914 641798
rect 311014 641698 311138 641798
rect 311238 641698 311362 641798
rect 311462 641698 311586 641798
rect 311686 641698 311810 641798
rect 311910 641698 312034 641798
rect 312134 641698 312258 641798
rect 312358 641698 312482 641798
rect 312582 641698 312706 641798
rect 312806 641698 312930 641798
rect 313030 641698 313154 641798
rect 313254 641698 313378 641798
rect 313478 641698 313602 641798
rect 313702 641698 313826 641798
rect 313926 641698 314050 641798
rect 314150 641698 314274 641798
rect 314374 641698 314498 641798
rect 314598 641698 314722 641798
rect 314822 641698 314946 641798
rect 315046 641698 315170 641798
rect 315270 641698 315394 641798
rect 315494 641698 315618 641798
rect 315718 641698 315842 641798
rect 315942 641698 315966 641798
rect 309306 641664 315966 641698
rect 335576 642714 342236 642744
rect 335576 642614 335616 642714
rect 335716 642614 335840 642714
rect 335940 642614 336064 642714
rect 336164 642614 336288 642714
rect 336388 642614 336512 642714
rect 336612 642614 336736 642714
rect 336836 642614 336960 642714
rect 337060 642614 337184 642714
rect 337284 642614 337408 642714
rect 337508 642614 337632 642714
rect 337732 642614 337856 642714
rect 337956 642614 338080 642714
rect 338180 642614 338304 642714
rect 338404 642614 338528 642714
rect 338628 642614 338752 642714
rect 338852 642614 338976 642714
rect 339076 642614 339200 642714
rect 339300 642614 339424 642714
rect 339524 642614 339648 642714
rect 339748 642614 339872 642714
rect 339972 642614 340096 642714
rect 340196 642614 340320 642714
rect 340420 642614 340544 642714
rect 340644 642614 340768 642714
rect 340868 642614 340992 642714
rect 341092 642614 341216 642714
rect 341316 642614 341440 642714
rect 341540 642614 341664 642714
rect 341764 642614 341888 642714
rect 341988 642614 342112 642714
rect 342212 642614 342236 642714
rect 335576 642490 342236 642614
rect 335576 642390 335616 642490
rect 335716 642390 335840 642490
rect 335940 642390 336064 642490
rect 336164 642390 336288 642490
rect 336388 642390 336512 642490
rect 336612 642390 336736 642490
rect 336836 642390 336960 642490
rect 337060 642390 337184 642490
rect 337284 642390 337408 642490
rect 337508 642390 337632 642490
rect 337732 642390 337856 642490
rect 337956 642390 338080 642490
rect 338180 642390 338304 642490
rect 338404 642390 338528 642490
rect 338628 642390 338752 642490
rect 338852 642390 338976 642490
rect 339076 642390 339200 642490
rect 339300 642390 339424 642490
rect 339524 642390 339648 642490
rect 339748 642390 339872 642490
rect 339972 642390 340096 642490
rect 340196 642390 340320 642490
rect 340420 642390 340544 642490
rect 340644 642390 340768 642490
rect 340868 642390 340992 642490
rect 341092 642390 341216 642490
rect 341316 642390 341440 642490
rect 341540 642390 341664 642490
rect 341764 642390 341888 642490
rect 341988 642390 342112 642490
rect 342212 642390 342236 642490
rect 335576 642266 342236 642390
rect 335576 642166 335616 642266
rect 335716 642166 335840 642266
rect 335940 642166 336064 642266
rect 336164 642166 336288 642266
rect 336388 642166 336512 642266
rect 336612 642166 336736 642266
rect 336836 642166 336960 642266
rect 337060 642166 337184 642266
rect 337284 642166 337408 642266
rect 337508 642166 337632 642266
rect 337732 642166 337856 642266
rect 337956 642166 338080 642266
rect 338180 642166 338304 642266
rect 338404 642166 338528 642266
rect 338628 642166 338752 642266
rect 338852 642166 338976 642266
rect 339076 642166 339200 642266
rect 339300 642166 339424 642266
rect 339524 642166 339648 642266
rect 339748 642166 339872 642266
rect 339972 642166 340096 642266
rect 340196 642166 340320 642266
rect 340420 642166 340544 642266
rect 340644 642166 340768 642266
rect 340868 642166 340992 642266
rect 341092 642166 341216 642266
rect 341316 642166 341440 642266
rect 341540 642166 341664 642266
rect 341764 642166 341888 642266
rect 341988 642166 342112 642266
rect 342212 642166 342236 642266
rect 335576 642042 342236 642166
rect 335576 641942 335616 642042
rect 335716 641942 335840 642042
rect 335940 641942 336064 642042
rect 336164 641942 336288 642042
rect 336388 641942 336512 642042
rect 336612 641942 336736 642042
rect 336836 641942 336960 642042
rect 337060 641942 337184 642042
rect 337284 641942 337408 642042
rect 337508 641942 337632 642042
rect 337732 641942 337856 642042
rect 337956 641942 338080 642042
rect 338180 641942 338304 642042
rect 338404 641942 338528 642042
rect 338628 641942 338752 642042
rect 338852 641942 338976 642042
rect 339076 641942 339200 642042
rect 339300 641942 339424 642042
rect 339524 641942 339648 642042
rect 339748 641942 339872 642042
rect 339972 641942 340096 642042
rect 340196 641942 340320 642042
rect 340420 641942 340544 642042
rect 340644 641942 340768 642042
rect 340868 641942 340992 642042
rect 341092 641942 341216 642042
rect 341316 641942 341440 642042
rect 341540 641942 341664 642042
rect 341764 641942 341888 642042
rect 341988 641942 342112 642042
rect 342212 641942 342236 642042
rect 335576 641818 342236 641942
rect 335576 641718 335616 641818
rect 335716 641718 335840 641818
rect 335940 641718 336064 641818
rect 336164 641718 336288 641818
rect 336388 641718 336512 641818
rect 336612 641718 336736 641818
rect 336836 641718 336960 641818
rect 337060 641718 337184 641818
rect 337284 641718 337408 641818
rect 337508 641718 337632 641818
rect 337732 641718 337856 641818
rect 337956 641718 338080 641818
rect 338180 641718 338304 641818
rect 338404 641718 338528 641818
rect 338628 641718 338752 641818
rect 338852 641718 338976 641818
rect 339076 641718 339200 641818
rect 339300 641718 339424 641818
rect 339524 641718 339648 641818
rect 339748 641718 339872 641818
rect 339972 641718 340096 641818
rect 340196 641718 340320 641818
rect 340420 641718 340544 641818
rect 340644 641718 340768 641818
rect 340868 641718 340992 641818
rect 341092 641718 341216 641818
rect 341316 641718 341440 641818
rect 341540 641718 341664 641818
rect 341764 641718 341888 641818
rect 341988 641718 342112 641818
rect 342212 641718 342236 641818
rect 335576 641684 342236 641718
rect 297820 637996 298880 638020
rect 297820 637896 297850 637996
rect 297950 637896 298074 637996
rect 298174 637896 298298 637996
rect 298398 637896 298522 637996
rect 298622 637896 298746 637996
rect 298846 637896 298880 637996
rect 297820 637772 298880 637896
rect 297820 637672 297850 637772
rect 297950 637672 298074 637772
rect 298174 637672 298298 637772
rect 298398 637672 298522 637772
rect 298622 637672 298746 637772
rect 298846 637672 298880 637772
rect 297820 637548 298880 637672
rect 297820 637448 297850 637548
rect 297950 637448 298074 637548
rect 298174 637448 298298 637548
rect 298398 637448 298522 637548
rect 298622 637448 298746 637548
rect 298846 637448 298880 637548
rect 297820 637324 298880 637448
rect 297820 637224 297850 637324
rect 297950 637224 298074 637324
rect 298174 637224 298298 637324
rect 298398 637224 298522 637324
rect 298622 637224 298746 637324
rect 298846 637224 298880 637324
rect 297820 637100 298880 637224
rect 297820 637000 297850 637100
rect 297950 637000 298074 637100
rect 298174 637000 298298 637100
rect 298398 637000 298522 637100
rect 298622 637000 298746 637100
rect 298846 637000 298880 637100
rect 297820 636876 298880 637000
rect 297820 636776 297850 636876
rect 297950 636776 298074 636876
rect 298174 636776 298298 636876
rect 298398 636776 298522 636876
rect 298622 636776 298746 636876
rect 298846 636776 298880 636876
rect 297820 636652 298880 636776
rect 297820 636552 297850 636652
rect 297950 636552 298074 636652
rect 298174 636552 298298 636652
rect 298398 636552 298522 636652
rect 298622 636552 298746 636652
rect 298846 636552 298880 636652
rect 297820 636428 298880 636552
rect 297820 636328 297850 636428
rect 297950 636328 298074 636428
rect 298174 636328 298298 636428
rect 298398 636328 298522 636428
rect 298622 636328 298746 636428
rect 298846 636328 298880 636428
rect 297820 636204 298880 636328
rect 297820 636104 297850 636204
rect 297950 636104 298074 636204
rect 298174 636104 298298 636204
rect 298398 636104 298522 636204
rect 298622 636104 298746 636204
rect 298846 636104 298880 636204
rect 297820 635980 298880 636104
rect 297820 635880 297850 635980
rect 297950 635880 298074 635980
rect 298174 635880 298298 635980
rect 298398 635880 298522 635980
rect 298622 635880 298746 635980
rect 298846 635880 298880 635980
rect 297820 635756 298880 635880
rect 297820 635656 297850 635756
rect 297950 635656 298074 635756
rect 298174 635656 298298 635756
rect 298398 635656 298522 635756
rect 298622 635656 298746 635756
rect 298846 635656 298880 635756
rect 297820 635532 298880 635656
rect 297820 635432 297850 635532
rect 297950 635432 298074 635532
rect 298174 635432 298298 635532
rect 298398 635432 298522 635532
rect 298622 635432 298746 635532
rect 298846 635432 298880 635532
rect 297820 635308 298880 635432
rect 297820 635208 297850 635308
rect 297950 635208 298074 635308
rect 298174 635208 298298 635308
rect 298398 635208 298522 635308
rect 298622 635208 298746 635308
rect 298846 635208 298880 635308
rect 297820 635084 298880 635208
rect 297820 634984 297850 635084
rect 297950 634984 298074 635084
rect 298174 634984 298298 635084
rect 298398 634984 298522 635084
rect 298622 634984 298746 635084
rect 298846 634984 298880 635084
rect 297820 634860 298880 634984
rect 297820 634760 297850 634860
rect 297950 634760 298074 634860
rect 298174 634760 298298 634860
rect 298398 634760 298522 634860
rect 298622 634760 298746 634860
rect 298846 634760 298880 634860
rect 297820 634636 298880 634760
rect 297820 634536 297850 634636
rect 297950 634536 298074 634636
rect 298174 634536 298298 634636
rect 298398 634536 298522 634636
rect 298622 634536 298746 634636
rect 298846 634536 298880 634636
rect 297820 634412 298880 634536
rect 297820 634312 297850 634412
rect 297950 634312 298074 634412
rect 298174 634312 298298 634412
rect 298398 634312 298522 634412
rect 298622 634312 298746 634412
rect 298846 634312 298880 634412
rect 297820 634188 298880 634312
rect 297820 634088 297850 634188
rect 297950 634088 298074 634188
rect 298174 634088 298298 634188
rect 298398 634088 298522 634188
rect 298622 634088 298746 634188
rect 298846 634088 298880 634188
rect 297820 633964 298880 634088
rect 297820 633864 297850 633964
rect 297950 633864 298074 633964
rect 298174 633864 298298 633964
rect 298398 633864 298522 633964
rect 298622 633864 298746 633964
rect 298846 633864 298880 633964
rect 297820 633740 298880 633864
rect 297820 633640 297850 633740
rect 297950 633640 298074 633740
rect 298174 633640 298298 633740
rect 298398 633640 298522 633740
rect 298622 633640 298746 633740
rect 298846 633640 298880 633740
rect 297820 633516 298880 633640
rect 297820 633416 297850 633516
rect 297950 633416 298074 633516
rect 298174 633416 298298 633516
rect 298398 633416 298522 633516
rect 298622 633416 298746 633516
rect 298846 633416 298880 633516
rect 297820 633292 298880 633416
rect 297820 633192 297850 633292
rect 297950 633192 298074 633292
rect 298174 633192 298298 633292
rect 298398 633192 298522 633292
rect 298622 633192 298746 633292
rect 298846 633192 298880 633292
rect 297820 633068 298880 633192
rect 297820 632968 297850 633068
rect 297950 632968 298074 633068
rect 298174 632968 298298 633068
rect 298398 632968 298522 633068
rect 298622 632968 298746 633068
rect 298846 632968 298880 633068
rect 297820 632844 298880 632968
rect 297820 632744 297850 632844
rect 297950 632744 298074 632844
rect 298174 632744 298298 632844
rect 298398 632744 298522 632844
rect 298622 632744 298746 632844
rect 298846 632744 298880 632844
rect 297820 632620 298880 632744
rect 297820 632520 297850 632620
rect 297950 632520 298074 632620
rect 298174 632520 298298 632620
rect 298398 632520 298522 632620
rect 298622 632520 298746 632620
rect 298846 632520 298880 632620
rect 297820 632396 298880 632520
rect 297820 632296 297850 632396
rect 297950 632296 298074 632396
rect 298174 632296 298298 632396
rect 298398 632296 298522 632396
rect 298622 632296 298746 632396
rect 298846 632296 298880 632396
rect 297820 632172 298880 632296
rect 297820 632072 297850 632172
rect 297950 632072 298074 632172
rect 298174 632072 298298 632172
rect 298398 632072 298522 632172
rect 298622 632072 298746 632172
rect 298846 632072 298880 632172
rect 297820 631948 298880 632072
rect 297820 631848 297850 631948
rect 297950 631848 298074 631948
rect 298174 631848 298298 631948
rect 298398 631848 298522 631948
rect 298622 631848 298746 631948
rect 298846 631848 298880 631948
rect 297820 631724 298880 631848
rect 297820 631624 297850 631724
rect 297950 631624 298074 631724
rect 298174 631624 298298 631724
rect 298398 631624 298522 631724
rect 298622 631624 298746 631724
rect 298846 631624 298880 631724
rect 297820 631500 298880 631624
rect 297820 631400 297850 631500
rect 297950 631400 298074 631500
rect 298174 631400 298298 631500
rect 298398 631400 298522 631500
rect 298622 631400 298746 631500
rect 298846 631400 298880 631500
rect 297820 631360 298880 631400
rect 342100 637996 343160 638020
rect 342100 637896 342130 637996
rect 342230 637896 342354 637996
rect 342454 637896 342578 637996
rect 342678 637896 342802 637996
rect 342902 637896 343026 637996
rect 343126 637896 343160 637996
rect 342100 637772 343160 637896
rect 342100 637672 342130 637772
rect 342230 637672 342354 637772
rect 342454 637672 342578 637772
rect 342678 637672 342802 637772
rect 342902 637672 343026 637772
rect 343126 637672 343160 637772
rect 342100 637548 343160 637672
rect 342100 637448 342130 637548
rect 342230 637448 342354 637548
rect 342454 637448 342578 637548
rect 342678 637448 342802 637548
rect 342902 637448 343026 637548
rect 343126 637448 343160 637548
rect 342100 637324 343160 637448
rect 342100 637224 342130 637324
rect 342230 637224 342354 637324
rect 342454 637224 342578 637324
rect 342678 637224 342802 637324
rect 342902 637224 343026 637324
rect 343126 637224 343160 637324
rect 342100 637100 343160 637224
rect 342100 637000 342130 637100
rect 342230 637000 342354 637100
rect 342454 637000 342578 637100
rect 342678 637000 342802 637100
rect 342902 637000 343026 637100
rect 343126 637000 343160 637100
rect 342100 636876 343160 637000
rect 342100 636776 342130 636876
rect 342230 636776 342354 636876
rect 342454 636776 342578 636876
rect 342678 636776 342802 636876
rect 342902 636776 343026 636876
rect 343126 636776 343160 636876
rect 342100 636652 343160 636776
rect 342100 636552 342130 636652
rect 342230 636552 342354 636652
rect 342454 636552 342578 636652
rect 342678 636552 342802 636652
rect 342902 636552 343026 636652
rect 343126 636552 343160 636652
rect 342100 636428 343160 636552
rect 342100 636328 342130 636428
rect 342230 636328 342354 636428
rect 342454 636328 342578 636428
rect 342678 636328 342802 636428
rect 342902 636328 343026 636428
rect 343126 636328 343160 636428
rect 342100 636204 343160 636328
rect 342100 636104 342130 636204
rect 342230 636104 342354 636204
rect 342454 636104 342578 636204
rect 342678 636104 342802 636204
rect 342902 636104 343026 636204
rect 343126 636104 343160 636204
rect 342100 635980 343160 636104
rect 342100 635880 342130 635980
rect 342230 635880 342354 635980
rect 342454 635880 342578 635980
rect 342678 635880 342802 635980
rect 342902 635880 343026 635980
rect 343126 635880 343160 635980
rect 342100 635756 343160 635880
rect 342100 635656 342130 635756
rect 342230 635656 342354 635756
rect 342454 635656 342578 635756
rect 342678 635656 342802 635756
rect 342902 635656 343026 635756
rect 343126 635656 343160 635756
rect 342100 635532 343160 635656
rect 342100 635432 342130 635532
rect 342230 635432 342354 635532
rect 342454 635432 342578 635532
rect 342678 635432 342802 635532
rect 342902 635432 343026 635532
rect 343126 635432 343160 635532
rect 342100 635308 343160 635432
rect 342100 635208 342130 635308
rect 342230 635208 342354 635308
rect 342454 635208 342578 635308
rect 342678 635208 342802 635308
rect 342902 635208 343026 635308
rect 343126 635208 343160 635308
rect 342100 635084 343160 635208
rect 342100 634984 342130 635084
rect 342230 634984 342354 635084
rect 342454 634984 342578 635084
rect 342678 634984 342802 635084
rect 342902 634984 343026 635084
rect 343126 634984 343160 635084
rect 342100 634860 343160 634984
rect 342100 634760 342130 634860
rect 342230 634760 342354 634860
rect 342454 634760 342578 634860
rect 342678 634760 342802 634860
rect 342902 634760 343026 634860
rect 343126 634760 343160 634860
rect 342100 634636 343160 634760
rect 342100 634536 342130 634636
rect 342230 634536 342354 634636
rect 342454 634536 342578 634636
rect 342678 634536 342802 634636
rect 342902 634536 343026 634636
rect 343126 634536 343160 634636
rect 342100 634412 343160 634536
rect 342100 634312 342130 634412
rect 342230 634312 342354 634412
rect 342454 634312 342578 634412
rect 342678 634312 342802 634412
rect 342902 634312 343026 634412
rect 343126 634312 343160 634412
rect 342100 634188 343160 634312
rect 342100 634088 342130 634188
rect 342230 634088 342354 634188
rect 342454 634088 342578 634188
rect 342678 634088 342802 634188
rect 342902 634088 343026 634188
rect 343126 634088 343160 634188
rect 342100 633964 343160 634088
rect 342100 633864 342130 633964
rect 342230 633864 342354 633964
rect 342454 633864 342578 633964
rect 342678 633864 342802 633964
rect 342902 633864 343026 633964
rect 343126 633864 343160 633964
rect 342100 633740 343160 633864
rect 342100 633640 342130 633740
rect 342230 633640 342354 633740
rect 342454 633640 342578 633740
rect 342678 633640 342802 633740
rect 342902 633640 343026 633740
rect 343126 633640 343160 633740
rect 342100 633516 343160 633640
rect 342100 633416 342130 633516
rect 342230 633416 342354 633516
rect 342454 633416 342578 633516
rect 342678 633416 342802 633516
rect 342902 633416 343026 633516
rect 343126 633416 343160 633516
rect 342100 633292 343160 633416
rect 342100 633192 342130 633292
rect 342230 633192 342354 633292
rect 342454 633192 342578 633292
rect 342678 633192 342802 633292
rect 342902 633192 343026 633292
rect 343126 633192 343160 633292
rect 342100 633068 343160 633192
rect 342100 632968 342130 633068
rect 342230 632968 342354 633068
rect 342454 632968 342578 633068
rect 342678 632968 342802 633068
rect 342902 632968 343026 633068
rect 343126 632968 343160 633068
rect 342100 632844 343160 632968
rect 342100 632744 342130 632844
rect 342230 632744 342354 632844
rect 342454 632744 342578 632844
rect 342678 632744 342802 632844
rect 342902 632744 343026 632844
rect 343126 632744 343160 632844
rect 342100 632620 343160 632744
rect 342100 632520 342130 632620
rect 342230 632520 342354 632620
rect 342454 632520 342578 632620
rect 342678 632520 342802 632620
rect 342902 632520 343026 632620
rect 343126 632520 343160 632620
rect 342100 632396 343160 632520
rect 342100 632296 342130 632396
rect 342230 632296 342354 632396
rect 342454 632296 342578 632396
rect 342678 632296 342802 632396
rect 342902 632296 343026 632396
rect 343126 632296 343160 632396
rect 342100 632172 343160 632296
rect 342100 632072 342130 632172
rect 342230 632072 342354 632172
rect 342454 632072 342578 632172
rect 342678 632072 342802 632172
rect 342902 632072 343026 632172
rect 343126 632072 343160 632172
rect 342100 631948 343160 632072
rect 342100 631848 342130 631948
rect 342230 631848 342354 631948
rect 342454 631848 342578 631948
rect 342678 631848 342802 631948
rect 342902 631848 343026 631948
rect 343126 631848 343160 631948
rect 342100 631724 343160 631848
rect 342100 631624 342130 631724
rect 342230 631624 342354 631724
rect 342454 631624 342578 631724
rect 342678 631624 342802 631724
rect 342902 631624 343026 631724
rect 343126 631624 343160 631724
rect 342100 631500 343160 631624
rect 342100 631400 342130 631500
rect 342230 631400 342354 631500
rect 342454 631400 342578 631500
rect 342678 631400 342802 631500
rect 342902 631400 343026 631500
rect 343126 631400 343160 631500
rect 342100 631360 343160 631400
rect 319383 628868 319617 628885
rect 319383 628668 319400 628868
rect 319600 628668 319617 628868
rect 319383 628651 319617 628668
rect 319817 628868 320051 628885
rect 319817 628668 319834 628868
rect 320034 628668 320051 628868
rect 319817 628651 320051 628668
rect 320251 628868 320485 628885
rect 320251 628668 320268 628868
rect 320468 628668 320485 628868
rect 320251 628651 320485 628668
rect 320685 628868 320919 628885
rect 320685 628668 320702 628868
rect 320902 628668 320919 628868
rect 320685 628651 320919 628668
rect 321119 628868 321353 628885
rect 321119 628668 321136 628868
rect 321336 628668 321353 628868
rect 321119 628651 321353 628668
rect 321553 628868 321787 628885
rect 321553 628668 321570 628868
rect 321770 628668 321787 628868
rect 321553 628651 321787 628668
rect 321987 628868 322221 628885
rect 321987 628668 322004 628868
rect 322204 628668 322221 628868
rect 321987 628651 322221 628668
rect 322421 628868 322655 628885
rect 322421 628668 322438 628868
rect 322638 628668 322655 628868
rect 322421 628651 322655 628668
rect 322855 628868 323089 628885
rect 322855 628668 322872 628868
rect 323072 628668 323089 628868
rect 322855 628651 323089 628668
rect 323289 628868 323523 628885
rect 323289 628668 323306 628868
rect 323506 628668 323523 628868
rect 323289 628651 323523 628668
rect 323723 628868 323957 628885
rect 323723 628668 323740 628868
rect 323940 628668 323957 628868
rect 323723 628651 323957 628668
rect 324123 628868 324357 628885
rect 324123 628668 324140 628868
rect 324340 628668 324357 628868
rect 324123 628651 324357 628668
rect 324523 628868 324757 628885
rect 324523 628668 324540 628868
rect 324740 628668 324757 628868
rect 324523 628651 324757 628668
rect 324923 628868 325157 628885
rect 324923 628668 324940 628868
rect 325140 628668 325157 628868
rect 324923 628651 325157 628668
rect 325323 628868 325557 628885
rect 325323 628668 325340 628868
rect 325540 628668 325557 628868
rect 325323 628651 325557 628668
rect 325723 628868 325957 628885
rect 325723 628668 325740 628868
rect 325940 628668 325957 628868
rect 325723 628651 325957 628668
rect 326123 628868 326357 628885
rect 326123 628668 326140 628868
rect 326340 628668 326357 628868
rect 326123 628651 326357 628668
rect 326523 628868 326757 628885
rect 326523 628668 326540 628868
rect 326740 628668 326757 628868
rect 326523 628651 326757 628668
rect 326923 628868 327157 628885
rect 326923 628668 326940 628868
rect 327140 628668 327157 628868
rect 326923 628651 327157 628668
rect 327323 628868 327557 628885
rect 327323 628668 327340 628868
rect 327540 628668 327557 628868
rect 327323 628651 327557 628668
rect 328923 628868 329157 628885
rect 328923 628668 328940 628868
rect 329140 628668 329157 628868
rect 328923 628651 329157 628668
rect 329323 628868 329557 628885
rect 329323 628668 329340 628868
rect 329540 628668 329557 628868
rect 329323 628651 329557 628668
rect 329723 628868 329957 628885
rect 329723 628668 329740 628868
rect 329940 628668 329957 628868
rect 329723 628651 329957 628668
rect 330123 628868 330357 628885
rect 330123 628668 330140 628868
rect 330340 628668 330357 628868
rect 330123 628651 330357 628668
rect 330523 628868 330757 628885
rect 330523 628668 330540 628868
rect 330740 628668 330757 628868
rect 330523 628651 330757 628668
rect 330923 628868 331157 628885
rect 330923 628668 330940 628868
rect 331140 628668 331157 628868
rect 330923 628651 331157 628668
rect 331323 628868 331557 628885
rect 331323 628668 331340 628868
rect 331540 628668 331557 628868
rect 331323 628651 331557 628668
rect 331723 628868 331957 628885
rect 331723 628668 331740 628868
rect 331940 628668 331957 628868
rect 331723 628651 331957 628668
rect 332123 628868 332357 628885
rect 332123 628668 332140 628868
rect 332340 628668 332357 628868
rect 332123 628651 332357 628668
rect 319383 628434 319617 628451
rect 319383 628234 319400 628434
rect 319600 628234 319617 628434
rect 319383 628217 319617 628234
rect 319817 628434 320051 628451
rect 319817 628234 319834 628434
rect 320034 628234 320051 628434
rect 319817 628217 320051 628234
rect 320251 628434 320485 628451
rect 320251 628234 320268 628434
rect 320468 628234 320485 628434
rect 320251 628217 320485 628234
rect 320685 628434 320919 628451
rect 320685 628234 320702 628434
rect 320902 628234 320919 628434
rect 320685 628217 320919 628234
rect 321119 628434 321353 628451
rect 321119 628234 321136 628434
rect 321336 628234 321353 628434
rect 321119 628217 321353 628234
rect 321553 628434 321787 628451
rect 321553 628234 321570 628434
rect 321770 628234 321787 628434
rect 321553 628217 321787 628234
rect 321987 628434 322221 628451
rect 321987 628234 322004 628434
rect 322204 628234 322221 628434
rect 321987 628217 322221 628234
rect 322421 628434 322655 628451
rect 322421 628234 322438 628434
rect 322638 628234 322655 628434
rect 322421 628217 322655 628234
rect 322855 628434 323089 628451
rect 322855 628234 322872 628434
rect 323072 628234 323089 628434
rect 322855 628217 323089 628234
rect 323289 628434 323523 628451
rect 323289 628234 323306 628434
rect 323506 628234 323523 628434
rect 323289 628217 323523 628234
rect 323723 628434 323957 628451
rect 323723 628234 323740 628434
rect 323940 628234 323957 628434
rect 323723 628217 323957 628234
rect 319383 628000 319617 628017
rect 319383 627800 319400 628000
rect 319600 627800 319617 628000
rect 319383 627783 319617 627800
rect 319817 628000 320051 628017
rect 319817 627800 319834 628000
rect 320034 627800 320051 628000
rect 319817 627783 320051 627800
rect 320251 628000 320485 628017
rect 320251 627800 320268 628000
rect 320468 627800 320485 628000
rect 320251 627783 320485 627800
rect 320685 628000 320919 628017
rect 320685 627800 320702 628000
rect 320902 627800 320919 628000
rect 320685 627783 320919 627800
rect 321119 628000 321353 628017
rect 321119 627800 321136 628000
rect 321336 627800 321353 628000
rect 321119 627783 321353 627800
rect 321553 628000 321787 628017
rect 321553 627800 321570 628000
rect 321770 627800 321787 628000
rect 321553 627783 321787 627800
rect 321987 628000 322221 628017
rect 321987 627800 322004 628000
rect 322204 627800 322221 628000
rect 321987 627783 322221 627800
rect 322421 628000 322655 628017
rect 322421 627800 322438 628000
rect 322638 627800 322655 628000
rect 322421 627783 322655 627800
rect 322855 628000 323089 628017
rect 322855 627800 322872 628000
rect 323072 627800 323089 628000
rect 322855 627783 323089 627800
rect 323289 628000 323523 628017
rect 323289 627800 323306 628000
rect 323506 627800 323523 628000
rect 323289 627783 323523 627800
rect 323723 628000 323957 628017
rect 323723 627800 323740 628000
rect 323940 627800 323957 628000
rect 323723 627783 323957 627800
rect 302960 626030 303550 626090
rect 302960 625970 302980 626030
rect 303040 625970 303100 626030
rect 303160 625970 303220 626030
rect 303280 625970 303340 626030
rect 303400 625970 303460 626030
rect 303520 625970 303550 626030
rect 302960 625910 303550 625970
rect 302960 625850 302980 625910
rect 303040 625850 303100 625910
rect 303160 625850 303220 625910
rect 303280 625850 303340 625910
rect 303400 625850 303460 625910
rect 303520 625850 303550 625910
rect 297820 624596 298878 624606
rect 297820 624496 297850 624596
rect 297950 624496 298074 624596
rect 298174 624496 298298 624596
rect 298398 624496 298522 624596
rect 298622 624496 298746 624596
rect 298846 624496 298878 624596
rect 297820 624372 298878 624496
rect 297820 624272 297850 624372
rect 297950 624272 298074 624372
rect 298174 624272 298298 624372
rect 298398 624272 298522 624372
rect 298622 624272 298746 624372
rect 298846 624272 298878 624372
rect 297820 624148 298878 624272
rect 297820 624048 297850 624148
rect 297950 624048 298074 624148
rect 298174 624048 298298 624148
rect 298398 624048 298522 624148
rect 298622 624048 298746 624148
rect 298846 624048 298878 624148
rect 297820 623924 298878 624048
rect 302960 624184 303550 625850
rect 302960 624114 302972 624184
rect 303032 624114 303044 624184
rect 303104 624114 303116 624184
rect 303176 624114 303188 624184
rect 303248 624114 303260 624184
rect 303320 624114 303332 624184
rect 303392 624114 303404 624184
rect 303464 624114 303476 624184
rect 303536 624114 303550 624184
rect 302960 624090 303550 624114
rect 302960 624020 302972 624090
rect 303032 624020 303044 624090
rect 303104 624020 303116 624090
rect 303176 624020 303188 624090
rect 303248 624020 303260 624090
rect 303320 624020 303332 624090
rect 303392 624020 303404 624090
rect 303464 624020 303476 624090
rect 303536 624020 303550 624090
rect 302960 624010 303550 624020
rect 342100 624596 343158 624606
rect 342100 624496 342130 624596
rect 342230 624496 342354 624596
rect 342454 624496 342578 624596
rect 342678 624496 342802 624596
rect 342902 624496 343026 624596
rect 343126 624496 343158 624596
rect 342100 624372 343158 624496
rect 342100 624272 342130 624372
rect 342230 624272 342354 624372
rect 342454 624272 342578 624372
rect 342678 624272 342802 624372
rect 342902 624272 343026 624372
rect 343126 624272 343158 624372
rect 342100 624148 343158 624272
rect 342100 624048 342130 624148
rect 342230 624048 342354 624148
rect 342454 624048 342578 624148
rect 342678 624048 342802 624148
rect 342902 624048 343026 624148
rect 343126 624048 343158 624148
rect 297820 623824 297850 623924
rect 297950 623824 298074 623924
rect 298174 623824 298298 623924
rect 298398 623824 298522 623924
rect 298622 623824 298746 623924
rect 298846 623824 298878 623924
rect 297820 623700 298878 623824
rect 297820 623600 297850 623700
rect 297950 623600 298074 623700
rect 298174 623600 298298 623700
rect 298398 623600 298522 623700
rect 298622 623600 298746 623700
rect 298846 623600 298878 623700
rect 297820 623476 298878 623600
rect 297820 623376 297850 623476
rect 297950 623376 298074 623476
rect 298174 623376 298298 623476
rect 298398 623376 298522 623476
rect 298622 623376 298746 623476
rect 298846 623376 298878 623476
rect 297820 623252 298878 623376
rect 297820 623152 297850 623252
rect 297950 623152 298074 623252
rect 298174 623152 298298 623252
rect 298398 623152 298522 623252
rect 298622 623152 298746 623252
rect 298846 623152 298878 623252
rect 297820 623028 298878 623152
rect 297820 622928 297850 623028
rect 297950 622928 298074 623028
rect 298174 622928 298298 623028
rect 298398 622928 298522 623028
rect 298622 622928 298746 623028
rect 298846 622928 298878 623028
rect 297820 622804 298878 622928
rect 297820 622704 297850 622804
rect 297950 622704 298074 622804
rect 298174 622704 298298 622804
rect 298398 622704 298522 622804
rect 298622 622704 298746 622804
rect 298846 622704 298878 622804
rect 297820 622580 298878 622704
rect 297820 622480 297850 622580
rect 297950 622480 298074 622580
rect 298174 622480 298298 622580
rect 298398 622480 298522 622580
rect 298622 622480 298746 622580
rect 298846 622480 298878 622580
rect 297820 622356 298878 622480
rect 297820 622256 297850 622356
rect 297950 622256 298074 622356
rect 298174 622256 298298 622356
rect 298398 622256 298522 622356
rect 298622 622256 298746 622356
rect 298846 622256 298878 622356
rect 297820 622132 298878 622256
rect 297820 622032 297850 622132
rect 297950 622032 298074 622132
rect 298174 622032 298298 622132
rect 298398 622032 298522 622132
rect 298622 622032 298746 622132
rect 298846 622032 298878 622132
rect 297820 621908 298878 622032
rect 297820 621808 297850 621908
rect 297950 621808 298074 621908
rect 298174 621808 298298 621908
rect 298398 621808 298522 621908
rect 298622 621808 298746 621908
rect 298846 621808 298878 621908
rect 297820 621684 298878 621808
rect 297820 621584 297850 621684
rect 297950 621584 298074 621684
rect 298174 621584 298298 621684
rect 298398 621584 298522 621684
rect 298622 621584 298746 621684
rect 298846 621584 298878 621684
rect 297820 621460 298878 621584
rect 297820 621360 297850 621460
rect 297950 621360 298074 621460
rect 298174 621360 298298 621460
rect 298398 621360 298522 621460
rect 298622 621360 298746 621460
rect 298846 621360 298878 621460
rect 297820 621236 298878 621360
rect 297820 621136 297850 621236
rect 297950 621136 298074 621236
rect 298174 621136 298298 621236
rect 298398 621136 298522 621236
rect 298622 621136 298746 621236
rect 298846 621136 298878 621236
rect 297820 621012 298878 621136
rect 297820 620912 297850 621012
rect 297950 620912 298074 621012
rect 298174 620912 298298 621012
rect 298398 620912 298522 621012
rect 298622 620912 298746 621012
rect 298846 620912 298878 621012
rect 297820 620788 298878 620912
rect 297820 620688 297850 620788
rect 297950 620688 298074 620788
rect 298174 620688 298298 620788
rect 298398 620688 298522 620788
rect 298622 620688 298746 620788
rect 298846 620688 298878 620788
rect 297820 620564 298878 620688
rect 297820 620464 297850 620564
rect 297950 620464 298074 620564
rect 298174 620464 298298 620564
rect 298398 620464 298522 620564
rect 298622 620464 298746 620564
rect 298846 620464 298878 620564
rect 297820 620340 298878 620464
rect 297820 620240 297850 620340
rect 297950 620240 298074 620340
rect 298174 620240 298298 620340
rect 298398 620240 298522 620340
rect 298622 620240 298746 620340
rect 298846 620240 298878 620340
rect 297820 620116 298878 620240
rect 297820 620016 297850 620116
rect 297950 620016 298074 620116
rect 298174 620016 298298 620116
rect 298398 620016 298522 620116
rect 298622 620016 298746 620116
rect 298846 620016 298878 620116
rect 297820 619892 298878 620016
rect 297820 619792 297850 619892
rect 297950 619792 298074 619892
rect 298174 619792 298298 619892
rect 298398 619792 298522 619892
rect 298622 619792 298746 619892
rect 298846 619792 298878 619892
rect 297820 619668 298878 619792
rect 297820 619568 297850 619668
rect 297950 619568 298074 619668
rect 298174 619568 298298 619668
rect 298398 619568 298522 619668
rect 298622 619568 298746 619668
rect 298846 619568 298878 619668
rect 297820 619444 298878 619568
rect 297820 619344 297850 619444
rect 297950 619344 298074 619444
rect 298174 619344 298298 619444
rect 298398 619344 298522 619444
rect 298622 619344 298746 619444
rect 298846 619344 298878 619444
rect 297820 619220 298878 619344
rect 297820 619120 297850 619220
rect 297950 619120 298074 619220
rect 298174 619120 298298 619220
rect 298398 619120 298522 619220
rect 298622 619120 298746 619220
rect 298846 619120 298878 619220
rect 297820 618996 298878 619120
rect 297820 618896 297850 618996
rect 297950 618896 298074 618996
rect 298174 618896 298298 618996
rect 298398 618896 298522 618996
rect 298622 618896 298746 618996
rect 298846 618896 298878 618996
rect 297820 618772 298878 618896
rect 297820 618672 297850 618772
rect 297950 618672 298074 618772
rect 298174 618672 298298 618772
rect 298398 618672 298522 618772
rect 298622 618672 298746 618772
rect 298846 618672 298878 618772
rect 297820 618548 298878 618672
rect 297820 618448 297850 618548
rect 297950 618448 298074 618548
rect 298174 618448 298298 618548
rect 298398 618448 298522 618548
rect 298622 618448 298746 618548
rect 298846 618448 298878 618548
rect 297820 618324 298878 618448
rect 297820 618224 297850 618324
rect 297950 618224 298074 618324
rect 298174 618224 298298 618324
rect 298398 618224 298522 618324
rect 298622 618224 298746 618324
rect 298846 618224 298878 618324
rect 297820 618100 298878 618224
rect 297820 618000 297850 618100
rect 297950 618000 298074 618100
rect 298174 618000 298298 618100
rect 298398 618000 298522 618100
rect 298622 618000 298746 618100
rect 298846 618000 298878 618100
rect 297820 617980 298878 618000
rect 342100 623924 343158 624048
rect 342100 623824 342130 623924
rect 342230 623824 342354 623924
rect 342454 623824 342578 623924
rect 342678 623824 342802 623924
rect 342902 623824 343026 623924
rect 343126 623824 343158 623924
rect 342100 623700 343158 623824
rect 342100 623600 342130 623700
rect 342230 623600 342354 623700
rect 342454 623600 342578 623700
rect 342678 623600 342802 623700
rect 342902 623600 343026 623700
rect 343126 623600 343158 623700
rect 342100 623476 343158 623600
rect 342100 623376 342130 623476
rect 342230 623376 342354 623476
rect 342454 623376 342578 623476
rect 342678 623376 342802 623476
rect 342902 623376 343026 623476
rect 343126 623376 343158 623476
rect 342100 623252 343158 623376
rect 342100 623152 342130 623252
rect 342230 623152 342354 623252
rect 342454 623152 342578 623252
rect 342678 623152 342802 623252
rect 342902 623152 343026 623252
rect 343126 623152 343158 623252
rect 342100 623028 343158 623152
rect 342100 622928 342130 623028
rect 342230 622928 342354 623028
rect 342454 622928 342578 623028
rect 342678 622928 342802 623028
rect 342902 622928 343026 623028
rect 343126 622928 343158 623028
rect 342100 622804 343158 622928
rect 342100 622704 342130 622804
rect 342230 622704 342354 622804
rect 342454 622704 342578 622804
rect 342678 622704 342802 622804
rect 342902 622704 343026 622804
rect 343126 622704 343158 622804
rect 342100 622580 343158 622704
rect 342100 622480 342130 622580
rect 342230 622480 342354 622580
rect 342454 622480 342578 622580
rect 342678 622480 342802 622580
rect 342902 622480 343026 622580
rect 343126 622480 343158 622580
rect 342100 622356 343158 622480
rect 342100 622256 342130 622356
rect 342230 622256 342354 622356
rect 342454 622256 342578 622356
rect 342678 622256 342802 622356
rect 342902 622256 343026 622356
rect 343126 622256 343158 622356
rect 342100 622132 343158 622256
rect 342100 622032 342130 622132
rect 342230 622032 342354 622132
rect 342454 622032 342578 622132
rect 342678 622032 342802 622132
rect 342902 622032 343026 622132
rect 343126 622032 343158 622132
rect 342100 621908 343158 622032
rect 342100 621808 342130 621908
rect 342230 621808 342354 621908
rect 342454 621808 342578 621908
rect 342678 621808 342802 621908
rect 342902 621808 343026 621908
rect 343126 621808 343158 621908
rect 342100 621684 343158 621808
rect 342100 621584 342130 621684
rect 342230 621584 342354 621684
rect 342454 621584 342578 621684
rect 342678 621584 342802 621684
rect 342902 621584 343026 621684
rect 343126 621584 343158 621684
rect 342100 621460 343158 621584
rect 342100 621360 342130 621460
rect 342230 621360 342354 621460
rect 342454 621360 342578 621460
rect 342678 621360 342802 621460
rect 342902 621360 343026 621460
rect 343126 621360 343158 621460
rect 342100 621236 343158 621360
rect 342100 621136 342130 621236
rect 342230 621136 342354 621236
rect 342454 621136 342578 621236
rect 342678 621136 342802 621236
rect 342902 621136 343026 621236
rect 343126 621136 343158 621236
rect 342100 621012 343158 621136
rect 342100 620912 342130 621012
rect 342230 620912 342354 621012
rect 342454 620912 342578 621012
rect 342678 620912 342802 621012
rect 342902 620912 343026 621012
rect 343126 620912 343158 621012
rect 342100 620788 343158 620912
rect 342100 620688 342130 620788
rect 342230 620688 342354 620788
rect 342454 620688 342578 620788
rect 342678 620688 342802 620788
rect 342902 620688 343026 620788
rect 343126 620688 343158 620788
rect 342100 620564 343158 620688
rect 342100 620464 342130 620564
rect 342230 620464 342354 620564
rect 342454 620464 342578 620564
rect 342678 620464 342802 620564
rect 342902 620464 343026 620564
rect 343126 620464 343158 620564
rect 342100 620340 343158 620464
rect 342100 620240 342130 620340
rect 342230 620240 342354 620340
rect 342454 620240 342578 620340
rect 342678 620240 342802 620340
rect 342902 620240 343026 620340
rect 343126 620240 343158 620340
rect 342100 620116 343158 620240
rect 342100 620016 342130 620116
rect 342230 620016 342354 620116
rect 342454 620016 342578 620116
rect 342678 620016 342802 620116
rect 342902 620016 343026 620116
rect 343126 620016 343158 620116
rect 342100 619892 343158 620016
rect 342100 619792 342130 619892
rect 342230 619792 342354 619892
rect 342454 619792 342578 619892
rect 342678 619792 342802 619892
rect 342902 619792 343026 619892
rect 343126 619792 343158 619892
rect 342100 619668 343158 619792
rect 342100 619568 342130 619668
rect 342230 619568 342354 619668
rect 342454 619568 342578 619668
rect 342678 619568 342802 619668
rect 342902 619568 343026 619668
rect 343126 619568 343158 619668
rect 342100 619444 343158 619568
rect 342100 619344 342130 619444
rect 342230 619344 342354 619444
rect 342454 619344 342578 619444
rect 342678 619344 342802 619444
rect 342902 619344 343026 619444
rect 343126 619344 343158 619444
rect 342100 619220 343158 619344
rect 342100 619120 342130 619220
rect 342230 619120 342354 619220
rect 342454 619120 342578 619220
rect 342678 619120 342802 619220
rect 342902 619120 343026 619220
rect 343126 619120 343158 619220
rect 342100 618996 343158 619120
rect 342100 618896 342130 618996
rect 342230 618896 342354 618996
rect 342454 618896 342578 618996
rect 342678 618896 342802 618996
rect 342902 618896 343026 618996
rect 343126 618896 343158 618996
rect 342100 618772 343158 618896
rect 342100 618672 342130 618772
rect 342230 618672 342354 618772
rect 342454 618672 342578 618772
rect 342678 618672 342802 618772
rect 342902 618672 343026 618772
rect 343126 618672 343158 618772
rect 342100 618548 343158 618672
rect 342100 618448 342130 618548
rect 342230 618448 342354 618548
rect 342454 618448 342578 618548
rect 342678 618448 342802 618548
rect 342902 618448 343026 618548
rect 343126 618448 343158 618548
rect 342100 618324 343158 618448
rect 342100 618224 342130 618324
rect 342230 618224 342354 618324
rect 342454 618224 342578 618324
rect 342678 618224 342802 618324
rect 342902 618224 343026 618324
rect 343126 618224 343158 618324
rect 342100 618100 343158 618224
rect 342100 618000 342130 618100
rect 342230 618000 342354 618100
rect 342454 618000 342578 618100
rect 342678 618000 342802 618100
rect 342902 618000 343026 618100
rect 343126 618000 343158 618100
rect 342100 617980 343158 618000
rect 298836 615474 305496 615504
rect 298836 615374 298876 615474
rect 298976 615374 299100 615474
rect 299200 615374 299324 615474
rect 299424 615374 299548 615474
rect 299648 615374 299772 615474
rect 299872 615374 299996 615474
rect 300096 615374 300220 615474
rect 300320 615374 300444 615474
rect 300544 615374 300668 615474
rect 300768 615374 300892 615474
rect 300992 615374 301116 615474
rect 301216 615374 301340 615474
rect 301440 615374 301564 615474
rect 301664 615374 301788 615474
rect 301888 615374 302012 615474
rect 302112 615374 302236 615474
rect 302336 615374 302460 615474
rect 302560 615374 302684 615474
rect 302784 615374 302908 615474
rect 303008 615374 303132 615474
rect 303232 615374 303356 615474
rect 303456 615374 303580 615474
rect 303680 615374 303804 615474
rect 303904 615374 304028 615474
rect 304128 615374 304252 615474
rect 304352 615374 304476 615474
rect 304576 615374 304700 615474
rect 304800 615374 304924 615474
rect 305024 615374 305148 615474
rect 305248 615374 305372 615474
rect 305472 615374 305496 615474
rect 298836 615250 305496 615374
rect 298836 615150 298876 615250
rect 298976 615150 299100 615250
rect 299200 615150 299324 615250
rect 299424 615150 299548 615250
rect 299648 615150 299772 615250
rect 299872 615150 299996 615250
rect 300096 615150 300220 615250
rect 300320 615150 300444 615250
rect 300544 615150 300668 615250
rect 300768 615150 300892 615250
rect 300992 615150 301116 615250
rect 301216 615150 301340 615250
rect 301440 615150 301564 615250
rect 301664 615150 301788 615250
rect 301888 615150 302012 615250
rect 302112 615150 302236 615250
rect 302336 615150 302460 615250
rect 302560 615150 302684 615250
rect 302784 615150 302908 615250
rect 303008 615150 303132 615250
rect 303232 615150 303356 615250
rect 303456 615150 303580 615250
rect 303680 615150 303804 615250
rect 303904 615150 304028 615250
rect 304128 615150 304252 615250
rect 304352 615150 304476 615250
rect 304576 615150 304700 615250
rect 304800 615150 304924 615250
rect 305024 615150 305148 615250
rect 305248 615150 305372 615250
rect 305472 615150 305496 615250
rect 298836 615026 305496 615150
rect 298836 614926 298876 615026
rect 298976 614926 299100 615026
rect 299200 614926 299324 615026
rect 299424 614926 299548 615026
rect 299648 614926 299772 615026
rect 299872 614926 299996 615026
rect 300096 614926 300220 615026
rect 300320 614926 300444 615026
rect 300544 614926 300668 615026
rect 300768 614926 300892 615026
rect 300992 614926 301116 615026
rect 301216 614926 301340 615026
rect 301440 614926 301564 615026
rect 301664 614926 301788 615026
rect 301888 614926 302012 615026
rect 302112 614926 302236 615026
rect 302336 614926 302460 615026
rect 302560 614926 302684 615026
rect 302784 614926 302908 615026
rect 303008 614926 303132 615026
rect 303232 614926 303356 615026
rect 303456 614926 303580 615026
rect 303680 614926 303804 615026
rect 303904 614926 304028 615026
rect 304128 614926 304252 615026
rect 304352 614926 304476 615026
rect 304576 614926 304700 615026
rect 304800 614926 304924 615026
rect 305024 614926 305148 615026
rect 305248 614926 305372 615026
rect 305472 614926 305496 615026
rect 298836 614802 305496 614926
rect 298836 614702 298876 614802
rect 298976 614702 299100 614802
rect 299200 614702 299324 614802
rect 299424 614702 299548 614802
rect 299648 614702 299772 614802
rect 299872 614702 299996 614802
rect 300096 614702 300220 614802
rect 300320 614702 300444 614802
rect 300544 614702 300668 614802
rect 300768 614702 300892 614802
rect 300992 614702 301116 614802
rect 301216 614702 301340 614802
rect 301440 614702 301564 614802
rect 301664 614702 301788 614802
rect 301888 614702 302012 614802
rect 302112 614702 302236 614802
rect 302336 614702 302460 614802
rect 302560 614702 302684 614802
rect 302784 614702 302908 614802
rect 303008 614702 303132 614802
rect 303232 614702 303356 614802
rect 303456 614702 303580 614802
rect 303680 614702 303804 614802
rect 303904 614702 304028 614802
rect 304128 614702 304252 614802
rect 304352 614702 304476 614802
rect 304576 614702 304700 614802
rect 304800 614702 304924 614802
rect 305024 614702 305148 614802
rect 305248 614702 305372 614802
rect 305472 614702 305496 614802
rect 298836 614578 305496 614702
rect 298836 614478 298876 614578
rect 298976 614478 299100 614578
rect 299200 614478 299324 614578
rect 299424 614478 299548 614578
rect 299648 614478 299772 614578
rect 299872 614478 299996 614578
rect 300096 614478 300220 614578
rect 300320 614478 300444 614578
rect 300544 614478 300668 614578
rect 300768 614478 300892 614578
rect 300992 614478 301116 614578
rect 301216 614478 301340 614578
rect 301440 614478 301564 614578
rect 301664 614478 301788 614578
rect 301888 614478 302012 614578
rect 302112 614478 302236 614578
rect 302336 614478 302460 614578
rect 302560 614478 302684 614578
rect 302784 614478 302908 614578
rect 303008 614478 303132 614578
rect 303232 614478 303356 614578
rect 303456 614478 303580 614578
rect 303680 614478 303804 614578
rect 303904 614478 304028 614578
rect 304128 614478 304252 614578
rect 304352 614478 304476 614578
rect 304576 614478 304700 614578
rect 304800 614478 304924 614578
rect 305024 614478 305148 614578
rect 305248 614478 305372 614578
rect 305472 614478 305496 614578
rect 298836 614444 305496 614478
rect 309306 615474 315966 615504
rect 309306 615374 309346 615474
rect 309446 615374 309570 615474
rect 309670 615374 309794 615474
rect 309894 615374 310018 615474
rect 310118 615374 310242 615474
rect 310342 615374 310466 615474
rect 310566 615374 310690 615474
rect 310790 615374 310914 615474
rect 311014 615374 311138 615474
rect 311238 615374 311362 615474
rect 311462 615374 311586 615474
rect 311686 615374 311810 615474
rect 311910 615374 312034 615474
rect 312134 615374 312258 615474
rect 312358 615374 312482 615474
rect 312582 615374 312706 615474
rect 312806 615374 312930 615474
rect 313030 615374 313154 615474
rect 313254 615374 313378 615474
rect 313478 615374 313602 615474
rect 313702 615374 313826 615474
rect 313926 615374 314050 615474
rect 314150 615374 314274 615474
rect 314374 615374 314498 615474
rect 314598 615374 314722 615474
rect 314822 615374 314946 615474
rect 315046 615374 315170 615474
rect 315270 615374 315394 615474
rect 315494 615374 315618 615474
rect 315718 615374 315842 615474
rect 315942 615374 315966 615474
rect 309306 615250 315966 615374
rect 309306 615150 309346 615250
rect 309446 615150 309570 615250
rect 309670 615150 309794 615250
rect 309894 615150 310018 615250
rect 310118 615150 310242 615250
rect 310342 615150 310466 615250
rect 310566 615150 310690 615250
rect 310790 615150 310914 615250
rect 311014 615150 311138 615250
rect 311238 615150 311362 615250
rect 311462 615150 311586 615250
rect 311686 615150 311810 615250
rect 311910 615150 312034 615250
rect 312134 615150 312258 615250
rect 312358 615150 312482 615250
rect 312582 615150 312706 615250
rect 312806 615150 312930 615250
rect 313030 615150 313154 615250
rect 313254 615150 313378 615250
rect 313478 615150 313602 615250
rect 313702 615150 313826 615250
rect 313926 615150 314050 615250
rect 314150 615150 314274 615250
rect 314374 615150 314498 615250
rect 314598 615150 314722 615250
rect 314822 615150 314946 615250
rect 315046 615150 315170 615250
rect 315270 615150 315394 615250
rect 315494 615150 315618 615250
rect 315718 615150 315842 615250
rect 315942 615150 315966 615250
rect 309306 615026 315966 615150
rect 309306 614926 309346 615026
rect 309446 614926 309570 615026
rect 309670 614926 309794 615026
rect 309894 614926 310018 615026
rect 310118 614926 310242 615026
rect 310342 614926 310466 615026
rect 310566 614926 310690 615026
rect 310790 614926 310914 615026
rect 311014 614926 311138 615026
rect 311238 614926 311362 615026
rect 311462 614926 311586 615026
rect 311686 614926 311810 615026
rect 311910 614926 312034 615026
rect 312134 614926 312258 615026
rect 312358 614926 312482 615026
rect 312582 614926 312706 615026
rect 312806 614926 312930 615026
rect 313030 614926 313154 615026
rect 313254 614926 313378 615026
rect 313478 614926 313602 615026
rect 313702 614926 313826 615026
rect 313926 614926 314050 615026
rect 314150 614926 314274 615026
rect 314374 614926 314498 615026
rect 314598 614926 314722 615026
rect 314822 614926 314946 615026
rect 315046 614926 315170 615026
rect 315270 614926 315394 615026
rect 315494 614926 315618 615026
rect 315718 614926 315842 615026
rect 315942 614926 315966 615026
rect 309306 614802 315966 614926
rect 309306 614702 309346 614802
rect 309446 614702 309570 614802
rect 309670 614702 309794 614802
rect 309894 614702 310018 614802
rect 310118 614702 310242 614802
rect 310342 614702 310466 614802
rect 310566 614702 310690 614802
rect 310790 614702 310914 614802
rect 311014 614702 311138 614802
rect 311238 614702 311362 614802
rect 311462 614702 311586 614802
rect 311686 614702 311810 614802
rect 311910 614702 312034 614802
rect 312134 614702 312258 614802
rect 312358 614702 312482 614802
rect 312582 614702 312706 614802
rect 312806 614702 312930 614802
rect 313030 614702 313154 614802
rect 313254 614702 313378 614802
rect 313478 614702 313602 614802
rect 313702 614702 313826 614802
rect 313926 614702 314050 614802
rect 314150 614702 314274 614802
rect 314374 614702 314498 614802
rect 314598 614702 314722 614802
rect 314822 614702 314946 614802
rect 315046 614702 315170 614802
rect 315270 614702 315394 614802
rect 315494 614702 315618 614802
rect 315718 614702 315842 614802
rect 315942 614702 315966 614802
rect 309306 614578 315966 614702
rect 309306 614478 309346 614578
rect 309446 614478 309570 614578
rect 309670 614478 309794 614578
rect 309894 614478 310018 614578
rect 310118 614478 310242 614578
rect 310342 614478 310466 614578
rect 310566 614478 310690 614578
rect 310790 614478 310914 614578
rect 311014 614478 311138 614578
rect 311238 614478 311362 614578
rect 311462 614478 311586 614578
rect 311686 614478 311810 614578
rect 311910 614478 312034 614578
rect 312134 614478 312258 614578
rect 312358 614478 312482 614578
rect 312582 614478 312706 614578
rect 312806 614478 312930 614578
rect 313030 614478 313154 614578
rect 313254 614478 313378 614578
rect 313478 614478 313602 614578
rect 313702 614478 313826 614578
rect 313926 614478 314050 614578
rect 314150 614478 314274 614578
rect 314374 614478 314498 614578
rect 314598 614478 314722 614578
rect 314822 614478 314946 614578
rect 315046 614478 315170 614578
rect 315270 614478 315394 614578
rect 315494 614478 315618 614578
rect 315718 614478 315842 614578
rect 315942 614478 315966 614578
rect 309306 614444 315966 614478
rect 335576 615494 342236 615524
rect 335576 615394 335616 615494
rect 335716 615394 335840 615494
rect 335940 615394 336064 615494
rect 336164 615394 336288 615494
rect 336388 615394 336512 615494
rect 336612 615394 336736 615494
rect 336836 615394 336960 615494
rect 337060 615394 337184 615494
rect 337284 615394 337408 615494
rect 337508 615394 337632 615494
rect 337732 615394 337856 615494
rect 337956 615394 338080 615494
rect 338180 615394 338304 615494
rect 338404 615394 338528 615494
rect 338628 615394 338752 615494
rect 338852 615394 338976 615494
rect 339076 615394 339200 615494
rect 339300 615394 339424 615494
rect 339524 615394 339648 615494
rect 339748 615394 339872 615494
rect 339972 615394 340096 615494
rect 340196 615394 340320 615494
rect 340420 615394 340544 615494
rect 340644 615394 340768 615494
rect 340868 615394 340992 615494
rect 341092 615394 341216 615494
rect 341316 615394 341440 615494
rect 341540 615394 341664 615494
rect 341764 615394 341888 615494
rect 341988 615394 342112 615494
rect 342212 615394 342236 615494
rect 335576 615270 342236 615394
rect 335576 615170 335616 615270
rect 335716 615170 335840 615270
rect 335940 615170 336064 615270
rect 336164 615170 336288 615270
rect 336388 615170 336512 615270
rect 336612 615170 336736 615270
rect 336836 615170 336960 615270
rect 337060 615170 337184 615270
rect 337284 615170 337408 615270
rect 337508 615170 337632 615270
rect 337732 615170 337856 615270
rect 337956 615170 338080 615270
rect 338180 615170 338304 615270
rect 338404 615170 338528 615270
rect 338628 615170 338752 615270
rect 338852 615170 338976 615270
rect 339076 615170 339200 615270
rect 339300 615170 339424 615270
rect 339524 615170 339648 615270
rect 339748 615170 339872 615270
rect 339972 615170 340096 615270
rect 340196 615170 340320 615270
rect 340420 615170 340544 615270
rect 340644 615170 340768 615270
rect 340868 615170 340992 615270
rect 341092 615170 341216 615270
rect 341316 615170 341440 615270
rect 341540 615170 341664 615270
rect 341764 615170 341888 615270
rect 341988 615170 342112 615270
rect 342212 615170 342236 615270
rect 335576 615046 342236 615170
rect 335576 614946 335616 615046
rect 335716 614946 335840 615046
rect 335940 614946 336064 615046
rect 336164 614946 336288 615046
rect 336388 614946 336512 615046
rect 336612 614946 336736 615046
rect 336836 614946 336960 615046
rect 337060 614946 337184 615046
rect 337284 614946 337408 615046
rect 337508 614946 337632 615046
rect 337732 614946 337856 615046
rect 337956 614946 338080 615046
rect 338180 614946 338304 615046
rect 338404 614946 338528 615046
rect 338628 614946 338752 615046
rect 338852 614946 338976 615046
rect 339076 614946 339200 615046
rect 339300 614946 339424 615046
rect 339524 614946 339648 615046
rect 339748 614946 339872 615046
rect 339972 614946 340096 615046
rect 340196 614946 340320 615046
rect 340420 614946 340544 615046
rect 340644 614946 340768 615046
rect 340868 614946 340992 615046
rect 341092 614946 341216 615046
rect 341316 614946 341440 615046
rect 341540 614946 341664 615046
rect 341764 614946 341888 615046
rect 341988 614946 342112 615046
rect 342212 614946 342236 615046
rect 335576 614822 342236 614946
rect 335576 614722 335616 614822
rect 335716 614722 335840 614822
rect 335940 614722 336064 614822
rect 336164 614722 336288 614822
rect 336388 614722 336512 614822
rect 336612 614722 336736 614822
rect 336836 614722 336960 614822
rect 337060 614722 337184 614822
rect 337284 614722 337408 614822
rect 337508 614722 337632 614822
rect 337732 614722 337856 614822
rect 337956 614722 338080 614822
rect 338180 614722 338304 614822
rect 338404 614722 338528 614822
rect 338628 614722 338752 614822
rect 338852 614722 338976 614822
rect 339076 614722 339200 614822
rect 339300 614722 339424 614822
rect 339524 614722 339648 614822
rect 339748 614722 339872 614822
rect 339972 614722 340096 614822
rect 340196 614722 340320 614822
rect 340420 614722 340544 614822
rect 340644 614722 340768 614822
rect 340868 614722 340992 614822
rect 341092 614722 341216 614822
rect 341316 614722 341440 614822
rect 341540 614722 341664 614822
rect 341764 614722 341888 614822
rect 341988 614722 342112 614822
rect 342212 614722 342236 614822
rect 335576 614598 342236 614722
rect 335576 614498 335616 614598
rect 335716 614498 335840 614598
rect 335940 614498 336064 614598
rect 336164 614498 336288 614598
rect 336388 614498 336512 614598
rect 336612 614498 336736 614598
rect 336836 614498 336960 614598
rect 337060 614498 337184 614598
rect 337284 614498 337408 614598
rect 337508 614498 337632 614598
rect 337732 614498 337856 614598
rect 337956 614498 338080 614598
rect 338180 614498 338304 614598
rect 338404 614498 338528 614598
rect 338628 614498 338752 614598
rect 338852 614498 338976 614598
rect 339076 614498 339200 614598
rect 339300 614498 339424 614598
rect 339524 614498 339648 614598
rect 339748 614498 339872 614598
rect 339972 614498 340096 614598
rect 340196 614498 340320 614598
rect 340420 614498 340544 614598
rect 340644 614498 340768 614598
rect 340868 614498 340992 614598
rect 341092 614498 341216 614598
rect 341316 614498 341440 614598
rect 341540 614498 341664 614598
rect 341764 614498 341888 614598
rect 341988 614498 342112 614598
rect 342212 614498 342236 614598
rect 335576 614464 342236 614498
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 298876 642594 298976 642694
rect 299100 642594 299200 642694
rect 299324 642594 299424 642694
rect 299548 642594 299648 642694
rect 299772 642594 299872 642694
rect 299996 642594 300096 642694
rect 300220 642594 300320 642694
rect 300444 642594 300544 642694
rect 300668 642594 300768 642694
rect 300892 642594 300992 642694
rect 301116 642594 301216 642694
rect 301340 642594 301440 642694
rect 301564 642594 301664 642694
rect 301788 642594 301888 642694
rect 302012 642594 302112 642694
rect 302236 642594 302336 642694
rect 302460 642594 302560 642694
rect 302684 642594 302784 642694
rect 302908 642594 303008 642694
rect 303132 642594 303232 642694
rect 303356 642594 303456 642694
rect 303580 642594 303680 642694
rect 303804 642594 303904 642694
rect 304028 642594 304128 642694
rect 304252 642594 304352 642694
rect 304476 642594 304576 642694
rect 304700 642594 304800 642694
rect 304924 642594 305024 642694
rect 305148 642594 305248 642694
rect 305372 642594 305472 642694
rect 298876 642370 298976 642470
rect 299100 642370 299200 642470
rect 299324 642370 299424 642470
rect 299548 642370 299648 642470
rect 299772 642370 299872 642470
rect 299996 642370 300096 642470
rect 300220 642370 300320 642470
rect 300444 642370 300544 642470
rect 300668 642370 300768 642470
rect 300892 642370 300992 642470
rect 301116 642370 301216 642470
rect 301340 642370 301440 642470
rect 301564 642370 301664 642470
rect 301788 642370 301888 642470
rect 302012 642370 302112 642470
rect 302236 642370 302336 642470
rect 302460 642370 302560 642470
rect 302684 642370 302784 642470
rect 302908 642370 303008 642470
rect 303132 642370 303232 642470
rect 303356 642370 303456 642470
rect 303580 642370 303680 642470
rect 303804 642370 303904 642470
rect 304028 642370 304128 642470
rect 304252 642370 304352 642470
rect 304476 642370 304576 642470
rect 304700 642370 304800 642470
rect 304924 642370 305024 642470
rect 305148 642370 305248 642470
rect 305372 642370 305472 642470
rect 298876 642146 298976 642246
rect 299100 642146 299200 642246
rect 299324 642146 299424 642246
rect 299548 642146 299648 642246
rect 299772 642146 299872 642246
rect 299996 642146 300096 642246
rect 300220 642146 300320 642246
rect 300444 642146 300544 642246
rect 300668 642146 300768 642246
rect 300892 642146 300992 642246
rect 301116 642146 301216 642246
rect 301340 642146 301440 642246
rect 301564 642146 301664 642246
rect 301788 642146 301888 642246
rect 302012 642146 302112 642246
rect 302236 642146 302336 642246
rect 302460 642146 302560 642246
rect 302684 642146 302784 642246
rect 302908 642146 303008 642246
rect 303132 642146 303232 642246
rect 303356 642146 303456 642246
rect 303580 642146 303680 642246
rect 303804 642146 303904 642246
rect 304028 642146 304128 642246
rect 304252 642146 304352 642246
rect 304476 642146 304576 642246
rect 304700 642146 304800 642246
rect 304924 642146 305024 642246
rect 305148 642146 305248 642246
rect 305372 642146 305472 642246
rect 298876 641922 298976 642022
rect 299100 641922 299200 642022
rect 299324 641922 299424 642022
rect 299548 641922 299648 642022
rect 299772 641922 299872 642022
rect 299996 641922 300096 642022
rect 300220 641922 300320 642022
rect 300444 641922 300544 642022
rect 300668 641922 300768 642022
rect 300892 641922 300992 642022
rect 301116 641922 301216 642022
rect 301340 641922 301440 642022
rect 301564 641922 301664 642022
rect 301788 641922 301888 642022
rect 302012 641922 302112 642022
rect 302236 641922 302336 642022
rect 302460 641922 302560 642022
rect 302684 641922 302784 642022
rect 302908 641922 303008 642022
rect 303132 641922 303232 642022
rect 303356 641922 303456 642022
rect 303580 641922 303680 642022
rect 303804 641922 303904 642022
rect 304028 641922 304128 642022
rect 304252 641922 304352 642022
rect 304476 641922 304576 642022
rect 304700 641922 304800 642022
rect 304924 641922 305024 642022
rect 305148 641922 305248 642022
rect 305372 641922 305472 642022
rect 298876 641698 298976 641798
rect 299100 641698 299200 641798
rect 299324 641698 299424 641798
rect 299548 641698 299648 641798
rect 299772 641698 299872 641798
rect 299996 641698 300096 641798
rect 300220 641698 300320 641798
rect 300444 641698 300544 641798
rect 300668 641698 300768 641798
rect 300892 641698 300992 641798
rect 301116 641698 301216 641798
rect 301340 641698 301440 641798
rect 301564 641698 301664 641798
rect 301788 641698 301888 641798
rect 302012 641698 302112 641798
rect 302236 641698 302336 641798
rect 302460 641698 302560 641798
rect 302684 641698 302784 641798
rect 302908 641698 303008 641798
rect 303132 641698 303232 641798
rect 303356 641698 303456 641798
rect 303580 641698 303680 641798
rect 303804 641698 303904 641798
rect 304028 641698 304128 641798
rect 304252 641698 304352 641798
rect 304476 641698 304576 641798
rect 304700 641698 304800 641798
rect 304924 641698 305024 641798
rect 305148 641698 305248 641798
rect 305372 641698 305472 641798
rect 309346 642594 309446 642694
rect 309570 642594 309670 642694
rect 309794 642594 309894 642694
rect 310018 642594 310118 642694
rect 310242 642594 310342 642694
rect 310466 642594 310566 642694
rect 310690 642594 310790 642694
rect 310914 642594 311014 642694
rect 311138 642594 311238 642694
rect 311362 642594 311462 642694
rect 311586 642594 311686 642694
rect 311810 642594 311910 642694
rect 312034 642594 312134 642694
rect 312258 642594 312358 642694
rect 312482 642594 312582 642694
rect 312706 642594 312806 642694
rect 312930 642594 313030 642694
rect 313154 642594 313254 642694
rect 313378 642594 313478 642694
rect 313602 642594 313702 642694
rect 313826 642594 313926 642694
rect 314050 642594 314150 642694
rect 314274 642594 314374 642694
rect 314498 642594 314598 642694
rect 314722 642594 314822 642694
rect 314946 642594 315046 642694
rect 315170 642594 315270 642694
rect 315394 642594 315494 642694
rect 315618 642594 315718 642694
rect 315842 642594 315942 642694
rect 309346 642370 309446 642470
rect 309570 642370 309670 642470
rect 309794 642370 309894 642470
rect 310018 642370 310118 642470
rect 310242 642370 310342 642470
rect 310466 642370 310566 642470
rect 310690 642370 310790 642470
rect 310914 642370 311014 642470
rect 311138 642370 311238 642470
rect 311362 642370 311462 642470
rect 311586 642370 311686 642470
rect 311810 642370 311910 642470
rect 312034 642370 312134 642470
rect 312258 642370 312358 642470
rect 312482 642370 312582 642470
rect 312706 642370 312806 642470
rect 312930 642370 313030 642470
rect 313154 642370 313254 642470
rect 313378 642370 313478 642470
rect 313602 642370 313702 642470
rect 313826 642370 313926 642470
rect 314050 642370 314150 642470
rect 314274 642370 314374 642470
rect 314498 642370 314598 642470
rect 314722 642370 314822 642470
rect 314946 642370 315046 642470
rect 315170 642370 315270 642470
rect 315394 642370 315494 642470
rect 315618 642370 315718 642470
rect 315842 642370 315942 642470
rect 309346 642146 309446 642246
rect 309570 642146 309670 642246
rect 309794 642146 309894 642246
rect 310018 642146 310118 642246
rect 310242 642146 310342 642246
rect 310466 642146 310566 642246
rect 310690 642146 310790 642246
rect 310914 642146 311014 642246
rect 311138 642146 311238 642246
rect 311362 642146 311462 642246
rect 311586 642146 311686 642246
rect 311810 642146 311910 642246
rect 312034 642146 312134 642246
rect 312258 642146 312358 642246
rect 312482 642146 312582 642246
rect 312706 642146 312806 642246
rect 312930 642146 313030 642246
rect 313154 642146 313254 642246
rect 313378 642146 313478 642246
rect 313602 642146 313702 642246
rect 313826 642146 313926 642246
rect 314050 642146 314150 642246
rect 314274 642146 314374 642246
rect 314498 642146 314598 642246
rect 314722 642146 314822 642246
rect 314946 642146 315046 642246
rect 315170 642146 315270 642246
rect 315394 642146 315494 642246
rect 315618 642146 315718 642246
rect 315842 642146 315942 642246
rect 309346 641922 309446 642022
rect 309570 641922 309670 642022
rect 309794 641922 309894 642022
rect 310018 641922 310118 642022
rect 310242 641922 310342 642022
rect 310466 641922 310566 642022
rect 310690 641922 310790 642022
rect 310914 641922 311014 642022
rect 311138 641922 311238 642022
rect 311362 641922 311462 642022
rect 311586 641922 311686 642022
rect 311810 641922 311910 642022
rect 312034 641922 312134 642022
rect 312258 641922 312358 642022
rect 312482 641922 312582 642022
rect 312706 641922 312806 642022
rect 312930 641922 313030 642022
rect 313154 641922 313254 642022
rect 313378 641922 313478 642022
rect 313602 641922 313702 642022
rect 313826 641922 313926 642022
rect 314050 641922 314150 642022
rect 314274 641922 314374 642022
rect 314498 641922 314598 642022
rect 314722 641922 314822 642022
rect 314946 641922 315046 642022
rect 315170 641922 315270 642022
rect 315394 641922 315494 642022
rect 315618 641922 315718 642022
rect 315842 641922 315942 642022
rect 309346 641698 309446 641798
rect 309570 641698 309670 641798
rect 309794 641698 309894 641798
rect 310018 641698 310118 641798
rect 310242 641698 310342 641798
rect 310466 641698 310566 641798
rect 310690 641698 310790 641798
rect 310914 641698 311014 641798
rect 311138 641698 311238 641798
rect 311362 641698 311462 641798
rect 311586 641698 311686 641798
rect 311810 641698 311910 641798
rect 312034 641698 312134 641798
rect 312258 641698 312358 641798
rect 312482 641698 312582 641798
rect 312706 641698 312806 641798
rect 312930 641698 313030 641798
rect 313154 641698 313254 641798
rect 313378 641698 313478 641798
rect 313602 641698 313702 641798
rect 313826 641698 313926 641798
rect 314050 641698 314150 641798
rect 314274 641698 314374 641798
rect 314498 641698 314598 641798
rect 314722 641698 314822 641798
rect 314946 641698 315046 641798
rect 315170 641698 315270 641798
rect 315394 641698 315494 641798
rect 315618 641698 315718 641798
rect 315842 641698 315942 641798
rect 335616 642614 335716 642714
rect 335840 642614 335940 642714
rect 336064 642614 336164 642714
rect 336288 642614 336388 642714
rect 336512 642614 336612 642714
rect 336736 642614 336836 642714
rect 336960 642614 337060 642714
rect 337184 642614 337284 642714
rect 337408 642614 337508 642714
rect 337632 642614 337732 642714
rect 337856 642614 337956 642714
rect 338080 642614 338180 642714
rect 338304 642614 338404 642714
rect 338528 642614 338628 642714
rect 338752 642614 338852 642714
rect 338976 642614 339076 642714
rect 339200 642614 339300 642714
rect 339424 642614 339524 642714
rect 339648 642614 339748 642714
rect 339872 642614 339972 642714
rect 340096 642614 340196 642714
rect 340320 642614 340420 642714
rect 340544 642614 340644 642714
rect 340768 642614 340868 642714
rect 340992 642614 341092 642714
rect 341216 642614 341316 642714
rect 341440 642614 341540 642714
rect 341664 642614 341764 642714
rect 341888 642614 341988 642714
rect 342112 642614 342212 642714
rect 335616 642390 335716 642490
rect 335840 642390 335940 642490
rect 336064 642390 336164 642490
rect 336288 642390 336388 642490
rect 336512 642390 336612 642490
rect 336736 642390 336836 642490
rect 336960 642390 337060 642490
rect 337184 642390 337284 642490
rect 337408 642390 337508 642490
rect 337632 642390 337732 642490
rect 337856 642390 337956 642490
rect 338080 642390 338180 642490
rect 338304 642390 338404 642490
rect 338528 642390 338628 642490
rect 338752 642390 338852 642490
rect 338976 642390 339076 642490
rect 339200 642390 339300 642490
rect 339424 642390 339524 642490
rect 339648 642390 339748 642490
rect 339872 642390 339972 642490
rect 340096 642390 340196 642490
rect 340320 642390 340420 642490
rect 340544 642390 340644 642490
rect 340768 642390 340868 642490
rect 340992 642390 341092 642490
rect 341216 642390 341316 642490
rect 341440 642390 341540 642490
rect 341664 642390 341764 642490
rect 341888 642390 341988 642490
rect 342112 642390 342212 642490
rect 335616 642166 335716 642266
rect 335840 642166 335940 642266
rect 336064 642166 336164 642266
rect 336288 642166 336388 642266
rect 336512 642166 336612 642266
rect 336736 642166 336836 642266
rect 336960 642166 337060 642266
rect 337184 642166 337284 642266
rect 337408 642166 337508 642266
rect 337632 642166 337732 642266
rect 337856 642166 337956 642266
rect 338080 642166 338180 642266
rect 338304 642166 338404 642266
rect 338528 642166 338628 642266
rect 338752 642166 338852 642266
rect 338976 642166 339076 642266
rect 339200 642166 339300 642266
rect 339424 642166 339524 642266
rect 339648 642166 339748 642266
rect 339872 642166 339972 642266
rect 340096 642166 340196 642266
rect 340320 642166 340420 642266
rect 340544 642166 340644 642266
rect 340768 642166 340868 642266
rect 340992 642166 341092 642266
rect 341216 642166 341316 642266
rect 341440 642166 341540 642266
rect 341664 642166 341764 642266
rect 341888 642166 341988 642266
rect 342112 642166 342212 642266
rect 335616 641942 335716 642042
rect 335840 641942 335940 642042
rect 336064 641942 336164 642042
rect 336288 641942 336388 642042
rect 336512 641942 336612 642042
rect 336736 641942 336836 642042
rect 336960 641942 337060 642042
rect 337184 641942 337284 642042
rect 337408 641942 337508 642042
rect 337632 641942 337732 642042
rect 337856 641942 337956 642042
rect 338080 641942 338180 642042
rect 338304 641942 338404 642042
rect 338528 641942 338628 642042
rect 338752 641942 338852 642042
rect 338976 641942 339076 642042
rect 339200 641942 339300 642042
rect 339424 641942 339524 642042
rect 339648 641942 339748 642042
rect 339872 641942 339972 642042
rect 340096 641942 340196 642042
rect 340320 641942 340420 642042
rect 340544 641942 340644 642042
rect 340768 641942 340868 642042
rect 340992 641942 341092 642042
rect 341216 641942 341316 642042
rect 341440 641942 341540 642042
rect 341664 641942 341764 642042
rect 341888 641942 341988 642042
rect 342112 641942 342212 642042
rect 335616 641718 335716 641818
rect 335840 641718 335940 641818
rect 336064 641718 336164 641818
rect 336288 641718 336388 641818
rect 336512 641718 336612 641818
rect 336736 641718 336836 641818
rect 336960 641718 337060 641818
rect 337184 641718 337284 641818
rect 337408 641718 337508 641818
rect 337632 641718 337732 641818
rect 337856 641718 337956 641818
rect 338080 641718 338180 641818
rect 338304 641718 338404 641818
rect 338528 641718 338628 641818
rect 338752 641718 338852 641818
rect 338976 641718 339076 641818
rect 339200 641718 339300 641818
rect 339424 641718 339524 641818
rect 339648 641718 339748 641818
rect 339872 641718 339972 641818
rect 340096 641718 340196 641818
rect 340320 641718 340420 641818
rect 340544 641718 340644 641818
rect 340768 641718 340868 641818
rect 340992 641718 341092 641818
rect 341216 641718 341316 641818
rect 341440 641718 341540 641818
rect 341664 641718 341764 641818
rect 341888 641718 341988 641818
rect 342112 641718 342212 641818
rect 297850 637896 297950 637996
rect 298074 637896 298174 637996
rect 298298 637896 298398 637996
rect 298522 637896 298622 637996
rect 298746 637896 298846 637996
rect 297850 637672 297950 637772
rect 298074 637672 298174 637772
rect 298298 637672 298398 637772
rect 298522 637672 298622 637772
rect 298746 637672 298846 637772
rect 297850 637448 297950 637548
rect 298074 637448 298174 637548
rect 298298 637448 298398 637548
rect 298522 637448 298622 637548
rect 298746 637448 298846 637548
rect 297850 637224 297950 637324
rect 298074 637224 298174 637324
rect 298298 637224 298398 637324
rect 298522 637224 298622 637324
rect 298746 637224 298846 637324
rect 297850 637000 297950 637100
rect 298074 637000 298174 637100
rect 298298 637000 298398 637100
rect 298522 637000 298622 637100
rect 298746 637000 298846 637100
rect 297850 636776 297950 636876
rect 298074 636776 298174 636876
rect 298298 636776 298398 636876
rect 298522 636776 298622 636876
rect 298746 636776 298846 636876
rect 297850 636552 297950 636652
rect 298074 636552 298174 636652
rect 298298 636552 298398 636652
rect 298522 636552 298622 636652
rect 298746 636552 298846 636652
rect 297850 636328 297950 636428
rect 298074 636328 298174 636428
rect 298298 636328 298398 636428
rect 298522 636328 298622 636428
rect 298746 636328 298846 636428
rect 297850 636104 297950 636204
rect 298074 636104 298174 636204
rect 298298 636104 298398 636204
rect 298522 636104 298622 636204
rect 298746 636104 298846 636204
rect 297850 635880 297950 635980
rect 298074 635880 298174 635980
rect 298298 635880 298398 635980
rect 298522 635880 298622 635980
rect 298746 635880 298846 635980
rect 297850 635656 297950 635756
rect 298074 635656 298174 635756
rect 298298 635656 298398 635756
rect 298522 635656 298622 635756
rect 298746 635656 298846 635756
rect 297850 635432 297950 635532
rect 298074 635432 298174 635532
rect 298298 635432 298398 635532
rect 298522 635432 298622 635532
rect 298746 635432 298846 635532
rect 297850 635208 297950 635308
rect 298074 635208 298174 635308
rect 298298 635208 298398 635308
rect 298522 635208 298622 635308
rect 298746 635208 298846 635308
rect 297850 634984 297950 635084
rect 298074 634984 298174 635084
rect 298298 634984 298398 635084
rect 298522 634984 298622 635084
rect 298746 634984 298846 635084
rect 297850 634760 297950 634860
rect 298074 634760 298174 634860
rect 298298 634760 298398 634860
rect 298522 634760 298622 634860
rect 298746 634760 298846 634860
rect 297850 634536 297950 634636
rect 298074 634536 298174 634636
rect 298298 634536 298398 634636
rect 298522 634536 298622 634636
rect 298746 634536 298846 634636
rect 297850 634312 297950 634412
rect 298074 634312 298174 634412
rect 298298 634312 298398 634412
rect 298522 634312 298622 634412
rect 298746 634312 298846 634412
rect 297850 634088 297950 634188
rect 298074 634088 298174 634188
rect 298298 634088 298398 634188
rect 298522 634088 298622 634188
rect 298746 634088 298846 634188
rect 297850 633864 297950 633964
rect 298074 633864 298174 633964
rect 298298 633864 298398 633964
rect 298522 633864 298622 633964
rect 298746 633864 298846 633964
rect 297850 633640 297950 633740
rect 298074 633640 298174 633740
rect 298298 633640 298398 633740
rect 298522 633640 298622 633740
rect 298746 633640 298846 633740
rect 297850 633416 297950 633516
rect 298074 633416 298174 633516
rect 298298 633416 298398 633516
rect 298522 633416 298622 633516
rect 298746 633416 298846 633516
rect 297850 633192 297950 633292
rect 298074 633192 298174 633292
rect 298298 633192 298398 633292
rect 298522 633192 298622 633292
rect 298746 633192 298846 633292
rect 297850 632968 297950 633068
rect 298074 632968 298174 633068
rect 298298 632968 298398 633068
rect 298522 632968 298622 633068
rect 298746 632968 298846 633068
rect 297850 632744 297950 632844
rect 298074 632744 298174 632844
rect 298298 632744 298398 632844
rect 298522 632744 298622 632844
rect 298746 632744 298846 632844
rect 297850 632520 297950 632620
rect 298074 632520 298174 632620
rect 298298 632520 298398 632620
rect 298522 632520 298622 632620
rect 298746 632520 298846 632620
rect 297850 632296 297950 632396
rect 298074 632296 298174 632396
rect 298298 632296 298398 632396
rect 298522 632296 298622 632396
rect 298746 632296 298846 632396
rect 297850 632072 297950 632172
rect 298074 632072 298174 632172
rect 298298 632072 298398 632172
rect 298522 632072 298622 632172
rect 298746 632072 298846 632172
rect 297850 631848 297950 631948
rect 298074 631848 298174 631948
rect 298298 631848 298398 631948
rect 298522 631848 298622 631948
rect 298746 631848 298846 631948
rect 297850 631624 297950 631724
rect 298074 631624 298174 631724
rect 298298 631624 298398 631724
rect 298522 631624 298622 631724
rect 298746 631624 298846 631724
rect 297850 631400 297950 631500
rect 298074 631400 298174 631500
rect 298298 631400 298398 631500
rect 298522 631400 298622 631500
rect 298746 631400 298846 631500
rect 342130 637896 342230 637996
rect 342354 637896 342454 637996
rect 342578 637896 342678 637996
rect 342802 637896 342902 637996
rect 343026 637896 343126 637996
rect 342130 637672 342230 637772
rect 342354 637672 342454 637772
rect 342578 637672 342678 637772
rect 342802 637672 342902 637772
rect 343026 637672 343126 637772
rect 342130 637448 342230 637548
rect 342354 637448 342454 637548
rect 342578 637448 342678 637548
rect 342802 637448 342902 637548
rect 343026 637448 343126 637548
rect 342130 637224 342230 637324
rect 342354 637224 342454 637324
rect 342578 637224 342678 637324
rect 342802 637224 342902 637324
rect 343026 637224 343126 637324
rect 342130 637000 342230 637100
rect 342354 637000 342454 637100
rect 342578 637000 342678 637100
rect 342802 637000 342902 637100
rect 343026 637000 343126 637100
rect 342130 636776 342230 636876
rect 342354 636776 342454 636876
rect 342578 636776 342678 636876
rect 342802 636776 342902 636876
rect 343026 636776 343126 636876
rect 342130 636552 342230 636652
rect 342354 636552 342454 636652
rect 342578 636552 342678 636652
rect 342802 636552 342902 636652
rect 343026 636552 343126 636652
rect 342130 636328 342230 636428
rect 342354 636328 342454 636428
rect 342578 636328 342678 636428
rect 342802 636328 342902 636428
rect 343026 636328 343126 636428
rect 342130 636104 342230 636204
rect 342354 636104 342454 636204
rect 342578 636104 342678 636204
rect 342802 636104 342902 636204
rect 343026 636104 343126 636204
rect 342130 635880 342230 635980
rect 342354 635880 342454 635980
rect 342578 635880 342678 635980
rect 342802 635880 342902 635980
rect 343026 635880 343126 635980
rect 342130 635656 342230 635756
rect 342354 635656 342454 635756
rect 342578 635656 342678 635756
rect 342802 635656 342902 635756
rect 343026 635656 343126 635756
rect 342130 635432 342230 635532
rect 342354 635432 342454 635532
rect 342578 635432 342678 635532
rect 342802 635432 342902 635532
rect 343026 635432 343126 635532
rect 342130 635208 342230 635308
rect 342354 635208 342454 635308
rect 342578 635208 342678 635308
rect 342802 635208 342902 635308
rect 343026 635208 343126 635308
rect 342130 634984 342230 635084
rect 342354 634984 342454 635084
rect 342578 634984 342678 635084
rect 342802 634984 342902 635084
rect 343026 634984 343126 635084
rect 342130 634760 342230 634860
rect 342354 634760 342454 634860
rect 342578 634760 342678 634860
rect 342802 634760 342902 634860
rect 343026 634760 343126 634860
rect 342130 634536 342230 634636
rect 342354 634536 342454 634636
rect 342578 634536 342678 634636
rect 342802 634536 342902 634636
rect 343026 634536 343126 634636
rect 342130 634312 342230 634412
rect 342354 634312 342454 634412
rect 342578 634312 342678 634412
rect 342802 634312 342902 634412
rect 343026 634312 343126 634412
rect 342130 634088 342230 634188
rect 342354 634088 342454 634188
rect 342578 634088 342678 634188
rect 342802 634088 342902 634188
rect 343026 634088 343126 634188
rect 342130 633864 342230 633964
rect 342354 633864 342454 633964
rect 342578 633864 342678 633964
rect 342802 633864 342902 633964
rect 343026 633864 343126 633964
rect 342130 633640 342230 633740
rect 342354 633640 342454 633740
rect 342578 633640 342678 633740
rect 342802 633640 342902 633740
rect 343026 633640 343126 633740
rect 342130 633416 342230 633516
rect 342354 633416 342454 633516
rect 342578 633416 342678 633516
rect 342802 633416 342902 633516
rect 343026 633416 343126 633516
rect 342130 633192 342230 633292
rect 342354 633192 342454 633292
rect 342578 633192 342678 633292
rect 342802 633192 342902 633292
rect 343026 633192 343126 633292
rect 342130 632968 342230 633068
rect 342354 632968 342454 633068
rect 342578 632968 342678 633068
rect 342802 632968 342902 633068
rect 343026 632968 343126 633068
rect 342130 632744 342230 632844
rect 342354 632744 342454 632844
rect 342578 632744 342678 632844
rect 342802 632744 342902 632844
rect 343026 632744 343126 632844
rect 342130 632520 342230 632620
rect 342354 632520 342454 632620
rect 342578 632520 342678 632620
rect 342802 632520 342902 632620
rect 343026 632520 343126 632620
rect 342130 632296 342230 632396
rect 342354 632296 342454 632396
rect 342578 632296 342678 632396
rect 342802 632296 342902 632396
rect 343026 632296 343126 632396
rect 342130 632072 342230 632172
rect 342354 632072 342454 632172
rect 342578 632072 342678 632172
rect 342802 632072 342902 632172
rect 343026 632072 343126 632172
rect 342130 631848 342230 631948
rect 342354 631848 342454 631948
rect 342578 631848 342678 631948
rect 342802 631848 342902 631948
rect 343026 631848 343126 631948
rect 342130 631624 342230 631724
rect 342354 631624 342454 631724
rect 342578 631624 342678 631724
rect 342802 631624 342902 631724
rect 343026 631624 343126 631724
rect 342130 631400 342230 631500
rect 342354 631400 342454 631500
rect 342578 631400 342678 631500
rect 342802 631400 342902 631500
rect 343026 631400 343126 631500
rect 319400 628668 319600 628868
rect 319834 628668 320034 628868
rect 320268 628668 320468 628868
rect 320702 628668 320902 628868
rect 321136 628668 321336 628868
rect 321570 628668 321770 628868
rect 322004 628668 322204 628868
rect 322438 628668 322638 628868
rect 322872 628668 323072 628868
rect 323306 628668 323506 628868
rect 323740 628668 323940 628868
rect 324140 628668 324340 628868
rect 324540 628668 324740 628868
rect 324940 628668 325140 628868
rect 325340 628668 325540 628868
rect 325740 628668 325940 628868
rect 326140 628668 326340 628868
rect 326540 628668 326740 628868
rect 326940 628668 327140 628868
rect 327340 628668 327540 628868
rect 328940 628668 329140 628868
rect 329340 628668 329540 628868
rect 329740 628668 329940 628868
rect 330140 628668 330340 628868
rect 330540 628668 330740 628868
rect 330940 628668 331140 628868
rect 331340 628668 331540 628868
rect 331740 628668 331940 628868
rect 332140 628668 332340 628868
rect 319400 628234 319600 628434
rect 319834 628234 320034 628434
rect 320268 628234 320468 628434
rect 320702 628234 320902 628434
rect 321136 628234 321336 628434
rect 321570 628234 321770 628434
rect 322004 628234 322204 628434
rect 322438 628234 322638 628434
rect 322872 628234 323072 628434
rect 323306 628234 323506 628434
rect 323740 628234 323940 628434
rect 319400 627800 319600 628000
rect 319834 627800 320034 628000
rect 320268 627800 320468 628000
rect 320702 627800 320902 628000
rect 321136 627800 321336 628000
rect 321570 627800 321770 628000
rect 322004 627800 322204 628000
rect 322438 627800 322638 628000
rect 322872 627800 323072 628000
rect 323306 627800 323506 628000
rect 323740 627800 323940 628000
rect 302980 625970 303040 626030
rect 303100 625970 303160 626030
rect 303220 625970 303280 626030
rect 303340 625970 303400 626030
rect 303460 625970 303520 626030
rect 302980 625850 303040 625910
rect 303100 625850 303160 625910
rect 303220 625850 303280 625910
rect 303340 625850 303400 625910
rect 303460 625850 303520 625910
rect 297850 624496 297950 624596
rect 298074 624496 298174 624596
rect 298298 624496 298398 624596
rect 298522 624496 298622 624596
rect 298746 624496 298846 624596
rect 297850 624272 297950 624372
rect 298074 624272 298174 624372
rect 298298 624272 298398 624372
rect 298522 624272 298622 624372
rect 298746 624272 298846 624372
rect 297850 624048 297950 624148
rect 298074 624048 298174 624148
rect 298298 624048 298398 624148
rect 298522 624048 298622 624148
rect 298746 624048 298846 624148
rect 342130 624496 342230 624596
rect 342354 624496 342454 624596
rect 342578 624496 342678 624596
rect 342802 624496 342902 624596
rect 343026 624496 343126 624596
rect 342130 624272 342230 624372
rect 342354 624272 342454 624372
rect 342578 624272 342678 624372
rect 342802 624272 342902 624372
rect 343026 624272 343126 624372
rect 342130 624048 342230 624148
rect 342354 624048 342454 624148
rect 342578 624048 342678 624148
rect 342802 624048 342902 624148
rect 343026 624048 343126 624148
rect 297850 623824 297950 623924
rect 298074 623824 298174 623924
rect 298298 623824 298398 623924
rect 298522 623824 298622 623924
rect 298746 623824 298846 623924
rect 297850 623600 297950 623700
rect 298074 623600 298174 623700
rect 298298 623600 298398 623700
rect 298522 623600 298622 623700
rect 298746 623600 298846 623700
rect 297850 623376 297950 623476
rect 298074 623376 298174 623476
rect 298298 623376 298398 623476
rect 298522 623376 298622 623476
rect 298746 623376 298846 623476
rect 297850 623152 297950 623252
rect 298074 623152 298174 623252
rect 298298 623152 298398 623252
rect 298522 623152 298622 623252
rect 298746 623152 298846 623252
rect 297850 622928 297950 623028
rect 298074 622928 298174 623028
rect 298298 622928 298398 623028
rect 298522 622928 298622 623028
rect 298746 622928 298846 623028
rect 297850 622704 297950 622804
rect 298074 622704 298174 622804
rect 298298 622704 298398 622804
rect 298522 622704 298622 622804
rect 298746 622704 298846 622804
rect 297850 622480 297950 622580
rect 298074 622480 298174 622580
rect 298298 622480 298398 622580
rect 298522 622480 298622 622580
rect 298746 622480 298846 622580
rect 297850 622256 297950 622356
rect 298074 622256 298174 622356
rect 298298 622256 298398 622356
rect 298522 622256 298622 622356
rect 298746 622256 298846 622356
rect 297850 622032 297950 622132
rect 298074 622032 298174 622132
rect 298298 622032 298398 622132
rect 298522 622032 298622 622132
rect 298746 622032 298846 622132
rect 297850 621808 297950 621908
rect 298074 621808 298174 621908
rect 298298 621808 298398 621908
rect 298522 621808 298622 621908
rect 298746 621808 298846 621908
rect 297850 621584 297950 621684
rect 298074 621584 298174 621684
rect 298298 621584 298398 621684
rect 298522 621584 298622 621684
rect 298746 621584 298846 621684
rect 297850 621360 297950 621460
rect 298074 621360 298174 621460
rect 298298 621360 298398 621460
rect 298522 621360 298622 621460
rect 298746 621360 298846 621460
rect 297850 621136 297950 621236
rect 298074 621136 298174 621236
rect 298298 621136 298398 621236
rect 298522 621136 298622 621236
rect 298746 621136 298846 621236
rect 297850 620912 297950 621012
rect 298074 620912 298174 621012
rect 298298 620912 298398 621012
rect 298522 620912 298622 621012
rect 298746 620912 298846 621012
rect 297850 620688 297950 620788
rect 298074 620688 298174 620788
rect 298298 620688 298398 620788
rect 298522 620688 298622 620788
rect 298746 620688 298846 620788
rect 297850 620464 297950 620564
rect 298074 620464 298174 620564
rect 298298 620464 298398 620564
rect 298522 620464 298622 620564
rect 298746 620464 298846 620564
rect 297850 620240 297950 620340
rect 298074 620240 298174 620340
rect 298298 620240 298398 620340
rect 298522 620240 298622 620340
rect 298746 620240 298846 620340
rect 297850 620016 297950 620116
rect 298074 620016 298174 620116
rect 298298 620016 298398 620116
rect 298522 620016 298622 620116
rect 298746 620016 298846 620116
rect 297850 619792 297950 619892
rect 298074 619792 298174 619892
rect 298298 619792 298398 619892
rect 298522 619792 298622 619892
rect 298746 619792 298846 619892
rect 297850 619568 297950 619668
rect 298074 619568 298174 619668
rect 298298 619568 298398 619668
rect 298522 619568 298622 619668
rect 298746 619568 298846 619668
rect 297850 619344 297950 619444
rect 298074 619344 298174 619444
rect 298298 619344 298398 619444
rect 298522 619344 298622 619444
rect 298746 619344 298846 619444
rect 297850 619120 297950 619220
rect 298074 619120 298174 619220
rect 298298 619120 298398 619220
rect 298522 619120 298622 619220
rect 298746 619120 298846 619220
rect 297850 618896 297950 618996
rect 298074 618896 298174 618996
rect 298298 618896 298398 618996
rect 298522 618896 298622 618996
rect 298746 618896 298846 618996
rect 297850 618672 297950 618772
rect 298074 618672 298174 618772
rect 298298 618672 298398 618772
rect 298522 618672 298622 618772
rect 298746 618672 298846 618772
rect 297850 618448 297950 618548
rect 298074 618448 298174 618548
rect 298298 618448 298398 618548
rect 298522 618448 298622 618548
rect 298746 618448 298846 618548
rect 297850 618224 297950 618324
rect 298074 618224 298174 618324
rect 298298 618224 298398 618324
rect 298522 618224 298622 618324
rect 298746 618224 298846 618324
rect 297850 618000 297950 618100
rect 298074 618000 298174 618100
rect 298298 618000 298398 618100
rect 298522 618000 298622 618100
rect 298746 618000 298846 618100
rect 342130 623824 342230 623924
rect 342354 623824 342454 623924
rect 342578 623824 342678 623924
rect 342802 623824 342902 623924
rect 343026 623824 343126 623924
rect 342130 623600 342230 623700
rect 342354 623600 342454 623700
rect 342578 623600 342678 623700
rect 342802 623600 342902 623700
rect 343026 623600 343126 623700
rect 342130 623376 342230 623476
rect 342354 623376 342454 623476
rect 342578 623376 342678 623476
rect 342802 623376 342902 623476
rect 343026 623376 343126 623476
rect 342130 623152 342230 623252
rect 342354 623152 342454 623252
rect 342578 623152 342678 623252
rect 342802 623152 342902 623252
rect 343026 623152 343126 623252
rect 342130 622928 342230 623028
rect 342354 622928 342454 623028
rect 342578 622928 342678 623028
rect 342802 622928 342902 623028
rect 343026 622928 343126 623028
rect 342130 622704 342230 622804
rect 342354 622704 342454 622804
rect 342578 622704 342678 622804
rect 342802 622704 342902 622804
rect 343026 622704 343126 622804
rect 342130 622480 342230 622580
rect 342354 622480 342454 622580
rect 342578 622480 342678 622580
rect 342802 622480 342902 622580
rect 343026 622480 343126 622580
rect 342130 622256 342230 622356
rect 342354 622256 342454 622356
rect 342578 622256 342678 622356
rect 342802 622256 342902 622356
rect 343026 622256 343126 622356
rect 342130 622032 342230 622132
rect 342354 622032 342454 622132
rect 342578 622032 342678 622132
rect 342802 622032 342902 622132
rect 343026 622032 343126 622132
rect 342130 621808 342230 621908
rect 342354 621808 342454 621908
rect 342578 621808 342678 621908
rect 342802 621808 342902 621908
rect 343026 621808 343126 621908
rect 342130 621584 342230 621684
rect 342354 621584 342454 621684
rect 342578 621584 342678 621684
rect 342802 621584 342902 621684
rect 343026 621584 343126 621684
rect 342130 621360 342230 621460
rect 342354 621360 342454 621460
rect 342578 621360 342678 621460
rect 342802 621360 342902 621460
rect 343026 621360 343126 621460
rect 342130 621136 342230 621236
rect 342354 621136 342454 621236
rect 342578 621136 342678 621236
rect 342802 621136 342902 621236
rect 343026 621136 343126 621236
rect 342130 620912 342230 621012
rect 342354 620912 342454 621012
rect 342578 620912 342678 621012
rect 342802 620912 342902 621012
rect 343026 620912 343126 621012
rect 342130 620688 342230 620788
rect 342354 620688 342454 620788
rect 342578 620688 342678 620788
rect 342802 620688 342902 620788
rect 343026 620688 343126 620788
rect 342130 620464 342230 620564
rect 342354 620464 342454 620564
rect 342578 620464 342678 620564
rect 342802 620464 342902 620564
rect 343026 620464 343126 620564
rect 342130 620240 342230 620340
rect 342354 620240 342454 620340
rect 342578 620240 342678 620340
rect 342802 620240 342902 620340
rect 343026 620240 343126 620340
rect 342130 620016 342230 620116
rect 342354 620016 342454 620116
rect 342578 620016 342678 620116
rect 342802 620016 342902 620116
rect 343026 620016 343126 620116
rect 342130 619792 342230 619892
rect 342354 619792 342454 619892
rect 342578 619792 342678 619892
rect 342802 619792 342902 619892
rect 343026 619792 343126 619892
rect 342130 619568 342230 619668
rect 342354 619568 342454 619668
rect 342578 619568 342678 619668
rect 342802 619568 342902 619668
rect 343026 619568 343126 619668
rect 342130 619344 342230 619444
rect 342354 619344 342454 619444
rect 342578 619344 342678 619444
rect 342802 619344 342902 619444
rect 343026 619344 343126 619444
rect 342130 619120 342230 619220
rect 342354 619120 342454 619220
rect 342578 619120 342678 619220
rect 342802 619120 342902 619220
rect 343026 619120 343126 619220
rect 342130 618896 342230 618996
rect 342354 618896 342454 618996
rect 342578 618896 342678 618996
rect 342802 618896 342902 618996
rect 343026 618896 343126 618996
rect 342130 618672 342230 618772
rect 342354 618672 342454 618772
rect 342578 618672 342678 618772
rect 342802 618672 342902 618772
rect 343026 618672 343126 618772
rect 342130 618448 342230 618548
rect 342354 618448 342454 618548
rect 342578 618448 342678 618548
rect 342802 618448 342902 618548
rect 343026 618448 343126 618548
rect 342130 618224 342230 618324
rect 342354 618224 342454 618324
rect 342578 618224 342678 618324
rect 342802 618224 342902 618324
rect 343026 618224 343126 618324
rect 342130 618000 342230 618100
rect 342354 618000 342454 618100
rect 342578 618000 342678 618100
rect 342802 618000 342902 618100
rect 343026 618000 343126 618100
rect 298876 615374 298976 615474
rect 299100 615374 299200 615474
rect 299324 615374 299424 615474
rect 299548 615374 299648 615474
rect 299772 615374 299872 615474
rect 299996 615374 300096 615474
rect 300220 615374 300320 615474
rect 300444 615374 300544 615474
rect 300668 615374 300768 615474
rect 300892 615374 300992 615474
rect 301116 615374 301216 615474
rect 301340 615374 301440 615474
rect 301564 615374 301664 615474
rect 301788 615374 301888 615474
rect 302012 615374 302112 615474
rect 302236 615374 302336 615474
rect 302460 615374 302560 615474
rect 302684 615374 302784 615474
rect 302908 615374 303008 615474
rect 303132 615374 303232 615474
rect 303356 615374 303456 615474
rect 303580 615374 303680 615474
rect 303804 615374 303904 615474
rect 304028 615374 304128 615474
rect 304252 615374 304352 615474
rect 304476 615374 304576 615474
rect 304700 615374 304800 615474
rect 304924 615374 305024 615474
rect 305148 615374 305248 615474
rect 305372 615374 305472 615474
rect 298876 615150 298976 615250
rect 299100 615150 299200 615250
rect 299324 615150 299424 615250
rect 299548 615150 299648 615250
rect 299772 615150 299872 615250
rect 299996 615150 300096 615250
rect 300220 615150 300320 615250
rect 300444 615150 300544 615250
rect 300668 615150 300768 615250
rect 300892 615150 300992 615250
rect 301116 615150 301216 615250
rect 301340 615150 301440 615250
rect 301564 615150 301664 615250
rect 301788 615150 301888 615250
rect 302012 615150 302112 615250
rect 302236 615150 302336 615250
rect 302460 615150 302560 615250
rect 302684 615150 302784 615250
rect 302908 615150 303008 615250
rect 303132 615150 303232 615250
rect 303356 615150 303456 615250
rect 303580 615150 303680 615250
rect 303804 615150 303904 615250
rect 304028 615150 304128 615250
rect 304252 615150 304352 615250
rect 304476 615150 304576 615250
rect 304700 615150 304800 615250
rect 304924 615150 305024 615250
rect 305148 615150 305248 615250
rect 305372 615150 305472 615250
rect 298876 614926 298976 615026
rect 299100 614926 299200 615026
rect 299324 614926 299424 615026
rect 299548 614926 299648 615026
rect 299772 614926 299872 615026
rect 299996 614926 300096 615026
rect 300220 614926 300320 615026
rect 300444 614926 300544 615026
rect 300668 614926 300768 615026
rect 300892 614926 300992 615026
rect 301116 614926 301216 615026
rect 301340 614926 301440 615026
rect 301564 614926 301664 615026
rect 301788 614926 301888 615026
rect 302012 614926 302112 615026
rect 302236 614926 302336 615026
rect 302460 614926 302560 615026
rect 302684 614926 302784 615026
rect 302908 614926 303008 615026
rect 303132 614926 303232 615026
rect 303356 614926 303456 615026
rect 303580 614926 303680 615026
rect 303804 614926 303904 615026
rect 304028 614926 304128 615026
rect 304252 614926 304352 615026
rect 304476 614926 304576 615026
rect 304700 614926 304800 615026
rect 304924 614926 305024 615026
rect 305148 614926 305248 615026
rect 305372 614926 305472 615026
rect 298876 614702 298976 614802
rect 299100 614702 299200 614802
rect 299324 614702 299424 614802
rect 299548 614702 299648 614802
rect 299772 614702 299872 614802
rect 299996 614702 300096 614802
rect 300220 614702 300320 614802
rect 300444 614702 300544 614802
rect 300668 614702 300768 614802
rect 300892 614702 300992 614802
rect 301116 614702 301216 614802
rect 301340 614702 301440 614802
rect 301564 614702 301664 614802
rect 301788 614702 301888 614802
rect 302012 614702 302112 614802
rect 302236 614702 302336 614802
rect 302460 614702 302560 614802
rect 302684 614702 302784 614802
rect 302908 614702 303008 614802
rect 303132 614702 303232 614802
rect 303356 614702 303456 614802
rect 303580 614702 303680 614802
rect 303804 614702 303904 614802
rect 304028 614702 304128 614802
rect 304252 614702 304352 614802
rect 304476 614702 304576 614802
rect 304700 614702 304800 614802
rect 304924 614702 305024 614802
rect 305148 614702 305248 614802
rect 305372 614702 305472 614802
rect 298876 614478 298976 614578
rect 299100 614478 299200 614578
rect 299324 614478 299424 614578
rect 299548 614478 299648 614578
rect 299772 614478 299872 614578
rect 299996 614478 300096 614578
rect 300220 614478 300320 614578
rect 300444 614478 300544 614578
rect 300668 614478 300768 614578
rect 300892 614478 300992 614578
rect 301116 614478 301216 614578
rect 301340 614478 301440 614578
rect 301564 614478 301664 614578
rect 301788 614478 301888 614578
rect 302012 614478 302112 614578
rect 302236 614478 302336 614578
rect 302460 614478 302560 614578
rect 302684 614478 302784 614578
rect 302908 614478 303008 614578
rect 303132 614478 303232 614578
rect 303356 614478 303456 614578
rect 303580 614478 303680 614578
rect 303804 614478 303904 614578
rect 304028 614478 304128 614578
rect 304252 614478 304352 614578
rect 304476 614478 304576 614578
rect 304700 614478 304800 614578
rect 304924 614478 305024 614578
rect 305148 614478 305248 614578
rect 305372 614478 305472 614578
rect 309346 615374 309446 615474
rect 309570 615374 309670 615474
rect 309794 615374 309894 615474
rect 310018 615374 310118 615474
rect 310242 615374 310342 615474
rect 310466 615374 310566 615474
rect 310690 615374 310790 615474
rect 310914 615374 311014 615474
rect 311138 615374 311238 615474
rect 311362 615374 311462 615474
rect 311586 615374 311686 615474
rect 311810 615374 311910 615474
rect 312034 615374 312134 615474
rect 312258 615374 312358 615474
rect 312482 615374 312582 615474
rect 312706 615374 312806 615474
rect 312930 615374 313030 615474
rect 313154 615374 313254 615474
rect 313378 615374 313478 615474
rect 313602 615374 313702 615474
rect 313826 615374 313926 615474
rect 314050 615374 314150 615474
rect 314274 615374 314374 615474
rect 314498 615374 314598 615474
rect 314722 615374 314822 615474
rect 314946 615374 315046 615474
rect 315170 615374 315270 615474
rect 315394 615374 315494 615474
rect 315618 615374 315718 615474
rect 315842 615374 315942 615474
rect 309346 615150 309446 615250
rect 309570 615150 309670 615250
rect 309794 615150 309894 615250
rect 310018 615150 310118 615250
rect 310242 615150 310342 615250
rect 310466 615150 310566 615250
rect 310690 615150 310790 615250
rect 310914 615150 311014 615250
rect 311138 615150 311238 615250
rect 311362 615150 311462 615250
rect 311586 615150 311686 615250
rect 311810 615150 311910 615250
rect 312034 615150 312134 615250
rect 312258 615150 312358 615250
rect 312482 615150 312582 615250
rect 312706 615150 312806 615250
rect 312930 615150 313030 615250
rect 313154 615150 313254 615250
rect 313378 615150 313478 615250
rect 313602 615150 313702 615250
rect 313826 615150 313926 615250
rect 314050 615150 314150 615250
rect 314274 615150 314374 615250
rect 314498 615150 314598 615250
rect 314722 615150 314822 615250
rect 314946 615150 315046 615250
rect 315170 615150 315270 615250
rect 315394 615150 315494 615250
rect 315618 615150 315718 615250
rect 315842 615150 315942 615250
rect 309346 614926 309446 615026
rect 309570 614926 309670 615026
rect 309794 614926 309894 615026
rect 310018 614926 310118 615026
rect 310242 614926 310342 615026
rect 310466 614926 310566 615026
rect 310690 614926 310790 615026
rect 310914 614926 311014 615026
rect 311138 614926 311238 615026
rect 311362 614926 311462 615026
rect 311586 614926 311686 615026
rect 311810 614926 311910 615026
rect 312034 614926 312134 615026
rect 312258 614926 312358 615026
rect 312482 614926 312582 615026
rect 312706 614926 312806 615026
rect 312930 614926 313030 615026
rect 313154 614926 313254 615026
rect 313378 614926 313478 615026
rect 313602 614926 313702 615026
rect 313826 614926 313926 615026
rect 314050 614926 314150 615026
rect 314274 614926 314374 615026
rect 314498 614926 314598 615026
rect 314722 614926 314822 615026
rect 314946 614926 315046 615026
rect 315170 614926 315270 615026
rect 315394 614926 315494 615026
rect 315618 614926 315718 615026
rect 315842 614926 315942 615026
rect 309346 614702 309446 614802
rect 309570 614702 309670 614802
rect 309794 614702 309894 614802
rect 310018 614702 310118 614802
rect 310242 614702 310342 614802
rect 310466 614702 310566 614802
rect 310690 614702 310790 614802
rect 310914 614702 311014 614802
rect 311138 614702 311238 614802
rect 311362 614702 311462 614802
rect 311586 614702 311686 614802
rect 311810 614702 311910 614802
rect 312034 614702 312134 614802
rect 312258 614702 312358 614802
rect 312482 614702 312582 614802
rect 312706 614702 312806 614802
rect 312930 614702 313030 614802
rect 313154 614702 313254 614802
rect 313378 614702 313478 614802
rect 313602 614702 313702 614802
rect 313826 614702 313926 614802
rect 314050 614702 314150 614802
rect 314274 614702 314374 614802
rect 314498 614702 314598 614802
rect 314722 614702 314822 614802
rect 314946 614702 315046 614802
rect 315170 614702 315270 614802
rect 315394 614702 315494 614802
rect 315618 614702 315718 614802
rect 315842 614702 315942 614802
rect 309346 614478 309446 614578
rect 309570 614478 309670 614578
rect 309794 614478 309894 614578
rect 310018 614478 310118 614578
rect 310242 614478 310342 614578
rect 310466 614478 310566 614578
rect 310690 614478 310790 614578
rect 310914 614478 311014 614578
rect 311138 614478 311238 614578
rect 311362 614478 311462 614578
rect 311586 614478 311686 614578
rect 311810 614478 311910 614578
rect 312034 614478 312134 614578
rect 312258 614478 312358 614578
rect 312482 614478 312582 614578
rect 312706 614478 312806 614578
rect 312930 614478 313030 614578
rect 313154 614478 313254 614578
rect 313378 614478 313478 614578
rect 313602 614478 313702 614578
rect 313826 614478 313926 614578
rect 314050 614478 314150 614578
rect 314274 614478 314374 614578
rect 314498 614478 314598 614578
rect 314722 614478 314822 614578
rect 314946 614478 315046 614578
rect 315170 614478 315270 614578
rect 315394 614478 315494 614578
rect 315618 614478 315718 614578
rect 315842 614478 315942 614578
rect 335616 615394 335716 615494
rect 335840 615394 335940 615494
rect 336064 615394 336164 615494
rect 336288 615394 336388 615494
rect 336512 615394 336612 615494
rect 336736 615394 336836 615494
rect 336960 615394 337060 615494
rect 337184 615394 337284 615494
rect 337408 615394 337508 615494
rect 337632 615394 337732 615494
rect 337856 615394 337956 615494
rect 338080 615394 338180 615494
rect 338304 615394 338404 615494
rect 338528 615394 338628 615494
rect 338752 615394 338852 615494
rect 338976 615394 339076 615494
rect 339200 615394 339300 615494
rect 339424 615394 339524 615494
rect 339648 615394 339748 615494
rect 339872 615394 339972 615494
rect 340096 615394 340196 615494
rect 340320 615394 340420 615494
rect 340544 615394 340644 615494
rect 340768 615394 340868 615494
rect 340992 615394 341092 615494
rect 341216 615394 341316 615494
rect 341440 615394 341540 615494
rect 341664 615394 341764 615494
rect 341888 615394 341988 615494
rect 342112 615394 342212 615494
rect 335616 615170 335716 615270
rect 335840 615170 335940 615270
rect 336064 615170 336164 615270
rect 336288 615170 336388 615270
rect 336512 615170 336612 615270
rect 336736 615170 336836 615270
rect 336960 615170 337060 615270
rect 337184 615170 337284 615270
rect 337408 615170 337508 615270
rect 337632 615170 337732 615270
rect 337856 615170 337956 615270
rect 338080 615170 338180 615270
rect 338304 615170 338404 615270
rect 338528 615170 338628 615270
rect 338752 615170 338852 615270
rect 338976 615170 339076 615270
rect 339200 615170 339300 615270
rect 339424 615170 339524 615270
rect 339648 615170 339748 615270
rect 339872 615170 339972 615270
rect 340096 615170 340196 615270
rect 340320 615170 340420 615270
rect 340544 615170 340644 615270
rect 340768 615170 340868 615270
rect 340992 615170 341092 615270
rect 341216 615170 341316 615270
rect 341440 615170 341540 615270
rect 341664 615170 341764 615270
rect 341888 615170 341988 615270
rect 342112 615170 342212 615270
rect 335616 614946 335716 615046
rect 335840 614946 335940 615046
rect 336064 614946 336164 615046
rect 336288 614946 336388 615046
rect 336512 614946 336612 615046
rect 336736 614946 336836 615046
rect 336960 614946 337060 615046
rect 337184 614946 337284 615046
rect 337408 614946 337508 615046
rect 337632 614946 337732 615046
rect 337856 614946 337956 615046
rect 338080 614946 338180 615046
rect 338304 614946 338404 615046
rect 338528 614946 338628 615046
rect 338752 614946 338852 615046
rect 338976 614946 339076 615046
rect 339200 614946 339300 615046
rect 339424 614946 339524 615046
rect 339648 614946 339748 615046
rect 339872 614946 339972 615046
rect 340096 614946 340196 615046
rect 340320 614946 340420 615046
rect 340544 614946 340644 615046
rect 340768 614946 340868 615046
rect 340992 614946 341092 615046
rect 341216 614946 341316 615046
rect 341440 614946 341540 615046
rect 341664 614946 341764 615046
rect 341888 614946 341988 615046
rect 342112 614946 342212 615046
rect 335616 614722 335716 614822
rect 335840 614722 335940 614822
rect 336064 614722 336164 614822
rect 336288 614722 336388 614822
rect 336512 614722 336612 614822
rect 336736 614722 336836 614822
rect 336960 614722 337060 614822
rect 337184 614722 337284 614822
rect 337408 614722 337508 614822
rect 337632 614722 337732 614822
rect 337856 614722 337956 614822
rect 338080 614722 338180 614822
rect 338304 614722 338404 614822
rect 338528 614722 338628 614822
rect 338752 614722 338852 614822
rect 338976 614722 339076 614822
rect 339200 614722 339300 614822
rect 339424 614722 339524 614822
rect 339648 614722 339748 614822
rect 339872 614722 339972 614822
rect 340096 614722 340196 614822
rect 340320 614722 340420 614822
rect 340544 614722 340644 614822
rect 340768 614722 340868 614822
rect 340992 614722 341092 614822
rect 341216 614722 341316 614822
rect 341440 614722 341540 614822
rect 341664 614722 341764 614822
rect 341888 614722 341988 614822
rect 342112 614722 342212 614822
rect 335616 614498 335716 614598
rect 335840 614498 335940 614598
rect 336064 614498 336164 614598
rect 336288 614498 336388 614598
rect 336512 614498 336612 614598
rect 336736 614498 336836 614598
rect 336960 614498 337060 614598
rect 337184 614498 337284 614598
rect 337408 614498 337508 614598
rect 337632 614498 337732 614598
rect 337856 614498 337956 614598
rect 338080 614498 338180 614598
rect 338304 614498 338404 614598
rect 338528 614498 338628 614598
rect 338752 614498 338852 614598
rect 338976 614498 339076 614598
rect 339200 614498 339300 614598
rect 339424 614498 339524 614598
rect 339648 614498 339748 614598
rect 339872 614498 339972 614598
rect 340096 614498 340196 614598
rect 340320 614498 340420 614598
rect 340544 614498 340644 614598
rect 340768 614498 340868 614598
rect 340992 614498 341092 614598
rect 341216 614498 341316 614598
rect 341440 614498 341540 614598
rect 341664 614498 341764 614598
rect 341888 614498 341988 614598
rect 342112 614498 342212 614598
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 690577 173094 704800
rect -800 680242 1700 685242
rect 170894 684353 170922 690577
rect 173066 684353 173094 690577
rect 170894 683764 173094 684353
rect 173394 690577 175594 704800
rect 175894 702300 180894 704800
rect 173394 684353 173422 690577
rect 175566 684353 175594 690577
rect 173394 683764 175594 684353
rect -800 643842 1660 648642
rect -800 633842 1660 638642
rect 217294 626176 222294 704800
rect 222594 690610 224794 704800
rect 222594 684386 222622 690610
rect 224766 684386 224794 690610
rect 222594 683913 224794 684386
rect 225094 694292 227294 704800
rect 227594 694292 232594 704800
rect 225094 692092 232594 694292
rect 225094 683913 227294 692092
rect 217294 626112 217344 626176
rect 217408 626112 217472 626176
rect 217536 626112 217600 626176
rect 217664 626112 217728 626176
rect 217792 626112 217856 626176
rect 217920 626112 217984 626176
rect 218048 626112 218112 626176
rect 218176 626112 218240 626176
rect 218304 626112 218368 626176
rect 218432 626112 218496 626176
rect 218560 626112 218624 626176
rect 218688 626112 218752 626176
rect 218816 626112 218880 626176
rect 218944 626112 219008 626176
rect 219072 626112 219136 626176
rect 219200 626112 219264 626176
rect 219328 626112 219392 626176
rect 219456 626112 219520 626176
rect 219584 626112 219648 626176
rect 219712 626112 219776 626176
rect 219840 626112 219904 626176
rect 219968 626112 220032 626176
rect 220096 626112 220160 626176
rect 220224 626112 220288 626176
rect 220352 626112 220416 626176
rect 220480 626112 220544 626176
rect 220608 626112 220672 626176
rect 220736 626112 220800 626176
rect 220864 626112 220928 626176
rect 220992 626112 221056 626176
rect 221120 626112 221184 626176
rect 221248 626112 221312 626176
rect 221376 626112 221440 626176
rect 221504 626112 221568 626176
rect 221632 626112 221696 626176
rect 221760 626112 221824 626176
rect 221888 626112 221952 626176
rect 222016 626112 222080 626176
rect 222144 626112 222294 626176
rect 217294 626048 222294 626112
rect 217294 625984 217344 626048
rect 217408 625984 217472 626048
rect 217536 625984 217600 626048
rect 217664 625984 217728 626048
rect 217792 625984 217856 626048
rect 217920 625984 217984 626048
rect 218048 625984 218112 626048
rect 218176 625984 218240 626048
rect 218304 625984 218368 626048
rect 218432 625984 218496 626048
rect 218560 625984 218624 626048
rect 218688 625984 218752 626048
rect 218816 625984 218880 626048
rect 218944 625984 219008 626048
rect 219072 625984 219136 626048
rect 219200 625984 219264 626048
rect 219328 625984 219392 626048
rect 219456 625984 219520 626048
rect 219584 625984 219648 626048
rect 219712 625984 219776 626048
rect 219840 625984 219904 626048
rect 219968 625984 220032 626048
rect 220096 625984 220160 626048
rect 220224 625984 220288 626048
rect 220352 625984 220416 626048
rect 220480 625984 220544 626048
rect 220608 625984 220672 626048
rect 220736 625984 220800 626048
rect 220864 625984 220928 626048
rect 220992 625984 221056 626048
rect 221120 625984 221184 626048
rect 221248 625984 221312 626048
rect 221376 625984 221440 626048
rect 221504 625984 221568 626048
rect 221632 625984 221696 626048
rect 221760 625984 221824 626048
rect 221888 625984 221952 626048
rect 222016 625984 222080 626048
rect 222144 625984 222294 626048
rect 217294 625920 222294 625984
rect 217294 625856 217344 625920
rect 217408 625856 217472 625920
rect 217536 625856 217600 625920
rect 217664 625856 217728 625920
rect 217792 625856 217856 625920
rect 217920 625856 217984 625920
rect 218048 625856 218112 625920
rect 218176 625856 218240 625920
rect 218304 625856 218368 625920
rect 218432 625856 218496 625920
rect 218560 625856 218624 625920
rect 218688 625856 218752 625920
rect 218816 625856 218880 625920
rect 218944 625856 219008 625920
rect 219072 625856 219136 625920
rect 219200 625856 219264 625920
rect 219328 625856 219392 625920
rect 219456 625856 219520 625920
rect 219584 625856 219648 625920
rect 219712 625856 219776 625920
rect 219840 625856 219904 625920
rect 219968 625856 220032 625920
rect 220096 625856 220160 625920
rect 220224 625856 220288 625920
rect 220352 625856 220416 625920
rect 220480 625856 220544 625920
rect 220608 625856 220672 625920
rect 220736 625856 220800 625920
rect 220864 625856 220928 625920
rect 220992 625856 221056 625920
rect 221120 625856 221184 625920
rect 221248 625856 221312 625920
rect 221376 625856 221440 625920
rect 221504 625856 221568 625920
rect 221632 625856 221696 625920
rect 221760 625856 221824 625920
rect 221888 625856 221952 625920
rect 222016 625856 222080 625920
rect 222144 625856 222294 625920
rect 217294 625792 222294 625856
rect 217294 625728 217344 625792
rect 217408 625728 217472 625792
rect 217536 625728 217600 625792
rect 217664 625728 217728 625792
rect 217792 625728 217856 625792
rect 217920 625728 217984 625792
rect 218048 625728 218112 625792
rect 218176 625728 218240 625792
rect 218304 625728 218368 625792
rect 218432 625728 218496 625792
rect 218560 625728 218624 625792
rect 218688 625728 218752 625792
rect 218816 625728 218880 625792
rect 218944 625728 219008 625792
rect 219072 625728 219136 625792
rect 219200 625728 219264 625792
rect 219328 625728 219392 625792
rect 219456 625728 219520 625792
rect 219584 625728 219648 625792
rect 219712 625728 219776 625792
rect 219840 625728 219904 625792
rect 219968 625728 220032 625792
rect 220096 625728 220160 625792
rect 220224 625728 220288 625792
rect 220352 625728 220416 625792
rect 220480 625728 220544 625792
rect 220608 625728 220672 625792
rect 220736 625728 220800 625792
rect 220864 625728 220928 625792
rect 220992 625728 221056 625792
rect 221120 625728 221184 625792
rect 221248 625728 221312 625792
rect 221376 625728 221440 625792
rect 221504 625728 221568 625792
rect 221632 625728 221696 625792
rect 221760 625728 221824 625792
rect 221888 625728 221952 625792
rect 222016 625728 222080 625792
rect 222144 625728 222294 625792
rect 217294 625700 222294 625728
rect 227594 626176 232594 692092
rect 227594 626112 227640 626176
rect 227704 626112 227768 626176
rect 227832 626112 227896 626176
rect 227960 626112 228024 626176
rect 228088 626112 228152 626176
rect 228216 626112 228280 626176
rect 228344 626112 228408 626176
rect 228472 626112 228536 626176
rect 228600 626112 228664 626176
rect 228728 626112 228792 626176
rect 228856 626112 228920 626176
rect 228984 626112 229048 626176
rect 229112 626112 229176 626176
rect 229240 626112 229304 626176
rect 229368 626112 229432 626176
rect 229496 626112 229560 626176
rect 229624 626112 229688 626176
rect 229752 626112 229816 626176
rect 229880 626112 229944 626176
rect 230008 626112 230072 626176
rect 230136 626112 230200 626176
rect 230264 626112 230328 626176
rect 230392 626112 230456 626176
rect 230520 626112 230584 626176
rect 230648 626112 230712 626176
rect 230776 626112 230840 626176
rect 230904 626112 230968 626176
rect 231032 626112 231096 626176
rect 231160 626112 231224 626176
rect 231288 626112 231352 626176
rect 231416 626112 231480 626176
rect 231544 626112 231608 626176
rect 231672 626112 231736 626176
rect 231800 626112 231864 626176
rect 231928 626112 231992 626176
rect 232056 626112 232120 626176
rect 232184 626112 232248 626176
rect 232312 626112 232376 626176
rect 232440 626112 232594 626176
rect 227594 626048 232594 626112
rect 227594 625984 227640 626048
rect 227704 625984 227768 626048
rect 227832 625984 227896 626048
rect 227960 625984 228024 626048
rect 228088 625984 228152 626048
rect 228216 625984 228280 626048
rect 228344 625984 228408 626048
rect 228472 625984 228536 626048
rect 228600 625984 228664 626048
rect 228728 625984 228792 626048
rect 228856 625984 228920 626048
rect 228984 625984 229048 626048
rect 229112 625984 229176 626048
rect 229240 625984 229304 626048
rect 229368 625984 229432 626048
rect 229496 625984 229560 626048
rect 229624 625984 229688 626048
rect 229752 625984 229816 626048
rect 229880 625984 229944 626048
rect 230008 625984 230072 626048
rect 230136 625984 230200 626048
rect 230264 625984 230328 626048
rect 230392 625984 230456 626048
rect 230520 625984 230584 626048
rect 230648 625984 230712 626048
rect 230776 625984 230840 626048
rect 230904 625984 230968 626048
rect 231032 625984 231096 626048
rect 231160 625984 231224 626048
rect 231288 625984 231352 626048
rect 231416 625984 231480 626048
rect 231544 625984 231608 626048
rect 231672 625984 231736 626048
rect 231800 625984 231864 626048
rect 231928 625984 231992 626048
rect 232056 625984 232120 626048
rect 232184 625984 232248 626048
rect 232312 625984 232376 626048
rect 232440 625984 232594 626048
rect 227594 625920 232594 625984
rect 227594 625856 227640 625920
rect 227704 625856 227768 625920
rect 227832 625856 227896 625920
rect 227960 625856 228024 625920
rect 228088 625856 228152 625920
rect 228216 625856 228280 625920
rect 228344 625856 228408 625920
rect 228472 625856 228536 625920
rect 228600 625856 228664 625920
rect 228728 625856 228792 625920
rect 228856 625856 228920 625920
rect 228984 625856 229048 625920
rect 229112 625856 229176 625920
rect 229240 625856 229304 625920
rect 229368 625856 229432 625920
rect 229496 625856 229560 625920
rect 229624 625856 229688 625920
rect 229752 625856 229816 625920
rect 229880 625856 229944 625920
rect 230008 625856 230072 625920
rect 230136 625856 230200 625920
rect 230264 625856 230328 625920
rect 230392 625856 230456 625920
rect 230520 625856 230584 625920
rect 230648 625856 230712 625920
rect 230776 625856 230840 625920
rect 230904 625856 230968 625920
rect 231032 625856 231096 625920
rect 231160 625856 231224 625920
rect 231288 625856 231352 625920
rect 231416 625856 231480 625920
rect 231544 625856 231608 625920
rect 231672 625856 231736 625920
rect 231800 625856 231864 625920
rect 231928 625856 231992 625920
rect 232056 625856 232120 625920
rect 232184 625856 232248 625920
rect 232312 625856 232376 625920
rect 232440 625856 232594 625920
rect 227594 625792 232594 625856
rect 227594 625728 227640 625792
rect 227704 625728 227768 625792
rect 227832 625728 227896 625792
rect 227960 625728 228024 625792
rect 228088 625728 228152 625792
rect 228216 625728 228280 625792
rect 228344 625728 228408 625792
rect 228472 625728 228536 625792
rect 228600 625728 228664 625792
rect 228728 625728 228792 625792
rect 228856 625728 228920 625792
rect 228984 625728 229048 625792
rect 229112 625728 229176 625792
rect 229240 625728 229304 625792
rect 229368 625728 229432 625792
rect 229496 625728 229560 625792
rect 229624 625728 229688 625792
rect 229752 625728 229816 625792
rect 229880 625728 229944 625792
rect 230008 625728 230072 625792
rect 230136 625728 230200 625792
rect 230264 625728 230328 625792
rect 230392 625728 230456 625792
rect 230520 625728 230584 625792
rect 230648 625728 230712 625792
rect 230776 625728 230840 625792
rect 230904 625728 230968 625792
rect 231032 625728 231096 625792
rect 231160 625728 231224 625792
rect 231288 625728 231352 625792
rect 231416 625728 231480 625792
rect 231544 625728 231608 625792
rect 231672 625728 231736 625792
rect 231800 625728 231864 625792
rect 231928 625728 231992 625792
rect 232056 625728 232120 625792
rect 232184 625728 232248 625792
rect 232312 625728 232376 625792
rect 232440 625728 232594 625792
rect 227594 625700 232594 625728
rect 288920 690084 295576 690584
rect 288920 684340 289800 690084
rect 294584 684340 295576 690084
rect 288920 650584 295576 684340
rect 318994 683600 323994 704800
rect 324294 690593 326494 704800
rect 326794 694292 328994 704800
rect 329294 694292 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 326794 692092 334294 694292
rect 324294 684369 324322 690593
rect 326466 684369 326494 690593
rect 324294 684038 326494 684369
rect 329294 683600 334294 692092
rect 510594 690560 515394 704800
rect 510594 684336 510602 690560
rect 515386 684336 515394 690560
rect 288920 644840 289920 650584
rect 294704 644840 295576 650584
rect 288920 637184 295576 644840
rect 298820 650584 315980 651400
rect 298820 644840 298920 650584
rect 303704 644840 304920 650584
rect 309704 644840 310920 650584
rect 315704 644840 315980 650584
rect 318994 650200 334400 683600
rect 510594 651406 515394 684336
rect 298820 642694 315980 644840
rect 298820 642594 298876 642694
rect 298976 642594 299100 642694
rect 299200 642594 299324 642694
rect 299424 642594 299548 642694
rect 299648 642594 299772 642694
rect 299872 642594 299996 642694
rect 300096 642594 300220 642694
rect 300320 642594 300444 642694
rect 300544 642594 300668 642694
rect 300768 642594 300892 642694
rect 300992 642594 301116 642694
rect 301216 642594 301340 642694
rect 301440 642594 301564 642694
rect 301664 642594 301788 642694
rect 301888 642594 302012 642694
rect 302112 642594 302236 642694
rect 302336 642594 302460 642694
rect 302560 642594 302684 642694
rect 302784 642594 302908 642694
rect 303008 642594 303132 642694
rect 303232 642594 303356 642694
rect 303456 642594 303580 642694
rect 303680 642594 303804 642694
rect 303904 642594 304028 642694
rect 304128 642594 304252 642694
rect 304352 642594 304476 642694
rect 304576 642594 304700 642694
rect 304800 642594 304924 642694
rect 305024 642594 305148 642694
rect 305248 642594 305372 642694
rect 305472 642594 309346 642694
rect 309446 642594 309570 642694
rect 309670 642594 309794 642694
rect 309894 642594 310018 642694
rect 310118 642594 310242 642694
rect 310342 642594 310466 642694
rect 310566 642594 310690 642694
rect 310790 642594 310914 642694
rect 311014 642594 311138 642694
rect 311238 642594 311362 642694
rect 311462 642594 311586 642694
rect 311686 642594 311810 642694
rect 311910 642594 312034 642694
rect 312134 642594 312258 642694
rect 312358 642594 312482 642694
rect 312582 642594 312706 642694
rect 312806 642594 312930 642694
rect 313030 642594 313154 642694
rect 313254 642594 313378 642694
rect 313478 642594 313602 642694
rect 313702 642594 313826 642694
rect 313926 642594 314050 642694
rect 314150 642594 314274 642694
rect 314374 642594 314498 642694
rect 314598 642594 314722 642694
rect 314822 642594 314946 642694
rect 315046 642594 315170 642694
rect 315270 642594 315394 642694
rect 315494 642594 315618 642694
rect 315718 642594 315842 642694
rect 315942 642594 315980 642694
rect 298820 642470 315980 642594
rect 298820 642370 298876 642470
rect 298976 642370 299100 642470
rect 299200 642370 299324 642470
rect 299424 642370 299548 642470
rect 299648 642370 299772 642470
rect 299872 642370 299996 642470
rect 300096 642370 300220 642470
rect 300320 642370 300444 642470
rect 300544 642370 300668 642470
rect 300768 642370 300892 642470
rect 300992 642370 301116 642470
rect 301216 642370 301340 642470
rect 301440 642370 301564 642470
rect 301664 642370 301788 642470
rect 301888 642370 302012 642470
rect 302112 642370 302236 642470
rect 302336 642370 302460 642470
rect 302560 642370 302684 642470
rect 302784 642370 302908 642470
rect 303008 642370 303132 642470
rect 303232 642370 303356 642470
rect 303456 642370 303580 642470
rect 303680 642370 303804 642470
rect 303904 642370 304028 642470
rect 304128 642370 304252 642470
rect 304352 642370 304476 642470
rect 304576 642370 304700 642470
rect 304800 642370 304924 642470
rect 305024 642370 305148 642470
rect 305248 642370 305372 642470
rect 305472 642370 309346 642470
rect 309446 642370 309570 642470
rect 309670 642370 309794 642470
rect 309894 642370 310018 642470
rect 310118 642370 310242 642470
rect 310342 642370 310466 642470
rect 310566 642370 310690 642470
rect 310790 642370 310914 642470
rect 311014 642370 311138 642470
rect 311238 642370 311362 642470
rect 311462 642370 311586 642470
rect 311686 642370 311810 642470
rect 311910 642370 312034 642470
rect 312134 642370 312258 642470
rect 312358 642370 312482 642470
rect 312582 642370 312706 642470
rect 312806 642370 312930 642470
rect 313030 642370 313154 642470
rect 313254 642370 313378 642470
rect 313478 642370 313602 642470
rect 313702 642370 313826 642470
rect 313926 642370 314050 642470
rect 314150 642370 314274 642470
rect 314374 642370 314498 642470
rect 314598 642370 314722 642470
rect 314822 642370 314946 642470
rect 315046 642370 315170 642470
rect 315270 642370 315394 642470
rect 315494 642370 315618 642470
rect 315718 642370 315842 642470
rect 315942 642370 315980 642470
rect 298820 642246 315980 642370
rect 298820 642146 298876 642246
rect 298976 642146 299100 642246
rect 299200 642146 299324 642246
rect 299424 642146 299548 642246
rect 299648 642146 299772 642246
rect 299872 642146 299996 642246
rect 300096 642146 300220 642246
rect 300320 642146 300444 642246
rect 300544 642146 300668 642246
rect 300768 642146 300892 642246
rect 300992 642146 301116 642246
rect 301216 642146 301340 642246
rect 301440 642146 301564 642246
rect 301664 642146 301788 642246
rect 301888 642146 302012 642246
rect 302112 642146 302236 642246
rect 302336 642146 302460 642246
rect 302560 642146 302684 642246
rect 302784 642146 302908 642246
rect 303008 642146 303132 642246
rect 303232 642146 303356 642246
rect 303456 642146 303580 642246
rect 303680 642146 303804 642246
rect 303904 642146 304028 642246
rect 304128 642146 304252 642246
rect 304352 642146 304476 642246
rect 304576 642146 304700 642246
rect 304800 642146 304924 642246
rect 305024 642146 305148 642246
rect 305248 642146 305372 642246
rect 305472 642146 309346 642246
rect 309446 642146 309570 642246
rect 309670 642146 309794 642246
rect 309894 642146 310018 642246
rect 310118 642146 310242 642246
rect 310342 642146 310466 642246
rect 310566 642146 310690 642246
rect 310790 642146 310914 642246
rect 311014 642146 311138 642246
rect 311238 642146 311362 642246
rect 311462 642146 311586 642246
rect 311686 642146 311810 642246
rect 311910 642146 312034 642246
rect 312134 642146 312258 642246
rect 312358 642146 312482 642246
rect 312582 642146 312706 642246
rect 312806 642146 312930 642246
rect 313030 642146 313154 642246
rect 313254 642146 313378 642246
rect 313478 642146 313602 642246
rect 313702 642146 313826 642246
rect 313926 642146 314050 642246
rect 314150 642146 314274 642246
rect 314374 642146 314498 642246
rect 314598 642146 314722 642246
rect 314822 642146 314946 642246
rect 315046 642146 315170 642246
rect 315270 642146 315394 642246
rect 315494 642146 315618 642246
rect 315718 642146 315842 642246
rect 315942 642146 315980 642246
rect 298820 642022 315980 642146
rect 298820 641922 298876 642022
rect 298976 641922 299100 642022
rect 299200 641922 299324 642022
rect 299424 641922 299548 642022
rect 299648 641922 299772 642022
rect 299872 641922 299996 642022
rect 300096 641922 300220 642022
rect 300320 641922 300444 642022
rect 300544 641922 300668 642022
rect 300768 641922 300892 642022
rect 300992 641922 301116 642022
rect 301216 641922 301340 642022
rect 301440 641922 301564 642022
rect 301664 641922 301788 642022
rect 301888 641922 302012 642022
rect 302112 641922 302236 642022
rect 302336 641922 302460 642022
rect 302560 641922 302684 642022
rect 302784 641922 302908 642022
rect 303008 641922 303132 642022
rect 303232 641922 303356 642022
rect 303456 641922 303580 642022
rect 303680 641922 303804 642022
rect 303904 641922 304028 642022
rect 304128 641922 304252 642022
rect 304352 641922 304476 642022
rect 304576 641922 304700 642022
rect 304800 641922 304924 642022
rect 305024 641922 305148 642022
rect 305248 641922 305372 642022
rect 305472 641922 309346 642022
rect 309446 641922 309570 642022
rect 309670 641922 309794 642022
rect 309894 641922 310018 642022
rect 310118 641922 310242 642022
rect 310342 641922 310466 642022
rect 310566 641922 310690 642022
rect 310790 641922 310914 642022
rect 311014 641922 311138 642022
rect 311238 641922 311362 642022
rect 311462 641922 311586 642022
rect 311686 641922 311810 642022
rect 311910 641922 312034 642022
rect 312134 641922 312258 642022
rect 312358 641922 312482 642022
rect 312582 641922 312706 642022
rect 312806 641922 312930 642022
rect 313030 641922 313154 642022
rect 313254 641922 313378 642022
rect 313478 641922 313602 642022
rect 313702 641922 313826 642022
rect 313926 641922 314050 642022
rect 314150 641922 314274 642022
rect 314374 641922 314498 642022
rect 314598 641922 314722 642022
rect 314822 641922 314946 642022
rect 315046 641922 315170 642022
rect 315270 641922 315394 642022
rect 315494 641922 315618 642022
rect 315718 641922 315842 642022
rect 315942 641922 315980 642022
rect 298820 641798 315980 641922
rect 298820 641698 298876 641798
rect 298976 641698 299100 641798
rect 299200 641698 299324 641798
rect 299424 641698 299548 641798
rect 299648 641698 299772 641798
rect 299872 641698 299996 641798
rect 300096 641698 300220 641798
rect 300320 641698 300444 641798
rect 300544 641698 300668 641798
rect 300768 641698 300892 641798
rect 300992 641698 301116 641798
rect 301216 641698 301340 641798
rect 301440 641698 301564 641798
rect 301664 641698 301788 641798
rect 301888 641698 302012 641798
rect 302112 641698 302236 641798
rect 302336 641698 302460 641798
rect 302560 641698 302684 641798
rect 302784 641698 302908 641798
rect 303008 641698 303132 641798
rect 303232 641698 303356 641798
rect 303456 641698 303580 641798
rect 303680 641698 303804 641798
rect 303904 641698 304028 641798
rect 304128 641698 304252 641798
rect 304352 641698 304476 641798
rect 304576 641698 304700 641798
rect 304800 641698 304924 641798
rect 305024 641698 305148 641798
rect 305248 641698 305372 641798
rect 305472 641698 309346 641798
rect 309446 641698 309570 641798
rect 309670 641698 309794 641798
rect 309894 641698 310018 641798
rect 310118 641698 310242 641798
rect 310342 641698 310466 641798
rect 310566 641698 310690 641798
rect 310790 641698 310914 641798
rect 311014 641698 311138 641798
rect 311238 641698 311362 641798
rect 311462 641698 311586 641798
rect 311686 641698 311810 641798
rect 311910 641698 312034 641798
rect 312134 641698 312258 641798
rect 312358 641698 312482 641798
rect 312582 641698 312706 641798
rect 312806 641698 312930 641798
rect 313030 641698 313154 641798
rect 313254 641698 313378 641798
rect 313478 641698 313602 641798
rect 313702 641698 313826 641798
rect 313926 641698 314050 641798
rect 314150 641698 314274 641798
rect 314374 641698 314498 641798
rect 314598 641698 314722 641798
rect 314822 641698 314946 641798
rect 315046 641698 315170 641798
rect 315270 641698 315394 641798
rect 315494 641698 315618 641798
rect 315718 641698 315842 641798
rect 315942 641698 315980 641798
rect 298820 641660 315980 641698
rect 288920 631440 289920 637184
rect 294704 631440 295576 637184
rect 288920 623784 295576 631440
rect 297820 637996 298880 638020
rect 297820 637896 297850 637996
rect 297950 637896 298074 637996
rect 298174 637896 298298 637996
rect 298398 637896 298522 637996
rect 298622 637896 298746 637996
rect 298846 637896 298880 637996
rect 297820 637772 298880 637896
rect 297820 637672 297850 637772
rect 297950 637672 298074 637772
rect 298174 637672 298298 637772
rect 298398 637672 298522 637772
rect 298622 637672 298746 637772
rect 298846 637672 298880 637772
rect 297820 637548 298880 637672
rect 297820 637448 297850 637548
rect 297950 637448 298074 637548
rect 298174 637448 298298 637548
rect 298398 637448 298522 637548
rect 298622 637448 298746 637548
rect 298846 637448 298880 637548
rect 297820 637324 298880 637448
rect 297820 637224 297850 637324
rect 297950 637224 298074 637324
rect 298174 637224 298298 637324
rect 298398 637224 298522 637324
rect 298622 637224 298746 637324
rect 298846 637224 298880 637324
rect 297820 637100 298880 637224
rect 297820 637000 297850 637100
rect 297950 637000 298074 637100
rect 298174 637000 298298 637100
rect 298398 637000 298522 637100
rect 298622 637000 298746 637100
rect 298846 637000 298880 637100
rect 297820 636876 298880 637000
rect 297820 636776 297850 636876
rect 297950 636776 298074 636876
rect 298174 636776 298298 636876
rect 298398 636776 298522 636876
rect 298622 636776 298746 636876
rect 298846 636776 298880 636876
rect 297820 636652 298880 636776
rect 297820 636552 297850 636652
rect 297950 636552 298074 636652
rect 298174 636552 298298 636652
rect 298398 636552 298522 636652
rect 298622 636552 298746 636652
rect 298846 636552 298880 636652
rect 297820 636428 298880 636552
rect 297820 636328 297850 636428
rect 297950 636328 298074 636428
rect 298174 636328 298298 636428
rect 298398 636328 298522 636428
rect 298622 636328 298746 636428
rect 298846 636328 298880 636428
rect 297820 636204 298880 636328
rect 297820 636104 297850 636204
rect 297950 636104 298074 636204
rect 298174 636104 298298 636204
rect 298398 636104 298522 636204
rect 298622 636104 298746 636204
rect 298846 636104 298880 636204
rect 297820 635980 298880 636104
rect 297820 635880 297850 635980
rect 297950 635880 298074 635980
rect 298174 635880 298298 635980
rect 298398 635880 298522 635980
rect 298622 635880 298746 635980
rect 298846 635880 298880 635980
rect 297820 635756 298880 635880
rect 297820 635656 297850 635756
rect 297950 635656 298074 635756
rect 298174 635656 298298 635756
rect 298398 635656 298522 635756
rect 298622 635656 298746 635756
rect 298846 635656 298880 635756
rect 297820 635532 298880 635656
rect 297820 635432 297850 635532
rect 297950 635432 298074 635532
rect 298174 635432 298298 635532
rect 298398 635432 298522 635532
rect 298622 635432 298746 635532
rect 298846 635432 298880 635532
rect 297820 635308 298880 635432
rect 297820 635208 297850 635308
rect 297950 635208 298074 635308
rect 298174 635208 298298 635308
rect 298398 635208 298522 635308
rect 298622 635208 298746 635308
rect 298846 635208 298880 635308
rect 297820 635084 298880 635208
rect 297820 634984 297850 635084
rect 297950 634984 298074 635084
rect 298174 634984 298298 635084
rect 298398 634984 298522 635084
rect 298622 634984 298746 635084
rect 298846 634984 298880 635084
rect 297820 634860 298880 634984
rect 297820 634760 297850 634860
rect 297950 634760 298074 634860
rect 298174 634760 298298 634860
rect 298398 634760 298522 634860
rect 298622 634760 298746 634860
rect 298846 634760 298880 634860
rect 297820 634636 298880 634760
rect 297820 634536 297850 634636
rect 297950 634536 298074 634636
rect 298174 634536 298298 634636
rect 298398 634536 298522 634636
rect 298622 634536 298746 634636
rect 298846 634536 298880 634636
rect 297820 634412 298880 634536
rect 297820 634312 297850 634412
rect 297950 634312 298074 634412
rect 298174 634312 298298 634412
rect 298398 634312 298522 634412
rect 298622 634312 298746 634412
rect 298846 634312 298880 634412
rect 297820 634188 298880 634312
rect 297820 634088 297850 634188
rect 297950 634088 298074 634188
rect 298174 634088 298298 634188
rect 298398 634088 298522 634188
rect 298622 634088 298746 634188
rect 298846 634088 298880 634188
rect 297820 633964 298880 634088
rect 297820 633864 297850 633964
rect 297950 633864 298074 633964
rect 298174 633864 298298 633964
rect 298398 633864 298522 633964
rect 298622 633864 298746 633964
rect 298846 633864 298880 633964
rect 297820 633740 298880 633864
rect 297820 633640 297850 633740
rect 297950 633640 298074 633740
rect 298174 633640 298298 633740
rect 298398 633640 298522 633740
rect 298622 633640 298746 633740
rect 298846 633640 298880 633740
rect 297820 633516 298880 633640
rect 297820 633416 297850 633516
rect 297950 633416 298074 633516
rect 298174 633416 298298 633516
rect 298398 633416 298522 633516
rect 298622 633416 298746 633516
rect 298846 633416 298880 633516
rect 297820 633292 298880 633416
rect 297820 633192 297850 633292
rect 297950 633192 298074 633292
rect 298174 633192 298298 633292
rect 298398 633192 298522 633292
rect 298622 633192 298746 633292
rect 298846 633192 298880 633292
rect 297820 633068 298880 633192
rect 297820 632968 297850 633068
rect 297950 632968 298074 633068
rect 298174 632968 298298 633068
rect 298398 632968 298522 633068
rect 298622 632968 298746 633068
rect 298846 632968 298880 633068
rect 297820 632844 298880 632968
rect 297820 632744 297850 632844
rect 297950 632744 298074 632844
rect 298174 632744 298298 632844
rect 298398 632744 298522 632844
rect 298622 632744 298746 632844
rect 298846 632744 298880 632844
rect 297820 632620 298880 632744
rect 297820 632520 297850 632620
rect 297950 632520 298074 632620
rect 298174 632520 298298 632620
rect 298398 632520 298522 632620
rect 298622 632520 298746 632620
rect 298846 632520 298880 632620
rect 297820 632396 298880 632520
rect 297820 632296 297850 632396
rect 297950 632296 298074 632396
rect 298174 632296 298298 632396
rect 298398 632296 298522 632396
rect 298622 632296 298746 632396
rect 298846 632296 298880 632396
rect 297820 632172 298880 632296
rect 297820 632072 297850 632172
rect 297950 632072 298074 632172
rect 298174 632072 298298 632172
rect 298398 632072 298522 632172
rect 298622 632072 298746 632172
rect 298846 632072 298880 632172
rect 297820 631948 298880 632072
rect 297820 631848 297850 631948
rect 297950 631848 298074 631948
rect 298174 631848 298298 631948
rect 298398 631848 298522 631948
rect 298622 631848 298746 631948
rect 298846 631848 298880 631948
rect 297820 631724 298880 631848
rect 297820 631624 297850 631724
rect 297950 631624 298074 631724
rect 298174 631624 298298 631724
rect 298398 631624 298522 631724
rect 298622 631624 298746 631724
rect 298846 631624 298880 631724
rect 297820 631500 298880 631624
rect 297820 631400 297850 631500
rect 297950 631400 298074 631500
rect 298174 631400 298298 631500
rect 298398 631400 298522 631500
rect 298622 631400 298746 631500
rect 298846 631400 298880 631500
rect 297820 631360 298880 631400
rect 319000 628868 334400 650200
rect 335580 650904 342400 651380
rect 335580 645160 336480 650904
rect 341264 645160 342400 650904
rect 335580 642744 342400 645160
rect 510602 650961 515394 651406
rect 515386 645217 515394 650961
rect 510602 644744 515394 645217
rect 335576 642714 342400 642744
rect 335576 642614 335616 642714
rect 335716 642614 335840 642714
rect 335940 642614 336064 642714
rect 336164 642614 336288 642714
rect 336388 642614 336512 642714
rect 336612 642614 336736 642714
rect 336836 642614 336960 642714
rect 337060 642614 337184 642714
rect 337284 642614 337408 642714
rect 337508 642614 337632 642714
rect 337732 642614 337856 642714
rect 337956 642614 338080 642714
rect 338180 642614 338304 642714
rect 338404 642614 338528 642714
rect 338628 642614 338752 642714
rect 338852 642614 338976 642714
rect 339076 642614 339200 642714
rect 339300 642614 339424 642714
rect 339524 642614 339648 642714
rect 339748 642614 339872 642714
rect 339972 642614 340096 642714
rect 340196 642614 340320 642714
rect 340420 642614 340544 642714
rect 340644 642614 340768 642714
rect 340868 642614 340992 642714
rect 341092 642614 341216 642714
rect 341316 642614 341440 642714
rect 341540 642614 341664 642714
rect 341764 642614 341888 642714
rect 341988 642614 342112 642714
rect 342212 642614 342400 642714
rect 335576 642490 342400 642614
rect 335576 642390 335616 642490
rect 335716 642390 335840 642490
rect 335940 642390 336064 642490
rect 336164 642390 336288 642490
rect 336388 642390 336512 642490
rect 336612 642390 336736 642490
rect 336836 642390 336960 642490
rect 337060 642390 337184 642490
rect 337284 642390 337408 642490
rect 337508 642390 337632 642490
rect 337732 642390 337856 642490
rect 337956 642390 338080 642490
rect 338180 642390 338304 642490
rect 338404 642390 338528 642490
rect 338628 642390 338752 642490
rect 338852 642390 338976 642490
rect 339076 642390 339200 642490
rect 339300 642390 339424 642490
rect 339524 642390 339648 642490
rect 339748 642390 339872 642490
rect 339972 642390 340096 642490
rect 340196 642390 340320 642490
rect 340420 642390 340544 642490
rect 340644 642390 340768 642490
rect 340868 642390 340992 642490
rect 341092 642390 341216 642490
rect 341316 642390 341440 642490
rect 341540 642390 341664 642490
rect 341764 642390 341888 642490
rect 341988 642390 342112 642490
rect 342212 642390 342400 642490
rect 335576 642266 342400 642390
rect 335576 642166 335616 642266
rect 335716 642166 335840 642266
rect 335940 642166 336064 642266
rect 336164 642166 336288 642266
rect 336388 642166 336512 642266
rect 336612 642166 336736 642266
rect 336836 642166 336960 642266
rect 337060 642166 337184 642266
rect 337284 642166 337408 642266
rect 337508 642166 337632 642266
rect 337732 642166 337856 642266
rect 337956 642166 338080 642266
rect 338180 642166 338304 642266
rect 338404 642166 338528 642266
rect 338628 642166 338752 642266
rect 338852 642166 338976 642266
rect 339076 642166 339200 642266
rect 339300 642166 339424 642266
rect 339524 642166 339648 642266
rect 339748 642166 339872 642266
rect 339972 642166 340096 642266
rect 340196 642166 340320 642266
rect 340420 642166 340544 642266
rect 340644 642166 340768 642266
rect 340868 642166 340992 642266
rect 341092 642166 341216 642266
rect 341316 642166 341440 642266
rect 341540 642166 341664 642266
rect 341764 642166 341888 642266
rect 341988 642166 342112 642266
rect 342212 642166 342400 642266
rect 335576 642042 342400 642166
rect 335576 641942 335616 642042
rect 335716 641942 335840 642042
rect 335940 641942 336064 642042
rect 336164 641942 336288 642042
rect 336388 641942 336512 642042
rect 336612 641942 336736 642042
rect 336836 641942 336960 642042
rect 337060 641942 337184 642042
rect 337284 641942 337408 642042
rect 337508 641942 337632 642042
rect 337732 641942 337856 642042
rect 337956 641942 338080 642042
rect 338180 641942 338304 642042
rect 338404 641942 338528 642042
rect 338628 641942 338752 642042
rect 338852 641942 338976 642042
rect 339076 641942 339200 642042
rect 339300 641942 339424 642042
rect 339524 641942 339648 642042
rect 339748 641942 339872 642042
rect 339972 641942 340096 642042
rect 340196 641942 340320 642042
rect 340420 641942 340544 642042
rect 340644 641942 340768 642042
rect 340868 641942 340992 642042
rect 341092 641942 341216 642042
rect 341316 641942 341440 642042
rect 341540 641942 341664 642042
rect 341764 641942 341888 642042
rect 341988 641942 342112 642042
rect 342212 641942 342400 642042
rect 335576 641818 342400 641942
rect 335576 641718 335616 641818
rect 335716 641718 335840 641818
rect 335940 641718 336064 641818
rect 336164 641718 336288 641818
rect 336388 641718 336512 641818
rect 336612 641718 336736 641818
rect 336836 641718 336960 641818
rect 337060 641718 337184 641818
rect 337284 641718 337408 641818
rect 337508 641718 337632 641818
rect 337732 641718 337856 641818
rect 337956 641718 338080 641818
rect 338180 641718 338304 641818
rect 338404 641718 338528 641818
rect 338628 641718 338752 641818
rect 338852 641718 338976 641818
rect 339076 641718 339200 641818
rect 339300 641718 339424 641818
rect 339524 641718 339648 641818
rect 339748 641718 339872 641818
rect 339972 641718 340096 641818
rect 340196 641718 340320 641818
rect 340420 641718 340544 641818
rect 340644 641718 340768 641818
rect 340868 641718 340992 641818
rect 341092 641718 341216 641818
rect 341316 641718 341440 641818
rect 341540 641718 341664 641818
rect 341764 641718 341888 641818
rect 341988 641718 342112 641818
rect 342212 641718 342400 641818
rect 335576 641684 342400 641718
rect 335580 641660 342400 641684
rect 342100 637996 343160 638020
rect 342100 637896 342130 637996
rect 342230 637896 342354 637996
rect 342454 637896 342578 637996
rect 342678 637896 342802 637996
rect 342902 637896 343026 637996
rect 343126 637896 343160 637996
rect 342100 637772 343160 637896
rect 342100 637672 342130 637772
rect 342230 637672 342354 637772
rect 342454 637672 342578 637772
rect 342678 637672 342802 637772
rect 342902 637672 343026 637772
rect 343126 637672 343160 637772
rect 342100 637548 343160 637672
rect 342100 637448 342130 637548
rect 342230 637448 342354 637548
rect 342454 637448 342578 637548
rect 342678 637448 342802 637548
rect 342902 637448 343026 637548
rect 343126 637448 343160 637548
rect 342100 637324 343160 637448
rect 342100 637224 342130 637324
rect 342230 637224 342354 637324
rect 342454 637224 342578 637324
rect 342678 637224 342802 637324
rect 342902 637224 343026 637324
rect 343126 637224 343160 637324
rect 342100 637100 343160 637224
rect 342100 637000 342130 637100
rect 342230 637000 342354 637100
rect 342454 637000 342578 637100
rect 342678 637000 342802 637100
rect 342902 637000 343026 637100
rect 343126 637000 343160 637100
rect 342100 636876 343160 637000
rect 342100 636776 342130 636876
rect 342230 636776 342354 636876
rect 342454 636776 342578 636876
rect 342678 636776 342802 636876
rect 342902 636776 343026 636876
rect 343126 636776 343160 636876
rect 342100 636652 343160 636776
rect 342100 636552 342130 636652
rect 342230 636552 342354 636652
rect 342454 636552 342578 636652
rect 342678 636552 342802 636652
rect 342902 636552 343026 636652
rect 343126 636552 343160 636652
rect 342100 636428 343160 636552
rect 342100 636328 342130 636428
rect 342230 636328 342354 636428
rect 342454 636328 342578 636428
rect 342678 636328 342802 636428
rect 342902 636328 343026 636428
rect 343126 636328 343160 636428
rect 342100 636204 343160 636328
rect 342100 636104 342130 636204
rect 342230 636104 342354 636204
rect 342454 636104 342578 636204
rect 342678 636104 342802 636204
rect 342902 636104 343026 636204
rect 343126 636104 343160 636204
rect 342100 635980 343160 636104
rect 342100 635880 342130 635980
rect 342230 635880 342354 635980
rect 342454 635880 342578 635980
rect 342678 635880 342802 635980
rect 342902 635880 343026 635980
rect 343126 635880 343160 635980
rect 342100 635756 343160 635880
rect 342100 635656 342130 635756
rect 342230 635656 342354 635756
rect 342454 635656 342578 635756
rect 342678 635656 342802 635756
rect 342902 635656 343026 635756
rect 343126 635656 343160 635756
rect 342100 635532 343160 635656
rect 342100 635432 342130 635532
rect 342230 635432 342354 635532
rect 342454 635432 342578 635532
rect 342678 635432 342802 635532
rect 342902 635432 343026 635532
rect 343126 635432 343160 635532
rect 342100 635308 343160 635432
rect 342100 635208 342130 635308
rect 342230 635208 342354 635308
rect 342454 635208 342578 635308
rect 342678 635208 342802 635308
rect 342902 635208 343026 635308
rect 343126 635208 343160 635308
rect 342100 635084 343160 635208
rect 342100 634984 342130 635084
rect 342230 634984 342354 635084
rect 342454 634984 342578 635084
rect 342678 634984 342802 635084
rect 342902 634984 343026 635084
rect 343126 634984 343160 635084
rect 342100 634860 343160 634984
rect 342100 634760 342130 634860
rect 342230 634760 342354 634860
rect 342454 634760 342578 634860
rect 342678 634760 342802 634860
rect 342902 634760 343026 634860
rect 343126 634760 343160 634860
rect 342100 634636 343160 634760
rect 342100 634536 342130 634636
rect 342230 634536 342354 634636
rect 342454 634536 342578 634636
rect 342678 634536 342802 634636
rect 342902 634536 343026 634636
rect 343126 634536 343160 634636
rect 342100 634412 343160 634536
rect 342100 634312 342130 634412
rect 342230 634312 342354 634412
rect 342454 634312 342578 634412
rect 342678 634312 342802 634412
rect 342902 634312 343026 634412
rect 343126 634312 343160 634412
rect 342100 634188 343160 634312
rect 342100 634088 342130 634188
rect 342230 634088 342354 634188
rect 342454 634088 342578 634188
rect 342678 634088 342802 634188
rect 342902 634088 343026 634188
rect 343126 634088 343160 634188
rect 342100 633964 343160 634088
rect 342100 633864 342130 633964
rect 342230 633864 342354 633964
rect 342454 633864 342578 633964
rect 342678 633864 342802 633964
rect 342902 633864 343026 633964
rect 343126 633864 343160 633964
rect 342100 633740 343160 633864
rect 342100 633640 342130 633740
rect 342230 633640 342354 633740
rect 342454 633640 342578 633740
rect 342678 633640 342802 633740
rect 342902 633640 343026 633740
rect 343126 633640 343160 633740
rect 342100 633516 343160 633640
rect 342100 633416 342130 633516
rect 342230 633416 342354 633516
rect 342454 633416 342578 633516
rect 342678 633416 342802 633516
rect 342902 633416 343026 633516
rect 343126 633416 343160 633516
rect 342100 633292 343160 633416
rect 342100 633192 342130 633292
rect 342230 633192 342354 633292
rect 342454 633192 342578 633292
rect 342678 633192 342802 633292
rect 342902 633192 343026 633292
rect 343126 633192 343160 633292
rect 342100 633068 343160 633192
rect 342100 632968 342130 633068
rect 342230 632968 342354 633068
rect 342454 632968 342578 633068
rect 342678 632968 342802 633068
rect 342902 632968 343026 633068
rect 343126 632968 343160 633068
rect 342100 632844 343160 632968
rect 342100 632744 342130 632844
rect 342230 632744 342354 632844
rect 342454 632744 342578 632844
rect 342678 632744 342802 632844
rect 342902 632744 343026 632844
rect 343126 632744 343160 632844
rect 342100 632620 343160 632744
rect 342100 632520 342130 632620
rect 342230 632520 342354 632620
rect 342454 632520 342578 632620
rect 342678 632520 342802 632620
rect 342902 632520 343026 632620
rect 343126 632520 343160 632620
rect 342100 632396 343160 632520
rect 342100 632296 342130 632396
rect 342230 632296 342354 632396
rect 342454 632296 342578 632396
rect 342678 632296 342802 632396
rect 342902 632296 343026 632396
rect 343126 632296 343160 632396
rect 342100 632172 343160 632296
rect 342100 632072 342130 632172
rect 342230 632072 342354 632172
rect 342454 632072 342578 632172
rect 342678 632072 342802 632172
rect 342902 632072 343026 632172
rect 343126 632072 343160 632172
rect 342100 631948 343160 632072
rect 342100 631848 342130 631948
rect 342230 631848 342354 631948
rect 342454 631848 342578 631948
rect 342678 631848 342802 631948
rect 342902 631848 343026 631948
rect 343126 631848 343160 631948
rect 342100 631724 343160 631848
rect 342100 631624 342130 631724
rect 342230 631624 342354 631724
rect 342454 631624 342578 631724
rect 342678 631624 342802 631724
rect 342902 631624 343026 631724
rect 343126 631624 343160 631724
rect 342100 631500 343160 631624
rect 342100 631400 342130 631500
rect 342230 631400 342354 631500
rect 342454 631400 342578 631500
rect 342678 631400 342802 631500
rect 342902 631400 343026 631500
rect 343126 631400 343160 631500
rect 342100 631360 343160 631400
rect 510594 637561 515394 644744
rect 510594 631817 510602 637561
rect 515386 631817 515394 637561
rect 319000 628668 319400 628868
rect 319600 628668 319834 628868
rect 320034 628668 320268 628868
rect 320468 628668 320702 628868
rect 320902 628668 321136 628868
rect 321336 628668 321570 628868
rect 321770 628668 322004 628868
rect 322204 628668 322438 628868
rect 322638 628668 322872 628868
rect 323072 628668 323306 628868
rect 323506 628668 323740 628868
rect 323940 628668 324140 628868
rect 324340 628668 324540 628868
rect 324740 628668 324940 628868
rect 325140 628668 325340 628868
rect 325540 628668 325740 628868
rect 325940 628668 326140 628868
rect 326340 628668 326540 628868
rect 326740 628668 326940 628868
rect 327140 628668 327340 628868
rect 327540 628668 328940 628868
rect 329140 628668 329340 628868
rect 329540 628668 329740 628868
rect 329940 628668 330140 628868
rect 330340 628668 330540 628868
rect 330740 628668 330940 628868
rect 331140 628668 331340 628868
rect 331540 628668 331740 628868
rect 331940 628668 332140 628868
rect 332340 628668 334400 628868
rect 319000 628434 334400 628668
rect 319000 628234 319400 628434
rect 319600 628234 319834 628434
rect 320034 628234 320268 628434
rect 320468 628234 320702 628434
rect 320902 628234 321136 628434
rect 321336 628234 321570 628434
rect 321770 628234 322004 628434
rect 322204 628234 322438 628434
rect 322638 628234 322872 628434
rect 323072 628234 323306 628434
rect 323506 628234 323740 628434
rect 323940 628234 334400 628434
rect 319000 628000 334400 628234
rect 319000 627800 319400 628000
rect 319600 627800 319834 628000
rect 320034 627800 320268 628000
rect 320468 627800 320702 628000
rect 320902 627800 321136 628000
rect 321336 627800 321570 628000
rect 321770 627800 322004 628000
rect 322204 627800 322438 628000
rect 322638 627800 322872 628000
rect 323072 627800 323306 628000
rect 323506 627800 323740 628000
rect 323940 627800 334400 628000
rect 319000 627600 334400 627800
rect 297792 626176 303552 626240
rect 297792 626112 297856 626176
rect 297920 626112 297984 626176
rect 298048 626112 298112 626176
rect 298176 626112 298240 626176
rect 298304 626112 298368 626176
rect 298432 626112 298496 626176
rect 298560 626112 298624 626176
rect 298688 626112 298752 626176
rect 298816 626112 298880 626176
rect 298944 626112 303552 626176
rect 297792 626048 303552 626112
rect 297792 625984 297856 626048
rect 297920 625984 297984 626048
rect 298048 625984 298112 626048
rect 298176 625984 298240 626048
rect 298304 625984 298368 626048
rect 298432 625984 298496 626048
rect 298560 625984 298624 626048
rect 298688 625984 298752 626048
rect 298816 625984 298880 626048
rect 298944 626030 303552 626048
rect 298944 625984 302980 626030
rect 297792 625970 302980 625984
rect 303040 625970 303100 626030
rect 303160 625970 303220 626030
rect 303280 625970 303340 626030
rect 303400 625970 303460 626030
rect 303520 625970 303552 626030
rect 297792 625920 303552 625970
rect 297792 625856 297856 625920
rect 297920 625856 297984 625920
rect 298048 625856 298112 625920
rect 298176 625856 298240 625920
rect 298304 625856 298368 625920
rect 298432 625856 298496 625920
rect 298560 625856 298624 625920
rect 298688 625856 298752 625920
rect 298816 625856 298880 625920
rect 298944 625910 303552 625920
rect 298944 625856 302980 625910
rect 297792 625850 302980 625856
rect 303040 625850 303100 625910
rect 303160 625850 303220 625910
rect 303280 625850 303340 625910
rect 303400 625850 303460 625910
rect 303520 625850 303552 625910
rect 297792 625792 303552 625850
rect 297792 625728 297856 625792
rect 297920 625728 297984 625792
rect 298048 625728 298112 625792
rect 298176 625728 298240 625792
rect 298304 625728 298368 625792
rect 298432 625728 298496 625792
rect 298560 625728 298624 625792
rect 298688 625728 298752 625792
rect 298816 625728 298880 625792
rect 298944 625728 303552 625792
rect 297792 625664 303552 625728
rect 510594 624606 515394 631817
rect 297820 624600 298878 624606
rect 342100 624600 343186 624606
rect 288920 618040 289920 623784
rect 294704 618040 295576 623784
rect 288920 610764 295576 618040
rect 297720 624596 298880 624600
rect 297720 624496 297850 624596
rect 297950 624496 298074 624596
rect 298174 624496 298298 624596
rect 298398 624496 298522 624596
rect 298622 624496 298746 624596
rect 298846 624496 298880 624596
rect 297720 624372 298880 624496
rect 297720 624272 297850 624372
rect 297950 624272 298074 624372
rect 298174 624272 298298 624372
rect 298398 624272 298522 624372
rect 298622 624272 298746 624372
rect 298846 624272 298880 624372
rect 297720 624148 298880 624272
rect 297720 624048 297850 624148
rect 297950 624048 298074 624148
rect 298174 624048 298298 624148
rect 298398 624048 298522 624148
rect 298622 624048 298746 624148
rect 298846 624048 298880 624148
rect 297720 623924 298880 624048
rect 297720 623824 297850 623924
rect 297950 623824 298074 623924
rect 298174 623824 298298 623924
rect 298398 623824 298522 623924
rect 298622 623824 298746 623924
rect 298846 623824 298880 623924
rect 297720 623700 298880 623824
rect 297720 623600 297850 623700
rect 297950 623600 298074 623700
rect 298174 623600 298298 623700
rect 298398 623600 298522 623700
rect 298622 623600 298746 623700
rect 298846 623600 298880 623700
rect 297720 623476 298880 623600
rect 297720 623376 297850 623476
rect 297950 623376 298074 623476
rect 298174 623376 298298 623476
rect 298398 623376 298522 623476
rect 298622 623376 298746 623476
rect 298846 623376 298880 623476
rect 297720 623252 298880 623376
rect 297720 623152 297850 623252
rect 297950 623152 298074 623252
rect 298174 623152 298298 623252
rect 298398 623152 298522 623252
rect 298622 623152 298746 623252
rect 298846 623152 298880 623252
rect 297720 623028 298880 623152
rect 297720 622928 297850 623028
rect 297950 622928 298074 623028
rect 298174 622928 298298 623028
rect 298398 622928 298522 623028
rect 298622 622928 298746 623028
rect 298846 622928 298880 623028
rect 297720 622804 298880 622928
rect 297720 622704 297850 622804
rect 297950 622704 298074 622804
rect 298174 622704 298298 622804
rect 298398 622704 298522 622804
rect 298622 622704 298746 622804
rect 298846 622704 298880 622804
rect 297720 622580 298880 622704
rect 297720 622480 297850 622580
rect 297950 622480 298074 622580
rect 298174 622480 298298 622580
rect 298398 622480 298522 622580
rect 298622 622480 298746 622580
rect 298846 622480 298880 622580
rect 297720 622356 298880 622480
rect 297720 622256 297850 622356
rect 297950 622256 298074 622356
rect 298174 622256 298298 622356
rect 298398 622256 298522 622356
rect 298622 622256 298746 622356
rect 298846 622256 298880 622356
rect 297720 622132 298880 622256
rect 297720 622032 297850 622132
rect 297950 622032 298074 622132
rect 298174 622032 298298 622132
rect 298398 622032 298522 622132
rect 298622 622032 298746 622132
rect 298846 622032 298880 622132
rect 297720 621908 298880 622032
rect 297720 621808 297850 621908
rect 297950 621808 298074 621908
rect 298174 621808 298298 621908
rect 298398 621808 298522 621908
rect 298622 621808 298746 621908
rect 298846 621808 298880 621908
rect 297720 621684 298880 621808
rect 297720 621584 297850 621684
rect 297950 621584 298074 621684
rect 298174 621584 298298 621684
rect 298398 621584 298522 621684
rect 298622 621584 298746 621684
rect 298846 621584 298880 621684
rect 297720 621460 298880 621584
rect 297720 621360 297850 621460
rect 297950 621360 298074 621460
rect 298174 621360 298298 621460
rect 298398 621360 298522 621460
rect 298622 621360 298746 621460
rect 298846 621360 298880 621460
rect 297720 621236 298880 621360
rect 297720 621136 297850 621236
rect 297950 621136 298074 621236
rect 298174 621136 298298 621236
rect 298398 621136 298522 621236
rect 298622 621136 298746 621236
rect 298846 621136 298880 621236
rect 297720 621012 298880 621136
rect 297720 620912 297850 621012
rect 297950 620912 298074 621012
rect 298174 620912 298298 621012
rect 298398 620912 298522 621012
rect 298622 620912 298746 621012
rect 298846 620912 298880 621012
rect 297720 620788 298880 620912
rect 297720 620688 297850 620788
rect 297950 620688 298074 620788
rect 298174 620688 298298 620788
rect 298398 620688 298522 620788
rect 298622 620688 298746 620788
rect 298846 620688 298880 620788
rect 297720 620564 298880 620688
rect 297720 620464 297850 620564
rect 297950 620464 298074 620564
rect 298174 620464 298298 620564
rect 298398 620464 298522 620564
rect 298622 620464 298746 620564
rect 298846 620464 298880 620564
rect 297720 620340 298880 620464
rect 297720 620240 297850 620340
rect 297950 620240 298074 620340
rect 298174 620240 298298 620340
rect 298398 620240 298522 620340
rect 298622 620240 298746 620340
rect 298846 620240 298880 620340
rect 297720 620116 298880 620240
rect 297720 620016 297850 620116
rect 297950 620016 298074 620116
rect 298174 620016 298298 620116
rect 298398 620016 298522 620116
rect 298622 620016 298746 620116
rect 298846 620016 298880 620116
rect 297720 619892 298880 620016
rect 297720 619792 297850 619892
rect 297950 619792 298074 619892
rect 298174 619792 298298 619892
rect 298398 619792 298522 619892
rect 298622 619792 298746 619892
rect 298846 619792 298880 619892
rect 297720 619668 298880 619792
rect 297720 619568 297850 619668
rect 297950 619568 298074 619668
rect 298174 619568 298298 619668
rect 298398 619568 298522 619668
rect 298622 619568 298746 619668
rect 298846 619568 298880 619668
rect 297720 619444 298880 619568
rect 297720 619344 297850 619444
rect 297950 619344 298074 619444
rect 298174 619344 298298 619444
rect 298398 619344 298522 619444
rect 298622 619344 298746 619444
rect 298846 619344 298880 619444
rect 297720 619220 298880 619344
rect 297720 619120 297850 619220
rect 297950 619120 298074 619220
rect 298174 619120 298298 619220
rect 298398 619120 298522 619220
rect 298622 619120 298746 619220
rect 298846 619120 298880 619220
rect 297720 618996 298880 619120
rect 297720 618896 297850 618996
rect 297950 618896 298074 618996
rect 298174 618896 298298 618996
rect 298398 618896 298522 618996
rect 298622 618896 298746 618996
rect 298846 618896 298880 618996
rect 297720 618772 298880 618896
rect 297720 618672 297850 618772
rect 297950 618672 298074 618772
rect 298174 618672 298298 618772
rect 298398 618672 298522 618772
rect 298622 618672 298746 618772
rect 298846 618672 298880 618772
rect 297720 618548 298880 618672
rect 297720 618448 297850 618548
rect 297950 618448 298074 618548
rect 298174 618448 298298 618548
rect 298398 618448 298522 618548
rect 298622 618448 298746 618548
rect 298846 618448 298880 618548
rect 297720 618324 298880 618448
rect 297720 618224 297850 618324
rect 297950 618224 298074 618324
rect 298174 618224 298298 618324
rect 298398 618224 298522 618324
rect 298622 618224 298746 618324
rect 298846 618224 298880 618324
rect 297720 618100 298880 618224
rect 297720 618000 297850 618100
rect 297950 618000 298074 618100
rect 298174 618000 298298 618100
rect 298398 618000 298522 618100
rect 298622 618000 298746 618100
rect 298846 618000 298880 618100
rect 297720 617944 298880 618000
rect 342000 624596 343186 624600
rect 342000 624496 342130 624596
rect 342230 624496 342354 624596
rect 342454 624496 342578 624596
rect 342678 624496 342802 624596
rect 342902 624496 343026 624596
rect 343126 624496 343186 624596
rect 342000 624372 343186 624496
rect 342000 624272 342130 624372
rect 342230 624272 342354 624372
rect 342454 624272 342578 624372
rect 342678 624272 342802 624372
rect 342902 624272 343026 624372
rect 343126 624272 343186 624372
rect 342000 624148 343186 624272
rect 342000 624048 342130 624148
rect 342230 624048 342354 624148
rect 342454 624048 342578 624148
rect 342678 624048 342802 624148
rect 342902 624048 343026 624148
rect 343126 624048 343186 624148
rect 342000 623924 343186 624048
rect 342000 623824 342130 623924
rect 342230 623824 342354 623924
rect 342454 623824 342578 623924
rect 342678 623824 342802 623924
rect 342902 623824 343026 623924
rect 343126 623824 343186 623924
rect 342000 623700 343186 623824
rect 342000 623600 342130 623700
rect 342230 623600 342354 623700
rect 342454 623600 342578 623700
rect 342678 623600 342802 623700
rect 342902 623600 343026 623700
rect 343126 623600 343186 623700
rect 342000 623476 343186 623600
rect 342000 623376 342130 623476
rect 342230 623376 342354 623476
rect 342454 623376 342578 623476
rect 342678 623376 342802 623476
rect 342902 623376 343026 623476
rect 343126 623376 343186 623476
rect 342000 623252 343186 623376
rect 342000 623152 342130 623252
rect 342230 623152 342354 623252
rect 342454 623152 342578 623252
rect 342678 623152 342802 623252
rect 342902 623152 343026 623252
rect 343126 623152 343186 623252
rect 342000 623028 343186 623152
rect 342000 622928 342130 623028
rect 342230 622928 342354 623028
rect 342454 622928 342578 623028
rect 342678 622928 342802 623028
rect 342902 622928 343026 623028
rect 343126 622928 343186 623028
rect 342000 622804 343186 622928
rect 342000 622704 342130 622804
rect 342230 622704 342354 622804
rect 342454 622704 342578 622804
rect 342678 622704 342802 622804
rect 342902 622704 343026 622804
rect 343126 622704 343186 622804
rect 342000 622580 343186 622704
rect 342000 622480 342130 622580
rect 342230 622480 342354 622580
rect 342454 622480 342578 622580
rect 342678 622480 342802 622580
rect 342902 622480 343026 622580
rect 343126 622480 343186 622580
rect 342000 622356 343186 622480
rect 342000 622256 342130 622356
rect 342230 622256 342354 622356
rect 342454 622256 342578 622356
rect 342678 622256 342802 622356
rect 342902 622256 343026 622356
rect 343126 622256 343186 622356
rect 342000 622132 343186 622256
rect 342000 622032 342130 622132
rect 342230 622032 342354 622132
rect 342454 622032 342578 622132
rect 342678 622032 342802 622132
rect 342902 622032 343026 622132
rect 343126 622032 343186 622132
rect 342000 621908 343186 622032
rect 342000 621808 342130 621908
rect 342230 621808 342354 621908
rect 342454 621808 342578 621908
rect 342678 621808 342802 621908
rect 342902 621808 343026 621908
rect 343126 621808 343186 621908
rect 342000 621684 343186 621808
rect 342000 621584 342130 621684
rect 342230 621584 342354 621684
rect 342454 621584 342578 621684
rect 342678 621584 342802 621684
rect 342902 621584 343026 621684
rect 343126 621584 343186 621684
rect 342000 621460 343186 621584
rect 342000 621360 342130 621460
rect 342230 621360 342354 621460
rect 342454 621360 342578 621460
rect 342678 621360 342802 621460
rect 342902 621360 343026 621460
rect 343126 621360 343186 621460
rect 342000 621236 343186 621360
rect 342000 621136 342130 621236
rect 342230 621136 342354 621236
rect 342454 621136 342578 621236
rect 342678 621136 342802 621236
rect 342902 621136 343026 621236
rect 343126 621136 343186 621236
rect 342000 621012 343186 621136
rect 342000 620912 342130 621012
rect 342230 620912 342354 621012
rect 342454 620912 342578 621012
rect 342678 620912 342802 621012
rect 342902 620912 343026 621012
rect 343126 620912 343186 621012
rect 342000 620788 343186 620912
rect 342000 620688 342130 620788
rect 342230 620688 342354 620788
rect 342454 620688 342578 620788
rect 342678 620688 342802 620788
rect 342902 620688 343026 620788
rect 343126 620688 343186 620788
rect 342000 620564 343186 620688
rect 342000 620464 342130 620564
rect 342230 620464 342354 620564
rect 342454 620464 342578 620564
rect 342678 620464 342802 620564
rect 342902 620464 343026 620564
rect 343126 620464 343186 620564
rect 342000 620340 343186 620464
rect 342000 620240 342130 620340
rect 342230 620240 342354 620340
rect 342454 620240 342578 620340
rect 342678 620240 342802 620340
rect 342902 620240 343026 620340
rect 343126 620240 343186 620340
rect 342000 620116 343186 620240
rect 342000 620016 342130 620116
rect 342230 620016 342354 620116
rect 342454 620016 342578 620116
rect 342678 620016 342802 620116
rect 342902 620016 343026 620116
rect 343126 620016 343186 620116
rect 342000 619892 343186 620016
rect 342000 619792 342130 619892
rect 342230 619792 342354 619892
rect 342454 619792 342578 619892
rect 342678 619792 342802 619892
rect 342902 619792 343026 619892
rect 343126 619792 343186 619892
rect 342000 619668 343186 619792
rect 342000 619568 342130 619668
rect 342230 619568 342354 619668
rect 342454 619568 342578 619668
rect 342678 619568 342802 619668
rect 342902 619568 343026 619668
rect 343126 619568 343186 619668
rect 342000 619444 343186 619568
rect 342000 619344 342130 619444
rect 342230 619344 342354 619444
rect 342454 619344 342578 619444
rect 342678 619344 342802 619444
rect 342902 619344 343026 619444
rect 343126 619344 343186 619444
rect 342000 619220 343186 619344
rect 342000 619120 342130 619220
rect 342230 619120 342354 619220
rect 342454 619120 342578 619220
rect 342678 619120 342802 619220
rect 342902 619120 343026 619220
rect 343126 619120 343186 619220
rect 342000 618996 343186 619120
rect 342000 618896 342130 618996
rect 342230 618896 342354 618996
rect 342454 618896 342578 618996
rect 342678 618896 342802 618996
rect 342902 618896 343026 618996
rect 343126 618896 343186 618996
rect 342000 618772 343186 618896
rect 342000 618672 342130 618772
rect 342230 618672 342354 618772
rect 342454 618672 342578 618772
rect 342678 618672 342802 618772
rect 342902 618672 343026 618772
rect 343126 618672 343186 618772
rect 342000 618548 343186 618672
rect 342000 618448 342130 618548
rect 342230 618448 342354 618548
rect 342454 618448 342578 618548
rect 342678 618448 342802 618548
rect 342902 618448 343026 618548
rect 343126 618448 343186 618548
rect 342000 618324 343186 618448
rect 342000 618224 342130 618324
rect 342230 618224 342354 618324
rect 342454 618224 342578 618324
rect 342678 618224 342802 618324
rect 342902 618224 343026 618324
rect 343126 618224 343186 618324
rect 342000 618100 343186 618224
rect 342000 618000 342130 618100
rect 342230 618000 342354 618100
rect 342454 618000 342578 618100
rect 342678 618000 342802 618100
rect 342902 618000 343026 618100
rect 343126 618000 343186 618100
rect 342000 617944 343186 618000
rect 510602 624161 515394 624606
rect 515386 618417 515394 624161
rect 510602 617944 515394 618417
rect 288920 605020 289920 610764
rect 294704 605020 295576 610764
rect 288920 604520 295576 605020
rect 298820 615474 315960 615520
rect 298820 615374 298876 615474
rect 298976 615374 299100 615474
rect 299200 615374 299324 615474
rect 299424 615374 299548 615474
rect 299648 615374 299772 615474
rect 299872 615374 299996 615474
rect 300096 615374 300220 615474
rect 300320 615374 300444 615474
rect 300544 615374 300668 615474
rect 300768 615374 300892 615474
rect 300992 615374 301116 615474
rect 301216 615374 301340 615474
rect 301440 615374 301564 615474
rect 301664 615374 301788 615474
rect 301888 615374 302012 615474
rect 302112 615374 302236 615474
rect 302336 615374 302460 615474
rect 302560 615374 302684 615474
rect 302784 615374 302908 615474
rect 303008 615374 303132 615474
rect 303232 615374 303356 615474
rect 303456 615374 303580 615474
rect 303680 615374 303804 615474
rect 303904 615374 304028 615474
rect 304128 615374 304252 615474
rect 304352 615374 304476 615474
rect 304576 615374 304700 615474
rect 304800 615374 304924 615474
rect 305024 615374 305148 615474
rect 305248 615374 305372 615474
rect 305472 615374 309346 615474
rect 309446 615374 309570 615474
rect 309670 615374 309794 615474
rect 309894 615374 310018 615474
rect 310118 615374 310242 615474
rect 310342 615374 310466 615474
rect 310566 615374 310690 615474
rect 310790 615374 310914 615474
rect 311014 615374 311138 615474
rect 311238 615374 311362 615474
rect 311462 615374 311586 615474
rect 311686 615374 311810 615474
rect 311910 615374 312034 615474
rect 312134 615374 312258 615474
rect 312358 615374 312482 615474
rect 312582 615374 312706 615474
rect 312806 615374 312930 615474
rect 313030 615374 313154 615474
rect 313254 615374 313378 615474
rect 313478 615374 313602 615474
rect 313702 615374 313826 615474
rect 313926 615374 314050 615474
rect 314150 615374 314274 615474
rect 314374 615374 314498 615474
rect 314598 615374 314722 615474
rect 314822 615374 314946 615474
rect 315046 615374 315170 615474
rect 315270 615374 315394 615474
rect 315494 615374 315618 615474
rect 315718 615374 315842 615474
rect 315942 615374 315960 615474
rect 298820 615250 315960 615374
rect 298820 615150 298876 615250
rect 298976 615150 299100 615250
rect 299200 615150 299324 615250
rect 299424 615150 299548 615250
rect 299648 615150 299772 615250
rect 299872 615150 299996 615250
rect 300096 615150 300220 615250
rect 300320 615150 300444 615250
rect 300544 615150 300668 615250
rect 300768 615150 300892 615250
rect 300992 615150 301116 615250
rect 301216 615150 301340 615250
rect 301440 615150 301564 615250
rect 301664 615150 301788 615250
rect 301888 615150 302012 615250
rect 302112 615150 302236 615250
rect 302336 615150 302460 615250
rect 302560 615150 302684 615250
rect 302784 615150 302908 615250
rect 303008 615150 303132 615250
rect 303232 615150 303356 615250
rect 303456 615150 303580 615250
rect 303680 615150 303804 615250
rect 303904 615150 304028 615250
rect 304128 615150 304252 615250
rect 304352 615150 304476 615250
rect 304576 615150 304700 615250
rect 304800 615150 304924 615250
rect 305024 615150 305148 615250
rect 305248 615150 305372 615250
rect 305472 615150 309346 615250
rect 309446 615150 309570 615250
rect 309670 615150 309794 615250
rect 309894 615150 310018 615250
rect 310118 615150 310242 615250
rect 310342 615150 310466 615250
rect 310566 615150 310690 615250
rect 310790 615150 310914 615250
rect 311014 615150 311138 615250
rect 311238 615150 311362 615250
rect 311462 615150 311586 615250
rect 311686 615150 311810 615250
rect 311910 615150 312034 615250
rect 312134 615150 312258 615250
rect 312358 615150 312482 615250
rect 312582 615150 312706 615250
rect 312806 615150 312930 615250
rect 313030 615150 313154 615250
rect 313254 615150 313378 615250
rect 313478 615150 313602 615250
rect 313702 615150 313826 615250
rect 313926 615150 314050 615250
rect 314150 615150 314274 615250
rect 314374 615150 314498 615250
rect 314598 615150 314722 615250
rect 314822 615150 314946 615250
rect 315046 615150 315170 615250
rect 315270 615150 315394 615250
rect 315494 615150 315618 615250
rect 315718 615150 315842 615250
rect 315942 615150 315960 615250
rect 298820 615026 315960 615150
rect 298820 614926 298876 615026
rect 298976 614926 299100 615026
rect 299200 614926 299324 615026
rect 299424 614926 299548 615026
rect 299648 614926 299772 615026
rect 299872 614926 299996 615026
rect 300096 614926 300220 615026
rect 300320 614926 300444 615026
rect 300544 614926 300668 615026
rect 300768 614926 300892 615026
rect 300992 614926 301116 615026
rect 301216 614926 301340 615026
rect 301440 614926 301564 615026
rect 301664 614926 301788 615026
rect 301888 614926 302012 615026
rect 302112 614926 302236 615026
rect 302336 614926 302460 615026
rect 302560 614926 302684 615026
rect 302784 614926 302908 615026
rect 303008 614926 303132 615026
rect 303232 614926 303356 615026
rect 303456 614926 303580 615026
rect 303680 614926 303804 615026
rect 303904 614926 304028 615026
rect 304128 614926 304252 615026
rect 304352 614926 304476 615026
rect 304576 614926 304700 615026
rect 304800 614926 304924 615026
rect 305024 614926 305148 615026
rect 305248 614926 305372 615026
rect 305472 614926 309346 615026
rect 309446 614926 309570 615026
rect 309670 614926 309794 615026
rect 309894 614926 310018 615026
rect 310118 614926 310242 615026
rect 310342 614926 310466 615026
rect 310566 614926 310690 615026
rect 310790 614926 310914 615026
rect 311014 614926 311138 615026
rect 311238 614926 311362 615026
rect 311462 614926 311586 615026
rect 311686 614926 311810 615026
rect 311910 614926 312034 615026
rect 312134 614926 312258 615026
rect 312358 614926 312482 615026
rect 312582 614926 312706 615026
rect 312806 614926 312930 615026
rect 313030 614926 313154 615026
rect 313254 614926 313378 615026
rect 313478 614926 313602 615026
rect 313702 614926 313826 615026
rect 313926 614926 314050 615026
rect 314150 614926 314274 615026
rect 314374 614926 314498 615026
rect 314598 614926 314722 615026
rect 314822 614926 314946 615026
rect 315046 614926 315170 615026
rect 315270 614926 315394 615026
rect 315494 614926 315618 615026
rect 315718 614926 315842 615026
rect 315942 614926 315960 615026
rect 298820 614802 315960 614926
rect 298820 614702 298876 614802
rect 298976 614702 299100 614802
rect 299200 614702 299324 614802
rect 299424 614702 299548 614802
rect 299648 614702 299772 614802
rect 299872 614702 299996 614802
rect 300096 614702 300220 614802
rect 300320 614702 300444 614802
rect 300544 614702 300668 614802
rect 300768 614702 300892 614802
rect 300992 614702 301116 614802
rect 301216 614702 301340 614802
rect 301440 614702 301564 614802
rect 301664 614702 301788 614802
rect 301888 614702 302012 614802
rect 302112 614702 302236 614802
rect 302336 614702 302460 614802
rect 302560 614702 302684 614802
rect 302784 614702 302908 614802
rect 303008 614702 303132 614802
rect 303232 614702 303356 614802
rect 303456 614702 303580 614802
rect 303680 614702 303804 614802
rect 303904 614702 304028 614802
rect 304128 614702 304252 614802
rect 304352 614702 304476 614802
rect 304576 614702 304700 614802
rect 304800 614702 304924 614802
rect 305024 614702 305148 614802
rect 305248 614702 305372 614802
rect 305472 614702 309346 614802
rect 309446 614702 309570 614802
rect 309670 614702 309794 614802
rect 309894 614702 310018 614802
rect 310118 614702 310242 614802
rect 310342 614702 310466 614802
rect 310566 614702 310690 614802
rect 310790 614702 310914 614802
rect 311014 614702 311138 614802
rect 311238 614702 311362 614802
rect 311462 614702 311586 614802
rect 311686 614702 311810 614802
rect 311910 614702 312034 614802
rect 312134 614702 312258 614802
rect 312358 614702 312482 614802
rect 312582 614702 312706 614802
rect 312806 614702 312930 614802
rect 313030 614702 313154 614802
rect 313254 614702 313378 614802
rect 313478 614702 313602 614802
rect 313702 614702 313826 614802
rect 313926 614702 314050 614802
rect 314150 614702 314274 614802
rect 314374 614702 314498 614802
rect 314598 614702 314722 614802
rect 314822 614702 314946 614802
rect 315046 614702 315170 614802
rect 315270 614702 315394 614802
rect 315494 614702 315618 614802
rect 315718 614702 315842 614802
rect 315942 614702 315960 614802
rect 298820 614578 315960 614702
rect 298820 614478 298876 614578
rect 298976 614478 299100 614578
rect 299200 614478 299324 614578
rect 299424 614478 299548 614578
rect 299648 614478 299772 614578
rect 299872 614478 299996 614578
rect 300096 614478 300220 614578
rect 300320 614478 300444 614578
rect 300544 614478 300668 614578
rect 300768 614478 300892 614578
rect 300992 614478 301116 614578
rect 301216 614478 301340 614578
rect 301440 614478 301564 614578
rect 301664 614478 301788 614578
rect 301888 614478 302012 614578
rect 302112 614478 302236 614578
rect 302336 614478 302460 614578
rect 302560 614478 302684 614578
rect 302784 614478 302908 614578
rect 303008 614478 303132 614578
rect 303232 614478 303356 614578
rect 303456 614478 303580 614578
rect 303680 614478 303804 614578
rect 303904 614478 304028 614578
rect 304128 614478 304252 614578
rect 304352 614478 304476 614578
rect 304576 614478 304700 614578
rect 304800 614478 304924 614578
rect 305024 614478 305148 614578
rect 305248 614478 305372 614578
rect 305472 614478 309346 614578
rect 309446 614478 309570 614578
rect 309670 614478 309794 614578
rect 309894 614478 310018 614578
rect 310118 614478 310242 614578
rect 310342 614478 310466 614578
rect 310566 614478 310690 614578
rect 310790 614478 310914 614578
rect 311014 614478 311138 614578
rect 311238 614478 311362 614578
rect 311462 614478 311586 614578
rect 311686 614478 311810 614578
rect 311910 614478 312034 614578
rect 312134 614478 312258 614578
rect 312358 614478 312482 614578
rect 312582 614478 312706 614578
rect 312806 614478 312930 614578
rect 313030 614478 313154 614578
rect 313254 614478 313378 614578
rect 313478 614478 313602 614578
rect 313702 614478 313826 614578
rect 313926 614478 314050 614578
rect 314150 614478 314274 614578
rect 314374 614478 314498 614578
rect 314598 614478 314722 614578
rect 314822 614478 314946 614578
rect 315046 614478 315170 614578
rect 315270 614478 315394 614578
rect 315494 614478 315618 614578
rect 315718 614478 315842 614578
rect 315942 614478 315960 614578
rect 298820 613100 315960 614478
rect 298820 611080 315980 613100
rect 298820 605336 298920 611080
rect 303704 605336 304920 611080
rect 309704 605336 310920 611080
rect 315704 605336 315980 611080
rect 298820 604520 315980 605336
rect 316960 597324 330680 616840
rect 335560 615494 342400 615540
rect 335560 615394 335616 615494
rect 335716 615394 335840 615494
rect 335940 615394 336064 615494
rect 336164 615394 336288 615494
rect 336388 615394 336512 615494
rect 336612 615394 336736 615494
rect 336836 615394 336960 615494
rect 337060 615394 337184 615494
rect 337284 615394 337408 615494
rect 337508 615394 337632 615494
rect 337732 615394 337856 615494
rect 337956 615394 338080 615494
rect 338180 615394 338304 615494
rect 338404 615394 338528 615494
rect 338628 615394 338752 615494
rect 338852 615394 338976 615494
rect 339076 615394 339200 615494
rect 339300 615394 339424 615494
rect 339524 615394 339648 615494
rect 339748 615394 339872 615494
rect 339972 615394 340096 615494
rect 340196 615394 340320 615494
rect 340420 615394 340544 615494
rect 340644 615394 340768 615494
rect 340868 615394 340992 615494
rect 341092 615394 341216 615494
rect 341316 615394 341440 615494
rect 341540 615394 341664 615494
rect 341764 615394 341888 615494
rect 341988 615394 342112 615494
rect 342212 615394 342400 615494
rect 335560 615270 342400 615394
rect 335560 615170 335616 615270
rect 335716 615170 335840 615270
rect 335940 615170 336064 615270
rect 336164 615170 336288 615270
rect 336388 615170 336512 615270
rect 336612 615170 336736 615270
rect 336836 615170 336960 615270
rect 337060 615170 337184 615270
rect 337284 615170 337408 615270
rect 337508 615170 337632 615270
rect 337732 615170 337856 615270
rect 337956 615170 338080 615270
rect 338180 615170 338304 615270
rect 338404 615170 338528 615270
rect 338628 615170 338752 615270
rect 338852 615170 338976 615270
rect 339076 615170 339200 615270
rect 339300 615170 339424 615270
rect 339524 615170 339648 615270
rect 339748 615170 339872 615270
rect 339972 615170 340096 615270
rect 340196 615170 340320 615270
rect 340420 615170 340544 615270
rect 340644 615170 340768 615270
rect 340868 615170 340992 615270
rect 341092 615170 341216 615270
rect 341316 615170 341440 615270
rect 341540 615170 341664 615270
rect 341764 615170 341888 615270
rect 341988 615170 342112 615270
rect 342212 615170 342400 615270
rect 335560 615046 342400 615170
rect 335560 614946 335616 615046
rect 335716 614946 335840 615046
rect 335940 614946 336064 615046
rect 336164 614946 336288 615046
rect 336388 614946 336512 615046
rect 336612 614946 336736 615046
rect 336836 614946 336960 615046
rect 337060 614946 337184 615046
rect 337284 614946 337408 615046
rect 337508 614946 337632 615046
rect 337732 614946 337856 615046
rect 337956 614946 338080 615046
rect 338180 614946 338304 615046
rect 338404 614946 338528 615046
rect 338628 614946 338752 615046
rect 338852 614946 338976 615046
rect 339076 614946 339200 615046
rect 339300 614946 339424 615046
rect 339524 614946 339648 615046
rect 339748 614946 339872 615046
rect 339972 614946 340096 615046
rect 340196 614946 340320 615046
rect 340420 614946 340544 615046
rect 340644 614946 340768 615046
rect 340868 614946 340992 615046
rect 341092 614946 341216 615046
rect 341316 614946 341440 615046
rect 341540 614946 341664 615046
rect 341764 614946 341888 615046
rect 341988 614946 342112 615046
rect 342212 614946 342400 615046
rect 335560 614822 342400 614946
rect 335560 614722 335616 614822
rect 335716 614722 335840 614822
rect 335940 614722 336064 614822
rect 336164 614722 336288 614822
rect 336388 614722 336512 614822
rect 336612 614722 336736 614822
rect 336836 614722 336960 614822
rect 337060 614722 337184 614822
rect 337284 614722 337408 614822
rect 337508 614722 337632 614822
rect 337732 614722 337856 614822
rect 337956 614722 338080 614822
rect 338180 614722 338304 614822
rect 338404 614722 338528 614822
rect 338628 614722 338752 614822
rect 338852 614722 338976 614822
rect 339076 614722 339200 614822
rect 339300 614722 339424 614822
rect 339524 614722 339648 614822
rect 339748 614722 339872 614822
rect 339972 614722 340096 614822
rect 340196 614722 340320 614822
rect 340420 614722 340544 614822
rect 340644 614722 340768 614822
rect 340868 614722 340992 614822
rect 341092 614722 341216 614822
rect 341316 614722 341440 614822
rect 341540 614722 341664 614822
rect 341764 614722 341888 614822
rect 341988 614722 342112 614822
rect 342212 614722 342400 614822
rect 335560 614598 342400 614722
rect 335560 614498 335616 614598
rect 335716 614498 335840 614598
rect 335940 614498 336064 614598
rect 336164 614498 336288 614598
rect 336388 614498 336512 614598
rect 336612 614498 336736 614598
rect 336836 614498 336960 614598
rect 337060 614498 337184 614598
rect 337284 614498 337408 614598
rect 337508 614498 337632 614598
rect 337732 614498 337856 614598
rect 337956 614498 338080 614598
rect 338180 614498 338304 614598
rect 338404 614498 338528 614598
rect 338628 614498 338752 614598
rect 338852 614498 338976 614598
rect 339076 614498 339200 614598
rect 339300 614498 339424 614598
rect 339524 614498 339648 614598
rect 339748 614498 339872 614598
rect 339972 614498 340096 614598
rect 340196 614498 340320 614598
rect 340420 614498 340544 614598
rect 340644 614498 340768 614598
rect 340868 614498 340992 614598
rect 341092 614498 341216 614598
rect 341316 614498 341440 614598
rect 341540 614498 341664 614598
rect 341764 614498 341888 614598
rect 341988 614498 342112 614598
rect 342212 614498 342400 614598
rect 335560 614464 342400 614498
rect 335580 611084 342400 614464
rect 510594 611200 515394 617944
rect 335580 605340 336480 611084
rect 341264 605340 342400 611084
rect 335580 604720 342400 605340
rect 510602 610761 515394 611200
rect 515386 605017 515394 610761
rect 510602 604544 515394 605017
rect 520594 690560 525394 704800
rect 566594 702300 571594 704800
rect 520594 684336 520602 690560
rect 525386 684336 525394 690560
rect 520594 650961 525394 684336
rect 582300 677984 584800 682984
rect 520594 645217 520602 650961
rect 525386 645217 525394 650961
rect 520594 637561 525394 645217
rect 560050 644576 584800 644584
rect 560050 639792 560582 644576
rect 566726 639792 584800 644576
rect 560050 639784 584800 639792
rect 520594 631817 520602 637561
rect 525386 631817 525394 637561
rect 520594 624161 525394 631817
rect 560050 634576 584800 634584
rect 560050 629792 560582 634576
rect 566726 629792 584800 634576
rect 560050 629784 584800 629792
rect 520594 618417 520602 624161
rect 525386 618417 525394 624161
rect 520594 610761 525394 618417
rect 520594 605017 520602 610761
rect 525386 605017 525394 610761
rect 520594 604544 525394 605017
rect 316960 591580 317480 597324
rect 322264 591580 325480 597324
rect 330264 591580 330680 597324
rect 316960 591080 330680 591580
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 339960 511642 340072 571500
rect -800 511530 340072 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect 340967 463692 341079 571500
rect -800 463580 341079 463692
rect -800 462486 17711 462510
rect -800 462422 13897 462486
rect 13961 462422 13977 462486
rect 14041 462422 14057 462486
rect 14121 462422 14137 462486
rect 14201 462422 14217 462486
rect 14281 462422 14297 462486
rect 14361 462422 14377 462486
rect 14441 462422 14457 462486
rect 14521 462422 14537 462486
rect 14601 462422 14617 462486
rect 14681 462422 14697 462486
rect 14761 462422 14777 462486
rect 14841 462422 14857 462486
rect 14921 462422 14937 462486
rect 15001 462422 15017 462486
rect 15081 462422 15097 462486
rect 15161 462422 15177 462486
rect 15241 462422 15257 462486
rect 15321 462422 15337 462486
rect 15401 462422 15417 462486
rect 15481 462422 15497 462486
rect 15561 462422 15577 462486
rect 15641 462422 15657 462486
rect 15721 462422 15737 462486
rect 15801 462422 15817 462486
rect 15881 462422 15897 462486
rect 15961 462422 15977 462486
rect 16041 462422 16057 462486
rect 16121 462422 16137 462486
rect 16201 462422 16217 462486
rect 16281 462422 16297 462486
rect 16361 462422 16377 462486
rect 16441 462422 16457 462486
rect 16521 462422 16537 462486
rect 16601 462422 16617 462486
rect 16681 462422 16697 462486
rect 16761 462422 16777 462486
rect 16841 462422 16857 462486
rect 16921 462422 16937 462486
rect 17001 462422 17017 462486
rect 17081 462422 17097 462486
rect 17161 462422 17177 462486
rect 17241 462422 17257 462486
rect 17321 462422 17337 462486
rect 17401 462422 17417 462486
rect 17481 462422 17497 462486
rect 17561 462422 17711 462486
rect -800 462398 17711 462422
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect 341738 420470 341850 571500
rect -800 420358 341850 420470
rect -800 419264 17694 419288
rect -800 419200 13911 419264
rect 13975 419200 13991 419264
rect 14055 419200 14071 419264
rect 14135 419200 14151 419264
rect 14215 419200 14231 419264
rect 14295 419200 14311 419264
rect 14375 419200 14391 419264
rect 14455 419200 14471 419264
rect 14535 419200 14551 419264
rect 14615 419200 14631 419264
rect 14695 419200 14711 419264
rect 14775 419200 14791 419264
rect 14855 419200 14871 419264
rect 14935 419200 14951 419264
rect 15015 419200 15031 419264
rect 15095 419200 15111 419264
rect 15175 419200 15191 419264
rect 15255 419200 15271 419264
rect 15335 419200 15351 419264
rect 15415 419200 15431 419264
rect 15495 419200 15511 419264
rect 15575 419200 15591 419264
rect 15655 419200 15671 419264
rect 15735 419200 15751 419264
rect 15815 419200 15831 419264
rect 15895 419200 15911 419264
rect 15975 419200 15991 419264
rect 16055 419200 16071 419264
rect 16135 419200 16151 419264
rect 16215 419200 16231 419264
rect 16295 419200 16311 419264
rect 16375 419200 16391 419264
rect 16455 419200 16471 419264
rect 16535 419200 16551 419264
rect 16615 419200 16631 419264
rect 16695 419200 16711 419264
rect 16775 419200 16791 419264
rect 16855 419200 16871 419264
rect 16935 419200 16951 419264
rect 17015 419200 17031 419264
rect 17095 419200 17111 419264
rect 17175 419200 17191 419264
rect 17255 419200 17271 419264
rect 17335 419200 17351 419264
rect 17415 419200 17431 419264
rect 17495 419200 17511 419264
rect 17575 419200 17694 419264
rect -800 419176 17694 419200
rect 533497 405408 533609 573580
rect 537376 454558 537488 573580
rect 539494 498980 539606 573580
rect 555452 555354 584800 555362
rect 555452 550570 556255 555354
rect 562319 550570 584800 555354
rect 555452 550562 584800 550570
rect 555452 545354 584800 545362
rect 555452 540570 556255 545354
rect 562319 540570 584800 545354
rect 555452 540562 584800 540570
rect 573371 500138 584800 500162
rect 573371 500074 573553 500138
rect 573617 500074 573633 500138
rect 573697 500074 573713 500138
rect 573777 500074 573793 500138
rect 573857 500074 573873 500138
rect 573937 500074 573953 500138
rect 574017 500074 574033 500138
rect 574097 500074 574113 500138
rect 574177 500074 574193 500138
rect 574257 500074 574273 500138
rect 574337 500074 574353 500138
rect 574417 500074 574433 500138
rect 574497 500074 574513 500138
rect 574577 500074 574593 500138
rect 574657 500074 574673 500138
rect 574737 500074 574753 500138
rect 574817 500074 574833 500138
rect 574897 500074 574913 500138
rect 574977 500074 574993 500138
rect 575057 500074 575073 500138
rect 575137 500074 575153 500138
rect 575217 500074 575233 500138
rect 575297 500074 575313 500138
rect 575377 500074 575393 500138
rect 575457 500074 575473 500138
rect 575537 500074 575553 500138
rect 575617 500074 575633 500138
rect 575697 500074 575713 500138
rect 575777 500074 575793 500138
rect 575857 500074 575873 500138
rect 575937 500074 575953 500138
rect 576017 500074 576033 500138
rect 576097 500074 576113 500138
rect 576177 500074 576193 500138
rect 576257 500074 576273 500138
rect 576337 500074 576353 500138
rect 576417 500074 576433 500138
rect 576497 500074 576513 500138
rect 576577 500074 576593 500138
rect 576657 500074 576673 500138
rect 576737 500074 584800 500138
rect 573371 500050 584800 500074
rect 539494 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 573405 455716 584800 455740
rect 573405 455652 573591 455716
rect 573655 455652 573671 455716
rect 573735 455652 573751 455716
rect 573815 455652 573831 455716
rect 573895 455652 573911 455716
rect 573975 455652 573991 455716
rect 574055 455652 574071 455716
rect 574135 455652 574151 455716
rect 574215 455652 574231 455716
rect 574295 455652 574311 455716
rect 574375 455652 574391 455716
rect 574455 455652 574471 455716
rect 574535 455652 574551 455716
rect 574615 455652 574631 455716
rect 574695 455652 574711 455716
rect 574775 455652 574791 455716
rect 574855 455652 574871 455716
rect 574935 455652 574951 455716
rect 575015 455652 575031 455716
rect 575095 455652 575111 455716
rect 575175 455652 575191 455716
rect 575255 455652 575271 455716
rect 575335 455652 575351 455716
rect 575415 455652 575431 455716
rect 575495 455652 575511 455716
rect 575575 455652 575591 455716
rect 575655 455652 575671 455716
rect 575735 455652 575751 455716
rect 575815 455652 575831 455716
rect 575895 455652 575911 455716
rect 575975 455652 575991 455716
rect 576055 455652 576071 455716
rect 576135 455652 576151 455716
rect 576215 455652 576231 455716
rect 576295 455652 576311 455716
rect 576375 455652 576391 455716
rect 576455 455652 576471 455716
rect 576535 455652 576551 455716
rect 576615 455652 576631 455716
rect 576695 455652 584800 455716
rect 573405 455628 584800 455652
rect 537376 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 533497 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 13406 196222 584800 196230
rect 13406 191438 13997 196222
rect 17421 191438 573605 196222
rect 576629 191438 584800 196222
rect 13406 191430 584800 191438
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 170922 684353 173066 690577
rect 173422 684353 175566 690577
rect 222622 684386 224766 690610
rect 217344 626112 217408 626176
rect 217472 626112 217536 626176
rect 217600 626112 217664 626176
rect 217728 626112 217792 626176
rect 217856 626112 217920 626176
rect 217984 626112 218048 626176
rect 218112 626112 218176 626176
rect 218240 626112 218304 626176
rect 218368 626112 218432 626176
rect 218496 626112 218560 626176
rect 218624 626112 218688 626176
rect 218752 626112 218816 626176
rect 218880 626112 218944 626176
rect 219008 626112 219072 626176
rect 219136 626112 219200 626176
rect 219264 626112 219328 626176
rect 219392 626112 219456 626176
rect 219520 626112 219584 626176
rect 219648 626112 219712 626176
rect 219776 626112 219840 626176
rect 219904 626112 219968 626176
rect 220032 626112 220096 626176
rect 220160 626112 220224 626176
rect 220288 626112 220352 626176
rect 220416 626112 220480 626176
rect 220544 626112 220608 626176
rect 220672 626112 220736 626176
rect 220800 626112 220864 626176
rect 220928 626112 220992 626176
rect 221056 626112 221120 626176
rect 221184 626112 221248 626176
rect 221312 626112 221376 626176
rect 221440 626112 221504 626176
rect 221568 626112 221632 626176
rect 221696 626112 221760 626176
rect 221824 626112 221888 626176
rect 221952 626112 222016 626176
rect 222080 626112 222144 626176
rect 217344 625984 217408 626048
rect 217472 625984 217536 626048
rect 217600 625984 217664 626048
rect 217728 625984 217792 626048
rect 217856 625984 217920 626048
rect 217984 625984 218048 626048
rect 218112 625984 218176 626048
rect 218240 625984 218304 626048
rect 218368 625984 218432 626048
rect 218496 625984 218560 626048
rect 218624 625984 218688 626048
rect 218752 625984 218816 626048
rect 218880 625984 218944 626048
rect 219008 625984 219072 626048
rect 219136 625984 219200 626048
rect 219264 625984 219328 626048
rect 219392 625984 219456 626048
rect 219520 625984 219584 626048
rect 219648 625984 219712 626048
rect 219776 625984 219840 626048
rect 219904 625984 219968 626048
rect 220032 625984 220096 626048
rect 220160 625984 220224 626048
rect 220288 625984 220352 626048
rect 220416 625984 220480 626048
rect 220544 625984 220608 626048
rect 220672 625984 220736 626048
rect 220800 625984 220864 626048
rect 220928 625984 220992 626048
rect 221056 625984 221120 626048
rect 221184 625984 221248 626048
rect 221312 625984 221376 626048
rect 221440 625984 221504 626048
rect 221568 625984 221632 626048
rect 221696 625984 221760 626048
rect 221824 625984 221888 626048
rect 221952 625984 222016 626048
rect 222080 625984 222144 626048
rect 217344 625856 217408 625920
rect 217472 625856 217536 625920
rect 217600 625856 217664 625920
rect 217728 625856 217792 625920
rect 217856 625856 217920 625920
rect 217984 625856 218048 625920
rect 218112 625856 218176 625920
rect 218240 625856 218304 625920
rect 218368 625856 218432 625920
rect 218496 625856 218560 625920
rect 218624 625856 218688 625920
rect 218752 625856 218816 625920
rect 218880 625856 218944 625920
rect 219008 625856 219072 625920
rect 219136 625856 219200 625920
rect 219264 625856 219328 625920
rect 219392 625856 219456 625920
rect 219520 625856 219584 625920
rect 219648 625856 219712 625920
rect 219776 625856 219840 625920
rect 219904 625856 219968 625920
rect 220032 625856 220096 625920
rect 220160 625856 220224 625920
rect 220288 625856 220352 625920
rect 220416 625856 220480 625920
rect 220544 625856 220608 625920
rect 220672 625856 220736 625920
rect 220800 625856 220864 625920
rect 220928 625856 220992 625920
rect 221056 625856 221120 625920
rect 221184 625856 221248 625920
rect 221312 625856 221376 625920
rect 221440 625856 221504 625920
rect 221568 625856 221632 625920
rect 221696 625856 221760 625920
rect 221824 625856 221888 625920
rect 221952 625856 222016 625920
rect 222080 625856 222144 625920
rect 217344 625728 217408 625792
rect 217472 625728 217536 625792
rect 217600 625728 217664 625792
rect 217728 625728 217792 625792
rect 217856 625728 217920 625792
rect 217984 625728 218048 625792
rect 218112 625728 218176 625792
rect 218240 625728 218304 625792
rect 218368 625728 218432 625792
rect 218496 625728 218560 625792
rect 218624 625728 218688 625792
rect 218752 625728 218816 625792
rect 218880 625728 218944 625792
rect 219008 625728 219072 625792
rect 219136 625728 219200 625792
rect 219264 625728 219328 625792
rect 219392 625728 219456 625792
rect 219520 625728 219584 625792
rect 219648 625728 219712 625792
rect 219776 625728 219840 625792
rect 219904 625728 219968 625792
rect 220032 625728 220096 625792
rect 220160 625728 220224 625792
rect 220288 625728 220352 625792
rect 220416 625728 220480 625792
rect 220544 625728 220608 625792
rect 220672 625728 220736 625792
rect 220800 625728 220864 625792
rect 220928 625728 220992 625792
rect 221056 625728 221120 625792
rect 221184 625728 221248 625792
rect 221312 625728 221376 625792
rect 221440 625728 221504 625792
rect 221568 625728 221632 625792
rect 221696 625728 221760 625792
rect 221824 625728 221888 625792
rect 221952 625728 222016 625792
rect 222080 625728 222144 625792
rect 227640 626112 227704 626176
rect 227768 626112 227832 626176
rect 227896 626112 227960 626176
rect 228024 626112 228088 626176
rect 228152 626112 228216 626176
rect 228280 626112 228344 626176
rect 228408 626112 228472 626176
rect 228536 626112 228600 626176
rect 228664 626112 228728 626176
rect 228792 626112 228856 626176
rect 228920 626112 228984 626176
rect 229048 626112 229112 626176
rect 229176 626112 229240 626176
rect 229304 626112 229368 626176
rect 229432 626112 229496 626176
rect 229560 626112 229624 626176
rect 229688 626112 229752 626176
rect 229816 626112 229880 626176
rect 229944 626112 230008 626176
rect 230072 626112 230136 626176
rect 230200 626112 230264 626176
rect 230328 626112 230392 626176
rect 230456 626112 230520 626176
rect 230584 626112 230648 626176
rect 230712 626112 230776 626176
rect 230840 626112 230904 626176
rect 230968 626112 231032 626176
rect 231096 626112 231160 626176
rect 231224 626112 231288 626176
rect 231352 626112 231416 626176
rect 231480 626112 231544 626176
rect 231608 626112 231672 626176
rect 231736 626112 231800 626176
rect 231864 626112 231928 626176
rect 231992 626112 232056 626176
rect 232120 626112 232184 626176
rect 232248 626112 232312 626176
rect 232376 626112 232440 626176
rect 227640 625984 227704 626048
rect 227768 625984 227832 626048
rect 227896 625984 227960 626048
rect 228024 625984 228088 626048
rect 228152 625984 228216 626048
rect 228280 625984 228344 626048
rect 228408 625984 228472 626048
rect 228536 625984 228600 626048
rect 228664 625984 228728 626048
rect 228792 625984 228856 626048
rect 228920 625984 228984 626048
rect 229048 625984 229112 626048
rect 229176 625984 229240 626048
rect 229304 625984 229368 626048
rect 229432 625984 229496 626048
rect 229560 625984 229624 626048
rect 229688 625984 229752 626048
rect 229816 625984 229880 626048
rect 229944 625984 230008 626048
rect 230072 625984 230136 626048
rect 230200 625984 230264 626048
rect 230328 625984 230392 626048
rect 230456 625984 230520 626048
rect 230584 625984 230648 626048
rect 230712 625984 230776 626048
rect 230840 625984 230904 626048
rect 230968 625984 231032 626048
rect 231096 625984 231160 626048
rect 231224 625984 231288 626048
rect 231352 625984 231416 626048
rect 231480 625984 231544 626048
rect 231608 625984 231672 626048
rect 231736 625984 231800 626048
rect 231864 625984 231928 626048
rect 231992 625984 232056 626048
rect 232120 625984 232184 626048
rect 232248 625984 232312 626048
rect 232376 625984 232440 626048
rect 227640 625856 227704 625920
rect 227768 625856 227832 625920
rect 227896 625856 227960 625920
rect 228024 625856 228088 625920
rect 228152 625856 228216 625920
rect 228280 625856 228344 625920
rect 228408 625856 228472 625920
rect 228536 625856 228600 625920
rect 228664 625856 228728 625920
rect 228792 625856 228856 625920
rect 228920 625856 228984 625920
rect 229048 625856 229112 625920
rect 229176 625856 229240 625920
rect 229304 625856 229368 625920
rect 229432 625856 229496 625920
rect 229560 625856 229624 625920
rect 229688 625856 229752 625920
rect 229816 625856 229880 625920
rect 229944 625856 230008 625920
rect 230072 625856 230136 625920
rect 230200 625856 230264 625920
rect 230328 625856 230392 625920
rect 230456 625856 230520 625920
rect 230584 625856 230648 625920
rect 230712 625856 230776 625920
rect 230840 625856 230904 625920
rect 230968 625856 231032 625920
rect 231096 625856 231160 625920
rect 231224 625856 231288 625920
rect 231352 625856 231416 625920
rect 231480 625856 231544 625920
rect 231608 625856 231672 625920
rect 231736 625856 231800 625920
rect 231864 625856 231928 625920
rect 231992 625856 232056 625920
rect 232120 625856 232184 625920
rect 232248 625856 232312 625920
rect 232376 625856 232440 625920
rect 227640 625728 227704 625792
rect 227768 625728 227832 625792
rect 227896 625728 227960 625792
rect 228024 625728 228088 625792
rect 228152 625728 228216 625792
rect 228280 625728 228344 625792
rect 228408 625728 228472 625792
rect 228536 625728 228600 625792
rect 228664 625728 228728 625792
rect 228792 625728 228856 625792
rect 228920 625728 228984 625792
rect 229048 625728 229112 625792
rect 229176 625728 229240 625792
rect 229304 625728 229368 625792
rect 229432 625728 229496 625792
rect 229560 625728 229624 625792
rect 229688 625728 229752 625792
rect 229816 625728 229880 625792
rect 229944 625728 230008 625792
rect 230072 625728 230136 625792
rect 230200 625728 230264 625792
rect 230328 625728 230392 625792
rect 230456 625728 230520 625792
rect 230584 625728 230648 625792
rect 230712 625728 230776 625792
rect 230840 625728 230904 625792
rect 230968 625728 231032 625792
rect 231096 625728 231160 625792
rect 231224 625728 231288 625792
rect 231352 625728 231416 625792
rect 231480 625728 231544 625792
rect 231608 625728 231672 625792
rect 231736 625728 231800 625792
rect 231864 625728 231928 625792
rect 231992 625728 232056 625792
rect 232120 625728 232184 625792
rect 232248 625728 232312 625792
rect 232376 625728 232440 625792
rect 289800 684340 294584 690084
rect 324322 684369 326466 690593
rect 510602 684336 515386 690560
rect 289920 644840 294704 650584
rect 298920 644840 303704 650584
rect 304920 644840 309704 650584
rect 310920 644840 315704 650584
rect 298876 642594 298976 642694
rect 299100 642594 299200 642694
rect 299324 642594 299424 642694
rect 299548 642594 299648 642694
rect 299772 642594 299872 642694
rect 299996 642594 300096 642694
rect 300220 642594 300320 642694
rect 300444 642594 300544 642694
rect 300668 642594 300768 642694
rect 300892 642594 300992 642694
rect 301116 642594 301216 642694
rect 301340 642594 301440 642694
rect 301564 642594 301664 642694
rect 301788 642594 301888 642694
rect 302012 642594 302112 642694
rect 302236 642594 302336 642694
rect 302460 642594 302560 642694
rect 302684 642594 302784 642694
rect 302908 642594 303008 642694
rect 303132 642594 303232 642694
rect 303356 642594 303456 642694
rect 303580 642594 303680 642694
rect 303804 642594 303904 642694
rect 304028 642594 304128 642694
rect 304252 642594 304352 642694
rect 304476 642594 304576 642694
rect 304700 642594 304800 642694
rect 304924 642594 305024 642694
rect 305148 642594 305248 642694
rect 305372 642594 305472 642694
rect 309346 642594 309446 642694
rect 309570 642594 309670 642694
rect 309794 642594 309894 642694
rect 310018 642594 310118 642694
rect 310242 642594 310342 642694
rect 310466 642594 310566 642694
rect 310690 642594 310790 642694
rect 310914 642594 311014 642694
rect 311138 642594 311238 642694
rect 311362 642594 311462 642694
rect 311586 642594 311686 642694
rect 311810 642594 311910 642694
rect 312034 642594 312134 642694
rect 312258 642594 312358 642694
rect 312482 642594 312582 642694
rect 312706 642594 312806 642694
rect 312930 642594 313030 642694
rect 313154 642594 313254 642694
rect 313378 642594 313478 642694
rect 313602 642594 313702 642694
rect 313826 642594 313926 642694
rect 314050 642594 314150 642694
rect 314274 642594 314374 642694
rect 314498 642594 314598 642694
rect 314722 642594 314822 642694
rect 314946 642594 315046 642694
rect 315170 642594 315270 642694
rect 315394 642594 315494 642694
rect 315618 642594 315718 642694
rect 315842 642594 315942 642694
rect 298876 642370 298976 642470
rect 299100 642370 299200 642470
rect 299324 642370 299424 642470
rect 299548 642370 299648 642470
rect 299772 642370 299872 642470
rect 299996 642370 300096 642470
rect 300220 642370 300320 642470
rect 300444 642370 300544 642470
rect 300668 642370 300768 642470
rect 300892 642370 300992 642470
rect 301116 642370 301216 642470
rect 301340 642370 301440 642470
rect 301564 642370 301664 642470
rect 301788 642370 301888 642470
rect 302012 642370 302112 642470
rect 302236 642370 302336 642470
rect 302460 642370 302560 642470
rect 302684 642370 302784 642470
rect 302908 642370 303008 642470
rect 303132 642370 303232 642470
rect 303356 642370 303456 642470
rect 303580 642370 303680 642470
rect 303804 642370 303904 642470
rect 304028 642370 304128 642470
rect 304252 642370 304352 642470
rect 304476 642370 304576 642470
rect 304700 642370 304800 642470
rect 304924 642370 305024 642470
rect 305148 642370 305248 642470
rect 305372 642370 305472 642470
rect 309346 642370 309446 642470
rect 309570 642370 309670 642470
rect 309794 642370 309894 642470
rect 310018 642370 310118 642470
rect 310242 642370 310342 642470
rect 310466 642370 310566 642470
rect 310690 642370 310790 642470
rect 310914 642370 311014 642470
rect 311138 642370 311238 642470
rect 311362 642370 311462 642470
rect 311586 642370 311686 642470
rect 311810 642370 311910 642470
rect 312034 642370 312134 642470
rect 312258 642370 312358 642470
rect 312482 642370 312582 642470
rect 312706 642370 312806 642470
rect 312930 642370 313030 642470
rect 313154 642370 313254 642470
rect 313378 642370 313478 642470
rect 313602 642370 313702 642470
rect 313826 642370 313926 642470
rect 314050 642370 314150 642470
rect 314274 642370 314374 642470
rect 314498 642370 314598 642470
rect 314722 642370 314822 642470
rect 314946 642370 315046 642470
rect 315170 642370 315270 642470
rect 315394 642370 315494 642470
rect 315618 642370 315718 642470
rect 315842 642370 315942 642470
rect 298876 642146 298976 642246
rect 299100 642146 299200 642246
rect 299324 642146 299424 642246
rect 299548 642146 299648 642246
rect 299772 642146 299872 642246
rect 299996 642146 300096 642246
rect 300220 642146 300320 642246
rect 300444 642146 300544 642246
rect 300668 642146 300768 642246
rect 300892 642146 300992 642246
rect 301116 642146 301216 642246
rect 301340 642146 301440 642246
rect 301564 642146 301664 642246
rect 301788 642146 301888 642246
rect 302012 642146 302112 642246
rect 302236 642146 302336 642246
rect 302460 642146 302560 642246
rect 302684 642146 302784 642246
rect 302908 642146 303008 642246
rect 303132 642146 303232 642246
rect 303356 642146 303456 642246
rect 303580 642146 303680 642246
rect 303804 642146 303904 642246
rect 304028 642146 304128 642246
rect 304252 642146 304352 642246
rect 304476 642146 304576 642246
rect 304700 642146 304800 642246
rect 304924 642146 305024 642246
rect 305148 642146 305248 642246
rect 305372 642146 305472 642246
rect 309346 642146 309446 642246
rect 309570 642146 309670 642246
rect 309794 642146 309894 642246
rect 310018 642146 310118 642246
rect 310242 642146 310342 642246
rect 310466 642146 310566 642246
rect 310690 642146 310790 642246
rect 310914 642146 311014 642246
rect 311138 642146 311238 642246
rect 311362 642146 311462 642246
rect 311586 642146 311686 642246
rect 311810 642146 311910 642246
rect 312034 642146 312134 642246
rect 312258 642146 312358 642246
rect 312482 642146 312582 642246
rect 312706 642146 312806 642246
rect 312930 642146 313030 642246
rect 313154 642146 313254 642246
rect 313378 642146 313478 642246
rect 313602 642146 313702 642246
rect 313826 642146 313926 642246
rect 314050 642146 314150 642246
rect 314274 642146 314374 642246
rect 314498 642146 314598 642246
rect 314722 642146 314822 642246
rect 314946 642146 315046 642246
rect 315170 642146 315270 642246
rect 315394 642146 315494 642246
rect 315618 642146 315718 642246
rect 315842 642146 315942 642246
rect 298876 641922 298976 642022
rect 299100 641922 299200 642022
rect 299324 641922 299424 642022
rect 299548 641922 299648 642022
rect 299772 641922 299872 642022
rect 299996 641922 300096 642022
rect 300220 641922 300320 642022
rect 300444 641922 300544 642022
rect 300668 641922 300768 642022
rect 300892 641922 300992 642022
rect 301116 641922 301216 642022
rect 301340 641922 301440 642022
rect 301564 641922 301664 642022
rect 301788 641922 301888 642022
rect 302012 641922 302112 642022
rect 302236 641922 302336 642022
rect 302460 641922 302560 642022
rect 302684 641922 302784 642022
rect 302908 641922 303008 642022
rect 303132 641922 303232 642022
rect 303356 641922 303456 642022
rect 303580 641922 303680 642022
rect 303804 641922 303904 642022
rect 304028 641922 304128 642022
rect 304252 641922 304352 642022
rect 304476 641922 304576 642022
rect 304700 641922 304800 642022
rect 304924 641922 305024 642022
rect 305148 641922 305248 642022
rect 305372 641922 305472 642022
rect 309346 641922 309446 642022
rect 309570 641922 309670 642022
rect 309794 641922 309894 642022
rect 310018 641922 310118 642022
rect 310242 641922 310342 642022
rect 310466 641922 310566 642022
rect 310690 641922 310790 642022
rect 310914 641922 311014 642022
rect 311138 641922 311238 642022
rect 311362 641922 311462 642022
rect 311586 641922 311686 642022
rect 311810 641922 311910 642022
rect 312034 641922 312134 642022
rect 312258 641922 312358 642022
rect 312482 641922 312582 642022
rect 312706 641922 312806 642022
rect 312930 641922 313030 642022
rect 313154 641922 313254 642022
rect 313378 641922 313478 642022
rect 313602 641922 313702 642022
rect 313826 641922 313926 642022
rect 314050 641922 314150 642022
rect 314274 641922 314374 642022
rect 314498 641922 314598 642022
rect 314722 641922 314822 642022
rect 314946 641922 315046 642022
rect 315170 641922 315270 642022
rect 315394 641922 315494 642022
rect 315618 641922 315718 642022
rect 315842 641922 315942 642022
rect 298876 641698 298976 641798
rect 299100 641698 299200 641798
rect 299324 641698 299424 641798
rect 299548 641698 299648 641798
rect 299772 641698 299872 641798
rect 299996 641698 300096 641798
rect 300220 641698 300320 641798
rect 300444 641698 300544 641798
rect 300668 641698 300768 641798
rect 300892 641698 300992 641798
rect 301116 641698 301216 641798
rect 301340 641698 301440 641798
rect 301564 641698 301664 641798
rect 301788 641698 301888 641798
rect 302012 641698 302112 641798
rect 302236 641698 302336 641798
rect 302460 641698 302560 641798
rect 302684 641698 302784 641798
rect 302908 641698 303008 641798
rect 303132 641698 303232 641798
rect 303356 641698 303456 641798
rect 303580 641698 303680 641798
rect 303804 641698 303904 641798
rect 304028 641698 304128 641798
rect 304252 641698 304352 641798
rect 304476 641698 304576 641798
rect 304700 641698 304800 641798
rect 304924 641698 305024 641798
rect 305148 641698 305248 641798
rect 305372 641698 305472 641798
rect 309346 641698 309446 641798
rect 309570 641698 309670 641798
rect 309794 641698 309894 641798
rect 310018 641698 310118 641798
rect 310242 641698 310342 641798
rect 310466 641698 310566 641798
rect 310690 641698 310790 641798
rect 310914 641698 311014 641798
rect 311138 641698 311238 641798
rect 311362 641698 311462 641798
rect 311586 641698 311686 641798
rect 311810 641698 311910 641798
rect 312034 641698 312134 641798
rect 312258 641698 312358 641798
rect 312482 641698 312582 641798
rect 312706 641698 312806 641798
rect 312930 641698 313030 641798
rect 313154 641698 313254 641798
rect 313378 641698 313478 641798
rect 313602 641698 313702 641798
rect 313826 641698 313926 641798
rect 314050 641698 314150 641798
rect 314274 641698 314374 641798
rect 314498 641698 314598 641798
rect 314722 641698 314822 641798
rect 314946 641698 315046 641798
rect 315170 641698 315270 641798
rect 315394 641698 315494 641798
rect 315618 641698 315718 641798
rect 315842 641698 315942 641798
rect 289920 631440 294704 637184
rect 297850 637896 297950 637996
rect 298074 637896 298174 637996
rect 298298 637896 298398 637996
rect 298522 637896 298622 637996
rect 298746 637896 298846 637996
rect 297850 637672 297950 637772
rect 298074 637672 298174 637772
rect 298298 637672 298398 637772
rect 298522 637672 298622 637772
rect 298746 637672 298846 637772
rect 297850 637448 297950 637548
rect 298074 637448 298174 637548
rect 298298 637448 298398 637548
rect 298522 637448 298622 637548
rect 298746 637448 298846 637548
rect 297850 637224 297950 637324
rect 298074 637224 298174 637324
rect 298298 637224 298398 637324
rect 298522 637224 298622 637324
rect 298746 637224 298846 637324
rect 297850 637000 297950 637100
rect 298074 637000 298174 637100
rect 298298 637000 298398 637100
rect 298522 637000 298622 637100
rect 298746 637000 298846 637100
rect 297850 636776 297950 636876
rect 298074 636776 298174 636876
rect 298298 636776 298398 636876
rect 298522 636776 298622 636876
rect 298746 636776 298846 636876
rect 297850 636552 297950 636652
rect 298074 636552 298174 636652
rect 298298 636552 298398 636652
rect 298522 636552 298622 636652
rect 298746 636552 298846 636652
rect 297850 636328 297950 636428
rect 298074 636328 298174 636428
rect 298298 636328 298398 636428
rect 298522 636328 298622 636428
rect 298746 636328 298846 636428
rect 297850 636104 297950 636204
rect 298074 636104 298174 636204
rect 298298 636104 298398 636204
rect 298522 636104 298622 636204
rect 298746 636104 298846 636204
rect 297850 635880 297950 635980
rect 298074 635880 298174 635980
rect 298298 635880 298398 635980
rect 298522 635880 298622 635980
rect 298746 635880 298846 635980
rect 297850 635656 297950 635756
rect 298074 635656 298174 635756
rect 298298 635656 298398 635756
rect 298522 635656 298622 635756
rect 298746 635656 298846 635756
rect 297850 635432 297950 635532
rect 298074 635432 298174 635532
rect 298298 635432 298398 635532
rect 298522 635432 298622 635532
rect 298746 635432 298846 635532
rect 297850 635208 297950 635308
rect 298074 635208 298174 635308
rect 298298 635208 298398 635308
rect 298522 635208 298622 635308
rect 298746 635208 298846 635308
rect 297850 634984 297950 635084
rect 298074 634984 298174 635084
rect 298298 634984 298398 635084
rect 298522 634984 298622 635084
rect 298746 634984 298846 635084
rect 297850 634760 297950 634860
rect 298074 634760 298174 634860
rect 298298 634760 298398 634860
rect 298522 634760 298622 634860
rect 298746 634760 298846 634860
rect 297850 634536 297950 634636
rect 298074 634536 298174 634636
rect 298298 634536 298398 634636
rect 298522 634536 298622 634636
rect 298746 634536 298846 634636
rect 297850 634312 297950 634412
rect 298074 634312 298174 634412
rect 298298 634312 298398 634412
rect 298522 634312 298622 634412
rect 298746 634312 298846 634412
rect 297850 634088 297950 634188
rect 298074 634088 298174 634188
rect 298298 634088 298398 634188
rect 298522 634088 298622 634188
rect 298746 634088 298846 634188
rect 297850 633864 297950 633964
rect 298074 633864 298174 633964
rect 298298 633864 298398 633964
rect 298522 633864 298622 633964
rect 298746 633864 298846 633964
rect 297850 633640 297950 633740
rect 298074 633640 298174 633740
rect 298298 633640 298398 633740
rect 298522 633640 298622 633740
rect 298746 633640 298846 633740
rect 297850 633416 297950 633516
rect 298074 633416 298174 633516
rect 298298 633416 298398 633516
rect 298522 633416 298622 633516
rect 298746 633416 298846 633516
rect 297850 633192 297950 633292
rect 298074 633192 298174 633292
rect 298298 633192 298398 633292
rect 298522 633192 298622 633292
rect 298746 633192 298846 633292
rect 297850 632968 297950 633068
rect 298074 632968 298174 633068
rect 298298 632968 298398 633068
rect 298522 632968 298622 633068
rect 298746 632968 298846 633068
rect 297850 632744 297950 632844
rect 298074 632744 298174 632844
rect 298298 632744 298398 632844
rect 298522 632744 298622 632844
rect 298746 632744 298846 632844
rect 297850 632520 297950 632620
rect 298074 632520 298174 632620
rect 298298 632520 298398 632620
rect 298522 632520 298622 632620
rect 298746 632520 298846 632620
rect 297850 632296 297950 632396
rect 298074 632296 298174 632396
rect 298298 632296 298398 632396
rect 298522 632296 298622 632396
rect 298746 632296 298846 632396
rect 297850 632072 297950 632172
rect 298074 632072 298174 632172
rect 298298 632072 298398 632172
rect 298522 632072 298622 632172
rect 298746 632072 298846 632172
rect 297850 631848 297950 631948
rect 298074 631848 298174 631948
rect 298298 631848 298398 631948
rect 298522 631848 298622 631948
rect 298746 631848 298846 631948
rect 297850 631624 297950 631724
rect 298074 631624 298174 631724
rect 298298 631624 298398 631724
rect 298522 631624 298622 631724
rect 298746 631624 298846 631724
rect 297850 631400 297950 631500
rect 298074 631400 298174 631500
rect 298298 631400 298398 631500
rect 298522 631400 298622 631500
rect 298746 631400 298846 631500
rect 336480 645160 341264 650904
rect 510602 645217 515386 650961
rect 335616 642614 335716 642714
rect 335840 642614 335940 642714
rect 336064 642614 336164 642714
rect 336288 642614 336388 642714
rect 336512 642614 336612 642714
rect 336736 642614 336836 642714
rect 336960 642614 337060 642714
rect 337184 642614 337284 642714
rect 337408 642614 337508 642714
rect 337632 642614 337732 642714
rect 337856 642614 337956 642714
rect 338080 642614 338180 642714
rect 338304 642614 338404 642714
rect 338528 642614 338628 642714
rect 338752 642614 338852 642714
rect 338976 642614 339076 642714
rect 339200 642614 339300 642714
rect 339424 642614 339524 642714
rect 339648 642614 339748 642714
rect 339872 642614 339972 642714
rect 340096 642614 340196 642714
rect 340320 642614 340420 642714
rect 340544 642614 340644 642714
rect 340768 642614 340868 642714
rect 340992 642614 341092 642714
rect 341216 642614 341316 642714
rect 341440 642614 341540 642714
rect 341664 642614 341764 642714
rect 341888 642614 341988 642714
rect 342112 642614 342212 642714
rect 335616 642390 335716 642490
rect 335840 642390 335940 642490
rect 336064 642390 336164 642490
rect 336288 642390 336388 642490
rect 336512 642390 336612 642490
rect 336736 642390 336836 642490
rect 336960 642390 337060 642490
rect 337184 642390 337284 642490
rect 337408 642390 337508 642490
rect 337632 642390 337732 642490
rect 337856 642390 337956 642490
rect 338080 642390 338180 642490
rect 338304 642390 338404 642490
rect 338528 642390 338628 642490
rect 338752 642390 338852 642490
rect 338976 642390 339076 642490
rect 339200 642390 339300 642490
rect 339424 642390 339524 642490
rect 339648 642390 339748 642490
rect 339872 642390 339972 642490
rect 340096 642390 340196 642490
rect 340320 642390 340420 642490
rect 340544 642390 340644 642490
rect 340768 642390 340868 642490
rect 340992 642390 341092 642490
rect 341216 642390 341316 642490
rect 341440 642390 341540 642490
rect 341664 642390 341764 642490
rect 341888 642390 341988 642490
rect 342112 642390 342212 642490
rect 335616 642166 335716 642266
rect 335840 642166 335940 642266
rect 336064 642166 336164 642266
rect 336288 642166 336388 642266
rect 336512 642166 336612 642266
rect 336736 642166 336836 642266
rect 336960 642166 337060 642266
rect 337184 642166 337284 642266
rect 337408 642166 337508 642266
rect 337632 642166 337732 642266
rect 337856 642166 337956 642266
rect 338080 642166 338180 642266
rect 338304 642166 338404 642266
rect 338528 642166 338628 642266
rect 338752 642166 338852 642266
rect 338976 642166 339076 642266
rect 339200 642166 339300 642266
rect 339424 642166 339524 642266
rect 339648 642166 339748 642266
rect 339872 642166 339972 642266
rect 340096 642166 340196 642266
rect 340320 642166 340420 642266
rect 340544 642166 340644 642266
rect 340768 642166 340868 642266
rect 340992 642166 341092 642266
rect 341216 642166 341316 642266
rect 341440 642166 341540 642266
rect 341664 642166 341764 642266
rect 341888 642166 341988 642266
rect 342112 642166 342212 642266
rect 335616 641942 335716 642042
rect 335840 641942 335940 642042
rect 336064 641942 336164 642042
rect 336288 641942 336388 642042
rect 336512 641942 336612 642042
rect 336736 641942 336836 642042
rect 336960 641942 337060 642042
rect 337184 641942 337284 642042
rect 337408 641942 337508 642042
rect 337632 641942 337732 642042
rect 337856 641942 337956 642042
rect 338080 641942 338180 642042
rect 338304 641942 338404 642042
rect 338528 641942 338628 642042
rect 338752 641942 338852 642042
rect 338976 641942 339076 642042
rect 339200 641942 339300 642042
rect 339424 641942 339524 642042
rect 339648 641942 339748 642042
rect 339872 641942 339972 642042
rect 340096 641942 340196 642042
rect 340320 641942 340420 642042
rect 340544 641942 340644 642042
rect 340768 641942 340868 642042
rect 340992 641942 341092 642042
rect 341216 641942 341316 642042
rect 341440 641942 341540 642042
rect 341664 641942 341764 642042
rect 341888 641942 341988 642042
rect 342112 641942 342212 642042
rect 335616 641718 335716 641818
rect 335840 641718 335940 641818
rect 336064 641718 336164 641818
rect 336288 641718 336388 641818
rect 336512 641718 336612 641818
rect 336736 641718 336836 641818
rect 336960 641718 337060 641818
rect 337184 641718 337284 641818
rect 337408 641718 337508 641818
rect 337632 641718 337732 641818
rect 337856 641718 337956 641818
rect 338080 641718 338180 641818
rect 338304 641718 338404 641818
rect 338528 641718 338628 641818
rect 338752 641718 338852 641818
rect 338976 641718 339076 641818
rect 339200 641718 339300 641818
rect 339424 641718 339524 641818
rect 339648 641718 339748 641818
rect 339872 641718 339972 641818
rect 340096 641718 340196 641818
rect 340320 641718 340420 641818
rect 340544 641718 340644 641818
rect 340768 641718 340868 641818
rect 340992 641718 341092 641818
rect 341216 641718 341316 641818
rect 341440 641718 341540 641818
rect 341664 641718 341764 641818
rect 341888 641718 341988 641818
rect 342112 641718 342212 641818
rect 342130 637896 342230 637996
rect 342354 637896 342454 637996
rect 342578 637896 342678 637996
rect 342802 637896 342902 637996
rect 343026 637896 343126 637996
rect 342130 637672 342230 637772
rect 342354 637672 342454 637772
rect 342578 637672 342678 637772
rect 342802 637672 342902 637772
rect 343026 637672 343126 637772
rect 342130 637448 342230 637548
rect 342354 637448 342454 637548
rect 342578 637448 342678 637548
rect 342802 637448 342902 637548
rect 343026 637448 343126 637548
rect 342130 637224 342230 637324
rect 342354 637224 342454 637324
rect 342578 637224 342678 637324
rect 342802 637224 342902 637324
rect 343026 637224 343126 637324
rect 342130 637000 342230 637100
rect 342354 637000 342454 637100
rect 342578 637000 342678 637100
rect 342802 637000 342902 637100
rect 343026 637000 343126 637100
rect 342130 636776 342230 636876
rect 342354 636776 342454 636876
rect 342578 636776 342678 636876
rect 342802 636776 342902 636876
rect 343026 636776 343126 636876
rect 342130 636552 342230 636652
rect 342354 636552 342454 636652
rect 342578 636552 342678 636652
rect 342802 636552 342902 636652
rect 343026 636552 343126 636652
rect 342130 636328 342230 636428
rect 342354 636328 342454 636428
rect 342578 636328 342678 636428
rect 342802 636328 342902 636428
rect 343026 636328 343126 636428
rect 342130 636104 342230 636204
rect 342354 636104 342454 636204
rect 342578 636104 342678 636204
rect 342802 636104 342902 636204
rect 343026 636104 343126 636204
rect 342130 635880 342230 635980
rect 342354 635880 342454 635980
rect 342578 635880 342678 635980
rect 342802 635880 342902 635980
rect 343026 635880 343126 635980
rect 342130 635656 342230 635756
rect 342354 635656 342454 635756
rect 342578 635656 342678 635756
rect 342802 635656 342902 635756
rect 343026 635656 343126 635756
rect 342130 635432 342230 635532
rect 342354 635432 342454 635532
rect 342578 635432 342678 635532
rect 342802 635432 342902 635532
rect 343026 635432 343126 635532
rect 342130 635208 342230 635308
rect 342354 635208 342454 635308
rect 342578 635208 342678 635308
rect 342802 635208 342902 635308
rect 343026 635208 343126 635308
rect 342130 634984 342230 635084
rect 342354 634984 342454 635084
rect 342578 634984 342678 635084
rect 342802 634984 342902 635084
rect 343026 634984 343126 635084
rect 342130 634760 342230 634860
rect 342354 634760 342454 634860
rect 342578 634760 342678 634860
rect 342802 634760 342902 634860
rect 343026 634760 343126 634860
rect 342130 634536 342230 634636
rect 342354 634536 342454 634636
rect 342578 634536 342678 634636
rect 342802 634536 342902 634636
rect 343026 634536 343126 634636
rect 342130 634312 342230 634412
rect 342354 634312 342454 634412
rect 342578 634312 342678 634412
rect 342802 634312 342902 634412
rect 343026 634312 343126 634412
rect 342130 634088 342230 634188
rect 342354 634088 342454 634188
rect 342578 634088 342678 634188
rect 342802 634088 342902 634188
rect 343026 634088 343126 634188
rect 342130 633864 342230 633964
rect 342354 633864 342454 633964
rect 342578 633864 342678 633964
rect 342802 633864 342902 633964
rect 343026 633864 343126 633964
rect 342130 633640 342230 633740
rect 342354 633640 342454 633740
rect 342578 633640 342678 633740
rect 342802 633640 342902 633740
rect 343026 633640 343126 633740
rect 342130 633416 342230 633516
rect 342354 633416 342454 633516
rect 342578 633416 342678 633516
rect 342802 633416 342902 633516
rect 343026 633416 343126 633516
rect 342130 633192 342230 633292
rect 342354 633192 342454 633292
rect 342578 633192 342678 633292
rect 342802 633192 342902 633292
rect 343026 633192 343126 633292
rect 342130 632968 342230 633068
rect 342354 632968 342454 633068
rect 342578 632968 342678 633068
rect 342802 632968 342902 633068
rect 343026 632968 343126 633068
rect 342130 632744 342230 632844
rect 342354 632744 342454 632844
rect 342578 632744 342678 632844
rect 342802 632744 342902 632844
rect 343026 632744 343126 632844
rect 342130 632520 342230 632620
rect 342354 632520 342454 632620
rect 342578 632520 342678 632620
rect 342802 632520 342902 632620
rect 343026 632520 343126 632620
rect 342130 632296 342230 632396
rect 342354 632296 342454 632396
rect 342578 632296 342678 632396
rect 342802 632296 342902 632396
rect 343026 632296 343126 632396
rect 342130 632072 342230 632172
rect 342354 632072 342454 632172
rect 342578 632072 342678 632172
rect 342802 632072 342902 632172
rect 343026 632072 343126 632172
rect 342130 631848 342230 631948
rect 342354 631848 342454 631948
rect 342578 631848 342678 631948
rect 342802 631848 342902 631948
rect 343026 631848 343126 631948
rect 342130 631624 342230 631724
rect 342354 631624 342454 631724
rect 342578 631624 342678 631724
rect 342802 631624 342902 631724
rect 343026 631624 343126 631724
rect 342130 631400 342230 631500
rect 342354 631400 342454 631500
rect 342578 631400 342678 631500
rect 342802 631400 342902 631500
rect 343026 631400 343126 631500
rect 510602 631817 515386 637561
rect 319400 628668 319600 628868
rect 319834 628668 320034 628868
rect 320268 628668 320468 628868
rect 320702 628668 320902 628868
rect 321136 628668 321336 628868
rect 321570 628668 321770 628868
rect 322004 628668 322204 628868
rect 322438 628668 322638 628868
rect 322872 628668 323072 628868
rect 323306 628668 323506 628868
rect 323740 628668 323940 628868
rect 324140 628668 324340 628868
rect 324540 628668 324740 628868
rect 324940 628668 325140 628868
rect 325340 628668 325540 628868
rect 325740 628668 325940 628868
rect 326140 628668 326340 628868
rect 326540 628668 326740 628868
rect 326940 628668 327140 628868
rect 327340 628668 327540 628868
rect 328940 628668 329140 628868
rect 329340 628668 329540 628868
rect 329740 628668 329940 628868
rect 330140 628668 330340 628868
rect 330540 628668 330740 628868
rect 330940 628668 331140 628868
rect 331340 628668 331540 628868
rect 331740 628668 331940 628868
rect 332140 628668 332340 628868
rect 319400 628234 319600 628434
rect 319834 628234 320034 628434
rect 320268 628234 320468 628434
rect 320702 628234 320902 628434
rect 321136 628234 321336 628434
rect 321570 628234 321770 628434
rect 322004 628234 322204 628434
rect 322438 628234 322638 628434
rect 322872 628234 323072 628434
rect 323306 628234 323506 628434
rect 323740 628234 323940 628434
rect 319400 627800 319600 628000
rect 319834 627800 320034 628000
rect 320268 627800 320468 628000
rect 320702 627800 320902 628000
rect 321136 627800 321336 628000
rect 321570 627800 321770 628000
rect 322004 627800 322204 628000
rect 322438 627800 322638 628000
rect 322872 627800 323072 628000
rect 323306 627800 323506 628000
rect 323740 627800 323940 628000
rect 297856 626112 297920 626176
rect 297984 626112 298048 626176
rect 298112 626112 298176 626176
rect 298240 626112 298304 626176
rect 298368 626112 298432 626176
rect 298496 626112 298560 626176
rect 298624 626112 298688 626176
rect 298752 626112 298816 626176
rect 298880 626112 298944 626176
rect 297856 625984 297920 626048
rect 297984 625984 298048 626048
rect 298112 625984 298176 626048
rect 298240 625984 298304 626048
rect 298368 625984 298432 626048
rect 298496 625984 298560 626048
rect 298624 625984 298688 626048
rect 298752 625984 298816 626048
rect 298880 625984 298944 626048
rect 297856 625856 297920 625920
rect 297984 625856 298048 625920
rect 298112 625856 298176 625920
rect 298240 625856 298304 625920
rect 298368 625856 298432 625920
rect 298496 625856 298560 625920
rect 298624 625856 298688 625920
rect 298752 625856 298816 625920
rect 298880 625856 298944 625920
rect 297856 625728 297920 625792
rect 297984 625728 298048 625792
rect 298112 625728 298176 625792
rect 298240 625728 298304 625792
rect 298368 625728 298432 625792
rect 298496 625728 298560 625792
rect 298624 625728 298688 625792
rect 298752 625728 298816 625792
rect 298880 625728 298944 625792
rect 289920 618040 294704 623784
rect 297850 624496 297950 624596
rect 298074 624496 298174 624596
rect 298298 624496 298398 624596
rect 298522 624496 298622 624596
rect 298746 624496 298846 624596
rect 297850 624272 297950 624372
rect 298074 624272 298174 624372
rect 298298 624272 298398 624372
rect 298522 624272 298622 624372
rect 298746 624272 298846 624372
rect 297850 624048 297950 624148
rect 298074 624048 298174 624148
rect 298298 624048 298398 624148
rect 298522 624048 298622 624148
rect 298746 624048 298846 624148
rect 297850 623824 297950 623924
rect 298074 623824 298174 623924
rect 298298 623824 298398 623924
rect 298522 623824 298622 623924
rect 298746 623824 298846 623924
rect 297850 623600 297950 623700
rect 298074 623600 298174 623700
rect 298298 623600 298398 623700
rect 298522 623600 298622 623700
rect 298746 623600 298846 623700
rect 297850 623376 297950 623476
rect 298074 623376 298174 623476
rect 298298 623376 298398 623476
rect 298522 623376 298622 623476
rect 298746 623376 298846 623476
rect 297850 623152 297950 623252
rect 298074 623152 298174 623252
rect 298298 623152 298398 623252
rect 298522 623152 298622 623252
rect 298746 623152 298846 623252
rect 297850 622928 297950 623028
rect 298074 622928 298174 623028
rect 298298 622928 298398 623028
rect 298522 622928 298622 623028
rect 298746 622928 298846 623028
rect 297850 622704 297950 622804
rect 298074 622704 298174 622804
rect 298298 622704 298398 622804
rect 298522 622704 298622 622804
rect 298746 622704 298846 622804
rect 297850 622480 297950 622580
rect 298074 622480 298174 622580
rect 298298 622480 298398 622580
rect 298522 622480 298622 622580
rect 298746 622480 298846 622580
rect 297850 622256 297950 622356
rect 298074 622256 298174 622356
rect 298298 622256 298398 622356
rect 298522 622256 298622 622356
rect 298746 622256 298846 622356
rect 297850 622032 297950 622132
rect 298074 622032 298174 622132
rect 298298 622032 298398 622132
rect 298522 622032 298622 622132
rect 298746 622032 298846 622132
rect 297850 621808 297950 621908
rect 298074 621808 298174 621908
rect 298298 621808 298398 621908
rect 298522 621808 298622 621908
rect 298746 621808 298846 621908
rect 297850 621584 297950 621684
rect 298074 621584 298174 621684
rect 298298 621584 298398 621684
rect 298522 621584 298622 621684
rect 298746 621584 298846 621684
rect 297850 621360 297950 621460
rect 298074 621360 298174 621460
rect 298298 621360 298398 621460
rect 298522 621360 298622 621460
rect 298746 621360 298846 621460
rect 297850 621136 297950 621236
rect 298074 621136 298174 621236
rect 298298 621136 298398 621236
rect 298522 621136 298622 621236
rect 298746 621136 298846 621236
rect 297850 620912 297950 621012
rect 298074 620912 298174 621012
rect 298298 620912 298398 621012
rect 298522 620912 298622 621012
rect 298746 620912 298846 621012
rect 297850 620688 297950 620788
rect 298074 620688 298174 620788
rect 298298 620688 298398 620788
rect 298522 620688 298622 620788
rect 298746 620688 298846 620788
rect 297850 620464 297950 620564
rect 298074 620464 298174 620564
rect 298298 620464 298398 620564
rect 298522 620464 298622 620564
rect 298746 620464 298846 620564
rect 297850 620240 297950 620340
rect 298074 620240 298174 620340
rect 298298 620240 298398 620340
rect 298522 620240 298622 620340
rect 298746 620240 298846 620340
rect 297850 620016 297950 620116
rect 298074 620016 298174 620116
rect 298298 620016 298398 620116
rect 298522 620016 298622 620116
rect 298746 620016 298846 620116
rect 297850 619792 297950 619892
rect 298074 619792 298174 619892
rect 298298 619792 298398 619892
rect 298522 619792 298622 619892
rect 298746 619792 298846 619892
rect 297850 619568 297950 619668
rect 298074 619568 298174 619668
rect 298298 619568 298398 619668
rect 298522 619568 298622 619668
rect 298746 619568 298846 619668
rect 297850 619344 297950 619444
rect 298074 619344 298174 619444
rect 298298 619344 298398 619444
rect 298522 619344 298622 619444
rect 298746 619344 298846 619444
rect 297850 619120 297950 619220
rect 298074 619120 298174 619220
rect 298298 619120 298398 619220
rect 298522 619120 298622 619220
rect 298746 619120 298846 619220
rect 297850 618896 297950 618996
rect 298074 618896 298174 618996
rect 298298 618896 298398 618996
rect 298522 618896 298622 618996
rect 298746 618896 298846 618996
rect 297850 618672 297950 618772
rect 298074 618672 298174 618772
rect 298298 618672 298398 618772
rect 298522 618672 298622 618772
rect 298746 618672 298846 618772
rect 297850 618448 297950 618548
rect 298074 618448 298174 618548
rect 298298 618448 298398 618548
rect 298522 618448 298622 618548
rect 298746 618448 298846 618548
rect 297850 618224 297950 618324
rect 298074 618224 298174 618324
rect 298298 618224 298398 618324
rect 298522 618224 298622 618324
rect 298746 618224 298846 618324
rect 297850 618000 297950 618100
rect 298074 618000 298174 618100
rect 298298 618000 298398 618100
rect 298522 618000 298622 618100
rect 298746 618000 298846 618100
rect 342130 624496 342230 624596
rect 342354 624496 342454 624596
rect 342578 624496 342678 624596
rect 342802 624496 342902 624596
rect 343026 624496 343126 624596
rect 342130 624272 342230 624372
rect 342354 624272 342454 624372
rect 342578 624272 342678 624372
rect 342802 624272 342902 624372
rect 343026 624272 343126 624372
rect 342130 624048 342230 624148
rect 342354 624048 342454 624148
rect 342578 624048 342678 624148
rect 342802 624048 342902 624148
rect 343026 624048 343126 624148
rect 342130 623824 342230 623924
rect 342354 623824 342454 623924
rect 342578 623824 342678 623924
rect 342802 623824 342902 623924
rect 343026 623824 343126 623924
rect 342130 623600 342230 623700
rect 342354 623600 342454 623700
rect 342578 623600 342678 623700
rect 342802 623600 342902 623700
rect 343026 623600 343126 623700
rect 342130 623376 342230 623476
rect 342354 623376 342454 623476
rect 342578 623376 342678 623476
rect 342802 623376 342902 623476
rect 343026 623376 343126 623476
rect 342130 623152 342230 623252
rect 342354 623152 342454 623252
rect 342578 623152 342678 623252
rect 342802 623152 342902 623252
rect 343026 623152 343126 623252
rect 342130 622928 342230 623028
rect 342354 622928 342454 623028
rect 342578 622928 342678 623028
rect 342802 622928 342902 623028
rect 343026 622928 343126 623028
rect 342130 622704 342230 622804
rect 342354 622704 342454 622804
rect 342578 622704 342678 622804
rect 342802 622704 342902 622804
rect 343026 622704 343126 622804
rect 342130 622480 342230 622580
rect 342354 622480 342454 622580
rect 342578 622480 342678 622580
rect 342802 622480 342902 622580
rect 343026 622480 343126 622580
rect 342130 622256 342230 622356
rect 342354 622256 342454 622356
rect 342578 622256 342678 622356
rect 342802 622256 342902 622356
rect 343026 622256 343126 622356
rect 342130 622032 342230 622132
rect 342354 622032 342454 622132
rect 342578 622032 342678 622132
rect 342802 622032 342902 622132
rect 343026 622032 343126 622132
rect 342130 621808 342230 621908
rect 342354 621808 342454 621908
rect 342578 621808 342678 621908
rect 342802 621808 342902 621908
rect 343026 621808 343126 621908
rect 342130 621584 342230 621684
rect 342354 621584 342454 621684
rect 342578 621584 342678 621684
rect 342802 621584 342902 621684
rect 343026 621584 343126 621684
rect 342130 621360 342230 621460
rect 342354 621360 342454 621460
rect 342578 621360 342678 621460
rect 342802 621360 342902 621460
rect 343026 621360 343126 621460
rect 342130 621136 342230 621236
rect 342354 621136 342454 621236
rect 342578 621136 342678 621236
rect 342802 621136 342902 621236
rect 343026 621136 343126 621236
rect 342130 620912 342230 621012
rect 342354 620912 342454 621012
rect 342578 620912 342678 621012
rect 342802 620912 342902 621012
rect 343026 620912 343126 621012
rect 342130 620688 342230 620788
rect 342354 620688 342454 620788
rect 342578 620688 342678 620788
rect 342802 620688 342902 620788
rect 343026 620688 343126 620788
rect 342130 620464 342230 620564
rect 342354 620464 342454 620564
rect 342578 620464 342678 620564
rect 342802 620464 342902 620564
rect 343026 620464 343126 620564
rect 342130 620240 342230 620340
rect 342354 620240 342454 620340
rect 342578 620240 342678 620340
rect 342802 620240 342902 620340
rect 343026 620240 343126 620340
rect 342130 620016 342230 620116
rect 342354 620016 342454 620116
rect 342578 620016 342678 620116
rect 342802 620016 342902 620116
rect 343026 620016 343126 620116
rect 342130 619792 342230 619892
rect 342354 619792 342454 619892
rect 342578 619792 342678 619892
rect 342802 619792 342902 619892
rect 343026 619792 343126 619892
rect 342130 619568 342230 619668
rect 342354 619568 342454 619668
rect 342578 619568 342678 619668
rect 342802 619568 342902 619668
rect 343026 619568 343126 619668
rect 342130 619344 342230 619444
rect 342354 619344 342454 619444
rect 342578 619344 342678 619444
rect 342802 619344 342902 619444
rect 343026 619344 343126 619444
rect 342130 619120 342230 619220
rect 342354 619120 342454 619220
rect 342578 619120 342678 619220
rect 342802 619120 342902 619220
rect 343026 619120 343126 619220
rect 342130 618896 342230 618996
rect 342354 618896 342454 618996
rect 342578 618896 342678 618996
rect 342802 618896 342902 618996
rect 343026 618896 343126 618996
rect 342130 618672 342230 618772
rect 342354 618672 342454 618772
rect 342578 618672 342678 618772
rect 342802 618672 342902 618772
rect 343026 618672 343126 618772
rect 342130 618448 342230 618548
rect 342354 618448 342454 618548
rect 342578 618448 342678 618548
rect 342802 618448 342902 618548
rect 343026 618448 343126 618548
rect 342130 618224 342230 618324
rect 342354 618224 342454 618324
rect 342578 618224 342678 618324
rect 342802 618224 342902 618324
rect 343026 618224 343126 618324
rect 342130 618000 342230 618100
rect 342354 618000 342454 618100
rect 342578 618000 342678 618100
rect 342802 618000 342902 618100
rect 343026 618000 343126 618100
rect 510602 618417 515386 624161
rect 289920 605020 294704 610764
rect 298876 615374 298976 615474
rect 299100 615374 299200 615474
rect 299324 615374 299424 615474
rect 299548 615374 299648 615474
rect 299772 615374 299872 615474
rect 299996 615374 300096 615474
rect 300220 615374 300320 615474
rect 300444 615374 300544 615474
rect 300668 615374 300768 615474
rect 300892 615374 300992 615474
rect 301116 615374 301216 615474
rect 301340 615374 301440 615474
rect 301564 615374 301664 615474
rect 301788 615374 301888 615474
rect 302012 615374 302112 615474
rect 302236 615374 302336 615474
rect 302460 615374 302560 615474
rect 302684 615374 302784 615474
rect 302908 615374 303008 615474
rect 303132 615374 303232 615474
rect 303356 615374 303456 615474
rect 303580 615374 303680 615474
rect 303804 615374 303904 615474
rect 304028 615374 304128 615474
rect 304252 615374 304352 615474
rect 304476 615374 304576 615474
rect 304700 615374 304800 615474
rect 304924 615374 305024 615474
rect 305148 615374 305248 615474
rect 305372 615374 305472 615474
rect 309346 615374 309446 615474
rect 309570 615374 309670 615474
rect 309794 615374 309894 615474
rect 310018 615374 310118 615474
rect 310242 615374 310342 615474
rect 310466 615374 310566 615474
rect 310690 615374 310790 615474
rect 310914 615374 311014 615474
rect 311138 615374 311238 615474
rect 311362 615374 311462 615474
rect 311586 615374 311686 615474
rect 311810 615374 311910 615474
rect 312034 615374 312134 615474
rect 312258 615374 312358 615474
rect 312482 615374 312582 615474
rect 312706 615374 312806 615474
rect 312930 615374 313030 615474
rect 313154 615374 313254 615474
rect 313378 615374 313478 615474
rect 313602 615374 313702 615474
rect 313826 615374 313926 615474
rect 314050 615374 314150 615474
rect 314274 615374 314374 615474
rect 314498 615374 314598 615474
rect 314722 615374 314822 615474
rect 314946 615374 315046 615474
rect 315170 615374 315270 615474
rect 315394 615374 315494 615474
rect 315618 615374 315718 615474
rect 315842 615374 315942 615474
rect 298876 615150 298976 615250
rect 299100 615150 299200 615250
rect 299324 615150 299424 615250
rect 299548 615150 299648 615250
rect 299772 615150 299872 615250
rect 299996 615150 300096 615250
rect 300220 615150 300320 615250
rect 300444 615150 300544 615250
rect 300668 615150 300768 615250
rect 300892 615150 300992 615250
rect 301116 615150 301216 615250
rect 301340 615150 301440 615250
rect 301564 615150 301664 615250
rect 301788 615150 301888 615250
rect 302012 615150 302112 615250
rect 302236 615150 302336 615250
rect 302460 615150 302560 615250
rect 302684 615150 302784 615250
rect 302908 615150 303008 615250
rect 303132 615150 303232 615250
rect 303356 615150 303456 615250
rect 303580 615150 303680 615250
rect 303804 615150 303904 615250
rect 304028 615150 304128 615250
rect 304252 615150 304352 615250
rect 304476 615150 304576 615250
rect 304700 615150 304800 615250
rect 304924 615150 305024 615250
rect 305148 615150 305248 615250
rect 305372 615150 305472 615250
rect 309346 615150 309446 615250
rect 309570 615150 309670 615250
rect 309794 615150 309894 615250
rect 310018 615150 310118 615250
rect 310242 615150 310342 615250
rect 310466 615150 310566 615250
rect 310690 615150 310790 615250
rect 310914 615150 311014 615250
rect 311138 615150 311238 615250
rect 311362 615150 311462 615250
rect 311586 615150 311686 615250
rect 311810 615150 311910 615250
rect 312034 615150 312134 615250
rect 312258 615150 312358 615250
rect 312482 615150 312582 615250
rect 312706 615150 312806 615250
rect 312930 615150 313030 615250
rect 313154 615150 313254 615250
rect 313378 615150 313478 615250
rect 313602 615150 313702 615250
rect 313826 615150 313926 615250
rect 314050 615150 314150 615250
rect 314274 615150 314374 615250
rect 314498 615150 314598 615250
rect 314722 615150 314822 615250
rect 314946 615150 315046 615250
rect 315170 615150 315270 615250
rect 315394 615150 315494 615250
rect 315618 615150 315718 615250
rect 315842 615150 315942 615250
rect 298876 614926 298976 615026
rect 299100 614926 299200 615026
rect 299324 614926 299424 615026
rect 299548 614926 299648 615026
rect 299772 614926 299872 615026
rect 299996 614926 300096 615026
rect 300220 614926 300320 615026
rect 300444 614926 300544 615026
rect 300668 614926 300768 615026
rect 300892 614926 300992 615026
rect 301116 614926 301216 615026
rect 301340 614926 301440 615026
rect 301564 614926 301664 615026
rect 301788 614926 301888 615026
rect 302012 614926 302112 615026
rect 302236 614926 302336 615026
rect 302460 614926 302560 615026
rect 302684 614926 302784 615026
rect 302908 614926 303008 615026
rect 303132 614926 303232 615026
rect 303356 614926 303456 615026
rect 303580 614926 303680 615026
rect 303804 614926 303904 615026
rect 304028 614926 304128 615026
rect 304252 614926 304352 615026
rect 304476 614926 304576 615026
rect 304700 614926 304800 615026
rect 304924 614926 305024 615026
rect 305148 614926 305248 615026
rect 305372 614926 305472 615026
rect 309346 614926 309446 615026
rect 309570 614926 309670 615026
rect 309794 614926 309894 615026
rect 310018 614926 310118 615026
rect 310242 614926 310342 615026
rect 310466 614926 310566 615026
rect 310690 614926 310790 615026
rect 310914 614926 311014 615026
rect 311138 614926 311238 615026
rect 311362 614926 311462 615026
rect 311586 614926 311686 615026
rect 311810 614926 311910 615026
rect 312034 614926 312134 615026
rect 312258 614926 312358 615026
rect 312482 614926 312582 615026
rect 312706 614926 312806 615026
rect 312930 614926 313030 615026
rect 313154 614926 313254 615026
rect 313378 614926 313478 615026
rect 313602 614926 313702 615026
rect 313826 614926 313926 615026
rect 314050 614926 314150 615026
rect 314274 614926 314374 615026
rect 314498 614926 314598 615026
rect 314722 614926 314822 615026
rect 314946 614926 315046 615026
rect 315170 614926 315270 615026
rect 315394 614926 315494 615026
rect 315618 614926 315718 615026
rect 315842 614926 315942 615026
rect 298876 614702 298976 614802
rect 299100 614702 299200 614802
rect 299324 614702 299424 614802
rect 299548 614702 299648 614802
rect 299772 614702 299872 614802
rect 299996 614702 300096 614802
rect 300220 614702 300320 614802
rect 300444 614702 300544 614802
rect 300668 614702 300768 614802
rect 300892 614702 300992 614802
rect 301116 614702 301216 614802
rect 301340 614702 301440 614802
rect 301564 614702 301664 614802
rect 301788 614702 301888 614802
rect 302012 614702 302112 614802
rect 302236 614702 302336 614802
rect 302460 614702 302560 614802
rect 302684 614702 302784 614802
rect 302908 614702 303008 614802
rect 303132 614702 303232 614802
rect 303356 614702 303456 614802
rect 303580 614702 303680 614802
rect 303804 614702 303904 614802
rect 304028 614702 304128 614802
rect 304252 614702 304352 614802
rect 304476 614702 304576 614802
rect 304700 614702 304800 614802
rect 304924 614702 305024 614802
rect 305148 614702 305248 614802
rect 305372 614702 305472 614802
rect 309346 614702 309446 614802
rect 309570 614702 309670 614802
rect 309794 614702 309894 614802
rect 310018 614702 310118 614802
rect 310242 614702 310342 614802
rect 310466 614702 310566 614802
rect 310690 614702 310790 614802
rect 310914 614702 311014 614802
rect 311138 614702 311238 614802
rect 311362 614702 311462 614802
rect 311586 614702 311686 614802
rect 311810 614702 311910 614802
rect 312034 614702 312134 614802
rect 312258 614702 312358 614802
rect 312482 614702 312582 614802
rect 312706 614702 312806 614802
rect 312930 614702 313030 614802
rect 313154 614702 313254 614802
rect 313378 614702 313478 614802
rect 313602 614702 313702 614802
rect 313826 614702 313926 614802
rect 314050 614702 314150 614802
rect 314274 614702 314374 614802
rect 314498 614702 314598 614802
rect 314722 614702 314822 614802
rect 314946 614702 315046 614802
rect 315170 614702 315270 614802
rect 315394 614702 315494 614802
rect 315618 614702 315718 614802
rect 315842 614702 315942 614802
rect 298876 614478 298976 614578
rect 299100 614478 299200 614578
rect 299324 614478 299424 614578
rect 299548 614478 299648 614578
rect 299772 614478 299872 614578
rect 299996 614478 300096 614578
rect 300220 614478 300320 614578
rect 300444 614478 300544 614578
rect 300668 614478 300768 614578
rect 300892 614478 300992 614578
rect 301116 614478 301216 614578
rect 301340 614478 301440 614578
rect 301564 614478 301664 614578
rect 301788 614478 301888 614578
rect 302012 614478 302112 614578
rect 302236 614478 302336 614578
rect 302460 614478 302560 614578
rect 302684 614478 302784 614578
rect 302908 614478 303008 614578
rect 303132 614478 303232 614578
rect 303356 614478 303456 614578
rect 303580 614478 303680 614578
rect 303804 614478 303904 614578
rect 304028 614478 304128 614578
rect 304252 614478 304352 614578
rect 304476 614478 304576 614578
rect 304700 614478 304800 614578
rect 304924 614478 305024 614578
rect 305148 614478 305248 614578
rect 305372 614478 305472 614578
rect 309346 614478 309446 614578
rect 309570 614478 309670 614578
rect 309794 614478 309894 614578
rect 310018 614478 310118 614578
rect 310242 614478 310342 614578
rect 310466 614478 310566 614578
rect 310690 614478 310790 614578
rect 310914 614478 311014 614578
rect 311138 614478 311238 614578
rect 311362 614478 311462 614578
rect 311586 614478 311686 614578
rect 311810 614478 311910 614578
rect 312034 614478 312134 614578
rect 312258 614478 312358 614578
rect 312482 614478 312582 614578
rect 312706 614478 312806 614578
rect 312930 614478 313030 614578
rect 313154 614478 313254 614578
rect 313378 614478 313478 614578
rect 313602 614478 313702 614578
rect 313826 614478 313926 614578
rect 314050 614478 314150 614578
rect 314274 614478 314374 614578
rect 314498 614478 314598 614578
rect 314722 614478 314822 614578
rect 314946 614478 315046 614578
rect 315170 614478 315270 614578
rect 315394 614478 315494 614578
rect 315618 614478 315718 614578
rect 315842 614478 315942 614578
rect 298920 605336 303704 611080
rect 304920 605336 309704 611080
rect 310920 605336 315704 611080
rect 335616 615394 335716 615494
rect 335840 615394 335940 615494
rect 336064 615394 336164 615494
rect 336288 615394 336388 615494
rect 336512 615394 336612 615494
rect 336736 615394 336836 615494
rect 336960 615394 337060 615494
rect 337184 615394 337284 615494
rect 337408 615394 337508 615494
rect 337632 615394 337732 615494
rect 337856 615394 337956 615494
rect 338080 615394 338180 615494
rect 338304 615394 338404 615494
rect 338528 615394 338628 615494
rect 338752 615394 338852 615494
rect 338976 615394 339076 615494
rect 339200 615394 339300 615494
rect 339424 615394 339524 615494
rect 339648 615394 339748 615494
rect 339872 615394 339972 615494
rect 340096 615394 340196 615494
rect 340320 615394 340420 615494
rect 340544 615394 340644 615494
rect 340768 615394 340868 615494
rect 340992 615394 341092 615494
rect 341216 615394 341316 615494
rect 341440 615394 341540 615494
rect 341664 615394 341764 615494
rect 341888 615394 341988 615494
rect 342112 615394 342212 615494
rect 335616 615170 335716 615270
rect 335840 615170 335940 615270
rect 336064 615170 336164 615270
rect 336288 615170 336388 615270
rect 336512 615170 336612 615270
rect 336736 615170 336836 615270
rect 336960 615170 337060 615270
rect 337184 615170 337284 615270
rect 337408 615170 337508 615270
rect 337632 615170 337732 615270
rect 337856 615170 337956 615270
rect 338080 615170 338180 615270
rect 338304 615170 338404 615270
rect 338528 615170 338628 615270
rect 338752 615170 338852 615270
rect 338976 615170 339076 615270
rect 339200 615170 339300 615270
rect 339424 615170 339524 615270
rect 339648 615170 339748 615270
rect 339872 615170 339972 615270
rect 340096 615170 340196 615270
rect 340320 615170 340420 615270
rect 340544 615170 340644 615270
rect 340768 615170 340868 615270
rect 340992 615170 341092 615270
rect 341216 615170 341316 615270
rect 341440 615170 341540 615270
rect 341664 615170 341764 615270
rect 341888 615170 341988 615270
rect 342112 615170 342212 615270
rect 335616 614946 335716 615046
rect 335840 614946 335940 615046
rect 336064 614946 336164 615046
rect 336288 614946 336388 615046
rect 336512 614946 336612 615046
rect 336736 614946 336836 615046
rect 336960 614946 337060 615046
rect 337184 614946 337284 615046
rect 337408 614946 337508 615046
rect 337632 614946 337732 615046
rect 337856 614946 337956 615046
rect 338080 614946 338180 615046
rect 338304 614946 338404 615046
rect 338528 614946 338628 615046
rect 338752 614946 338852 615046
rect 338976 614946 339076 615046
rect 339200 614946 339300 615046
rect 339424 614946 339524 615046
rect 339648 614946 339748 615046
rect 339872 614946 339972 615046
rect 340096 614946 340196 615046
rect 340320 614946 340420 615046
rect 340544 614946 340644 615046
rect 340768 614946 340868 615046
rect 340992 614946 341092 615046
rect 341216 614946 341316 615046
rect 341440 614946 341540 615046
rect 341664 614946 341764 615046
rect 341888 614946 341988 615046
rect 342112 614946 342212 615046
rect 335616 614722 335716 614822
rect 335840 614722 335940 614822
rect 336064 614722 336164 614822
rect 336288 614722 336388 614822
rect 336512 614722 336612 614822
rect 336736 614722 336836 614822
rect 336960 614722 337060 614822
rect 337184 614722 337284 614822
rect 337408 614722 337508 614822
rect 337632 614722 337732 614822
rect 337856 614722 337956 614822
rect 338080 614722 338180 614822
rect 338304 614722 338404 614822
rect 338528 614722 338628 614822
rect 338752 614722 338852 614822
rect 338976 614722 339076 614822
rect 339200 614722 339300 614822
rect 339424 614722 339524 614822
rect 339648 614722 339748 614822
rect 339872 614722 339972 614822
rect 340096 614722 340196 614822
rect 340320 614722 340420 614822
rect 340544 614722 340644 614822
rect 340768 614722 340868 614822
rect 340992 614722 341092 614822
rect 341216 614722 341316 614822
rect 341440 614722 341540 614822
rect 341664 614722 341764 614822
rect 341888 614722 341988 614822
rect 342112 614722 342212 614822
rect 335616 614498 335716 614598
rect 335840 614498 335940 614598
rect 336064 614498 336164 614598
rect 336288 614498 336388 614598
rect 336512 614498 336612 614598
rect 336736 614498 336836 614598
rect 336960 614498 337060 614598
rect 337184 614498 337284 614598
rect 337408 614498 337508 614598
rect 337632 614498 337732 614598
rect 337856 614498 337956 614598
rect 338080 614498 338180 614598
rect 338304 614498 338404 614598
rect 338528 614498 338628 614598
rect 338752 614498 338852 614598
rect 338976 614498 339076 614598
rect 339200 614498 339300 614598
rect 339424 614498 339524 614598
rect 339648 614498 339748 614598
rect 339872 614498 339972 614598
rect 340096 614498 340196 614598
rect 340320 614498 340420 614598
rect 340544 614498 340644 614598
rect 340768 614498 340868 614598
rect 340992 614498 341092 614598
rect 341216 614498 341316 614598
rect 341440 614498 341540 614598
rect 341664 614498 341764 614598
rect 341888 614498 341988 614598
rect 342112 614498 342212 614598
rect 336480 605340 341264 611084
rect 510602 605017 515386 610761
rect 520602 684336 525386 690560
rect 520602 645217 525386 650961
rect 560582 639792 566726 644576
rect 520602 631817 525386 637561
rect 560582 629792 566726 634576
rect 520602 618417 525386 624161
rect 520602 605017 525386 610761
rect 317480 591580 322264 597324
rect 325480 591580 330264 597324
rect 13897 462422 13961 462486
rect 13977 462422 14041 462486
rect 14057 462422 14121 462486
rect 14137 462422 14201 462486
rect 14217 462422 14281 462486
rect 14297 462422 14361 462486
rect 14377 462422 14441 462486
rect 14457 462422 14521 462486
rect 14537 462422 14601 462486
rect 14617 462422 14681 462486
rect 14697 462422 14761 462486
rect 14777 462422 14841 462486
rect 14857 462422 14921 462486
rect 14937 462422 15001 462486
rect 15017 462422 15081 462486
rect 15097 462422 15161 462486
rect 15177 462422 15241 462486
rect 15257 462422 15321 462486
rect 15337 462422 15401 462486
rect 15417 462422 15481 462486
rect 15497 462422 15561 462486
rect 15577 462422 15641 462486
rect 15657 462422 15721 462486
rect 15737 462422 15801 462486
rect 15817 462422 15881 462486
rect 15897 462422 15961 462486
rect 15977 462422 16041 462486
rect 16057 462422 16121 462486
rect 16137 462422 16201 462486
rect 16217 462422 16281 462486
rect 16297 462422 16361 462486
rect 16377 462422 16441 462486
rect 16457 462422 16521 462486
rect 16537 462422 16601 462486
rect 16617 462422 16681 462486
rect 16697 462422 16761 462486
rect 16777 462422 16841 462486
rect 16857 462422 16921 462486
rect 16937 462422 17001 462486
rect 17017 462422 17081 462486
rect 17097 462422 17161 462486
rect 17177 462422 17241 462486
rect 17257 462422 17321 462486
rect 17337 462422 17401 462486
rect 17417 462422 17481 462486
rect 17497 462422 17561 462486
rect 13911 419200 13975 419264
rect 13991 419200 14055 419264
rect 14071 419200 14135 419264
rect 14151 419200 14215 419264
rect 14231 419200 14295 419264
rect 14311 419200 14375 419264
rect 14391 419200 14455 419264
rect 14471 419200 14535 419264
rect 14551 419200 14615 419264
rect 14631 419200 14695 419264
rect 14711 419200 14775 419264
rect 14791 419200 14855 419264
rect 14871 419200 14935 419264
rect 14951 419200 15015 419264
rect 15031 419200 15095 419264
rect 15111 419200 15175 419264
rect 15191 419200 15255 419264
rect 15271 419200 15335 419264
rect 15351 419200 15415 419264
rect 15431 419200 15495 419264
rect 15511 419200 15575 419264
rect 15591 419200 15655 419264
rect 15671 419200 15735 419264
rect 15751 419200 15815 419264
rect 15831 419200 15895 419264
rect 15911 419200 15975 419264
rect 15991 419200 16055 419264
rect 16071 419200 16135 419264
rect 16151 419200 16215 419264
rect 16231 419200 16295 419264
rect 16311 419200 16375 419264
rect 16391 419200 16455 419264
rect 16471 419200 16535 419264
rect 16551 419200 16615 419264
rect 16631 419200 16695 419264
rect 16711 419200 16775 419264
rect 16791 419200 16855 419264
rect 16871 419200 16935 419264
rect 16951 419200 17015 419264
rect 17031 419200 17095 419264
rect 17111 419200 17175 419264
rect 17191 419200 17255 419264
rect 17271 419200 17335 419264
rect 17351 419200 17415 419264
rect 17431 419200 17495 419264
rect 17511 419200 17575 419264
rect 556255 550570 562319 555354
rect 556255 540570 562319 545354
rect 573553 500074 573617 500138
rect 573633 500074 573697 500138
rect 573713 500074 573777 500138
rect 573793 500074 573857 500138
rect 573873 500074 573937 500138
rect 573953 500074 574017 500138
rect 574033 500074 574097 500138
rect 574113 500074 574177 500138
rect 574193 500074 574257 500138
rect 574273 500074 574337 500138
rect 574353 500074 574417 500138
rect 574433 500074 574497 500138
rect 574513 500074 574577 500138
rect 574593 500074 574657 500138
rect 574673 500074 574737 500138
rect 574753 500074 574817 500138
rect 574833 500074 574897 500138
rect 574913 500074 574977 500138
rect 574993 500074 575057 500138
rect 575073 500074 575137 500138
rect 575153 500074 575217 500138
rect 575233 500074 575297 500138
rect 575313 500074 575377 500138
rect 575393 500074 575457 500138
rect 575473 500074 575537 500138
rect 575553 500074 575617 500138
rect 575633 500074 575697 500138
rect 575713 500074 575777 500138
rect 575793 500074 575857 500138
rect 575873 500074 575937 500138
rect 575953 500074 576017 500138
rect 576033 500074 576097 500138
rect 576113 500074 576177 500138
rect 576193 500074 576257 500138
rect 576273 500074 576337 500138
rect 576353 500074 576417 500138
rect 576433 500074 576497 500138
rect 576513 500074 576577 500138
rect 576593 500074 576657 500138
rect 576673 500074 576737 500138
rect 573591 455652 573655 455716
rect 573671 455652 573735 455716
rect 573751 455652 573815 455716
rect 573831 455652 573895 455716
rect 573911 455652 573975 455716
rect 573991 455652 574055 455716
rect 574071 455652 574135 455716
rect 574151 455652 574215 455716
rect 574231 455652 574295 455716
rect 574311 455652 574375 455716
rect 574391 455652 574455 455716
rect 574471 455652 574535 455716
rect 574551 455652 574615 455716
rect 574631 455652 574695 455716
rect 574711 455652 574775 455716
rect 574791 455652 574855 455716
rect 574871 455652 574935 455716
rect 574951 455652 575015 455716
rect 575031 455652 575095 455716
rect 575111 455652 575175 455716
rect 575191 455652 575255 455716
rect 575271 455652 575335 455716
rect 575351 455652 575415 455716
rect 575431 455652 575495 455716
rect 575511 455652 575575 455716
rect 575591 455652 575655 455716
rect 575671 455652 575735 455716
rect 575751 455652 575815 455716
rect 575831 455652 575895 455716
rect 575911 455652 575975 455716
rect 575991 455652 576055 455716
rect 576071 455652 576135 455716
rect 576151 455652 576215 455716
rect 576231 455652 576295 455716
rect 576311 455652 576375 455716
rect 576391 455652 576455 455716
rect 576471 455652 576535 455716
rect 576551 455652 576615 455716
rect 576631 455652 576695 455716
rect 13997 191438 17421 196222
rect 573605 191438 576629 196222
<< metal4 >>
rect 170628 690610 526162 690737
rect 170628 690577 222622 690610
rect 170628 684353 170922 690577
rect 173066 684353 173422 690577
rect 175566 684386 222622 690577
rect 224766 690593 526162 690610
rect 224766 690084 324322 690593
rect 224766 684386 289800 690084
rect 175566 684353 289800 684386
rect 170628 684340 289800 684353
rect 294584 684369 324322 690084
rect 326466 690560 526162 690593
rect 326466 684369 510602 690560
rect 294584 684340 510602 684369
rect 170628 684336 510602 684340
rect 515386 684336 520602 690560
rect 525386 684336 526162 690560
rect 170628 684183 526162 684336
rect 343420 651400 525804 651406
rect 285800 650961 525804 651400
rect 285800 650904 510602 650961
rect 285800 650584 336480 650904
rect 285800 644840 289920 650584
rect 294704 644840 298920 650584
rect 303704 644840 304920 650584
rect 309704 644840 310920 650584
rect 315704 645160 336480 650584
rect 341264 645217 510602 650904
rect 515386 645217 520602 650961
rect 525386 645217 525804 650961
rect 341264 645160 525804 645217
rect 315704 644840 525804 645160
rect 285800 644744 525804 644840
rect 560425 644576 566979 644980
rect 335560 642719 342216 642724
rect 335560 642714 342217 642719
rect 298820 642699 305476 642704
rect 309290 642699 315946 642704
rect 298820 642694 305477 642699
rect 298820 642594 298876 642694
rect 298976 642594 299100 642694
rect 299200 642594 299324 642694
rect 299424 642594 299548 642694
rect 299648 642594 299772 642694
rect 299872 642594 299996 642694
rect 300096 642594 300220 642694
rect 300320 642594 300444 642694
rect 300544 642594 300668 642694
rect 300768 642594 300892 642694
rect 300992 642594 301116 642694
rect 301216 642594 301340 642694
rect 301440 642594 301564 642694
rect 301664 642594 301788 642694
rect 301888 642594 302012 642694
rect 302112 642594 302236 642694
rect 302336 642594 302460 642694
rect 302560 642594 302684 642694
rect 302784 642594 302908 642694
rect 303008 642594 303132 642694
rect 303232 642594 303356 642694
rect 303456 642594 303580 642694
rect 303680 642594 303804 642694
rect 303904 642594 304028 642694
rect 304128 642594 304252 642694
rect 304352 642594 304476 642694
rect 304576 642594 304700 642694
rect 304800 642594 304924 642694
rect 305024 642594 305148 642694
rect 305248 642594 305372 642694
rect 305472 642594 305477 642694
rect 298820 642589 305477 642594
rect 309290 642694 315947 642699
rect 309290 642594 309346 642694
rect 309446 642594 309570 642694
rect 309670 642594 309794 642694
rect 309894 642594 310018 642694
rect 310118 642594 310242 642694
rect 310342 642594 310466 642694
rect 310566 642594 310690 642694
rect 310790 642594 310914 642694
rect 311014 642594 311138 642694
rect 311238 642594 311362 642694
rect 311462 642594 311586 642694
rect 311686 642594 311810 642694
rect 311910 642594 312034 642694
rect 312134 642594 312258 642694
rect 312358 642594 312482 642694
rect 312582 642594 312706 642694
rect 312806 642594 312930 642694
rect 313030 642594 313154 642694
rect 313254 642594 313378 642694
rect 313478 642594 313602 642694
rect 313702 642594 313826 642694
rect 313926 642594 314050 642694
rect 314150 642594 314274 642694
rect 314374 642594 314498 642694
rect 314598 642594 314722 642694
rect 314822 642594 314946 642694
rect 315046 642594 315170 642694
rect 315270 642594 315394 642694
rect 315494 642594 315618 642694
rect 315718 642594 315842 642694
rect 315942 642594 315947 642694
rect 309290 642589 315947 642594
rect 335560 642614 335616 642714
rect 335716 642614 335840 642714
rect 335940 642614 336064 642714
rect 336164 642614 336288 642714
rect 336388 642614 336512 642714
rect 336612 642614 336736 642714
rect 336836 642614 336960 642714
rect 337060 642614 337184 642714
rect 337284 642614 337408 642714
rect 337508 642614 337632 642714
rect 337732 642614 337856 642714
rect 337956 642614 338080 642714
rect 338180 642614 338304 642714
rect 338404 642614 338528 642714
rect 338628 642614 338752 642714
rect 338852 642614 338976 642714
rect 339076 642614 339200 642714
rect 339300 642614 339424 642714
rect 339524 642614 339648 642714
rect 339748 642614 339872 642714
rect 339972 642614 340096 642714
rect 340196 642614 340320 642714
rect 340420 642614 340544 642714
rect 340644 642614 340768 642714
rect 340868 642614 340992 642714
rect 341092 642614 341216 642714
rect 341316 642614 341440 642714
rect 341540 642614 341664 642714
rect 341764 642614 341888 642714
rect 341988 642614 342112 642714
rect 342212 642614 342217 642714
rect 335560 642609 342217 642614
rect 298820 642475 305476 642589
rect 309290 642475 315946 642589
rect 335560 642495 342216 642609
rect 335560 642490 342217 642495
rect 298820 642470 305477 642475
rect 298820 642370 298876 642470
rect 298976 642370 299100 642470
rect 299200 642370 299324 642470
rect 299424 642370 299548 642470
rect 299648 642370 299772 642470
rect 299872 642370 299996 642470
rect 300096 642370 300220 642470
rect 300320 642370 300444 642470
rect 300544 642370 300668 642470
rect 300768 642370 300892 642470
rect 300992 642370 301116 642470
rect 301216 642370 301340 642470
rect 301440 642370 301564 642470
rect 301664 642370 301788 642470
rect 301888 642370 302012 642470
rect 302112 642370 302236 642470
rect 302336 642370 302460 642470
rect 302560 642370 302684 642470
rect 302784 642370 302908 642470
rect 303008 642370 303132 642470
rect 303232 642370 303356 642470
rect 303456 642370 303580 642470
rect 303680 642370 303804 642470
rect 303904 642370 304028 642470
rect 304128 642370 304252 642470
rect 304352 642370 304476 642470
rect 304576 642370 304700 642470
rect 304800 642370 304924 642470
rect 305024 642370 305148 642470
rect 305248 642370 305372 642470
rect 305472 642370 305477 642470
rect 298820 642365 305477 642370
rect 309290 642470 315947 642475
rect 309290 642370 309346 642470
rect 309446 642370 309570 642470
rect 309670 642370 309794 642470
rect 309894 642370 310018 642470
rect 310118 642370 310242 642470
rect 310342 642370 310466 642470
rect 310566 642370 310690 642470
rect 310790 642370 310914 642470
rect 311014 642370 311138 642470
rect 311238 642370 311362 642470
rect 311462 642370 311586 642470
rect 311686 642370 311810 642470
rect 311910 642370 312034 642470
rect 312134 642370 312258 642470
rect 312358 642370 312482 642470
rect 312582 642370 312706 642470
rect 312806 642370 312930 642470
rect 313030 642370 313154 642470
rect 313254 642370 313378 642470
rect 313478 642370 313602 642470
rect 313702 642370 313826 642470
rect 313926 642370 314050 642470
rect 314150 642370 314274 642470
rect 314374 642370 314498 642470
rect 314598 642370 314722 642470
rect 314822 642370 314946 642470
rect 315046 642370 315170 642470
rect 315270 642370 315394 642470
rect 315494 642370 315618 642470
rect 315718 642370 315842 642470
rect 315942 642370 315947 642470
rect 309290 642365 315947 642370
rect 335560 642390 335616 642490
rect 335716 642390 335840 642490
rect 335940 642390 336064 642490
rect 336164 642390 336288 642490
rect 336388 642390 336512 642490
rect 336612 642390 336736 642490
rect 336836 642390 336960 642490
rect 337060 642390 337184 642490
rect 337284 642390 337408 642490
rect 337508 642390 337632 642490
rect 337732 642390 337856 642490
rect 337956 642390 338080 642490
rect 338180 642390 338304 642490
rect 338404 642390 338528 642490
rect 338628 642390 338752 642490
rect 338852 642390 338976 642490
rect 339076 642390 339200 642490
rect 339300 642390 339424 642490
rect 339524 642390 339648 642490
rect 339748 642390 339872 642490
rect 339972 642390 340096 642490
rect 340196 642390 340320 642490
rect 340420 642390 340544 642490
rect 340644 642390 340768 642490
rect 340868 642390 340992 642490
rect 341092 642390 341216 642490
rect 341316 642390 341440 642490
rect 341540 642390 341664 642490
rect 341764 642390 341888 642490
rect 341988 642390 342112 642490
rect 342212 642390 342217 642490
rect 335560 642385 342217 642390
rect 298820 642251 305476 642365
rect 309290 642251 315946 642365
rect 335560 642271 342216 642385
rect 335560 642266 342217 642271
rect 298820 642246 305477 642251
rect 298820 642146 298876 642246
rect 298976 642146 299100 642246
rect 299200 642146 299324 642246
rect 299424 642146 299548 642246
rect 299648 642146 299772 642246
rect 299872 642146 299996 642246
rect 300096 642146 300220 642246
rect 300320 642146 300444 642246
rect 300544 642146 300668 642246
rect 300768 642146 300892 642246
rect 300992 642146 301116 642246
rect 301216 642146 301340 642246
rect 301440 642146 301564 642246
rect 301664 642146 301788 642246
rect 301888 642146 302012 642246
rect 302112 642146 302236 642246
rect 302336 642146 302460 642246
rect 302560 642146 302684 642246
rect 302784 642146 302908 642246
rect 303008 642146 303132 642246
rect 303232 642146 303356 642246
rect 303456 642146 303580 642246
rect 303680 642146 303804 642246
rect 303904 642146 304028 642246
rect 304128 642146 304252 642246
rect 304352 642146 304476 642246
rect 304576 642146 304700 642246
rect 304800 642146 304924 642246
rect 305024 642146 305148 642246
rect 305248 642146 305372 642246
rect 305472 642146 305477 642246
rect 298820 642141 305477 642146
rect 309290 642246 315947 642251
rect 309290 642146 309346 642246
rect 309446 642146 309570 642246
rect 309670 642146 309794 642246
rect 309894 642146 310018 642246
rect 310118 642146 310242 642246
rect 310342 642146 310466 642246
rect 310566 642146 310690 642246
rect 310790 642146 310914 642246
rect 311014 642146 311138 642246
rect 311238 642146 311362 642246
rect 311462 642146 311586 642246
rect 311686 642146 311810 642246
rect 311910 642146 312034 642246
rect 312134 642146 312258 642246
rect 312358 642146 312482 642246
rect 312582 642146 312706 642246
rect 312806 642146 312930 642246
rect 313030 642146 313154 642246
rect 313254 642146 313378 642246
rect 313478 642146 313602 642246
rect 313702 642146 313826 642246
rect 313926 642146 314050 642246
rect 314150 642146 314274 642246
rect 314374 642146 314498 642246
rect 314598 642146 314722 642246
rect 314822 642146 314946 642246
rect 315046 642146 315170 642246
rect 315270 642146 315394 642246
rect 315494 642146 315618 642246
rect 315718 642146 315842 642246
rect 315942 642146 315947 642246
rect 309290 642141 315947 642146
rect 335560 642166 335616 642266
rect 335716 642166 335840 642266
rect 335940 642166 336064 642266
rect 336164 642166 336288 642266
rect 336388 642166 336512 642266
rect 336612 642166 336736 642266
rect 336836 642166 336960 642266
rect 337060 642166 337184 642266
rect 337284 642166 337408 642266
rect 337508 642166 337632 642266
rect 337732 642166 337856 642266
rect 337956 642166 338080 642266
rect 338180 642166 338304 642266
rect 338404 642166 338528 642266
rect 338628 642166 338752 642266
rect 338852 642166 338976 642266
rect 339076 642166 339200 642266
rect 339300 642166 339424 642266
rect 339524 642166 339648 642266
rect 339748 642166 339872 642266
rect 339972 642166 340096 642266
rect 340196 642166 340320 642266
rect 340420 642166 340544 642266
rect 340644 642166 340768 642266
rect 340868 642166 340992 642266
rect 341092 642166 341216 642266
rect 341316 642166 341440 642266
rect 341540 642166 341664 642266
rect 341764 642166 341888 642266
rect 341988 642166 342112 642266
rect 342212 642166 342217 642266
rect 335560 642161 342217 642166
rect 298820 642027 305476 642141
rect 309290 642027 315946 642141
rect 335560 642047 342216 642161
rect 335560 642042 342217 642047
rect 298820 642022 305477 642027
rect 298820 641922 298876 642022
rect 298976 641922 299100 642022
rect 299200 641922 299324 642022
rect 299424 641922 299548 642022
rect 299648 641922 299772 642022
rect 299872 641922 299996 642022
rect 300096 641922 300220 642022
rect 300320 641922 300444 642022
rect 300544 641922 300668 642022
rect 300768 641922 300892 642022
rect 300992 641922 301116 642022
rect 301216 641922 301340 642022
rect 301440 641922 301564 642022
rect 301664 641922 301788 642022
rect 301888 641922 302012 642022
rect 302112 641922 302236 642022
rect 302336 641922 302460 642022
rect 302560 641922 302684 642022
rect 302784 641922 302908 642022
rect 303008 641922 303132 642022
rect 303232 641922 303356 642022
rect 303456 641922 303580 642022
rect 303680 641922 303804 642022
rect 303904 641922 304028 642022
rect 304128 641922 304252 642022
rect 304352 641922 304476 642022
rect 304576 641922 304700 642022
rect 304800 641922 304924 642022
rect 305024 641922 305148 642022
rect 305248 641922 305372 642022
rect 305472 641922 305477 642022
rect 298820 641917 305477 641922
rect 309290 642022 315947 642027
rect 309290 641922 309346 642022
rect 309446 641922 309570 642022
rect 309670 641922 309794 642022
rect 309894 641922 310018 642022
rect 310118 641922 310242 642022
rect 310342 641922 310466 642022
rect 310566 641922 310690 642022
rect 310790 641922 310914 642022
rect 311014 641922 311138 642022
rect 311238 641922 311362 642022
rect 311462 641922 311586 642022
rect 311686 641922 311810 642022
rect 311910 641922 312034 642022
rect 312134 641922 312258 642022
rect 312358 641922 312482 642022
rect 312582 641922 312706 642022
rect 312806 641922 312930 642022
rect 313030 641922 313154 642022
rect 313254 641922 313378 642022
rect 313478 641922 313602 642022
rect 313702 641922 313826 642022
rect 313926 641922 314050 642022
rect 314150 641922 314274 642022
rect 314374 641922 314498 642022
rect 314598 641922 314722 642022
rect 314822 641922 314946 642022
rect 315046 641922 315170 642022
rect 315270 641922 315394 642022
rect 315494 641922 315618 642022
rect 315718 641922 315842 642022
rect 315942 641922 315947 642022
rect 309290 641917 315947 641922
rect 335560 641942 335616 642042
rect 335716 641942 335840 642042
rect 335940 641942 336064 642042
rect 336164 641942 336288 642042
rect 336388 641942 336512 642042
rect 336612 641942 336736 642042
rect 336836 641942 336960 642042
rect 337060 641942 337184 642042
rect 337284 641942 337408 642042
rect 337508 641942 337632 642042
rect 337732 641942 337856 642042
rect 337956 641942 338080 642042
rect 338180 641942 338304 642042
rect 338404 641942 338528 642042
rect 338628 641942 338752 642042
rect 338852 641942 338976 642042
rect 339076 641942 339200 642042
rect 339300 641942 339424 642042
rect 339524 641942 339648 642042
rect 339748 641942 339872 642042
rect 339972 641942 340096 642042
rect 340196 641942 340320 642042
rect 340420 641942 340544 642042
rect 340644 641942 340768 642042
rect 340868 641942 340992 642042
rect 341092 641942 341216 642042
rect 341316 641942 341440 642042
rect 341540 641942 341664 642042
rect 341764 641942 341888 642042
rect 341988 641942 342112 642042
rect 342212 641942 342217 642042
rect 335560 641937 342217 641942
rect 298820 641803 305476 641917
rect 309290 641803 315946 641917
rect 335560 641823 342216 641937
rect 335560 641818 342217 641823
rect 298820 641798 305477 641803
rect 298820 641698 298876 641798
rect 298976 641698 299100 641798
rect 299200 641698 299324 641798
rect 299424 641698 299548 641798
rect 299648 641698 299772 641798
rect 299872 641698 299996 641798
rect 300096 641698 300220 641798
rect 300320 641698 300444 641798
rect 300544 641698 300668 641798
rect 300768 641698 300892 641798
rect 300992 641698 301116 641798
rect 301216 641698 301340 641798
rect 301440 641698 301564 641798
rect 301664 641698 301788 641798
rect 301888 641698 302012 641798
rect 302112 641698 302236 641798
rect 302336 641698 302460 641798
rect 302560 641698 302684 641798
rect 302784 641698 302908 641798
rect 303008 641698 303132 641798
rect 303232 641698 303356 641798
rect 303456 641698 303580 641798
rect 303680 641698 303804 641798
rect 303904 641698 304028 641798
rect 304128 641698 304252 641798
rect 304352 641698 304476 641798
rect 304576 641698 304700 641798
rect 304800 641698 304924 641798
rect 305024 641698 305148 641798
rect 305248 641698 305372 641798
rect 305472 641698 305477 641798
rect 298820 641693 305477 641698
rect 309290 641798 315947 641803
rect 309290 641698 309346 641798
rect 309446 641698 309570 641798
rect 309670 641698 309794 641798
rect 309894 641698 310018 641798
rect 310118 641698 310242 641798
rect 310342 641698 310466 641798
rect 310566 641698 310690 641798
rect 310790 641698 310914 641798
rect 311014 641698 311138 641798
rect 311238 641698 311362 641798
rect 311462 641698 311586 641798
rect 311686 641698 311810 641798
rect 311910 641698 312034 641798
rect 312134 641698 312258 641798
rect 312358 641698 312482 641798
rect 312582 641698 312706 641798
rect 312806 641698 312930 641798
rect 313030 641698 313154 641798
rect 313254 641698 313378 641798
rect 313478 641698 313602 641798
rect 313702 641698 313826 641798
rect 313926 641698 314050 641798
rect 314150 641698 314274 641798
rect 314374 641698 314498 641798
rect 314598 641698 314722 641798
rect 314822 641698 314946 641798
rect 315046 641698 315170 641798
rect 315270 641698 315394 641798
rect 315494 641698 315618 641798
rect 315718 641698 315842 641798
rect 315942 641698 315947 641798
rect 309290 641693 315947 641698
rect 335560 641718 335616 641818
rect 335716 641718 335840 641818
rect 335940 641718 336064 641818
rect 336164 641718 336288 641818
rect 336388 641718 336512 641818
rect 336612 641718 336736 641818
rect 336836 641718 336960 641818
rect 337060 641718 337184 641818
rect 337284 641718 337408 641818
rect 337508 641718 337632 641818
rect 337732 641718 337856 641818
rect 337956 641718 338080 641818
rect 338180 641718 338304 641818
rect 338404 641718 338528 641818
rect 338628 641718 338752 641818
rect 338852 641718 338976 641818
rect 339076 641718 339200 641818
rect 339300 641718 339424 641818
rect 339524 641718 339648 641818
rect 339748 641718 339872 641818
rect 339972 641718 340096 641818
rect 340196 641718 340320 641818
rect 340420 641718 340544 641818
rect 340644 641718 340768 641818
rect 340868 641718 340992 641818
rect 341092 641718 341216 641818
rect 341316 641718 341440 641818
rect 341540 641718 341664 641818
rect 341764 641718 341888 641818
rect 341988 641718 342112 641818
rect 342212 641718 342217 641818
rect 335560 641713 342217 641718
rect 298820 641664 305476 641693
rect 309290 641664 315946 641693
rect 335560 641684 342216 641713
rect 560425 639792 560582 644576
rect 566726 639792 566979 644576
rect 289020 637996 298880 638020
rect 342125 638000 342235 638001
rect 342349 638000 342459 638001
rect 342573 638000 342683 638001
rect 342797 638000 342907 638001
rect 343021 638000 343131 638001
rect 289020 637896 297850 637996
rect 297950 637896 298074 637996
rect 298174 637896 298298 637996
rect 298398 637896 298522 637996
rect 298622 637896 298746 637996
rect 298846 637896 298880 637996
rect 289020 637772 298880 637896
rect 289020 637672 297850 637772
rect 297950 637672 298074 637772
rect 298174 637672 298298 637772
rect 298398 637672 298522 637772
rect 298622 637672 298746 637772
rect 298846 637672 298880 637772
rect 289020 637548 298880 637672
rect 289020 637448 297850 637548
rect 297950 637448 298074 637548
rect 298174 637448 298298 637548
rect 298398 637448 298522 637548
rect 298622 637448 298746 637548
rect 298846 637448 298880 637548
rect 289020 637324 298880 637448
rect 289020 637224 297850 637324
rect 297950 637224 298074 637324
rect 298174 637224 298298 637324
rect 298398 637224 298522 637324
rect 298622 637224 298746 637324
rect 298846 637224 298880 637324
rect 289020 637184 298880 637224
rect 289020 631440 289920 637184
rect 294704 637100 298880 637184
rect 294704 637000 297850 637100
rect 297950 637000 298074 637100
rect 298174 637000 298298 637100
rect 298398 637000 298522 637100
rect 298622 637000 298746 637100
rect 298846 637000 298880 637100
rect 294704 636876 298880 637000
rect 294704 636776 297850 636876
rect 297950 636776 298074 636876
rect 298174 636776 298298 636876
rect 298398 636776 298522 636876
rect 298622 636776 298746 636876
rect 298846 636776 298880 636876
rect 294704 636652 298880 636776
rect 294704 636552 297850 636652
rect 297950 636552 298074 636652
rect 298174 636552 298298 636652
rect 298398 636552 298522 636652
rect 298622 636552 298746 636652
rect 298846 636552 298880 636652
rect 294704 636428 298880 636552
rect 294704 636328 297850 636428
rect 297950 636328 298074 636428
rect 298174 636328 298298 636428
rect 298398 636328 298522 636428
rect 298622 636328 298746 636428
rect 298846 636328 298880 636428
rect 294704 636204 298880 636328
rect 294704 636104 297850 636204
rect 297950 636104 298074 636204
rect 298174 636104 298298 636204
rect 298398 636104 298522 636204
rect 298622 636104 298746 636204
rect 298846 636104 298880 636204
rect 294704 635980 298880 636104
rect 294704 635880 297850 635980
rect 297950 635880 298074 635980
rect 298174 635880 298298 635980
rect 298398 635880 298522 635980
rect 298622 635880 298746 635980
rect 298846 635880 298880 635980
rect 294704 635756 298880 635880
rect 294704 635656 297850 635756
rect 297950 635656 298074 635756
rect 298174 635656 298298 635756
rect 298398 635656 298522 635756
rect 298622 635656 298746 635756
rect 298846 635656 298880 635756
rect 294704 635532 298880 635656
rect 294704 635432 297850 635532
rect 297950 635432 298074 635532
rect 298174 635432 298298 635532
rect 298398 635432 298522 635532
rect 298622 635432 298746 635532
rect 298846 635432 298880 635532
rect 294704 635308 298880 635432
rect 294704 635208 297850 635308
rect 297950 635208 298074 635308
rect 298174 635208 298298 635308
rect 298398 635208 298522 635308
rect 298622 635208 298746 635308
rect 298846 635208 298880 635308
rect 294704 635084 298880 635208
rect 294704 634984 297850 635084
rect 297950 634984 298074 635084
rect 298174 634984 298298 635084
rect 298398 634984 298522 635084
rect 298622 634984 298746 635084
rect 298846 634984 298880 635084
rect 294704 634860 298880 634984
rect 294704 634760 297850 634860
rect 297950 634760 298074 634860
rect 298174 634760 298298 634860
rect 298398 634760 298522 634860
rect 298622 634760 298746 634860
rect 298846 634760 298880 634860
rect 294704 634636 298880 634760
rect 294704 634536 297850 634636
rect 297950 634536 298074 634636
rect 298174 634536 298298 634636
rect 298398 634536 298522 634636
rect 298622 634536 298746 634636
rect 298846 634536 298880 634636
rect 294704 634412 298880 634536
rect 294704 634312 297850 634412
rect 297950 634312 298074 634412
rect 298174 634312 298298 634412
rect 298398 634312 298522 634412
rect 298622 634312 298746 634412
rect 298846 634312 298880 634412
rect 294704 634188 298880 634312
rect 294704 634088 297850 634188
rect 297950 634088 298074 634188
rect 298174 634088 298298 634188
rect 298398 634088 298522 634188
rect 298622 634088 298746 634188
rect 298846 634088 298880 634188
rect 294704 633964 298880 634088
rect 294704 633864 297850 633964
rect 297950 633864 298074 633964
rect 298174 633864 298298 633964
rect 298398 633864 298522 633964
rect 298622 633864 298746 633964
rect 298846 633864 298880 633964
rect 294704 633740 298880 633864
rect 294704 633640 297850 633740
rect 297950 633640 298074 633740
rect 298174 633640 298298 633740
rect 298398 633640 298522 633740
rect 298622 633640 298746 633740
rect 298846 633640 298880 633740
rect 294704 633516 298880 633640
rect 294704 633416 297850 633516
rect 297950 633416 298074 633516
rect 298174 633416 298298 633516
rect 298398 633416 298522 633516
rect 298622 633416 298746 633516
rect 298846 633416 298880 633516
rect 294704 633292 298880 633416
rect 294704 633192 297850 633292
rect 297950 633192 298074 633292
rect 298174 633192 298298 633292
rect 298398 633192 298522 633292
rect 298622 633192 298746 633292
rect 298846 633192 298880 633292
rect 294704 633068 298880 633192
rect 294704 632968 297850 633068
rect 297950 632968 298074 633068
rect 298174 632968 298298 633068
rect 298398 632968 298522 633068
rect 298622 632968 298746 633068
rect 298846 632968 298880 633068
rect 294704 632844 298880 632968
rect 294704 632744 297850 632844
rect 297950 632744 298074 632844
rect 298174 632744 298298 632844
rect 298398 632744 298522 632844
rect 298622 632744 298746 632844
rect 298846 632744 298880 632844
rect 294704 632620 298880 632744
rect 294704 632520 297850 632620
rect 297950 632520 298074 632620
rect 298174 632520 298298 632620
rect 298398 632520 298522 632620
rect 298622 632520 298746 632620
rect 298846 632520 298880 632620
rect 294704 632396 298880 632520
rect 294704 632296 297850 632396
rect 297950 632296 298074 632396
rect 298174 632296 298298 632396
rect 298398 632296 298522 632396
rect 298622 632296 298746 632396
rect 298846 632296 298880 632396
rect 294704 632172 298880 632296
rect 294704 632072 297850 632172
rect 297950 632072 298074 632172
rect 298174 632072 298298 632172
rect 298398 632072 298522 632172
rect 298622 632072 298746 632172
rect 298846 632072 298880 632172
rect 294704 631948 298880 632072
rect 294704 631848 297850 631948
rect 297950 631848 298074 631948
rect 298174 631848 298298 631948
rect 298398 631848 298522 631948
rect 298622 631848 298746 631948
rect 298846 631848 298880 631948
rect 294704 631724 298880 631848
rect 294704 631624 297850 631724
rect 297950 631624 298074 631724
rect 298174 631624 298298 631724
rect 298398 631624 298522 631724
rect 298622 631624 298746 631724
rect 298846 631624 298880 631724
rect 294704 631500 298880 631624
rect 294704 631440 297850 631500
rect 289020 631400 297850 631440
rect 297950 631400 298074 631500
rect 298174 631400 298298 631500
rect 298398 631400 298522 631500
rect 298622 631400 298746 631500
rect 298846 631400 298880 631500
rect 289020 631340 298880 631400
rect 341994 637996 525800 638000
rect 341994 637896 342130 637996
rect 342230 637896 342354 637996
rect 342454 637896 342578 637996
rect 342678 637896 342802 637996
rect 342902 637896 343026 637996
rect 343126 637896 525800 637996
rect 341994 637772 525800 637896
rect 341994 637672 342130 637772
rect 342230 637672 342354 637772
rect 342454 637672 342578 637772
rect 342678 637672 342802 637772
rect 342902 637672 343026 637772
rect 343126 637672 525800 637772
rect 341994 637561 525800 637672
rect 341994 637548 510602 637561
rect 341994 637448 342130 637548
rect 342230 637448 342354 637548
rect 342454 637448 342578 637548
rect 342678 637448 342802 637548
rect 342902 637448 343026 637548
rect 343126 637448 510602 637548
rect 341994 637324 510602 637448
rect 341994 637224 342130 637324
rect 342230 637224 342354 637324
rect 342454 637224 342578 637324
rect 342678 637224 342802 637324
rect 342902 637224 343026 637324
rect 343126 637224 510602 637324
rect 341994 637100 510602 637224
rect 341994 637000 342130 637100
rect 342230 637000 342354 637100
rect 342454 637000 342578 637100
rect 342678 637000 342802 637100
rect 342902 637000 343026 637100
rect 343126 637000 510602 637100
rect 341994 636876 510602 637000
rect 341994 636776 342130 636876
rect 342230 636776 342354 636876
rect 342454 636776 342578 636876
rect 342678 636776 342802 636876
rect 342902 636776 343026 636876
rect 343126 636776 510602 636876
rect 341994 636652 510602 636776
rect 341994 636552 342130 636652
rect 342230 636552 342354 636652
rect 342454 636552 342578 636652
rect 342678 636552 342802 636652
rect 342902 636552 343026 636652
rect 343126 636552 510602 636652
rect 341994 636428 510602 636552
rect 341994 636328 342130 636428
rect 342230 636328 342354 636428
rect 342454 636328 342578 636428
rect 342678 636328 342802 636428
rect 342902 636328 343026 636428
rect 343126 636328 510602 636428
rect 341994 636204 510602 636328
rect 341994 636104 342130 636204
rect 342230 636104 342354 636204
rect 342454 636104 342578 636204
rect 342678 636104 342802 636204
rect 342902 636104 343026 636204
rect 343126 636104 510602 636204
rect 341994 635980 510602 636104
rect 341994 635880 342130 635980
rect 342230 635880 342354 635980
rect 342454 635880 342578 635980
rect 342678 635880 342802 635980
rect 342902 635880 343026 635980
rect 343126 635880 510602 635980
rect 341994 635756 510602 635880
rect 341994 635656 342130 635756
rect 342230 635656 342354 635756
rect 342454 635656 342578 635756
rect 342678 635656 342802 635756
rect 342902 635656 343026 635756
rect 343126 635656 510602 635756
rect 341994 635532 510602 635656
rect 341994 635432 342130 635532
rect 342230 635432 342354 635532
rect 342454 635432 342578 635532
rect 342678 635432 342802 635532
rect 342902 635432 343026 635532
rect 343126 635432 510602 635532
rect 341994 635308 510602 635432
rect 341994 635208 342130 635308
rect 342230 635208 342354 635308
rect 342454 635208 342578 635308
rect 342678 635208 342802 635308
rect 342902 635208 343026 635308
rect 343126 635208 510602 635308
rect 341994 635084 510602 635208
rect 341994 634984 342130 635084
rect 342230 634984 342354 635084
rect 342454 634984 342578 635084
rect 342678 634984 342802 635084
rect 342902 634984 343026 635084
rect 343126 634984 510602 635084
rect 341994 634860 510602 634984
rect 341994 634760 342130 634860
rect 342230 634760 342354 634860
rect 342454 634760 342578 634860
rect 342678 634760 342802 634860
rect 342902 634760 343026 634860
rect 343126 634760 510602 634860
rect 341994 634636 510602 634760
rect 341994 634536 342130 634636
rect 342230 634536 342354 634636
rect 342454 634536 342578 634636
rect 342678 634536 342802 634636
rect 342902 634536 343026 634636
rect 343126 634536 510602 634636
rect 341994 634412 510602 634536
rect 341994 634312 342130 634412
rect 342230 634312 342354 634412
rect 342454 634312 342578 634412
rect 342678 634312 342802 634412
rect 342902 634312 343026 634412
rect 343126 634312 510602 634412
rect 341994 634188 510602 634312
rect 341994 634088 342130 634188
rect 342230 634088 342354 634188
rect 342454 634088 342578 634188
rect 342678 634088 342802 634188
rect 342902 634088 343026 634188
rect 343126 634088 510602 634188
rect 341994 633964 510602 634088
rect 341994 633864 342130 633964
rect 342230 633864 342354 633964
rect 342454 633864 342578 633964
rect 342678 633864 342802 633964
rect 342902 633864 343026 633964
rect 343126 633864 510602 633964
rect 341994 633740 510602 633864
rect 341994 633640 342130 633740
rect 342230 633640 342354 633740
rect 342454 633640 342578 633740
rect 342678 633640 342802 633740
rect 342902 633640 343026 633740
rect 343126 633640 510602 633740
rect 341994 633516 510602 633640
rect 341994 633416 342130 633516
rect 342230 633416 342354 633516
rect 342454 633416 342578 633516
rect 342678 633416 342802 633516
rect 342902 633416 343026 633516
rect 343126 633416 510602 633516
rect 341994 633292 510602 633416
rect 341994 633192 342130 633292
rect 342230 633192 342354 633292
rect 342454 633192 342578 633292
rect 342678 633192 342802 633292
rect 342902 633192 343026 633292
rect 343126 633192 510602 633292
rect 341994 633068 510602 633192
rect 341994 632968 342130 633068
rect 342230 632968 342354 633068
rect 342454 632968 342578 633068
rect 342678 632968 342802 633068
rect 342902 632968 343026 633068
rect 343126 632968 510602 633068
rect 341994 632844 510602 632968
rect 341994 632744 342130 632844
rect 342230 632744 342354 632844
rect 342454 632744 342578 632844
rect 342678 632744 342802 632844
rect 342902 632744 343026 632844
rect 343126 632744 510602 632844
rect 341994 632620 510602 632744
rect 341994 632520 342130 632620
rect 342230 632520 342354 632620
rect 342454 632520 342578 632620
rect 342678 632520 342802 632620
rect 342902 632520 343026 632620
rect 343126 632520 510602 632620
rect 341994 632396 510602 632520
rect 341994 632296 342130 632396
rect 342230 632296 342354 632396
rect 342454 632296 342578 632396
rect 342678 632296 342802 632396
rect 342902 632296 343026 632396
rect 343126 632296 510602 632396
rect 341994 632172 510602 632296
rect 341994 632072 342130 632172
rect 342230 632072 342354 632172
rect 342454 632072 342578 632172
rect 342678 632072 342802 632172
rect 342902 632072 343026 632172
rect 343126 632072 510602 632172
rect 341994 631948 510602 632072
rect 341994 631848 342130 631948
rect 342230 631848 342354 631948
rect 342454 631848 342578 631948
rect 342678 631848 342802 631948
rect 342902 631848 343026 631948
rect 343126 631848 510602 631948
rect 341994 631817 510602 631848
rect 515386 631817 520602 637561
rect 525386 631817 525800 637561
rect 341994 631724 525800 631817
rect 341994 631624 342130 631724
rect 342230 631624 342354 631724
rect 342454 631624 342578 631724
rect 342678 631624 342802 631724
rect 342902 631624 343026 631724
rect 343126 631624 525800 631724
rect 341994 631500 525800 631624
rect 341994 631400 342130 631500
rect 342230 631400 342354 631500
rect 342454 631400 342578 631500
rect 342678 631400 342802 631500
rect 342902 631400 343026 631500
rect 343126 631400 525800 631500
rect 341994 631344 525800 631400
rect 560425 634576 566979 639792
rect 560425 629792 560582 634576
rect 566726 629792 566979 634576
rect 319399 628868 319601 628869
rect 319399 628668 319400 628868
rect 319600 628668 319601 628868
rect 319399 628667 319601 628668
rect 319833 628868 320035 628869
rect 319833 628668 319834 628868
rect 320034 628668 320035 628868
rect 319833 628667 320035 628668
rect 320267 628868 320469 628869
rect 320267 628668 320268 628868
rect 320468 628668 320469 628868
rect 320267 628667 320469 628668
rect 320701 628868 320903 628869
rect 320701 628668 320702 628868
rect 320902 628668 320903 628868
rect 320701 628667 320903 628668
rect 321135 628868 321337 628869
rect 321135 628668 321136 628868
rect 321336 628668 321337 628868
rect 321135 628667 321337 628668
rect 321569 628868 321771 628869
rect 321569 628668 321570 628868
rect 321770 628668 321771 628868
rect 321569 628667 321771 628668
rect 322003 628868 322205 628869
rect 322003 628668 322004 628868
rect 322204 628668 322205 628868
rect 322003 628667 322205 628668
rect 322437 628868 322639 628869
rect 322437 628668 322438 628868
rect 322638 628668 322639 628868
rect 322437 628667 322639 628668
rect 322871 628868 323073 628869
rect 322871 628668 322872 628868
rect 323072 628668 323073 628868
rect 322871 628667 323073 628668
rect 323305 628868 323507 628869
rect 323305 628668 323306 628868
rect 323506 628668 323507 628868
rect 323305 628667 323507 628668
rect 323739 628868 323941 628869
rect 323739 628668 323740 628868
rect 323940 628668 323941 628868
rect 323739 628667 323941 628668
rect 324139 628868 324341 628869
rect 324139 628668 324140 628868
rect 324340 628668 324341 628868
rect 324139 628667 324341 628668
rect 324539 628868 324741 628869
rect 324539 628668 324540 628868
rect 324740 628668 324741 628868
rect 324539 628667 324741 628668
rect 324939 628868 325141 628869
rect 324939 628668 324940 628868
rect 325140 628668 325141 628868
rect 324939 628667 325141 628668
rect 325339 628868 325541 628869
rect 325339 628668 325340 628868
rect 325540 628668 325541 628868
rect 325339 628667 325541 628668
rect 325739 628868 325941 628869
rect 325739 628668 325740 628868
rect 325940 628668 325941 628868
rect 325739 628667 325941 628668
rect 326139 628868 326341 628869
rect 326139 628668 326140 628868
rect 326340 628668 326341 628868
rect 326139 628667 326341 628668
rect 326539 628868 326741 628869
rect 326539 628668 326540 628868
rect 326740 628668 326741 628868
rect 326539 628667 326741 628668
rect 326939 628868 327141 628869
rect 326939 628668 326940 628868
rect 327140 628668 327141 628868
rect 326939 628667 327141 628668
rect 327339 628868 327541 628869
rect 327339 628668 327340 628868
rect 327540 628668 327541 628868
rect 327339 628667 327541 628668
rect 328939 628868 329141 628869
rect 328939 628668 328940 628868
rect 329140 628668 329141 628868
rect 328939 628667 329141 628668
rect 329339 628868 329541 628869
rect 329339 628668 329340 628868
rect 329540 628668 329541 628868
rect 329339 628667 329541 628668
rect 329739 628868 329941 628869
rect 329739 628668 329740 628868
rect 329940 628668 329941 628868
rect 329739 628667 329941 628668
rect 330139 628868 330341 628869
rect 330139 628668 330140 628868
rect 330340 628668 330341 628868
rect 330139 628667 330341 628668
rect 330539 628868 330741 628869
rect 330539 628668 330540 628868
rect 330740 628668 330741 628868
rect 330539 628667 330741 628668
rect 330939 628868 331141 628869
rect 330939 628668 330940 628868
rect 331140 628668 331141 628868
rect 330939 628667 331141 628668
rect 331339 628868 331541 628869
rect 331339 628668 331340 628868
rect 331540 628668 331541 628868
rect 331339 628667 331541 628668
rect 331739 628868 331941 628869
rect 331739 628668 331740 628868
rect 331940 628668 331941 628868
rect 331739 628667 331941 628668
rect 332139 628868 332341 628869
rect 332139 628668 332140 628868
rect 332340 628668 332341 628868
rect 332139 628667 332341 628668
rect 319399 628434 319601 628435
rect 319399 628234 319400 628434
rect 319600 628234 319601 628434
rect 319399 628233 319601 628234
rect 319833 628434 320035 628435
rect 319833 628234 319834 628434
rect 320034 628234 320035 628434
rect 319833 628233 320035 628234
rect 320267 628434 320469 628435
rect 320267 628234 320268 628434
rect 320468 628234 320469 628434
rect 320267 628233 320469 628234
rect 320701 628434 320903 628435
rect 320701 628234 320702 628434
rect 320902 628234 320903 628434
rect 320701 628233 320903 628234
rect 321135 628434 321337 628435
rect 321135 628234 321136 628434
rect 321336 628234 321337 628434
rect 321135 628233 321337 628234
rect 321569 628434 321771 628435
rect 321569 628234 321570 628434
rect 321770 628234 321771 628434
rect 321569 628233 321771 628234
rect 322003 628434 322205 628435
rect 322003 628234 322004 628434
rect 322204 628234 322205 628434
rect 322003 628233 322205 628234
rect 322437 628434 322639 628435
rect 322437 628234 322438 628434
rect 322638 628234 322639 628434
rect 322437 628233 322639 628234
rect 322871 628434 323073 628435
rect 322871 628234 322872 628434
rect 323072 628234 323073 628434
rect 322871 628233 323073 628234
rect 323305 628434 323507 628435
rect 323305 628234 323306 628434
rect 323506 628234 323507 628434
rect 323305 628233 323507 628234
rect 323739 628434 323941 628435
rect 323739 628234 323740 628434
rect 323940 628234 323941 628434
rect 323739 628233 323941 628234
rect 319399 628000 319601 628001
rect 319399 627800 319400 628000
rect 319600 627800 319601 628000
rect 319399 627799 319601 627800
rect 319833 628000 320035 628001
rect 319833 627800 319834 628000
rect 320034 627800 320035 628000
rect 319833 627799 320035 627800
rect 320267 628000 320469 628001
rect 320267 627800 320268 628000
rect 320468 627800 320469 628000
rect 320267 627799 320469 627800
rect 320701 628000 320903 628001
rect 320701 627800 320702 628000
rect 320902 627800 320903 628000
rect 320701 627799 320903 627800
rect 321135 628000 321337 628001
rect 321135 627800 321136 628000
rect 321336 627800 321337 628000
rect 321135 627799 321337 627800
rect 321569 628000 321771 628001
rect 321569 627800 321570 628000
rect 321770 627800 321771 628000
rect 321569 627799 321771 627800
rect 322003 628000 322205 628001
rect 322003 627800 322004 628000
rect 322204 627800 322205 628000
rect 322003 627799 322205 627800
rect 322437 628000 322639 628001
rect 322437 627800 322438 628000
rect 322638 627800 322639 628000
rect 322437 627799 322639 627800
rect 322871 628000 323073 628001
rect 322871 627800 322872 628000
rect 323072 627800 323073 628000
rect 322871 627799 323073 627800
rect 323305 628000 323507 628001
rect 323305 627800 323306 628000
rect 323506 627800 323507 628000
rect 323305 627799 323507 627800
rect 323739 628000 323941 628001
rect 323739 627800 323740 628000
rect 323940 627800 323941 628000
rect 323739 627799 323941 627800
rect 217216 626176 299008 626240
rect 217216 626112 217344 626176
rect 217408 626112 217472 626176
rect 217536 626112 217600 626176
rect 217664 626112 217728 626176
rect 217792 626112 217856 626176
rect 217920 626112 217984 626176
rect 218048 626112 218112 626176
rect 218176 626112 218240 626176
rect 218304 626112 218368 626176
rect 218432 626112 218496 626176
rect 218560 626112 218624 626176
rect 218688 626112 218752 626176
rect 218816 626112 218880 626176
rect 218944 626112 219008 626176
rect 219072 626112 219136 626176
rect 219200 626112 219264 626176
rect 219328 626112 219392 626176
rect 219456 626112 219520 626176
rect 219584 626112 219648 626176
rect 219712 626112 219776 626176
rect 219840 626112 219904 626176
rect 219968 626112 220032 626176
rect 220096 626112 220160 626176
rect 220224 626112 220288 626176
rect 220352 626112 220416 626176
rect 220480 626112 220544 626176
rect 220608 626112 220672 626176
rect 220736 626112 220800 626176
rect 220864 626112 220928 626176
rect 220992 626112 221056 626176
rect 221120 626112 221184 626176
rect 221248 626112 221312 626176
rect 221376 626112 221440 626176
rect 221504 626112 221568 626176
rect 221632 626112 221696 626176
rect 221760 626112 221824 626176
rect 221888 626112 221952 626176
rect 222016 626112 222080 626176
rect 222144 626112 227640 626176
rect 227704 626112 227768 626176
rect 227832 626112 227896 626176
rect 227960 626112 228024 626176
rect 228088 626112 228152 626176
rect 228216 626112 228280 626176
rect 228344 626112 228408 626176
rect 228472 626112 228536 626176
rect 228600 626112 228664 626176
rect 228728 626112 228792 626176
rect 228856 626112 228920 626176
rect 228984 626112 229048 626176
rect 229112 626112 229176 626176
rect 229240 626112 229304 626176
rect 229368 626112 229432 626176
rect 229496 626112 229560 626176
rect 229624 626112 229688 626176
rect 229752 626112 229816 626176
rect 229880 626112 229944 626176
rect 230008 626112 230072 626176
rect 230136 626112 230200 626176
rect 230264 626112 230328 626176
rect 230392 626112 230456 626176
rect 230520 626112 230584 626176
rect 230648 626112 230712 626176
rect 230776 626112 230840 626176
rect 230904 626112 230968 626176
rect 231032 626112 231096 626176
rect 231160 626112 231224 626176
rect 231288 626112 231352 626176
rect 231416 626112 231480 626176
rect 231544 626112 231608 626176
rect 231672 626112 231736 626176
rect 231800 626112 231864 626176
rect 231928 626112 231992 626176
rect 232056 626112 232120 626176
rect 232184 626112 232248 626176
rect 232312 626112 232376 626176
rect 232440 626112 297856 626176
rect 297920 626112 297984 626176
rect 298048 626112 298112 626176
rect 298176 626112 298240 626176
rect 298304 626112 298368 626176
rect 298432 626112 298496 626176
rect 298560 626112 298624 626176
rect 298688 626112 298752 626176
rect 298816 626112 298880 626176
rect 298944 626112 299008 626176
rect 217216 626048 299008 626112
rect 217216 625984 217344 626048
rect 217408 625984 217472 626048
rect 217536 625984 217600 626048
rect 217664 625984 217728 626048
rect 217792 625984 217856 626048
rect 217920 625984 217984 626048
rect 218048 625984 218112 626048
rect 218176 625984 218240 626048
rect 218304 625984 218368 626048
rect 218432 625984 218496 626048
rect 218560 625984 218624 626048
rect 218688 625984 218752 626048
rect 218816 625984 218880 626048
rect 218944 625984 219008 626048
rect 219072 625984 219136 626048
rect 219200 625984 219264 626048
rect 219328 625984 219392 626048
rect 219456 625984 219520 626048
rect 219584 625984 219648 626048
rect 219712 625984 219776 626048
rect 219840 625984 219904 626048
rect 219968 625984 220032 626048
rect 220096 625984 220160 626048
rect 220224 625984 220288 626048
rect 220352 625984 220416 626048
rect 220480 625984 220544 626048
rect 220608 625984 220672 626048
rect 220736 625984 220800 626048
rect 220864 625984 220928 626048
rect 220992 625984 221056 626048
rect 221120 625984 221184 626048
rect 221248 625984 221312 626048
rect 221376 625984 221440 626048
rect 221504 625984 221568 626048
rect 221632 625984 221696 626048
rect 221760 625984 221824 626048
rect 221888 625984 221952 626048
rect 222016 625984 222080 626048
rect 222144 625984 227640 626048
rect 227704 625984 227768 626048
rect 227832 625984 227896 626048
rect 227960 625984 228024 626048
rect 228088 625984 228152 626048
rect 228216 625984 228280 626048
rect 228344 625984 228408 626048
rect 228472 625984 228536 626048
rect 228600 625984 228664 626048
rect 228728 625984 228792 626048
rect 228856 625984 228920 626048
rect 228984 625984 229048 626048
rect 229112 625984 229176 626048
rect 229240 625984 229304 626048
rect 229368 625984 229432 626048
rect 229496 625984 229560 626048
rect 229624 625984 229688 626048
rect 229752 625984 229816 626048
rect 229880 625984 229944 626048
rect 230008 625984 230072 626048
rect 230136 625984 230200 626048
rect 230264 625984 230328 626048
rect 230392 625984 230456 626048
rect 230520 625984 230584 626048
rect 230648 625984 230712 626048
rect 230776 625984 230840 626048
rect 230904 625984 230968 626048
rect 231032 625984 231096 626048
rect 231160 625984 231224 626048
rect 231288 625984 231352 626048
rect 231416 625984 231480 626048
rect 231544 625984 231608 626048
rect 231672 625984 231736 626048
rect 231800 625984 231864 626048
rect 231928 625984 231992 626048
rect 232056 625984 232120 626048
rect 232184 625984 232248 626048
rect 232312 625984 232376 626048
rect 232440 625984 297856 626048
rect 297920 625984 297984 626048
rect 298048 625984 298112 626048
rect 298176 625984 298240 626048
rect 298304 625984 298368 626048
rect 298432 625984 298496 626048
rect 298560 625984 298624 626048
rect 298688 625984 298752 626048
rect 298816 625984 298880 626048
rect 298944 625984 299008 626048
rect 217216 625920 299008 625984
rect 217216 625856 217344 625920
rect 217408 625856 217472 625920
rect 217536 625856 217600 625920
rect 217664 625856 217728 625920
rect 217792 625856 217856 625920
rect 217920 625856 217984 625920
rect 218048 625856 218112 625920
rect 218176 625856 218240 625920
rect 218304 625856 218368 625920
rect 218432 625856 218496 625920
rect 218560 625856 218624 625920
rect 218688 625856 218752 625920
rect 218816 625856 218880 625920
rect 218944 625856 219008 625920
rect 219072 625856 219136 625920
rect 219200 625856 219264 625920
rect 219328 625856 219392 625920
rect 219456 625856 219520 625920
rect 219584 625856 219648 625920
rect 219712 625856 219776 625920
rect 219840 625856 219904 625920
rect 219968 625856 220032 625920
rect 220096 625856 220160 625920
rect 220224 625856 220288 625920
rect 220352 625856 220416 625920
rect 220480 625856 220544 625920
rect 220608 625856 220672 625920
rect 220736 625856 220800 625920
rect 220864 625856 220928 625920
rect 220992 625856 221056 625920
rect 221120 625856 221184 625920
rect 221248 625856 221312 625920
rect 221376 625856 221440 625920
rect 221504 625856 221568 625920
rect 221632 625856 221696 625920
rect 221760 625856 221824 625920
rect 221888 625856 221952 625920
rect 222016 625856 222080 625920
rect 222144 625856 227640 625920
rect 227704 625856 227768 625920
rect 227832 625856 227896 625920
rect 227960 625856 228024 625920
rect 228088 625856 228152 625920
rect 228216 625856 228280 625920
rect 228344 625856 228408 625920
rect 228472 625856 228536 625920
rect 228600 625856 228664 625920
rect 228728 625856 228792 625920
rect 228856 625856 228920 625920
rect 228984 625856 229048 625920
rect 229112 625856 229176 625920
rect 229240 625856 229304 625920
rect 229368 625856 229432 625920
rect 229496 625856 229560 625920
rect 229624 625856 229688 625920
rect 229752 625856 229816 625920
rect 229880 625856 229944 625920
rect 230008 625856 230072 625920
rect 230136 625856 230200 625920
rect 230264 625856 230328 625920
rect 230392 625856 230456 625920
rect 230520 625856 230584 625920
rect 230648 625856 230712 625920
rect 230776 625856 230840 625920
rect 230904 625856 230968 625920
rect 231032 625856 231096 625920
rect 231160 625856 231224 625920
rect 231288 625856 231352 625920
rect 231416 625856 231480 625920
rect 231544 625856 231608 625920
rect 231672 625856 231736 625920
rect 231800 625856 231864 625920
rect 231928 625856 231992 625920
rect 232056 625856 232120 625920
rect 232184 625856 232248 625920
rect 232312 625856 232376 625920
rect 232440 625856 297856 625920
rect 297920 625856 297984 625920
rect 298048 625856 298112 625920
rect 298176 625856 298240 625920
rect 298304 625856 298368 625920
rect 298432 625856 298496 625920
rect 298560 625856 298624 625920
rect 298688 625856 298752 625920
rect 298816 625856 298880 625920
rect 298944 625856 299008 625920
rect 217216 625792 299008 625856
rect 217216 625728 217344 625792
rect 217408 625728 217472 625792
rect 217536 625728 217600 625792
rect 217664 625728 217728 625792
rect 217792 625728 217856 625792
rect 217920 625728 217984 625792
rect 218048 625728 218112 625792
rect 218176 625728 218240 625792
rect 218304 625728 218368 625792
rect 218432 625728 218496 625792
rect 218560 625728 218624 625792
rect 218688 625728 218752 625792
rect 218816 625728 218880 625792
rect 218944 625728 219008 625792
rect 219072 625728 219136 625792
rect 219200 625728 219264 625792
rect 219328 625728 219392 625792
rect 219456 625728 219520 625792
rect 219584 625728 219648 625792
rect 219712 625728 219776 625792
rect 219840 625728 219904 625792
rect 219968 625728 220032 625792
rect 220096 625728 220160 625792
rect 220224 625728 220288 625792
rect 220352 625728 220416 625792
rect 220480 625728 220544 625792
rect 220608 625728 220672 625792
rect 220736 625728 220800 625792
rect 220864 625728 220928 625792
rect 220992 625728 221056 625792
rect 221120 625728 221184 625792
rect 221248 625728 221312 625792
rect 221376 625728 221440 625792
rect 221504 625728 221568 625792
rect 221632 625728 221696 625792
rect 221760 625728 221824 625792
rect 221888 625728 221952 625792
rect 222016 625728 222080 625792
rect 222144 625728 227640 625792
rect 227704 625728 227768 625792
rect 227832 625728 227896 625792
rect 227960 625728 228024 625792
rect 228088 625728 228152 625792
rect 228216 625728 228280 625792
rect 228344 625728 228408 625792
rect 228472 625728 228536 625792
rect 228600 625728 228664 625792
rect 228728 625728 228792 625792
rect 228856 625728 228920 625792
rect 228984 625728 229048 625792
rect 229112 625728 229176 625792
rect 229240 625728 229304 625792
rect 229368 625728 229432 625792
rect 229496 625728 229560 625792
rect 229624 625728 229688 625792
rect 229752 625728 229816 625792
rect 229880 625728 229944 625792
rect 230008 625728 230072 625792
rect 230136 625728 230200 625792
rect 230264 625728 230328 625792
rect 230392 625728 230456 625792
rect 230520 625728 230584 625792
rect 230648 625728 230712 625792
rect 230776 625728 230840 625792
rect 230904 625728 230968 625792
rect 231032 625728 231096 625792
rect 231160 625728 231224 625792
rect 231288 625728 231352 625792
rect 231416 625728 231480 625792
rect 231544 625728 231608 625792
rect 231672 625728 231736 625792
rect 231800 625728 231864 625792
rect 231928 625728 231992 625792
rect 232056 625728 232120 625792
rect 232184 625728 232248 625792
rect 232312 625728 232376 625792
rect 232440 625728 297856 625792
rect 297920 625728 297984 625792
rect 298048 625728 298112 625792
rect 298176 625728 298240 625792
rect 298304 625728 298368 625792
rect 298432 625728 298496 625792
rect 298560 625728 298624 625792
rect 298688 625728 298752 625792
rect 298816 625728 298880 625792
rect 298944 625728 299008 625792
rect 217216 625664 299008 625728
rect 289020 624596 298880 624620
rect 289020 624496 297850 624596
rect 297950 624496 298074 624596
rect 298174 624496 298298 624596
rect 298398 624496 298522 624596
rect 298622 624496 298746 624596
rect 298846 624496 298880 624596
rect 289020 624372 298880 624496
rect 289020 624272 297850 624372
rect 297950 624272 298074 624372
rect 298174 624272 298298 624372
rect 298398 624272 298522 624372
rect 298622 624272 298746 624372
rect 298846 624272 298880 624372
rect 289020 624148 298880 624272
rect 289020 624048 297850 624148
rect 297950 624048 298074 624148
rect 298174 624048 298298 624148
rect 298398 624048 298522 624148
rect 298622 624048 298746 624148
rect 298846 624048 298880 624148
rect 289020 623924 298880 624048
rect 289020 623824 297850 623924
rect 297950 623824 298074 623924
rect 298174 623824 298298 623924
rect 298398 623824 298522 623924
rect 298622 623824 298746 623924
rect 298846 623824 298880 623924
rect 289020 623784 298880 623824
rect 289020 618040 289920 623784
rect 294704 623700 298880 623784
rect 294704 623600 297850 623700
rect 297950 623600 298074 623700
rect 298174 623600 298298 623700
rect 298398 623600 298522 623700
rect 298622 623600 298746 623700
rect 298846 623600 298880 623700
rect 294704 623476 298880 623600
rect 294704 623376 297850 623476
rect 297950 623376 298074 623476
rect 298174 623376 298298 623476
rect 298398 623376 298522 623476
rect 298622 623376 298746 623476
rect 298846 623376 298880 623476
rect 294704 623252 298880 623376
rect 294704 623152 297850 623252
rect 297950 623152 298074 623252
rect 298174 623152 298298 623252
rect 298398 623152 298522 623252
rect 298622 623152 298746 623252
rect 298846 623152 298880 623252
rect 294704 623028 298880 623152
rect 294704 622928 297850 623028
rect 297950 622928 298074 623028
rect 298174 622928 298298 623028
rect 298398 622928 298522 623028
rect 298622 622928 298746 623028
rect 298846 622928 298880 623028
rect 294704 622804 298880 622928
rect 294704 622704 297850 622804
rect 297950 622704 298074 622804
rect 298174 622704 298298 622804
rect 298398 622704 298522 622804
rect 298622 622704 298746 622804
rect 298846 622704 298880 622804
rect 294704 622580 298880 622704
rect 294704 622480 297850 622580
rect 297950 622480 298074 622580
rect 298174 622480 298298 622580
rect 298398 622480 298522 622580
rect 298622 622480 298746 622580
rect 298846 622480 298880 622580
rect 294704 622356 298880 622480
rect 294704 622256 297850 622356
rect 297950 622256 298074 622356
rect 298174 622256 298298 622356
rect 298398 622256 298522 622356
rect 298622 622256 298746 622356
rect 298846 622256 298880 622356
rect 294704 622132 298880 622256
rect 294704 622032 297850 622132
rect 297950 622032 298074 622132
rect 298174 622032 298298 622132
rect 298398 622032 298522 622132
rect 298622 622032 298746 622132
rect 298846 622032 298880 622132
rect 294704 621908 298880 622032
rect 294704 621808 297850 621908
rect 297950 621808 298074 621908
rect 298174 621808 298298 621908
rect 298398 621808 298522 621908
rect 298622 621808 298746 621908
rect 298846 621808 298880 621908
rect 294704 621684 298880 621808
rect 294704 621584 297850 621684
rect 297950 621584 298074 621684
rect 298174 621584 298298 621684
rect 298398 621584 298522 621684
rect 298622 621584 298746 621684
rect 298846 621584 298880 621684
rect 294704 621460 298880 621584
rect 294704 621360 297850 621460
rect 297950 621360 298074 621460
rect 298174 621360 298298 621460
rect 298398 621360 298522 621460
rect 298622 621360 298746 621460
rect 298846 621360 298880 621460
rect 294704 621236 298880 621360
rect 294704 621136 297850 621236
rect 297950 621136 298074 621236
rect 298174 621136 298298 621236
rect 298398 621136 298522 621236
rect 298622 621136 298746 621236
rect 298846 621136 298880 621236
rect 294704 621012 298880 621136
rect 294704 620912 297850 621012
rect 297950 620912 298074 621012
rect 298174 620912 298298 621012
rect 298398 620912 298522 621012
rect 298622 620912 298746 621012
rect 298846 620912 298880 621012
rect 294704 620788 298880 620912
rect 294704 620688 297850 620788
rect 297950 620688 298074 620788
rect 298174 620688 298298 620788
rect 298398 620688 298522 620788
rect 298622 620688 298746 620788
rect 298846 620688 298880 620788
rect 294704 620564 298880 620688
rect 294704 620464 297850 620564
rect 297950 620464 298074 620564
rect 298174 620464 298298 620564
rect 298398 620464 298522 620564
rect 298622 620464 298746 620564
rect 298846 620464 298880 620564
rect 294704 620340 298880 620464
rect 294704 620240 297850 620340
rect 297950 620240 298074 620340
rect 298174 620240 298298 620340
rect 298398 620240 298522 620340
rect 298622 620240 298746 620340
rect 298846 620240 298880 620340
rect 294704 620116 298880 620240
rect 294704 620016 297850 620116
rect 297950 620016 298074 620116
rect 298174 620016 298298 620116
rect 298398 620016 298522 620116
rect 298622 620016 298746 620116
rect 298846 620016 298880 620116
rect 294704 619892 298880 620016
rect 294704 619792 297850 619892
rect 297950 619792 298074 619892
rect 298174 619792 298298 619892
rect 298398 619792 298522 619892
rect 298622 619792 298746 619892
rect 298846 619792 298880 619892
rect 294704 619668 298880 619792
rect 294704 619568 297850 619668
rect 297950 619568 298074 619668
rect 298174 619568 298298 619668
rect 298398 619568 298522 619668
rect 298622 619568 298746 619668
rect 298846 619568 298880 619668
rect 294704 619444 298880 619568
rect 294704 619344 297850 619444
rect 297950 619344 298074 619444
rect 298174 619344 298298 619444
rect 298398 619344 298522 619444
rect 298622 619344 298746 619444
rect 298846 619344 298880 619444
rect 294704 619220 298880 619344
rect 294704 619120 297850 619220
rect 297950 619120 298074 619220
rect 298174 619120 298298 619220
rect 298398 619120 298522 619220
rect 298622 619120 298746 619220
rect 298846 619120 298880 619220
rect 294704 618996 298880 619120
rect 294704 618896 297850 618996
rect 297950 618896 298074 618996
rect 298174 618896 298298 618996
rect 298398 618896 298522 618996
rect 298622 618896 298746 618996
rect 298846 618896 298880 618996
rect 294704 618772 298880 618896
rect 294704 618672 297850 618772
rect 297950 618672 298074 618772
rect 298174 618672 298298 618772
rect 298398 618672 298522 618772
rect 298622 618672 298746 618772
rect 298846 618672 298880 618772
rect 294704 618548 298880 618672
rect 294704 618448 297850 618548
rect 297950 618448 298074 618548
rect 298174 618448 298298 618548
rect 298398 618448 298522 618548
rect 298622 618448 298746 618548
rect 298846 618448 298880 618548
rect 294704 618324 298880 618448
rect 294704 618224 297850 618324
rect 297950 618224 298074 618324
rect 298174 618224 298298 618324
rect 298398 618224 298522 618324
rect 298622 618224 298746 618324
rect 298846 618224 298880 618324
rect 294704 618100 298880 618224
rect 294704 618040 297850 618100
rect 289020 618000 297850 618040
rect 297950 618000 298074 618100
rect 298174 618000 298298 618100
rect 298398 618000 298522 618100
rect 298622 618000 298746 618100
rect 298846 618000 298880 618100
rect 289020 617940 298880 618000
rect 342000 624596 525804 624606
rect 342000 624496 342130 624596
rect 342230 624496 342354 624596
rect 342454 624496 342578 624596
rect 342678 624496 342802 624596
rect 342902 624496 343026 624596
rect 343126 624496 525804 624596
rect 342000 624372 525804 624496
rect 342000 624272 342130 624372
rect 342230 624272 342354 624372
rect 342454 624272 342578 624372
rect 342678 624272 342802 624372
rect 342902 624272 343026 624372
rect 343126 624272 525804 624372
rect 342000 624161 525804 624272
rect 342000 624148 510602 624161
rect 342000 624048 342130 624148
rect 342230 624048 342354 624148
rect 342454 624048 342578 624148
rect 342678 624048 342802 624148
rect 342902 624048 343026 624148
rect 343126 624048 510602 624148
rect 342000 623924 510602 624048
rect 342000 623824 342130 623924
rect 342230 623824 342354 623924
rect 342454 623824 342578 623924
rect 342678 623824 342802 623924
rect 342902 623824 343026 623924
rect 343126 623824 510602 623924
rect 342000 623700 510602 623824
rect 342000 623600 342130 623700
rect 342230 623600 342354 623700
rect 342454 623600 342578 623700
rect 342678 623600 342802 623700
rect 342902 623600 343026 623700
rect 343126 623600 510602 623700
rect 342000 623476 510602 623600
rect 342000 623376 342130 623476
rect 342230 623376 342354 623476
rect 342454 623376 342578 623476
rect 342678 623376 342802 623476
rect 342902 623376 343026 623476
rect 343126 623376 510602 623476
rect 342000 623252 510602 623376
rect 342000 623152 342130 623252
rect 342230 623152 342354 623252
rect 342454 623152 342578 623252
rect 342678 623152 342802 623252
rect 342902 623152 343026 623252
rect 343126 623152 510602 623252
rect 342000 623028 510602 623152
rect 342000 622928 342130 623028
rect 342230 622928 342354 623028
rect 342454 622928 342578 623028
rect 342678 622928 342802 623028
rect 342902 622928 343026 623028
rect 343126 622928 510602 623028
rect 342000 622804 510602 622928
rect 342000 622704 342130 622804
rect 342230 622704 342354 622804
rect 342454 622704 342578 622804
rect 342678 622704 342802 622804
rect 342902 622704 343026 622804
rect 343126 622704 510602 622804
rect 342000 622580 510602 622704
rect 342000 622480 342130 622580
rect 342230 622480 342354 622580
rect 342454 622480 342578 622580
rect 342678 622480 342802 622580
rect 342902 622480 343026 622580
rect 343126 622480 510602 622580
rect 342000 622356 510602 622480
rect 342000 622256 342130 622356
rect 342230 622256 342354 622356
rect 342454 622256 342578 622356
rect 342678 622256 342802 622356
rect 342902 622256 343026 622356
rect 343126 622256 510602 622356
rect 342000 622132 510602 622256
rect 342000 622032 342130 622132
rect 342230 622032 342354 622132
rect 342454 622032 342578 622132
rect 342678 622032 342802 622132
rect 342902 622032 343026 622132
rect 343126 622032 510602 622132
rect 342000 621908 510602 622032
rect 342000 621808 342130 621908
rect 342230 621808 342354 621908
rect 342454 621808 342578 621908
rect 342678 621808 342802 621908
rect 342902 621808 343026 621908
rect 343126 621808 510602 621908
rect 342000 621684 510602 621808
rect 342000 621584 342130 621684
rect 342230 621584 342354 621684
rect 342454 621584 342578 621684
rect 342678 621584 342802 621684
rect 342902 621584 343026 621684
rect 343126 621584 510602 621684
rect 342000 621460 510602 621584
rect 342000 621360 342130 621460
rect 342230 621360 342354 621460
rect 342454 621360 342578 621460
rect 342678 621360 342802 621460
rect 342902 621360 343026 621460
rect 343126 621360 510602 621460
rect 342000 621236 510602 621360
rect 342000 621136 342130 621236
rect 342230 621136 342354 621236
rect 342454 621136 342578 621236
rect 342678 621136 342802 621236
rect 342902 621136 343026 621236
rect 343126 621136 510602 621236
rect 342000 621012 510602 621136
rect 342000 620912 342130 621012
rect 342230 620912 342354 621012
rect 342454 620912 342578 621012
rect 342678 620912 342802 621012
rect 342902 620912 343026 621012
rect 343126 620912 510602 621012
rect 342000 620788 510602 620912
rect 342000 620688 342130 620788
rect 342230 620688 342354 620788
rect 342454 620688 342578 620788
rect 342678 620688 342802 620788
rect 342902 620688 343026 620788
rect 343126 620688 510602 620788
rect 342000 620564 510602 620688
rect 342000 620464 342130 620564
rect 342230 620464 342354 620564
rect 342454 620464 342578 620564
rect 342678 620464 342802 620564
rect 342902 620464 343026 620564
rect 343126 620464 510602 620564
rect 342000 620340 510602 620464
rect 342000 620240 342130 620340
rect 342230 620240 342354 620340
rect 342454 620240 342578 620340
rect 342678 620240 342802 620340
rect 342902 620240 343026 620340
rect 343126 620240 510602 620340
rect 342000 620116 510602 620240
rect 342000 620016 342130 620116
rect 342230 620016 342354 620116
rect 342454 620016 342578 620116
rect 342678 620016 342802 620116
rect 342902 620016 343026 620116
rect 343126 620016 510602 620116
rect 342000 619892 510602 620016
rect 342000 619792 342130 619892
rect 342230 619792 342354 619892
rect 342454 619792 342578 619892
rect 342678 619792 342802 619892
rect 342902 619792 343026 619892
rect 343126 619792 510602 619892
rect 342000 619668 510602 619792
rect 342000 619568 342130 619668
rect 342230 619568 342354 619668
rect 342454 619568 342578 619668
rect 342678 619568 342802 619668
rect 342902 619568 343026 619668
rect 343126 619568 510602 619668
rect 342000 619444 510602 619568
rect 342000 619344 342130 619444
rect 342230 619344 342354 619444
rect 342454 619344 342578 619444
rect 342678 619344 342802 619444
rect 342902 619344 343026 619444
rect 343126 619344 510602 619444
rect 342000 619220 510602 619344
rect 342000 619120 342130 619220
rect 342230 619120 342354 619220
rect 342454 619120 342578 619220
rect 342678 619120 342802 619220
rect 342902 619120 343026 619220
rect 343126 619120 510602 619220
rect 342000 618996 510602 619120
rect 342000 618896 342130 618996
rect 342230 618896 342354 618996
rect 342454 618896 342578 618996
rect 342678 618896 342802 618996
rect 342902 618896 343026 618996
rect 343126 618896 510602 618996
rect 342000 618772 510602 618896
rect 342000 618672 342130 618772
rect 342230 618672 342354 618772
rect 342454 618672 342578 618772
rect 342678 618672 342802 618772
rect 342902 618672 343026 618772
rect 343126 618672 510602 618772
rect 342000 618548 510602 618672
rect 342000 618448 342130 618548
rect 342230 618448 342354 618548
rect 342454 618448 342578 618548
rect 342678 618448 342802 618548
rect 342902 618448 343026 618548
rect 343126 618448 510602 618548
rect 342000 618417 510602 618448
rect 515386 618417 520602 624161
rect 525386 618417 525804 624161
rect 342000 618324 525804 618417
rect 342000 618224 342130 618324
rect 342230 618224 342354 618324
rect 342454 618224 342578 618324
rect 342678 618224 342802 618324
rect 342902 618224 343026 618324
rect 343126 618224 525804 618324
rect 342000 618100 525804 618224
rect 342000 618000 342130 618100
rect 342230 618000 342354 618100
rect 342454 618000 342578 618100
rect 342678 618000 342802 618100
rect 342902 618000 343026 618100
rect 343126 618000 525804 618100
rect 342000 617944 525804 618000
rect 335560 615499 342216 615504
rect 335560 615494 342217 615499
rect 298820 615479 305476 615484
rect 309290 615479 315946 615484
rect 298820 615474 305477 615479
rect 298820 615374 298876 615474
rect 298976 615374 299100 615474
rect 299200 615374 299324 615474
rect 299424 615374 299548 615474
rect 299648 615374 299772 615474
rect 299872 615374 299996 615474
rect 300096 615374 300220 615474
rect 300320 615374 300444 615474
rect 300544 615374 300668 615474
rect 300768 615374 300892 615474
rect 300992 615374 301116 615474
rect 301216 615374 301340 615474
rect 301440 615374 301564 615474
rect 301664 615374 301788 615474
rect 301888 615374 302012 615474
rect 302112 615374 302236 615474
rect 302336 615374 302460 615474
rect 302560 615374 302684 615474
rect 302784 615374 302908 615474
rect 303008 615374 303132 615474
rect 303232 615374 303356 615474
rect 303456 615374 303580 615474
rect 303680 615374 303804 615474
rect 303904 615374 304028 615474
rect 304128 615374 304252 615474
rect 304352 615374 304476 615474
rect 304576 615374 304700 615474
rect 304800 615374 304924 615474
rect 305024 615374 305148 615474
rect 305248 615374 305372 615474
rect 305472 615374 305477 615474
rect 298820 615369 305477 615374
rect 309290 615474 315947 615479
rect 309290 615374 309346 615474
rect 309446 615374 309570 615474
rect 309670 615374 309794 615474
rect 309894 615374 310018 615474
rect 310118 615374 310242 615474
rect 310342 615374 310466 615474
rect 310566 615374 310690 615474
rect 310790 615374 310914 615474
rect 311014 615374 311138 615474
rect 311238 615374 311362 615474
rect 311462 615374 311586 615474
rect 311686 615374 311810 615474
rect 311910 615374 312034 615474
rect 312134 615374 312258 615474
rect 312358 615374 312482 615474
rect 312582 615374 312706 615474
rect 312806 615374 312930 615474
rect 313030 615374 313154 615474
rect 313254 615374 313378 615474
rect 313478 615374 313602 615474
rect 313702 615374 313826 615474
rect 313926 615374 314050 615474
rect 314150 615374 314274 615474
rect 314374 615374 314498 615474
rect 314598 615374 314722 615474
rect 314822 615374 314946 615474
rect 315046 615374 315170 615474
rect 315270 615374 315394 615474
rect 315494 615374 315618 615474
rect 315718 615374 315842 615474
rect 315942 615374 315947 615474
rect 309290 615369 315947 615374
rect 335560 615394 335616 615494
rect 335716 615394 335840 615494
rect 335940 615394 336064 615494
rect 336164 615394 336288 615494
rect 336388 615394 336512 615494
rect 336612 615394 336736 615494
rect 336836 615394 336960 615494
rect 337060 615394 337184 615494
rect 337284 615394 337408 615494
rect 337508 615394 337632 615494
rect 337732 615394 337856 615494
rect 337956 615394 338080 615494
rect 338180 615394 338304 615494
rect 338404 615394 338528 615494
rect 338628 615394 338752 615494
rect 338852 615394 338976 615494
rect 339076 615394 339200 615494
rect 339300 615394 339424 615494
rect 339524 615394 339648 615494
rect 339748 615394 339872 615494
rect 339972 615394 340096 615494
rect 340196 615394 340320 615494
rect 340420 615394 340544 615494
rect 340644 615394 340768 615494
rect 340868 615394 340992 615494
rect 341092 615394 341216 615494
rect 341316 615394 341440 615494
rect 341540 615394 341664 615494
rect 341764 615394 341888 615494
rect 341988 615394 342112 615494
rect 342212 615394 342217 615494
rect 335560 615389 342217 615394
rect 298820 615255 305476 615369
rect 309290 615255 315946 615369
rect 335560 615275 342216 615389
rect 335560 615270 342217 615275
rect 298820 615250 305477 615255
rect 298820 615150 298876 615250
rect 298976 615150 299100 615250
rect 299200 615150 299324 615250
rect 299424 615150 299548 615250
rect 299648 615150 299772 615250
rect 299872 615150 299996 615250
rect 300096 615150 300220 615250
rect 300320 615150 300444 615250
rect 300544 615150 300668 615250
rect 300768 615150 300892 615250
rect 300992 615150 301116 615250
rect 301216 615150 301340 615250
rect 301440 615150 301564 615250
rect 301664 615150 301788 615250
rect 301888 615150 302012 615250
rect 302112 615150 302236 615250
rect 302336 615150 302460 615250
rect 302560 615150 302684 615250
rect 302784 615150 302908 615250
rect 303008 615150 303132 615250
rect 303232 615150 303356 615250
rect 303456 615150 303580 615250
rect 303680 615150 303804 615250
rect 303904 615150 304028 615250
rect 304128 615150 304252 615250
rect 304352 615150 304476 615250
rect 304576 615150 304700 615250
rect 304800 615150 304924 615250
rect 305024 615150 305148 615250
rect 305248 615150 305372 615250
rect 305472 615150 305477 615250
rect 298820 615145 305477 615150
rect 309290 615250 315947 615255
rect 309290 615150 309346 615250
rect 309446 615150 309570 615250
rect 309670 615150 309794 615250
rect 309894 615150 310018 615250
rect 310118 615150 310242 615250
rect 310342 615150 310466 615250
rect 310566 615150 310690 615250
rect 310790 615150 310914 615250
rect 311014 615150 311138 615250
rect 311238 615150 311362 615250
rect 311462 615150 311586 615250
rect 311686 615150 311810 615250
rect 311910 615150 312034 615250
rect 312134 615150 312258 615250
rect 312358 615150 312482 615250
rect 312582 615150 312706 615250
rect 312806 615150 312930 615250
rect 313030 615150 313154 615250
rect 313254 615150 313378 615250
rect 313478 615150 313602 615250
rect 313702 615150 313826 615250
rect 313926 615150 314050 615250
rect 314150 615150 314274 615250
rect 314374 615150 314498 615250
rect 314598 615150 314722 615250
rect 314822 615150 314946 615250
rect 315046 615150 315170 615250
rect 315270 615150 315394 615250
rect 315494 615150 315618 615250
rect 315718 615150 315842 615250
rect 315942 615150 315947 615250
rect 309290 615145 315947 615150
rect 335560 615170 335616 615270
rect 335716 615170 335840 615270
rect 335940 615170 336064 615270
rect 336164 615170 336288 615270
rect 336388 615170 336512 615270
rect 336612 615170 336736 615270
rect 336836 615170 336960 615270
rect 337060 615170 337184 615270
rect 337284 615170 337408 615270
rect 337508 615170 337632 615270
rect 337732 615170 337856 615270
rect 337956 615170 338080 615270
rect 338180 615170 338304 615270
rect 338404 615170 338528 615270
rect 338628 615170 338752 615270
rect 338852 615170 338976 615270
rect 339076 615170 339200 615270
rect 339300 615170 339424 615270
rect 339524 615170 339648 615270
rect 339748 615170 339872 615270
rect 339972 615170 340096 615270
rect 340196 615170 340320 615270
rect 340420 615170 340544 615270
rect 340644 615170 340768 615270
rect 340868 615170 340992 615270
rect 341092 615170 341216 615270
rect 341316 615170 341440 615270
rect 341540 615170 341664 615270
rect 341764 615170 341888 615270
rect 341988 615170 342112 615270
rect 342212 615170 342217 615270
rect 335560 615165 342217 615170
rect 298820 615031 305476 615145
rect 309290 615031 315946 615145
rect 335560 615051 342216 615165
rect 335560 615046 342217 615051
rect 298820 615026 305477 615031
rect 298820 614926 298876 615026
rect 298976 614926 299100 615026
rect 299200 614926 299324 615026
rect 299424 614926 299548 615026
rect 299648 614926 299772 615026
rect 299872 614926 299996 615026
rect 300096 614926 300220 615026
rect 300320 614926 300444 615026
rect 300544 614926 300668 615026
rect 300768 614926 300892 615026
rect 300992 614926 301116 615026
rect 301216 614926 301340 615026
rect 301440 614926 301564 615026
rect 301664 614926 301788 615026
rect 301888 614926 302012 615026
rect 302112 614926 302236 615026
rect 302336 614926 302460 615026
rect 302560 614926 302684 615026
rect 302784 614926 302908 615026
rect 303008 614926 303132 615026
rect 303232 614926 303356 615026
rect 303456 614926 303580 615026
rect 303680 614926 303804 615026
rect 303904 614926 304028 615026
rect 304128 614926 304252 615026
rect 304352 614926 304476 615026
rect 304576 614926 304700 615026
rect 304800 614926 304924 615026
rect 305024 614926 305148 615026
rect 305248 614926 305372 615026
rect 305472 614926 305477 615026
rect 298820 614921 305477 614926
rect 309290 615026 315947 615031
rect 309290 614926 309346 615026
rect 309446 614926 309570 615026
rect 309670 614926 309794 615026
rect 309894 614926 310018 615026
rect 310118 614926 310242 615026
rect 310342 614926 310466 615026
rect 310566 614926 310690 615026
rect 310790 614926 310914 615026
rect 311014 614926 311138 615026
rect 311238 614926 311362 615026
rect 311462 614926 311586 615026
rect 311686 614926 311810 615026
rect 311910 614926 312034 615026
rect 312134 614926 312258 615026
rect 312358 614926 312482 615026
rect 312582 614926 312706 615026
rect 312806 614926 312930 615026
rect 313030 614926 313154 615026
rect 313254 614926 313378 615026
rect 313478 614926 313602 615026
rect 313702 614926 313826 615026
rect 313926 614926 314050 615026
rect 314150 614926 314274 615026
rect 314374 614926 314498 615026
rect 314598 614926 314722 615026
rect 314822 614926 314946 615026
rect 315046 614926 315170 615026
rect 315270 614926 315394 615026
rect 315494 614926 315618 615026
rect 315718 614926 315842 615026
rect 315942 614926 315947 615026
rect 309290 614921 315947 614926
rect 335560 614946 335616 615046
rect 335716 614946 335840 615046
rect 335940 614946 336064 615046
rect 336164 614946 336288 615046
rect 336388 614946 336512 615046
rect 336612 614946 336736 615046
rect 336836 614946 336960 615046
rect 337060 614946 337184 615046
rect 337284 614946 337408 615046
rect 337508 614946 337632 615046
rect 337732 614946 337856 615046
rect 337956 614946 338080 615046
rect 338180 614946 338304 615046
rect 338404 614946 338528 615046
rect 338628 614946 338752 615046
rect 338852 614946 338976 615046
rect 339076 614946 339200 615046
rect 339300 614946 339424 615046
rect 339524 614946 339648 615046
rect 339748 614946 339872 615046
rect 339972 614946 340096 615046
rect 340196 614946 340320 615046
rect 340420 614946 340544 615046
rect 340644 614946 340768 615046
rect 340868 614946 340992 615046
rect 341092 614946 341216 615046
rect 341316 614946 341440 615046
rect 341540 614946 341664 615046
rect 341764 614946 341888 615046
rect 341988 614946 342112 615046
rect 342212 614946 342217 615046
rect 335560 614941 342217 614946
rect 298820 614807 305476 614921
rect 309290 614807 315946 614921
rect 335560 614827 342216 614941
rect 335560 614822 342217 614827
rect 298820 614802 305477 614807
rect 298820 614702 298876 614802
rect 298976 614702 299100 614802
rect 299200 614702 299324 614802
rect 299424 614702 299548 614802
rect 299648 614702 299772 614802
rect 299872 614702 299996 614802
rect 300096 614702 300220 614802
rect 300320 614702 300444 614802
rect 300544 614702 300668 614802
rect 300768 614702 300892 614802
rect 300992 614702 301116 614802
rect 301216 614702 301340 614802
rect 301440 614702 301564 614802
rect 301664 614702 301788 614802
rect 301888 614702 302012 614802
rect 302112 614702 302236 614802
rect 302336 614702 302460 614802
rect 302560 614702 302684 614802
rect 302784 614702 302908 614802
rect 303008 614702 303132 614802
rect 303232 614702 303356 614802
rect 303456 614702 303580 614802
rect 303680 614702 303804 614802
rect 303904 614702 304028 614802
rect 304128 614702 304252 614802
rect 304352 614702 304476 614802
rect 304576 614702 304700 614802
rect 304800 614702 304924 614802
rect 305024 614702 305148 614802
rect 305248 614702 305372 614802
rect 305472 614702 305477 614802
rect 298820 614697 305477 614702
rect 309290 614802 315947 614807
rect 309290 614702 309346 614802
rect 309446 614702 309570 614802
rect 309670 614702 309794 614802
rect 309894 614702 310018 614802
rect 310118 614702 310242 614802
rect 310342 614702 310466 614802
rect 310566 614702 310690 614802
rect 310790 614702 310914 614802
rect 311014 614702 311138 614802
rect 311238 614702 311362 614802
rect 311462 614702 311586 614802
rect 311686 614702 311810 614802
rect 311910 614702 312034 614802
rect 312134 614702 312258 614802
rect 312358 614702 312482 614802
rect 312582 614702 312706 614802
rect 312806 614702 312930 614802
rect 313030 614702 313154 614802
rect 313254 614702 313378 614802
rect 313478 614702 313602 614802
rect 313702 614702 313826 614802
rect 313926 614702 314050 614802
rect 314150 614702 314274 614802
rect 314374 614702 314498 614802
rect 314598 614702 314722 614802
rect 314822 614702 314946 614802
rect 315046 614702 315170 614802
rect 315270 614702 315394 614802
rect 315494 614702 315618 614802
rect 315718 614702 315842 614802
rect 315942 614702 315947 614802
rect 309290 614697 315947 614702
rect 335560 614722 335616 614822
rect 335716 614722 335840 614822
rect 335940 614722 336064 614822
rect 336164 614722 336288 614822
rect 336388 614722 336512 614822
rect 336612 614722 336736 614822
rect 336836 614722 336960 614822
rect 337060 614722 337184 614822
rect 337284 614722 337408 614822
rect 337508 614722 337632 614822
rect 337732 614722 337856 614822
rect 337956 614722 338080 614822
rect 338180 614722 338304 614822
rect 338404 614722 338528 614822
rect 338628 614722 338752 614822
rect 338852 614722 338976 614822
rect 339076 614722 339200 614822
rect 339300 614722 339424 614822
rect 339524 614722 339648 614822
rect 339748 614722 339872 614822
rect 339972 614722 340096 614822
rect 340196 614722 340320 614822
rect 340420 614722 340544 614822
rect 340644 614722 340768 614822
rect 340868 614722 340992 614822
rect 341092 614722 341216 614822
rect 341316 614722 341440 614822
rect 341540 614722 341664 614822
rect 341764 614722 341888 614822
rect 341988 614722 342112 614822
rect 342212 614722 342217 614822
rect 335560 614717 342217 614722
rect 298820 614583 305476 614697
rect 309290 614583 315946 614697
rect 335560 614603 342216 614717
rect 335560 614598 342217 614603
rect 298820 614578 305477 614583
rect 298820 614478 298876 614578
rect 298976 614478 299100 614578
rect 299200 614478 299324 614578
rect 299424 614478 299548 614578
rect 299648 614478 299772 614578
rect 299872 614478 299996 614578
rect 300096 614478 300220 614578
rect 300320 614478 300444 614578
rect 300544 614478 300668 614578
rect 300768 614478 300892 614578
rect 300992 614478 301116 614578
rect 301216 614478 301340 614578
rect 301440 614478 301564 614578
rect 301664 614478 301788 614578
rect 301888 614478 302012 614578
rect 302112 614478 302236 614578
rect 302336 614478 302460 614578
rect 302560 614478 302684 614578
rect 302784 614478 302908 614578
rect 303008 614478 303132 614578
rect 303232 614478 303356 614578
rect 303456 614478 303580 614578
rect 303680 614478 303804 614578
rect 303904 614478 304028 614578
rect 304128 614478 304252 614578
rect 304352 614478 304476 614578
rect 304576 614478 304700 614578
rect 304800 614478 304924 614578
rect 305024 614478 305148 614578
rect 305248 614478 305372 614578
rect 305472 614478 305477 614578
rect 298820 614473 305477 614478
rect 309290 614578 315947 614583
rect 309290 614478 309346 614578
rect 309446 614478 309570 614578
rect 309670 614478 309794 614578
rect 309894 614478 310018 614578
rect 310118 614478 310242 614578
rect 310342 614478 310466 614578
rect 310566 614478 310690 614578
rect 310790 614478 310914 614578
rect 311014 614478 311138 614578
rect 311238 614478 311362 614578
rect 311462 614478 311586 614578
rect 311686 614478 311810 614578
rect 311910 614478 312034 614578
rect 312134 614478 312258 614578
rect 312358 614478 312482 614578
rect 312582 614478 312706 614578
rect 312806 614478 312930 614578
rect 313030 614478 313154 614578
rect 313254 614478 313378 614578
rect 313478 614478 313602 614578
rect 313702 614478 313826 614578
rect 313926 614478 314050 614578
rect 314150 614478 314274 614578
rect 314374 614478 314498 614578
rect 314598 614478 314722 614578
rect 314822 614478 314946 614578
rect 315046 614478 315170 614578
rect 315270 614478 315394 614578
rect 315494 614478 315618 614578
rect 315718 614478 315842 614578
rect 315942 614478 315947 614578
rect 309290 614473 315947 614478
rect 335560 614498 335616 614598
rect 335716 614498 335840 614598
rect 335940 614498 336064 614598
rect 336164 614498 336288 614598
rect 336388 614498 336512 614598
rect 336612 614498 336736 614598
rect 336836 614498 336960 614598
rect 337060 614498 337184 614598
rect 337284 614498 337408 614598
rect 337508 614498 337632 614598
rect 337732 614498 337856 614598
rect 337956 614498 338080 614598
rect 338180 614498 338304 614598
rect 338404 614498 338528 614598
rect 338628 614498 338752 614598
rect 338852 614498 338976 614598
rect 339076 614498 339200 614598
rect 339300 614498 339424 614598
rect 339524 614498 339648 614598
rect 339748 614498 339872 614598
rect 339972 614498 340096 614598
rect 340196 614498 340320 614598
rect 340420 614498 340544 614598
rect 340644 614498 340768 614598
rect 340868 614498 340992 614598
rect 341092 614498 341216 614598
rect 341316 614498 341440 614598
rect 341540 614498 341664 614598
rect 341764 614498 341888 614598
rect 341988 614498 342112 614598
rect 342212 614498 342217 614598
rect 335560 614493 342217 614498
rect 298820 614444 305476 614473
rect 309290 614444 315946 614473
rect 335560 614464 342216 614493
rect 316300 611176 525804 611206
rect 285800 611084 525804 611176
rect 285800 611080 336480 611084
rect 285800 610764 298920 611080
rect 285800 605020 289920 610764
rect 294704 605336 298920 610764
rect 303704 605336 304920 611080
rect 309704 605336 310920 611080
rect 315704 605340 336480 611080
rect 341264 610761 525804 611084
rect 341264 605340 510602 610761
rect 315704 605336 510602 605340
rect 294704 605020 510602 605336
rect 285800 605017 510602 605020
rect 515386 605017 520602 610761
rect 525386 605017 525804 610761
rect 285800 604544 525804 605017
rect 285800 604520 316300 604544
rect 560425 597806 566979 629792
rect 316064 597324 566979 597806
rect 316064 591580 317480 597324
rect 322264 591580 325480 597324
rect 330264 591580 566979 597324
rect 316064 591240 566979 591580
rect 316060 591140 566980 591240
rect 556059 555354 562613 559520
rect 556059 550570 556255 555354
rect 562319 550570 562613 555354
rect 556059 545354 562613 550570
rect 556059 540570 556255 545354
rect 562319 540570 562613 545354
rect 556059 540155 562613 540570
rect 573464 500138 576816 500473
rect 573464 500074 573553 500138
rect 573617 500074 573633 500138
rect 573697 500074 573713 500138
rect 573777 500074 573793 500138
rect 573857 500074 573873 500138
rect 573937 500074 573953 500138
rect 574017 500074 574033 500138
rect 574097 500074 574113 500138
rect 574177 500074 574193 500138
rect 574257 500074 574273 500138
rect 574337 500074 574353 500138
rect 574417 500074 574433 500138
rect 574497 500074 574513 500138
rect 574577 500074 574593 500138
rect 574657 500074 574673 500138
rect 574737 500074 574753 500138
rect 574817 500074 574833 500138
rect 574897 500074 574913 500138
rect 574977 500074 574993 500138
rect 575057 500074 575073 500138
rect 575137 500074 575153 500138
rect 575217 500074 575233 500138
rect 575297 500074 575313 500138
rect 575377 500074 575393 500138
rect 575457 500074 575473 500138
rect 575537 500074 575553 500138
rect 575617 500074 575633 500138
rect 575697 500074 575713 500138
rect 575777 500074 575793 500138
rect 575857 500074 575873 500138
rect 575937 500074 575953 500138
rect 576017 500074 576033 500138
rect 576097 500074 576113 500138
rect 576177 500074 576193 500138
rect 576257 500074 576273 500138
rect 576337 500074 576353 500138
rect 576417 500074 576433 500138
rect 576497 500074 576513 500138
rect 576577 500074 576593 500138
rect 576657 500074 576673 500138
rect 576737 500074 576816 500138
rect 13814 462486 17684 462771
rect 13814 462422 13897 462486
rect 13961 462422 13977 462486
rect 14041 462422 14057 462486
rect 14121 462422 14137 462486
rect 14201 462422 14217 462486
rect 14281 462422 14297 462486
rect 14361 462422 14377 462486
rect 14441 462422 14457 462486
rect 14521 462422 14537 462486
rect 14601 462422 14617 462486
rect 14681 462422 14697 462486
rect 14761 462422 14777 462486
rect 14841 462422 14857 462486
rect 14921 462422 14937 462486
rect 15001 462422 15017 462486
rect 15081 462422 15097 462486
rect 15161 462422 15177 462486
rect 15241 462422 15257 462486
rect 15321 462422 15337 462486
rect 15401 462422 15417 462486
rect 15481 462422 15497 462486
rect 15561 462422 15577 462486
rect 15641 462422 15657 462486
rect 15721 462422 15737 462486
rect 15801 462422 15817 462486
rect 15881 462422 15897 462486
rect 15961 462422 15977 462486
rect 16041 462422 16057 462486
rect 16121 462422 16137 462486
rect 16201 462422 16217 462486
rect 16281 462422 16297 462486
rect 16361 462422 16377 462486
rect 16441 462422 16457 462486
rect 16521 462422 16537 462486
rect 16601 462422 16617 462486
rect 16681 462422 16697 462486
rect 16761 462422 16777 462486
rect 16841 462422 16857 462486
rect 16921 462422 16937 462486
rect 17001 462422 17017 462486
rect 17081 462422 17097 462486
rect 17161 462422 17177 462486
rect 17241 462422 17257 462486
rect 17321 462422 17337 462486
rect 17401 462422 17417 462486
rect 17481 462422 17497 462486
rect 17561 462422 17684 462486
rect 13814 419264 17684 462422
rect 13814 419200 13911 419264
rect 13975 419200 13991 419264
rect 14055 419200 14071 419264
rect 14135 419200 14151 419264
rect 14215 419200 14231 419264
rect 14295 419200 14311 419264
rect 14375 419200 14391 419264
rect 14455 419200 14471 419264
rect 14535 419200 14551 419264
rect 14615 419200 14631 419264
rect 14695 419200 14711 419264
rect 14775 419200 14791 419264
rect 14855 419200 14871 419264
rect 14935 419200 14951 419264
rect 15015 419200 15031 419264
rect 15095 419200 15111 419264
rect 15175 419200 15191 419264
rect 15255 419200 15271 419264
rect 15335 419200 15351 419264
rect 15415 419200 15431 419264
rect 15495 419200 15511 419264
rect 15575 419200 15591 419264
rect 15655 419200 15671 419264
rect 15735 419200 15751 419264
rect 15815 419200 15831 419264
rect 15895 419200 15911 419264
rect 15975 419200 15991 419264
rect 16055 419200 16071 419264
rect 16135 419200 16151 419264
rect 16215 419200 16231 419264
rect 16295 419200 16311 419264
rect 16375 419200 16391 419264
rect 16455 419200 16471 419264
rect 16535 419200 16551 419264
rect 16615 419200 16631 419264
rect 16695 419200 16711 419264
rect 16775 419200 16791 419264
rect 16855 419200 16871 419264
rect 16935 419200 16951 419264
rect 17015 419200 17031 419264
rect 17095 419200 17111 419264
rect 17175 419200 17191 419264
rect 17255 419200 17271 419264
rect 17335 419200 17351 419264
rect 17415 419200 17431 419264
rect 17495 419200 17511 419264
rect 17575 419200 17684 419264
rect 13814 227257 17684 419200
rect 573464 455716 576816 500074
rect 573464 455652 573591 455716
rect 573655 455652 573671 455716
rect 573735 455652 573751 455716
rect 573815 455652 573831 455716
rect 573895 455652 573911 455716
rect 573975 455652 573991 455716
rect 574055 455652 574071 455716
rect 574135 455652 574151 455716
rect 574215 455652 574231 455716
rect 574295 455652 574311 455716
rect 574375 455652 574391 455716
rect 574455 455652 574471 455716
rect 574535 455652 574551 455716
rect 574615 455652 574631 455716
rect 574695 455652 574711 455716
rect 574775 455652 574791 455716
rect 574855 455652 574871 455716
rect 574935 455652 574951 455716
rect 575015 455652 575031 455716
rect 575095 455652 575111 455716
rect 575175 455652 575191 455716
rect 575255 455652 575271 455716
rect 575335 455652 575351 455716
rect 575415 455652 575431 455716
rect 575495 455652 575511 455716
rect 575575 455652 575591 455716
rect 575655 455652 575671 455716
rect 575735 455652 575751 455716
rect 575815 455652 575831 455716
rect 575895 455652 575911 455716
rect 575975 455652 575991 455716
rect 576055 455652 576071 455716
rect 576135 455652 576151 455716
rect 576215 455652 576231 455716
rect 576295 455652 576311 455716
rect 576375 455652 576391 455716
rect 576455 455652 576471 455716
rect 576535 455652 576551 455716
rect 576615 455652 576631 455716
rect 576695 455652 576816 455716
rect 13811 196222 17688 227257
rect 13811 191438 13997 196222
rect 17421 191438 17688 196222
rect 13811 191098 17688 191438
rect 573464 196222 576816 455652
rect 573464 191438 573605 196222
rect 576629 191438 576816 196222
rect 573464 191191 576816 191438
use bandgaptop_flat  bandgaptop_flat_0
timestamp 1622084101
transform 1 0 322204 0 1 615506
box -24404 -1106 20956 27190
<< labels >>
flabel metal3 s 572152 640142 580220 644150 0 FreeSans 20000 0 0 0 VCCD1
flabel metal3 s 567038 550960 577302 554546 0 FreeSans 20000 0 0 0 VDDA1
flabel metal3 s 511190 664896 514962 676272 0 FreeSans 20000 90 0 0 VSSA1
flabel metal3 s 561703 191929 571721 195859 0 FreeSans 20000 0 0 0 VSSD1
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
