magic
tech sky130A
magscale 1 2
timestamp 1620596431
<< locali >>
rect 8400 -5000 8600 5300
rect 9500 -5000 9900 5200
rect 10800 -5000 11200 5200
rect 12100 -5000 12500 5200
rect 13300 -5000 13800 5300
rect 14600 5100 14800 5300
rect 14600 4300 14700 5100
rect 14600 -5000 14800 4300
<< viali >>
rect 14700 4300 14800 5100
<< metal1 >>
rect 11200 8800 11500 8900
rect 8000 8300 9000 8500
rect 8000 7800 8200 8300
rect 8400 7700 8600 8200
rect 8800 7800 9000 8300
rect 9600 8300 10600 8500
rect 9200 7700 9400 8200
rect 9600 7800 9800 8300
rect 8400 7500 9400 7700
rect 10000 7700 10200 8200
rect 10400 7800 10600 8300
rect 11200 8400 11300 8800
rect 11400 8400 11500 8800
rect 13600 8800 14600 8900
rect 13600 8500 13700 8800
rect 14500 8500 14600 8800
rect 10800 7700 11000 8200
rect 11200 7800 11500 8400
rect 11600 8300 12600 8500
rect 11600 7800 11800 8300
rect 10000 7500 11000 7700
rect 12000 7700 12200 8200
rect 12400 7800 12600 8300
rect 13200 8300 14600 8500
rect 12800 7700 13000 8200
rect 13200 7800 13400 8300
rect 12000 7500 13000 7700
rect 13600 7700 13800 8200
rect 14000 7800 14200 8300
rect 14400 7700 14600 8300
rect 13600 7500 14600 7700
rect 9200 7100 10200 7300
rect 7900 6300 8200 7000
rect 7900 6000 8000 6300
rect 8100 6000 8200 6300
rect 7900 5900 8200 6000
rect 8300 6200 8600 7000
rect 8800 6500 9000 7000
rect 9200 6600 9400 7100
rect 9600 6500 9800 7000
rect 10000 6600 10200 7100
rect 10800 7100 12200 7300
rect 12800 7100 14600 7300
rect 8800 6300 9800 6500
rect 10400 6500 10600 7000
rect 10800 6600 11000 7100
rect 11200 6900 11500 7000
rect 11200 6700 11300 6900
rect 11400 6700 11500 6900
rect 11200 6600 11500 6700
rect 11600 6500 11800 7000
rect 12000 6600 12200 7100
rect 10400 6300 11800 6500
rect 12400 6500 12600 7100
rect 12800 6600 13000 7100
rect 13200 6500 13400 7000
rect 13600 6600 13800 7100
rect 14000 6500 14200 7000
rect 14400 6600 14600 7100
rect 12400 6300 14200 6500
rect 8300 4300 9400 6200
rect 11200 6100 11500 6200
rect 11200 5800 11300 6100
rect 11400 5800 11500 6100
rect 11200 5500 11500 5800
rect 11000 5000 11700 5500
rect 14800 5200 15400 5300
rect 14600 5100 15400 5200
rect 10000 3900 14500 5000
rect 14600 4300 14700 5100
rect 14800 4300 15000 5100
rect 14600 4100 15000 4300
rect 15300 4100 15400 5100
rect 14800 3900 15400 4100
rect 10000 3700 14600 3900
rect 8700 -4700 14600 3700
<< via1 >>
rect 11300 8400 11400 8800
rect 13700 8500 14500 8800
rect 8000 6000 8100 6300
rect 11300 6700 11400 6900
rect 11300 5800 11400 6100
rect 15000 4100 15300 5100
<< metal2 >>
rect 7300 8800 11500 8900
rect 7300 8600 11300 8800
rect 7300 6300 7600 8600
rect 11200 8400 11300 8600
rect 11400 8400 11500 8800
rect 13600 8800 15400 8900
rect 13600 8500 13700 8800
rect 14500 8500 15400 8800
rect 13600 8400 15400 8500
rect 11200 8300 11500 8400
rect 11200 6900 11500 7000
rect 11200 6700 11300 6900
rect 11400 6700 11500 6900
rect 7300 6000 8000 6300
rect 8100 6000 8200 6300
rect 7300 5900 8200 6000
rect 11200 6100 11500 6700
rect 11200 5800 11300 6100
rect 11400 5800 11500 6100
rect 11200 5700 11500 5800
rect 14900 5100 15400 8400
rect 14900 4100 15000 5100
rect 15300 4100 15400 5100
rect 14900 4000 15400 4100
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_2
timestamp 1620596431
transform 1 0 8937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_3
timestamp 1620596431
transform 1 0 9337 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_4
timestamp 1620596431
transform 1 0 9737 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_1
timestamp 1620596431
transform 1 0 8537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_0
timestamp 1620596431
transform 1 0 8137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_8
timestamp 1620596431
transform 1 0 11337 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_5
timestamp 1620596431
transform 1 0 10137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_6
timestamp 1620596431
transform 1 0 10537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_7
timestamp 1620596431
transform 1 0 10937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_9
timestamp 1620596431
transform 1 0 11737 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_10
timestamp 1620596431
transform 1 0 12137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_11
timestamp 1620596431
transform 1 0 12537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_12
timestamp 1620596431
transform 1 0 12937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_14
timestamp 1620596431
transform 1 0 13737 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_15
timestamp 1620596431
transform 1 0 14137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_16
timestamp 1620596431
transform 1 0 14537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_13
timestamp 1620596431
transform 1 0 13337 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 7 1288
timestamp 1620596431
transform 1 0 8374 0 1 -5042
box 26 26 1314 1314
<< labels >>
flabel space 11300 7300 11400 7700 1 FreeSans 1600 0 0 0 R3
flabel space 8500 7000 8600 7600 1 FreeSans 1600 0 0 0 R1
flabel metal1 11200 8300 11400 8500 1 FreeSans 1600 0 0 0 Vb
port 1 n
flabel metal2 14900 6100 15400 6400 1 FreeSans 1600 0 0 0 GND!
port 3 n
flabel metal1 8700 5500 9000 5800 1 FreeSans 1600 0 0 0 Va
port 2 n
<< end >>
