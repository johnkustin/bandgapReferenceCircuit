magic
tech sky130A
timestamp 1621317379
<< error_p >>
rect 8083 -9980 8354 -9969
rect 8083 -9983 8340 -9980
rect 8083 -10453 8340 -10439
rect 8343 -10450 8354 -9980
<< pwell >>
rect 8295 -8851 8326 -8782
<< psubdiff >>
rect 8295 -8851 8326 -8782
<< locali >>
rect 8292 -5751 13442 -5651
rect 8292 -6401 13392 -6201
rect 8292 -7051 13392 -6851
rect 8292 -7701 13392 -7501
rect 8292 -8351 13442 -8101
rect 8292 -8781 13442 -8751
rect 8291 -8782 13442 -8781
rect 8291 -8790 8315 -8782
rect 8326 -8790 13442 -8782
rect 8291 -8851 13442 -8790
rect 8291 -8860 8315 -8851
<< metal1 >>
rect 8442 -7056 13292 -5801
rect 8442 -7466 10333 -7056
rect 10362 -7088 10714 -7085
rect 10362 -7434 10365 -7088
rect 10711 -7434 10714 -7088
rect 10362 -7437 10714 -7434
rect 10742 -7466 13292 -7056
rect 8442 -7734 13292 -7466
rect 8442 -8075 12943 -7734
rect 13281 -8075 13292 -7734
rect 8442 -8381 13292 -8075
rect 8442 -8722 12947 -8381
rect 13285 -8722 13292 -8381
rect 8442 -8723 13292 -8722
rect 8083 -9983 8340 -9980
rect 8083 -10453 8340 -10450
<< via1 >>
rect 10365 -7434 10711 -7088
rect 12943 -8075 13281 -7734
rect 12947 -8722 13285 -8381
<< metal2 >>
rect 10362 -7088 10714 -7085
rect 10362 -7434 10365 -7088
rect 10711 -7434 10714 -7088
rect 10362 -9326 10714 -7434
rect 12817 -7734 13291 -7709
rect 12817 -8075 12943 -7734
rect 13281 -8075 13291 -7734
rect 12817 -8381 13291 -8075
rect 12817 -8722 12947 -8381
rect 13285 -8722 13291 -8381
rect 12817 -9957 13291 -8722
rect 8083 -9983 8343 -9980
rect 8340 -10450 8343 -9983
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 644 0 7 644
timestamp 1621270775
transform 0 1 8271 -1 0 -5638
box 13 13 657 657
<< end >>
