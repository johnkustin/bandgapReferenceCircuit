magic
tech sky130A
magscale 1 2
timestamp 1621197215
<< error_p >>
rect -6521 6350 -6481 6950
rect -6461 6350 -6421 6950
rect -5802 6350 -5762 6950
rect -5742 6350 -5702 6950
rect -5083 6350 -5043 6950
rect -5023 6350 -4983 6950
rect -4364 6350 -4324 6950
rect -4304 6350 -4264 6950
rect -3645 6350 -3605 6950
rect -3585 6350 -3545 6950
rect -2926 6350 -2886 6950
rect -2866 6350 -2826 6950
rect -2207 6350 -2167 6950
rect -2147 6350 -2107 6950
rect -1488 6350 -1448 6950
rect -1428 6350 -1388 6950
rect -769 6350 -729 6950
rect -709 6350 -669 6950
rect -50 6350 -10 6950
rect 10 6350 50 6950
rect 669 6350 709 6950
rect 729 6350 769 6950
rect 1388 6350 1428 6950
rect 1448 6350 1488 6950
rect 2107 6350 2147 6950
rect 2167 6350 2207 6950
rect 2826 6350 2866 6950
rect 2886 6350 2926 6950
rect 3545 6350 3585 6950
rect 3605 6350 3645 6950
rect 4264 6350 4304 6950
rect 4324 6350 4364 6950
rect 4983 6350 5023 6950
rect 5043 6350 5083 6950
rect 5702 6350 5742 6950
rect 5762 6350 5802 6950
rect 6421 6350 6461 6950
rect 6481 6350 6521 6950
rect -6521 5650 -6481 6250
rect -6461 5650 -6421 6250
rect -5802 5650 -5762 6250
rect -5742 5650 -5702 6250
rect -5083 5650 -5043 6250
rect -5023 5650 -4983 6250
rect -4364 5650 -4324 6250
rect -4304 5650 -4264 6250
rect -3645 5650 -3605 6250
rect -3585 5650 -3545 6250
rect -2926 5650 -2886 6250
rect -2866 5650 -2826 6250
rect -2207 5650 -2167 6250
rect -2147 5650 -2107 6250
rect -1488 5650 -1448 6250
rect -1428 5650 -1388 6250
rect -769 5650 -729 6250
rect -709 5650 -669 6250
rect -50 5650 -10 6250
rect 10 5650 50 6250
rect 669 5650 709 6250
rect 729 5650 769 6250
rect 1388 5650 1428 6250
rect 1448 5650 1488 6250
rect 2107 5650 2147 6250
rect 2167 5650 2207 6250
rect 2826 5650 2866 6250
rect 2886 5650 2926 6250
rect 3545 5650 3585 6250
rect 3605 5650 3645 6250
rect 4264 5650 4304 6250
rect 4324 5650 4364 6250
rect 4983 5650 5023 6250
rect 5043 5650 5083 6250
rect 5702 5650 5742 6250
rect 5762 5650 5802 6250
rect 6421 5650 6461 6250
rect 6481 5650 6521 6250
rect -6521 4950 -6481 5550
rect -6461 4950 -6421 5550
rect -5802 4950 -5762 5550
rect -5742 4950 -5702 5550
rect -5083 4950 -5043 5550
rect -5023 4950 -4983 5550
rect -4364 4950 -4324 5550
rect -4304 4950 -4264 5550
rect -3645 4950 -3605 5550
rect -3585 4950 -3545 5550
rect -2926 4950 -2886 5550
rect -2866 4950 -2826 5550
rect -2207 4950 -2167 5550
rect -2147 4950 -2107 5550
rect -1488 4950 -1448 5550
rect -1428 4950 -1388 5550
rect -769 4950 -729 5550
rect -709 4950 -669 5550
rect -50 4950 -10 5550
rect 10 4950 50 5550
rect 669 4950 709 5550
rect 729 4950 769 5550
rect 1388 4950 1428 5550
rect 1448 4950 1488 5550
rect 2107 4950 2147 5550
rect 2167 4950 2207 5550
rect 2826 4950 2866 5550
rect 2886 4950 2926 5550
rect 3545 4950 3585 5550
rect 3605 4950 3645 5550
rect 4264 4950 4304 5550
rect 4324 4950 4364 5550
rect 4983 4950 5023 5550
rect 5043 4950 5083 5550
rect 5702 4950 5742 5550
rect 5762 4950 5802 5550
rect 6421 4950 6461 5550
rect 6481 4950 6521 5550
rect -6521 4250 -6481 4850
rect -6461 4250 -6421 4850
rect -5802 4250 -5762 4850
rect -5742 4250 -5702 4850
rect -5083 4250 -5043 4850
rect -5023 4250 -4983 4850
rect -4364 4250 -4324 4850
rect -4304 4250 -4264 4850
rect -3645 4250 -3605 4850
rect -3585 4250 -3545 4850
rect -2926 4250 -2886 4850
rect -2866 4250 -2826 4850
rect -2207 4250 -2167 4850
rect -2147 4250 -2107 4850
rect -1488 4250 -1448 4850
rect -1428 4250 -1388 4850
rect -769 4250 -729 4850
rect -709 4250 -669 4850
rect -50 4250 -10 4850
rect 10 4250 50 4850
rect 669 4250 709 4850
rect 729 4250 769 4850
rect 1388 4250 1428 4850
rect 1448 4250 1488 4850
rect 2107 4250 2147 4850
rect 2167 4250 2207 4850
rect 2826 4250 2866 4850
rect 2886 4250 2926 4850
rect 3545 4250 3585 4850
rect 3605 4250 3645 4850
rect 4264 4250 4304 4850
rect 4324 4250 4364 4850
rect 4983 4250 5023 4850
rect 5043 4250 5083 4850
rect 5702 4250 5742 4850
rect 5762 4250 5802 4850
rect 6421 4250 6461 4850
rect 6481 4250 6521 4850
rect -6521 3550 -6481 4150
rect -6461 3550 -6421 4150
rect -5802 3550 -5762 4150
rect -5742 3550 -5702 4150
rect -5083 3550 -5043 4150
rect -5023 3550 -4983 4150
rect -4364 3550 -4324 4150
rect -4304 3550 -4264 4150
rect -3645 3550 -3605 4150
rect -3585 3550 -3545 4150
rect -2926 3550 -2886 4150
rect -2866 3550 -2826 4150
rect -2207 3550 -2167 4150
rect -2147 3550 -2107 4150
rect -1488 3550 -1448 4150
rect -1428 3550 -1388 4150
rect -769 3550 -729 4150
rect -709 3550 -669 4150
rect -50 3550 -10 4150
rect 10 3550 50 4150
rect 669 3550 709 4150
rect 729 3550 769 4150
rect 1388 3550 1428 4150
rect 1448 3550 1488 4150
rect 2107 3550 2147 4150
rect 2167 3550 2207 4150
rect 2826 3550 2866 4150
rect 2886 3550 2926 4150
rect 3545 3550 3585 4150
rect 3605 3550 3645 4150
rect 4264 3550 4304 4150
rect 4324 3550 4364 4150
rect 4983 3550 5023 4150
rect 5043 3550 5083 4150
rect 5702 3550 5742 4150
rect 5762 3550 5802 4150
rect 6421 3550 6461 4150
rect 6481 3550 6521 4150
rect -6521 2850 -6481 3450
rect -6461 2850 -6421 3450
rect -5802 2850 -5762 3450
rect -5742 2850 -5702 3450
rect -5083 2850 -5043 3450
rect -5023 2850 -4983 3450
rect -4364 2850 -4324 3450
rect -4304 2850 -4264 3450
rect -3645 2850 -3605 3450
rect -3585 2850 -3545 3450
rect -2926 2850 -2886 3450
rect -2866 2850 -2826 3450
rect -2207 2850 -2167 3450
rect -2147 2850 -2107 3450
rect -1488 2850 -1448 3450
rect -1428 2850 -1388 3450
rect -769 2850 -729 3450
rect -709 2850 -669 3450
rect -50 2850 -10 3450
rect 10 2850 50 3450
rect 669 2850 709 3450
rect 729 2850 769 3450
rect 1388 2850 1428 3450
rect 1448 2850 1488 3450
rect 2107 2850 2147 3450
rect 2167 2850 2207 3450
rect 2826 2850 2866 3450
rect 2886 2850 2926 3450
rect 3545 2850 3585 3450
rect 3605 2850 3645 3450
rect 4264 2850 4304 3450
rect 4324 2850 4364 3450
rect 4983 2850 5023 3450
rect 5043 2850 5083 3450
rect 5702 2850 5742 3450
rect 5762 2850 5802 3450
rect 6421 2850 6461 3450
rect 6481 2850 6521 3450
rect -6521 2150 -6481 2750
rect -6461 2150 -6421 2750
rect -5802 2150 -5762 2750
rect -5742 2150 -5702 2750
rect -5083 2150 -5043 2750
rect -5023 2150 -4983 2750
rect -4364 2150 -4324 2750
rect -4304 2150 -4264 2750
rect -3645 2150 -3605 2750
rect -3585 2150 -3545 2750
rect -2926 2150 -2886 2750
rect -2866 2150 -2826 2750
rect -2207 2150 -2167 2750
rect -2147 2150 -2107 2750
rect -1488 2150 -1448 2750
rect -1428 2150 -1388 2750
rect -769 2150 -729 2750
rect -709 2150 -669 2750
rect -50 2150 -10 2750
rect 10 2150 50 2750
rect 669 2150 709 2750
rect 729 2150 769 2750
rect 1388 2150 1428 2750
rect 1448 2150 1488 2750
rect 2107 2150 2147 2750
rect 2167 2150 2207 2750
rect 2826 2150 2866 2750
rect 2886 2150 2926 2750
rect 3545 2150 3585 2750
rect 3605 2150 3645 2750
rect 4264 2150 4304 2750
rect 4324 2150 4364 2750
rect 4983 2150 5023 2750
rect 5043 2150 5083 2750
rect 5702 2150 5742 2750
rect 5762 2150 5802 2750
rect 6421 2150 6461 2750
rect 6481 2150 6521 2750
rect -6521 1450 -6481 2050
rect -6461 1450 -6421 2050
rect -5802 1450 -5762 2050
rect -5742 1450 -5702 2050
rect -5083 1450 -5043 2050
rect -5023 1450 -4983 2050
rect -4364 1450 -4324 2050
rect -4304 1450 -4264 2050
rect -3645 1450 -3605 2050
rect -3585 1450 -3545 2050
rect -2926 1450 -2886 2050
rect -2866 1450 -2826 2050
rect -2207 1450 -2167 2050
rect -2147 1450 -2107 2050
rect -1488 1450 -1448 2050
rect -1428 1450 -1388 2050
rect -769 1450 -729 2050
rect -709 1450 -669 2050
rect -50 1450 -10 2050
rect 10 1450 50 2050
rect 669 1450 709 2050
rect 729 1450 769 2050
rect 1388 1450 1428 2050
rect 1448 1450 1488 2050
rect 2107 1450 2147 2050
rect 2167 1450 2207 2050
rect 2826 1450 2866 2050
rect 2886 1450 2926 2050
rect 3545 1450 3585 2050
rect 3605 1450 3645 2050
rect 4264 1450 4304 2050
rect 4324 1450 4364 2050
rect 4983 1450 5023 2050
rect 5043 1450 5083 2050
rect 5702 1450 5742 2050
rect 5762 1450 5802 2050
rect 6421 1450 6461 2050
rect 6481 1450 6521 2050
rect -6521 750 -6481 1350
rect -6461 750 -6421 1350
rect -5802 750 -5762 1350
rect -5742 750 -5702 1350
rect -5083 750 -5043 1350
rect -5023 750 -4983 1350
rect -4364 750 -4324 1350
rect -4304 750 -4264 1350
rect -3645 750 -3605 1350
rect -3585 750 -3545 1350
rect -2926 750 -2886 1350
rect -2866 750 -2826 1350
rect -2207 750 -2167 1350
rect -2147 750 -2107 1350
rect -1488 750 -1448 1350
rect -1428 750 -1388 1350
rect -769 750 -729 1350
rect -709 750 -669 1350
rect -50 750 -10 1350
rect 10 750 50 1350
rect 669 750 709 1350
rect 729 750 769 1350
rect 1388 750 1428 1350
rect 1448 750 1488 1350
rect 2107 750 2147 1350
rect 2167 750 2207 1350
rect 2826 750 2866 1350
rect 2886 750 2926 1350
rect 3545 750 3585 1350
rect 3605 750 3645 1350
rect 4264 750 4304 1350
rect 4324 750 4364 1350
rect 4983 750 5023 1350
rect 5043 750 5083 1350
rect 5702 750 5742 1350
rect 5762 750 5802 1350
rect 6421 750 6461 1350
rect 6481 750 6521 1350
rect -6521 50 -6481 650
rect -6461 50 -6421 650
rect -5802 50 -5762 650
rect -5742 50 -5702 650
rect -5083 50 -5043 650
rect -5023 50 -4983 650
rect -4364 50 -4324 650
rect -4304 50 -4264 650
rect -3645 50 -3605 650
rect -3585 50 -3545 650
rect -2926 50 -2886 650
rect -2866 50 -2826 650
rect -2207 50 -2167 650
rect -2147 50 -2107 650
rect -1488 50 -1448 650
rect -1428 50 -1388 650
rect -769 50 -729 650
rect -709 50 -669 650
rect -50 50 -10 650
rect 10 50 50 650
rect 669 50 709 650
rect 729 50 769 650
rect 1388 50 1428 650
rect 1448 50 1488 650
rect 2107 50 2147 650
rect 2167 50 2207 650
rect 2826 50 2866 650
rect 2886 50 2926 650
rect 3545 50 3585 650
rect 3605 50 3645 650
rect 4264 50 4304 650
rect 4324 50 4364 650
rect 4983 50 5023 650
rect 5043 50 5083 650
rect 5702 50 5742 650
rect 5762 50 5802 650
rect 6421 50 6461 650
rect 6481 50 6521 650
rect -6521 -650 -6481 -50
rect -6461 -650 -6421 -50
rect -5802 -650 -5762 -50
rect -5742 -650 -5702 -50
rect -5083 -650 -5043 -50
rect -5023 -650 -4983 -50
rect -4364 -650 -4324 -50
rect -4304 -650 -4264 -50
rect -3645 -650 -3605 -50
rect -3585 -650 -3545 -50
rect -2926 -650 -2886 -50
rect -2866 -650 -2826 -50
rect -2207 -650 -2167 -50
rect -2147 -650 -2107 -50
rect -1488 -650 -1448 -50
rect -1428 -650 -1388 -50
rect -769 -650 -729 -50
rect -709 -650 -669 -50
rect -50 -650 -10 -50
rect 10 -650 50 -50
rect 669 -650 709 -50
rect 729 -650 769 -50
rect 1388 -650 1428 -50
rect 1448 -650 1488 -50
rect 2107 -650 2147 -50
rect 2167 -650 2207 -50
rect 2826 -650 2866 -50
rect 2886 -650 2926 -50
rect 3545 -650 3585 -50
rect 3605 -650 3645 -50
rect 4264 -650 4304 -50
rect 4324 -650 4364 -50
rect 4983 -650 5023 -50
rect 5043 -650 5083 -50
rect 5702 -650 5742 -50
rect 5762 -650 5802 -50
rect 6421 -650 6461 -50
rect 6481 -650 6521 -50
rect -6521 -1350 -6481 -750
rect -6461 -1350 -6421 -750
rect -5802 -1350 -5762 -750
rect -5742 -1350 -5702 -750
rect -5083 -1350 -5043 -750
rect -5023 -1350 -4983 -750
rect -4364 -1350 -4324 -750
rect -4304 -1350 -4264 -750
rect -3645 -1350 -3605 -750
rect -3585 -1350 -3545 -750
rect -2926 -1350 -2886 -750
rect -2866 -1350 -2826 -750
rect -2207 -1350 -2167 -750
rect -2147 -1350 -2107 -750
rect -1488 -1350 -1448 -750
rect -1428 -1350 -1388 -750
rect -769 -1350 -729 -750
rect -709 -1350 -669 -750
rect -50 -1350 -10 -750
rect 10 -1350 50 -750
rect 669 -1350 709 -750
rect 729 -1350 769 -750
rect 1388 -1350 1428 -750
rect 1448 -1350 1488 -750
rect 2107 -1350 2147 -750
rect 2167 -1350 2207 -750
rect 2826 -1350 2866 -750
rect 2886 -1350 2926 -750
rect 3545 -1350 3585 -750
rect 3605 -1350 3645 -750
rect 4264 -1350 4304 -750
rect 4324 -1350 4364 -750
rect 4983 -1350 5023 -750
rect 5043 -1350 5083 -750
rect 5702 -1350 5742 -750
rect 5762 -1350 5802 -750
rect 6421 -1350 6461 -750
rect 6481 -1350 6521 -750
rect -6521 -2050 -6481 -1450
rect -6461 -2050 -6421 -1450
rect -5802 -2050 -5762 -1450
rect -5742 -2050 -5702 -1450
rect -5083 -2050 -5043 -1450
rect -5023 -2050 -4983 -1450
rect -4364 -2050 -4324 -1450
rect -4304 -2050 -4264 -1450
rect -3645 -2050 -3605 -1450
rect -3585 -2050 -3545 -1450
rect -2926 -2050 -2886 -1450
rect -2866 -2050 -2826 -1450
rect -2207 -2050 -2167 -1450
rect -2147 -2050 -2107 -1450
rect -1488 -2050 -1448 -1450
rect -1428 -2050 -1388 -1450
rect -769 -2050 -729 -1450
rect -709 -2050 -669 -1450
rect -50 -2050 -10 -1450
rect 10 -2050 50 -1450
rect 669 -2050 709 -1450
rect 729 -2050 769 -1450
rect 1388 -2050 1428 -1450
rect 1448 -2050 1488 -1450
rect 2107 -2050 2147 -1450
rect 2167 -2050 2207 -1450
rect 2826 -2050 2866 -1450
rect 2886 -2050 2926 -1450
rect 3545 -2050 3585 -1450
rect 3605 -2050 3645 -1450
rect 4264 -2050 4304 -1450
rect 4324 -2050 4364 -1450
rect 4983 -2050 5023 -1450
rect 5043 -2050 5083 -1450
rect 5702 -2050 5742 -1450
rect 5762 -2050 5802 -1450
rect 6421 -2050 6461 -1450
rect 6481 -2050 6521 -1450
rect -6521 -2750 -6481 -2150
rect -6461 -2750 -6421 -2150
rect -5802 -2750 -5762 -2150
rect -5742 -2750 -5702 -2150
rect -5083 -2750 -5043 -2150
rect -5023 -2750 -4983 -2150
rect -4364 -2750 -4324 -2150
rect -4304 -2750 -4264 -2150
rect -3645 -2750 -3605 -2150
rect -3585 -2750 -3545 -2150
rect -2926 -2750 -2886 -2150
rect -2866 -2750 -2826 -2150
rect -2207 -2750 -2167 -2150
rect -2147 -2750 -2107 -2150
rect -1488 -2750 -1448 -2150
rect -1428 -2750 -1388 -2150
rect -769 -2750 -729 -2150
rect -709 -2750 -669 -2150
rect -50 -2750 -10 -2150
rect 10 -2750 50 -2150
rect 669 -2750 709 -2150
rect 729 -2750 769 -2150
rect 1388 -2750 1428 -2150
rect 1448 -2750 1488 -2150
rect 2107 -2750 2147 -2150
rect 2167 -2750 2207 -2150
rect 2826 -2750 2866 -2150
rect 2886 -2750 2926 -2150
rect 3545 -2750 3585 -2150
rect 3605 -2750 3645 -2150
rect 4264 -2750 4304 -2150
rect 4324 -2750 4364 -2150
rect 4983 -2750 5023 -2150
rect 5043 -2750 5083 -2150
rect 5702 -2750 5742 -2150
rect 5762 -2750 5802 -2150
rect 6421 -2750 6461 -2150
rect 6481 -2750 6521 -2150
rect -6521 -3450 -6481 -2850
rect -6461 -3450 -6421 -2850
rect -5802 -3450 -5762 -2850
rect -5742 -3450 -5702 -2850
rect -5083 -3450 -5043 -2850
rect -5023 -3450 -4983 -2850
rect -4364 -3450 -4324 -2850
rect -4304 -3450 -4264 -2850
rect -3645 -3450 -3605 -2850
rect -3585 -3450 -3545 -2850
rect -2926 -3450 -2886 -2850
rect -2866 -3450 -2826 -2850
rect -2207 -3450 -2167 -2850
rect -2147 -3450 -2107 -2850
rect -1488 -3450 -1448 -2850
rect -1428 -3450 -1388 -2850
rect -769 -3450 -729 -2850
rect -709 -3450 -669 -2850
rect -50 -3450 -10 -2850
rect 10 -3450 50 -2850
rect 669 -3450 709 -2850
rect 729 -3450 769 -2850
rect 1388 -3450 1428 -2850
rect 1448 -3450 1488 -2850
rect 2107 -3450 2147 -2850
rect 2167 -3450 2207 -2850
rect 2826 -3450 2866 -2850
rect 2886 -3450 2926 -2850
rect 3545 -3450 3585 -2850
rect 3605 -3450 3645 -2850
rect 4264 -3450 4304 -2850
rect 4324 -3450 4364 -2850
rect 4983 -3450 5023 -2850
rect 5043 -3450 5083 -2850
rect 5702 -3450 5742 -2850
rect 5762 -3450 5802 -2850
rect 6421 -3450 6461 -2850
rect 6481 -3450 6521 -2850
rect -6521 -4150 -6481 -3550
rect -6461 -4150 -6421 -3550
rect -5802 -4150 -5762 -3550
rect -5742 -4150 -5702 -3550
rect -5083 -4150 -5043 -3550
rect -5023 -4150 -4983 -3550
rect -4364 -4150 -4324 -3550
rect -4304 -4150 -4264 -3550
rect -3645 -4150 -3605 -3550
rect -3585 -4150 -3545 -3550
rect -2926 -4150 -2886 -3550
rect -2866 -4150 -2826 -3550
rect -2207 -4150 -2167 -3550
rect -2147 -4150 -2107 -3550
rect -1488 -4150 -1448 -3550
rect -1428 -4150 -1388 -3550
rect -769 -4150 -729 -3550
rect -709 -4150 -669 -3550
rect -50 -4150 -10 -3550
rect 10 -4150 50 -3550
rect 669 -4150 709 -3550
rect 729 -4150 769 -3550
rect 1388 -4150 1428 -3550
rect 1448 -4150 1488 -3550
rect 2107 -4150 2147 -3550
rect 2167 -4150 2207 -3550
rect 2826 -4150 2866 -3550
rect 2886 -4150 2926 -3550
rect 3545 -4150 3585 -3550
rect 3605 -4150 3645 -3550
rect 4264 -4150 4304 -3550
rect 4324 -4150 4364 -3550
rect 4983 -4150 5023 -3550
rect 5043 -4150 5083 -3550
rect 5702 -4150 5742 -3550
rect 5762 -4150 5802 -3550
rect 6421 -4150 6461 -3550
rect 6481 -4150 6521 -3550
rect -6521 -4850 -6481 -4250
rect -6461 -4850 -6421 -4250
rect -5802 -4850 -5762 -4250
rect -5742 -4850 -5702 -4250
rect -5083 -4850 -5043 -4250
rect -5023 -4850 -4983 -4250
rect -4364 -4850 -4324 -4250
rect -4304 -4850 -4264 -4250
rect -3645 -4850 -3605 -4250
rect -3585 -4850 -3545 -4250
rect -2926 -4850 -2886 -4250
rect -2866 -4850 -2826 -4250
rect -2207 -4850 -2167 -4250
rect -2147 -4850 -2107 -4250
rect -1488 -4850 -1448 -4250
rect -1428 -4850 -1388 -4250
rect -769 -4850 -729 -4250
rect -709 -4850 -669 -4250
rect -50 -4850 -10 -4250
rect 10 -4850 50 -4250
rect 669 -4850 709 -4250
rect 729 -4850 769 -4250
rect 1388 -4850 1428 -4250
rect 1448 -4850 1488 -4250
rect 2107 -4850 2147 -4250
rect 2167 -4850 2207 -4250
rect 2826 -4850 2866 -4250
rect 2886 -4850 2926 -4250
rect 3545 -4850 3585 -4250
rect 3605 -4850 3645 -4250
rect 4264 -4850 4304 -4250
rect 4324 -4850 4364 -4250
rect 4983 -4850 5023 -4250
rect 5043 -4850 5083 -4250
rect 5702 -4850 5742 -4250
rect 5762 -4850 5802 -4250
rect 6421 -4850 6461 -4250
rect 6481 -4850 6521 -4250
rect -6521 -5550 -6481 -4950
rect -6461 -5550 -6421 -4950
rect -5802 -5550 -5762 -4950
rect -5742 -5550 -5702 -4950
rect -5083 -5550 -5043 -4950
rect -5023 -5550 -4983 -4950
rect -4364 -5550 -4324 -4950
rect -4304 -5550 -4264 -4950
rect -3645 -5550 -3605 -4950
rect -3585 -5550 -3545 -4950
rect -2926 -5550 -2886 -4950
rect -2866 -5550 -2826 -4950
rect -2207 -5550 -2167 -4950
rect -2147 -5550 -2107 -4950
rect -1488 -5550 -1448 -4950
rect -1428 -5550 -1388 -4950
rect -769 -5550 -729 -4950
rect -709 -5550 -669 -4950
rect -50 -5550 -10 -4950
rect 10 -5550 50 -4950
rect 669 -5550 709 -4950
rect 729 -5550 769 -4950
rect 1388 -5550 1428 -4950
rect 1448 -5550 1488 -4950
rect 2107 -5550 2147 -4950
rect 2167 -5550 2207 -4950
rect 2826 -5550 2866 -4950
rect 2886 -5550 2926 -4950
rect 3545 -5550 3585 -4950
rect 3605 -5550 3645 -4950
rect 4264 -5550 4304 -4950
rect 4324 -5550 4364 -4950
rect 4983 -5550 5023 -4950
rect 5043 -5550 5083 -4950
rect 5702 -5550 5742 -4950
rect 5762 -5550 5802 -4950
rect 6421 -5550 6461 -4950
rect 6481 -5550 6521 -4950
rect -6521 -6250 -6481 -5650
rect -6461 -6250 -6421 -5650
rect -5802 -6250 -5762 -5650
rect -5742 -6250 -5702 -5650
rect -5083 -6250 -5043 -5650
rect -5023 -6250 -4983 -5650
rect -4364 -6250 -4324 -5650
rect -4304 -6250 -4264 -5650
rect -3645 -6250 -3605 -5650
rect -3585 -6250 -3545 -5650
rect -2926 -6250 -2886 -5650
rect -2866 -6250 -2826 -5650
rect -2207 -6250 -2167 -5650
rect -2147 -6250 -2107 -5650
rect -1488 -6250 -1448 -5650
rect -1428 -6250 -1388 -5650
rect -769 -6250 -729 -5650
rect -709 -6250 -669 -5650
rect -50 -6250 -10 -5650
rect 10 -6250 50 -5650
rect 669 -6250 709 -5650
rect 729 -6250 769 -5650
rect 1388 -6250 1428 -5650
rect 1448 -6250 1488 -5650
rect 2107 -6250 2147 -5650
rect 2167 -6250 2207 -5650
rect 2826 -6250 2866 -5650
rect 2886 -6250 2926 -5650
rect 3545 -6250 3585 -5650
rect 3605 -6250 3645 -5650
rect 4264 -6250 4304 -5650
rect 4324 -6250 4364 -5650
rect 4983 -6250 5023 -5650
rect 5043 -6250 5083 -5650
rect 5702 -6250 5742 -5650
rect 5762 -6250 5802 -5650
rect 6421 -6250 6461 -5650
rect 6481 -6250 6521 -5650
rect -6521 -6950 -6481 -6350
rect -6461 -6950 -6421 -6350
rect -5802 -6950 -5762 -6350
rect -5742 -6950 -5702 -6350
rect -5083 -6950 -5043 -6350
rect -5023 -6950 -4983 -6350
rect -4364 -6950 -4324 -6350
rect -4304 -6950 -4264 -6350
rect -3645 -6950 -3605 -6350
rect -3585 -6950 -3545 -6350
rect -2926 -6950 -2886 -6350
rect -2866 -6950 -2826 -6350
rect -2207 -6950 -2167 -6350
rect -2147 -6950 -2107 -6350
rect -1488 -6950 -1448 -6350
rect -1428 -6950 -1388 -6350
rect -769 -6950 -729 -6350
rect -709 -6950 -669 -6350
rect -50 -6950 -10 -6350
rect 10 -6950 50 -6350
rect 669 -6950 709 -6350
rect 729 -6950 769 -6350
rect 1388 -6950 1428 -6350
rect 1448 -6950 1488 -6350
rect 2107 -6950 2147 -6350
rect 2167 -6950 2207 -6350
rect 2826 -6950 2866 -6350
rect 2886 -6950 2926 -6350
rect 3545 -6950 3585 -6350
rect 3605 -6950 3645 -6350
rect 4264 -6950 4304 -6350
rect 4324 -6950 4364 -6350
rect 4983 -6950 5023 -6350
rect 5043 -6950 5083 -6350
rect 5702 -6950 5742 -6350
rect 5762 -6950 5802 -6350
rect 6421 -6950 6461 -6350
rect 6481 -6950 6521 -6350
<< metal3 >>
rect -7180 6922 -6481 6950
rect -7180 6378 -6565 6922
rect -6501 6378 -6481 6922
rect -7180 6350 -6481 6378
rect -6461 6922 -5762 6950
rect -6461 6378 -5846 6922
rect -5782 6378 -5762 6922
rect -6461 6350 -5762 6378
rect -5742 6922 -5043 6950
rect -5742 6378 -5127 6922
rect -5063 6378 -5043 6922
rect -5742 6350 -5043 6378
rect -5023 6922 -4324 6950
rect -5023 6378 -4408 6922
rect -4344 6378 -4324 6922
rect -5023 6350 -4324 6378
rect -4304 6922 -3605 6950
rect -4304 6378 -3689 6922
rect -3625 6378 -3605 6922
rect -4304 6350 -3605 6378
rect -3585 6922 -2886 6950
rect -3585 6378 -2970 6922
rect -2906 6378 -2886 6922
rect -3585 6350 -2886 6378
rect -2866 6922 -2167 6950
rect -2866 6378 -2251 6922
rect -2187 6378 -2167 6922
rect -2866 6350 -2167 6378
rect -2147 6922 -1448 6950
rect -2147 6378 -1532 6922
rect -1468 6378 -1448 6922
rect -2147 6350 -1448 6378
rect -1428 6922 -729 6950
rect -1428 6378 -813 6922
rect -749 6378 -729 6922
rect -1428 6350 -729 6378
rect -709 6922 -10 6950
rect -709 6378 -94 6922
rect -30 6378 -10 6922
rect -709 6350 -10 6378
rect 10 6922 709 6950
rect 10 6378 625 6922
rect 689 6378 709 6922
rect 10 6350 709 6378
rect 729 6922 1428 6950
rect 729 6378 1344 6922
rect 1408 6378 1428 6922
rect 729 6350 1428 6378
rect 1448 6922 2147 6950
rect 1448 6378 2063 6922
rect 2127 6378 2147 6922
rect 1448 6350 2147 6378
rect 2167 6922 2866 6950
rect 2167 6378 2782 6922
rect 2846 6378 2866 6922
rect 2167 6350 2866 6378
rect 2886 6922 3585 6950
rect 2886 6378 3501 6922
rect 3565 6378 3585 6922
rect 2886 6350 3585 6378
rect 3605 6922 4304 6950
rect 3605 6378 4220 6922
rect 4284 6378 4304 6922
rect 3605 6350 4304 6378
rect 4324 6922 5023 6950
rect 4324 6378 4939 6922
rect 5003 6378 5023 6922
rect 4324 6350 5023 6378
rect 5043 6922 5742 6950
rect 5043 6378 5658 6922
rect 5722 6378 5742 6922
rect 5043 6350 5742 6378
rect 5762 6922 6461 6950
rect 5762 6378 6377 6922
rect 6441 6378 6461 6922
rect 5762 6350 6461 6378
rect 6481 6922 7180 6950
rect 6481 6378 7096 6922
rect 7160 6378 7180 6922
rect 6481 6350 7180 6378
rect -7180 6222 -6481 6250
rect -7180 5678 -6565 6222
rect -6501 5678 -6481 6222
rect -7180 5650 -6481 5678
rect -6461 6222 -5762 6250
rect -6461 5678 -5846 6222
rect -5782 5678 -5762 6222
rect -6461 5650 -5762 5678
rect -5742 6222 -5043 6250
rect -5742 5678 -5127 6222
rect -5063 5678 -5043 6222
rect -5742 5650 -5043 5678
rect -5023 6222 -4324 6250
rect -5023 5678 -4408 6222
rect -4344 5678 -4324 6222
rect -5023 5650 -4324 5678
rect -4304 6222 -3605 6250
rect -4304 5678 -3689 6222
rect -3625 5678 -3605 6222
rect -4304 5650 -3605 5678
rect -3585 6222 -2886 6250
rect -3585 5678 -2970 6222
rect -2906 5678 -2886 6222
rect -3585 5650 -2886 5678
rect -2866 6222 -2167 6250
rect -2866 5678 -2251 6222
rect -2187 5678 -2167 6222
rect -2866 5650 -2167 5678
rect -2147 6222 -1448 6250
rect -2147 5678 -1532 6222
rect -1468 5678 -1448 6222
rect -2147 5650 -1448 5678
rect -1428 6222 -729 6250
rect -1428 5678 -813 6222
rect -749 5678 -729 6222
rect -1428 5650 -729 5678
rect -709 6222 -10 6250
rect -709 5678 -94 6222
rect -30 5678 -10 6222
rect -709 5650 -10 5678
rect 10 6222 709 6250
rect 10 5678 625 6222
rect 689 5678 709 6222
rect 10 5650 709 5678
rect 729 6222 1428 6250
rect 729 5678 1344 6222
rect 1408 5678 1428 6222
rect 729 5650 1428 5678
rect 1448 6222 2147 6250
rect 1448 5678 2063 6222
rect 2127 5678 2147 6222
rect 1448 5650 2147 5678
rect 2167 6222 2866 6250
rect 2167 5678 2782 6222
rect 2846 5678 2866 6222
rect 2167 5650 2866 5678
rect 2886 6222 3585 6250
rect 2886 5678 3501 6222
rect 3565 5678 3585 6222
rect 2886 5650 3585 5678
rect 3605 6222 4304 6250
rect 3605 5678 4220 6222
rect 4284 5678 4304 6222
rect 3605 5650 4304 5678
rect 4324 6222 5023 6250
rect 4324 5678 4939 6222
rect 5003 5678 5023 6222
rect 4324 5650 5023 5678
rect 5043 6222 5742 6250
rect 5043 5678 5658 6222
rect 5722 5678 5742 6222
rect 5043 5650 5742 5678
rect 5762 6222 6461 6250
rect 5762 5678 6377 6222
rect 6441 5678 6461 6222
rect 5762 5650 6461 5678
rect 6481 6222 7180 6250
rect 6481 5678 7096 6222
rect 7160 5678 7180 6222
rect 6481 5650 7180 5678
rect -7180 5522 -6481 5550
rect -7180 4978 -6565 5522
rect -6501 4978 -6481 5522
rect -7180 4950 -6481 4978
rect -6461 5522 -5762 5550
rect -6461 4978 -5846 5522
rect -5782 4978 -5762 5522
rect -6461 4950 -5762 4978
rect -5742 5522 -5043 5550
rect -5742 4978 -5127 5522
rect -5063 4978 -5043 5522
rect -5742 4950 -5043 4978
rect -5023 5522 -4324 5550
rect -5023 4978 -4408 5522
rect -4344 4978 -4324 5522
rect -5023 4950 -4324 4978
rect -4304 5522 -3605 5550
rect -4304 4978 -3689 5522
rect -3625 4978 -3605 5522
rect -4304 4950 -3605 4978
rect -3585 5522 -2886 5550
rect -3585 4978 -2970 5522
rect -2906 4978 -2886 5522
rect -3585 4950 -2886 4978
rect -2866 5522 -2167 5550
rect -2866 4978 -2251 5522
rect -2187 4978 -2167 5522
rect -2866 4950 -2167 4978
rect -2147 5522 -1448 5550
rect -2147 4978 -1532 5522
rect -1468 4978 -1448 5522
rect -2147 4950 -1448 4978
rect -1428 5522 -729 5550
rect -1428 4978 -813 5522
rect -749 4978 -729 5522
rect -1428 4950 -729 4978
rect -709 5522 -10 5550
rect -709 4978 -94 5522
rect -30 4978 -10 5522
rect -709 4950 -10 4978
rect 10 5522 709 5550
rect 10 4978 625 5522
rect 689 4978 709 5522
rect 10 4950 709 4978
rect 729 5522 1428 5550
rect 729 4978 1344 5522
rect 1408 4978 1428 5522
rect 729 4950 1428 4978
rect 1448 5522 2147 5550
rect 1448 4978 2063 5522
rect 2127 4978 2147 5522
rect 1448 4950 2147 4978
rect 2167 5522 2866 5550
rect 2167 4978 2782 5522
rect 2846 4978 2866 5522
rect 2167 4950 2866 4978
rect 2886 5522 3585 5550
rect 2886 4978 3501 5522
rect 3565 4978 3585 5522
rect 2886 4950 3585 4978
rect 3605 5522 4304 5550
rect 3605 4978 4220 5522
rect 4284 4978 4304 5522
rect 3605 4950 4304 4978
rect 4324 5522 5023 5550
rect 4324 4978 4939 5522
rect 5003 4978 5023 5522
rect 4324 4950 5023 4978
rect 5043 5522 5742 5550
rect 5043 4978 5658 5522
rect 5722 4978 5742 5522
rect 5043 4950 5742 4978
rect 5762 5522 6461 5550
rect 5762 4978 6377 5522
rect 6441 4978 6461 5522
rect 5762 4950 6461 4978
rect 6481 5522 7180 5550
rect 6481 4978 7096 5522
rect 7160 4978 7180 5522
rect 6481 4950 7180 4978
rect -7180 4822 -6481 4850
rect -7180 4278 -6565 4822
rect -6501 4278 -6481 4822
rect -7180 4250 -6481 4278
rect -6461 4822 -5762 4850
rect -6461 4278 -5846 4822
rect -5782 4278 -5762 4822
rect -6461 4250 -5762 4278
rect -5742 4822 -5043 4850
rect -5742 4278 -5127 4822
rect -5063 4278 -5043 4822
rect -5742 4250 -5043 4278
rect -5023 4822 -4324 4850
rect -5023 4278 -4408 4822
rect -4344 4278 -4324 4822
rect -5023 4250 -4324 4278
rect -4304 4822 -3605 4850
rect -4304 4278 -3689 4822
rect -3625 4278 -3605 4822
rect -4304 4250 -3605 4278
rect -3585 4822 -2886 4850
rect -3585 4278 -2970 4822
rect -2906 4278 -2886 4822
rect -3585 4250 -2886 4278
rect -2866 4822 -2167 4850
rect -2866 4278 -2251 4822
rect -2187 4278 -2167 4822
rect -2866 4250 -2167 4278
rect -2147 4822 -1448 4850
rect -2147 4278 -1532 4822
rect -1468 4278 -1448 4822
rect -2147 4250 -1448 4278
rect -1428 4822 -729 4850
rect -1428 4278 -813 4822
rect -749 4278 -729 4822
rect -1428 4250 -729 4278
rect -709 4822 -10 4850
rect -709 4278 -94 4822
rect -30 4278 -10 4822
rect -709 4250 -10 4278
rect 10 4822 709 4850
rect 10 4278 625 4822
rect 689 4278 709 4822
rect 10 4250 709 4278
rect 729 4822 1428 4850
rect 729 4278 1344 4822
rect 1408 4278 1428 4822
rect 729 4250 1428 4278
rect 1448 4822 2147 4850
rect 1448 4278 2063 4822
rect 2127 4278 2147 4822
rect 1448 4250 2147 4278
rect 2167 4822 2866 4850
rect 2167 4278 2782 4822
rect 2846 4278 2866 4822
rect 2167 4250 2866 4278
rect 2886 4822 3585 4850
rect 2886 4278 3501 4822
rect 3565 4278 3585 4822
rect 2886 4250 3585 4278
rect 3605 4822 4304 4850
rect 3605 4278 4220 4822
rect 4284 4278 4304 4822
rect 3605 4250 4304 4278
rect 4324 4822 5023 4850
rect 4324 4278 4939 4822
rect 5003 4278 5023 4822
rect 4324 4250 5023 4278
rect 5043 4822 5742 4850
rect 5043 4278 5658 4822
rect 5722 4278 5742 4822
rect 5043 4250 5742 4278
rect 5762 4822 6461 4850
rect 5762 4278 6377 4822
rect 6441 4278 6461 4822
rect 5762 4250 6461 4278
rect 6481 4822 7180 4850
rect 6481 4278 7096 4822
rect 7160 4278 7180 4822
rect 6481 4250 7180 4278
rect -7180 4122 -6481 4150
rect -7180 3578 -6565 4122
rect -6501 3578 -6481 4122
rect -7180 3550 -6481 3578
rect -6461 4122 -5762 4150
rect -6461 3578 -5846 4122
rect -5782 3578 -5762 4122
rect -6461 3550 -5762 3578
rect -5742 4122 -5043 4150
rect -5742 3578 -5127 4122
rect -5063 3578 -5043 4122
rect -5742 3550 -5043 3578
rect -5023 4122 -4324 4150
rect -5023 3578 -4408 4122
rect -4344 3578 -4324 4122
rect -5023 3550 -4324 3578
rect -4304 4122 -3605 4150
rect -4304 3578 -3689 4122
rect -3625 3578 -3605 4122
rect -4304 3550 -3605 3578
rect -3585 4122 -2886 4150
rect -3585 3578 -2970 4122
rect -2906 3578 -2886 4122
rect -3585 3550 -2886 3578
rect -2866 4122 -2167 4150
rect -2866 3578 -2251 4122
rect -2187 3578 -2167 4122
rect -2866 3550 -2167 3578
rect -2147 4122 -1448 4150
rect -2147 3578 -1532 4122
rect -1468 3578 -1448 4122
rect -2147 3550 -1448 3578
rect -1428 4122 -729 4150
rect -1428 3578 -813 4122
rect -749 3578 -729 4122
rect -1428 3550 -729 3578
rect -709 4122 -10 4150
rect -709 3578 -94 4122
rect -30 3578 -10 4122
rect -709 3550 -10 3578
rect 10 4122 709 4150
rect 10 3578 625 4122
rect 689 3578 709 4122
rect 10 3550 709 3578
rect 729 4122 1428 4150
rect 729 3578 1344 4122
rect 1408 3578 1428 4122
rect 729 3550 1428 3578
rect 1448 4122 2147 4150
rect 1448 3578 2063 4122
rect 2127 3578 2147 4122
rect 1448 3550 2147 3578
rect 2167 4122 2866 4150
rect 2167 3578 2782 4122
rect 2846 3578 2866 4122
rect 2167 3550 2866 3578
rect 2886 4122 3585 4150
rect 2886 3578 3501 4122
rect 3565 3578 3585 4122
rect 2886 3550 3585 3578
rect 3605 4122 4304 4150
rect 3605 3578 4220 4122
rect 4284 3578 4304 4122
rect 3605 3550 4304 3578
rect 4324 4122 5023 4150
rect 4324 3578 4939 4122
rect 5003 3578 5023 4122
rect 4324 3550 5023 3578
rect 5043 4122 5742 4150
rect 5043 3578 5658 4122
rect 5722 3578 5742 4122
rect 5043 3550 5742 3578
rect 5762 4122 6461 4150
rect 5762 3578 6377 4122
rect 6441 3578 6461 4122
rect 5762 3550 6461 3578
rect 6481 4122 7180 4150
rect 6481 3578 7096 4122
rect 7160 3578 7180 4122
rect 6481 3550 7180 3578
rect -7180 3422 -6481 3450
rect -7180 2878 -6565 3422
rect -6501 2878 -6481 3422
rect -7180 2850 -6481 2878
rect -6461 3422 -5762 3450
rect -6461 2878 -5846 3422
rect -5782 2878 -5762 3422
rect -6461 2850 -5762 2878
rect -5742 3422 -5043 3450
rect -5742 2878 -5127 3422
rect -5063 2878 -5043 3422
rect -5742 2850 -5043 2878
rect -5023 3422 -4324 3450
rect -5023 2878 -4408 3422
rect -4344 2878 -4324 3422
rect -5023 2850 -4324 2878
rect -4304 3422 -3605 3450
rect -4304 2878 -3689 3422
rect -3625 2878 -3605 3422
rect -4304 2850 -3605 2878
rect -3585 3422 -2886 3450
rect -3585 2878 -2970 3422
rect -2906 2878 -2886 3422
rect -3585 2850 -2886 2878
rect -2866 3422 -2167 3450
rect -2866 2878 -2251 3422
rect -2187 2878 -2167 3422
rect -2866 2850 -2167 2878
rect -2147 3422 -1448 3450
rect -2147 2878 -1532 3422
rect -1468 2878 -1448 3422
rect -2147 2850 -1448 2878
rect -1428 3422 -729 3450
rect -1428 2878 -813 3422
rect -749 2878 -729 3422
rect -1428 2850 -729 2878
rect -709 3422 -10 3450
rect -709 2878 -94 3422
rect -30 2878 -10 3422
rect -709 2850 -10 2878
rect 10 3422 709 3450
rect 10 2878 625 3422
rect 689 2878 709 3422
rect 10 2850 709 2878
rect 729 3422 1428 3450
rect 729 2878 1344 3422
rect 1408 2878 1428 3422
rect 729 2850 1428 2878
rect 1448 3422 2147 3450
rect 1448 2878 2063 3422
rect 2127 2878 2147 3422
rect 1448 2850 2147 2878
rect 2167 3422 2866 3450
rect 2167 2878 2782 3422
rect 2846 2878 2866 3422
rect 2167 2850 2866 2878
rect 2886 3422 3585 3450
rect 2886 2878 3501 3422
rect 3565 2878 3585 3422
rect 2886 2850 3585 2878
rect 3605 3422 4304 3450
rect 3605 2878 4220 3422
rect 4284 2878 4304 3422
rect 3605 2850 4304 2878
rect 4324 3422 5023 3450
rect 4324 2878 4939 3422
rect 5003 2878 5023 3422
rect 4324 2850 5023 2878
rect 5043 3422 5742 3450
rect 5043 2878 5658 3422
rect 5722 2878 5742 3422
rect 5043 2850 5742 2878
rect 5762 3422 6461 3450
rect 5762 2878 6377 3422
rect 6441 2878 6461 3422
rect 5762 2850 6461 2878
rect 6481 3422 7180 3450
rect 6481 2878 7096 3422
rect 7160 2878 7180 3422
rect 6481 2850 7180 2878
rect -7180 2722 -6481 2750
rect -7180 2178 -6565 2722
rect -6501 2178 -6481 2722
rect -7180 2150 -6481 2178
rect -6461 2722 -5762 2750
rect -6461 2178 -5846 2722
rect -5782 2178 -5762 2722
rect -6461 2150 -5762 2178
rect -5742 2722 -5043 2750
rect -5742 2178 -5127 2722
rect -5063 2178 -5043 2722
rect -5742 2150 -5043 2178
rect -5023 2722 -4324 2750
rect -5023 2178 -4408 2722
rect -4344 2178 -4324 2722
rect -5023 2150 -4324 2178
rect -4304 2722 -3605 2750
rect -4304 2178 -3689 2722
rect -3625 2178 -3605 2722
rect -4304 2150 -3605 2178
rect -3585 2722 -2886 2750
rect -3585 2178 -2970 2722
rect -2906 2178 -2886 2722
rect -3585 2150 -2886 2178
rect -2866 2722 -2167 2750
rect -2866 2178 -2251 2722
rect -2187 2178 -2167 2722
rect -2866 2150 -2167 2178
rect -2147 2722 -1448 2750
rect -2147 2178 -1532 2722
rect -1468 2178 -1448 2722
rect -2147 2150 -1448 2178
rect -1428 2722 -729 2750
rect -1428 2178 -813 2722
rect -749 2178 -729 2722
rect -1428 2150 -729 2178
rect -709 2722 -10 2750
rect -709 2178 -94 2722
rect -30 2178 -10 2722
rect -709 2150 -10 2178
rect 10 2722 709 2750
rect 10 2178 625 2722
rect 689 2178 709 2722
rect 10 2150 709 2178
rect 729 2722 1428 2750
rect 729 2178 1344 2722
rect 1408 2178 1428 2722
rect 729 2150 1428 2178
rect 1448 2722 2147 2750
rect 1448 2178 2063 2722
rect 2127 2178 2147 2722
rect 1448 2150 2147 2178
rect 2167 2722 2866 2750
rect 2167 2178 2782 2722
rect 2846 2178 2866 2722
rect 2167 2150 2866 2178
rect 2886 2722 3585 2750
rect 2886 2178 3501 2722
rect 3565 2178 3585 2722
rect 2886 2150 3585 2178
rect 3605 2722 4304 2750
rect 3605 2178 4220 2722
rect 4284 2178 4304 2722
rect 3605 2150 4304 2178
rect 4324 2722 5023 2750
rect 4324 2178 4939 2722
rect 5003 2178 5023 2722
rect 4324 2150 5023 2178
rect 5043 2722 5742 2750
rect 5043 2178 5658 2722
rect 5722 2178 5742 2722
rect 5043 2150 5742 2178
rect 5762 2722 6461 2750
rect 5762 2178 6377 2722
rect 6441 2178 6461 2722
rect 5762 2150 6461 2178
rect 6481 2722 7180 2750
rect 6481 2178 7096 2722
rect 7160 2178 7180 2722
rect 6481 2150 7180 2178
rect -7180 2022 -6481 2050
rect -7180 1478 -6565 2022
rect -6501 1478 -6481 2022
rect -7180 1450 -6481 1478
rect -6461 2022 -5762 2050
rect -6461 1478 -5846 2022
rect -5782 1478 -5762 2022
rect -6461 1450 -5762 1478
rect -5742 2022 -5043 2050
rect -5742 1478 -5127 2022
rect -5063 1478 -5043 2022
rect -5742 1450 -5043 1478
rect -5023 2022 -4324 2050
rect -5023 1478 -4408 2022
rect -4344 1478 -4324 2022
rect -5023 1450 -4324 1478
rect -4304 2022 -3605 2050
rect -4304 1478 -3689 2022
rect -3625 1478 -3605 2022
rect -4304 1450 -3605 1478
rect -3585 2022 -2886 2050
rect -3585 1478 -2970 2022
rect -2906 1478 -2886 2022
rect -3585 1450 -2886 1478
rect -2866 2022 -2167 2050
rect -2866 1478 -2251 2022
rect -2187 1478 -2167 2022
rect -2866 1450 -2167 1478
rect -2147 2022 -1448 2050
rect -2147 1478 -1532 2022
rect -1468 1478 -1448 2022
rect -2147 1450 -1448 1478
rect -1428 2022 -729 2050
rect -1428 1478 -813 2022
rect -749 1478 -729 2022
rect -1428 1450 -729 1478
rect -709 2022 -10 2050
rect -709 1478 -94 2022
rect -30 1478 -10 2022
rect -709 1450 -10 1478
rect 10 2022 709 2050
rect 10 1478 625 2022
rect 689 1478 709 2022
rect 10 1450 709 1478
rect 729 2022 1428 2050
rect 729 1478 1344 2022
rect 1408 1478 1428 2022
rect 729 1450 1428 1478
rect 1448 2022 2147 2050
rect 1448 1478 2063 2022
rect 2127 1478 2147 2022
rect 1448 1450 2147 1478
rect 2167 2022 2866 2050
rect 2167 1478 2782 2022
rect 2846 1478 2866 2022
rect 2167 1450 2866 1478
rect 2886 2022 3585 2050
rect 2886 1478 3501 2022
rect 3565 1478 3585 2022
rect 2886 1450 3585 1478
rect 3605 2022 4304 2050
rect 3605 1478 4220 2022
rect 4284 1478 4304 2022
rect 3605 1450 4304 1478
rect 4324 2022 5023 2050
rect 4324 1478 4939 2022
rect 5003 1478 5023 2022
rect 4324 1450 5023 1478
rect 5043 2022 5742 2050
rect 5043 1478 5658 2022
rect 5722 1478 5742 2022
rect 5043 1450 5742 1478
rect 5762 2022 6461 2050
rect 5762 1478 6377 2022
rect 6441 1478 6461 2022
rect 5762 1450 6461 1478
rect 6481 2022 7180 2050
rect 6481 1478 7096 2022
rect 7160 1478 7180 2022
rect 6481 1450 7180 1478
rect -7180 1322 -6481 1350
rect -7180 778 -6565 1322
rect -6501 778 -6481 1322
rect -7180 750 -6481 778
rect -6461 1322 -5762 1350
rect -6461 778 -5846 1322
rect -5782 778 -5762 1322
rect -6461 750 -5762 778
rect -5742 1322 -5043 1350
rect -5742 778 -5127 1322
rect -5063 778 -5043 1322
rect -5742 750 -5043 778
rect -5023 1322 -4324 1350
rect -5023 778 -4408 1322
rect -4344 778 -4324 1322
rect -5023 750 -4324 778
rect -4304 1322 -3605 1350
rect -4304 778 -3689 1322
rect -3625 778 -3605 1322
rect -4304 750 -3605 778
rect -3585 1322 -2886 1350
rect -3585 778 -2970 1322
rect -2906 778 -2886 1322
rect -3585 750 -2886 778
rect -2866 1322 -2167 1350
rect -2866 778 -2251 1322
rect -2187 778 -2167 1322
rect -2866 750 -2167 778
rect -2147 1322 -1448 1350
rect -2147 778 -1532 1322
rect -1468 778 -1448 1322
rect -2147 750 -1448 778
rect -1428 1322 -729 1350
rect -1428 778 -813 1322
rect -749 778 -729 1322
rect -1428 750 -729 778
rect -709 1322 -10 1350
rect -709 778 -94 1322
rect -30 778 -10 1322
rect -709 750 -10 778
rect 10 1322 709 1350
rect 10 778 625 1322
rect 689 778 709 1322
rect 10 750 709 778
rect 729 1322 1428 1350
rect 729 778 1344 1322
rect 1408 778 1428 1322
rect 729 750 1428 778
rect 1448 1322 2147 1350
rect 1448 778 2063 1322
rect 2127 778 2147 1322
rect 1448 750 2147 778
rect 2167 1322 2866 1350
rect 2167 778 2782 1322
rect 2846 778 2866 1322
rect 2167 750 2866 778
rect 2886 1322 3585 1350
rect 2886 778 3501 1322
rect 3565 778 3585 1322
rect 2886 750 3585 778
rect 3605 1322 4304 1350
rect 3605 778 4220 1322
rect 4284 778 4304 1322
rect 3605 750 4304 778
rect 4324 1322 5023 1350
rect 4324 778 4939 1322
rect 5003 778 5023 1322
rect 4324 750 5023 778
rect 5043 1322 5742 1350
rect 5043 778 5658 1322
rect 5722 778 5742 1322
rect 5043 750 5742 778
rect 5762 1322 6461 1350
rect 5762 778 6377 1322
rect 6441 778 6461 1322
rect 5762 750 6461 778
rect 6481 1322 7180 1350
rect 6481 778 7096 1322
rect 7160 778 7180 1322
rect 6481 750 7180 778
rect -7180 622 -6481 650
rect -7180 78 -6565 622
rect -6501 78 -6481 622
rect -7180 50 -6481 78
rect -6461 622 -5762 650
rect -6461 78 -5846 622
rect -5782 78 -5762 622
rect -6461 50 -5762 78
rect -5742 622 -5043 650
rect -5742 78 -5127 622
rect -5063 78 -5043 622
rect -5742 50 -5043 78
rect -5023 622 -4324 650
rect -5023 78 -4408 622
rect -4344 78 -4324 622
rect -5023 50 -4324 78
rect -4304 622 -3605 650
rect -4304 78 -3689 622
rect -3625 78 -3605 622
rect -4304 50 -3605 78
rect -3585 622 -2886 650
rect -3585 78 -2970 622
rect -2906 78 -2886 622
rect -3585 50 -2886 78
rect -2866 622 -2167 650
rect -2866 78 -2251 622
rect -2187 78 -2167 622
rect -2866 50 -2167 78
rect -2147 622 -1448 650
rect -2147 78 -1532 622
rect -1468 78 -1448 622
rect -2147 50 -1448 78
rect -1428 622 -729 650
rect -1428 78 -813 622
rect -749 78 -729 622
rect -1428 50 -729 78
rect -709 622 -10 650
rect -709 78 -94 622
rect -30 78 -10 622
rect -709 50 -10 78
rect 10 622 709 650
rect 10 78 625 622
rect 689 78 709 622
rect 10 50 709 78
rect 729 622 1428 650
rect 729 78 1344 622
rect 1408 78 1428 622
rect 729 50 1428 78
rect 1448 622 2147 650
rect 1448 78 2063 622
rect 2127 78 2147 622
rect 1448 50 2147 78
rect 2167 622 2866 650
rect 2167 78 2782 622
rect 2846 78 2866 622
rect 2167 50 2866 78
rect 2886 622 3585 650
rect 2886 78 3501 622
rect 3565 78 3585 622
rect 2886 50 3585 78
rect 3605 622 4304 650
rect 3605 78 4220 622
rect 4284 78 4304 622
rect 3605 50 4304 78
rect 4324 622 5023 650
rect 4324 78 4939 622
rect 5003 78 5023 622
rect 4324 50 5023 78
rect 5043 622 5742 650
rect 5043 78 5658 622
rect 5722 78 5742 622
rect 5043 50 5742 78
rect 5762 622 6461 650
rect 5762 78 6377 622
rect 6441 78 6461 622
rect 5762 50 6461 78
rect 6481 622 7180 650
rect 6481 78 7096 622
rect 7160 78 7180 622
rect 6481 50 7180 78
rect -7180 -78 -6481 -50
rect -7180 -622 -6565 -78
rect -6501 -622 -6481 -78
rect -7180 -650 -6481 -622
rect -6461 -78 -5762 -50
rect -6461 -622 -5846 -78
rect -5782 -622 -5762 -78
rect -6461 -650 -5762 -622
rect -5742 -78 -5043 -50
rect -5742 -622 -5127 -78
rect -5063 -622 -5043 -78
rect -5742 -650 -5043 -622
rect -5023 -78 -4324 -50
rect -5023 -622 -4408 -78
rect -4344 -622 -4324 -78
rect -5023 -650 -4324 -622
rect -4304 -78 -3605 -50
rect -4304 -622 -3689 -78
rect -3625 -622 -3605 -78
rect -4304 -650 -3605 -622
rect -3585 -78 -2886 -50
rect -3585 -622 -2970 -78
rect -2906 -622 -2886 -78
rect -3585 -650 -2886 -622
rect -2866 -78 -2167 -50
rect -2866 -622 -2251 -78
rect -2187 -622 -2167 -78
rect -2866 -650 -2167 -622
rect -2147 -78 -1448 -50
rect -2147 -622 -1532 -78
rect -1468 -622 -1448 -78
rect -2147 -650 -1448 -622
rect -1428 -78 -729 -50
rect -1428 -622 -813 -78
rect -749 -622 -729 -78
rect -1428 -650 -729 -622
rect -709 -78 -10 -50
rect -709 -622 -94 -78
rect -30 -622 -10 -78
rect -709 -650 -10 -622
rect 10 -78 709 -50
rect 10 -622 625 -78
rect 689 -622 709 -78
rect 10 -650 709 -622
rect 729 -78 1428 -50
rect 729 -622 1344 -78
rect 1408 -622 1428 -78
rect 729 -650 1428 -622
rect 1448 -78 2147 -50
rect 1448 -622 2063 -78
rect 2127 -622 2147 -78
rect 1448 -650 2147 -622
rect 2167 -78 2866 -50
rect 2167 -622 2782 -78
rect 2846 -622 2866 -78
rect 2167 -650 2866 -622
rect 2886 -78 3585 -50
rect 2886 -622 3501 -78
rect 3565 -622 3585 -78
rect 2886 -650 3585 -622
rect 3605 -78 4304 -50
rect 3605 -622 4220 -78
rect 4284 -622 4304 -78
rect 3605 -650 4304 -622
rect 4324 -78 5023 -50
rect 4324 -622 4939 -78
rect 5003 -622 5023 -78
rect 4324 -650 5023 -622
rect 5043 -78 5742 -50
rect 5043 -622 5658 -78
rect 5722 -622 5742 -78
rect 5043 -650 5742 -622
rect 5762 -78 6461 -50
rect 5762 -622 6377 -78
rect 6441 -622 6461 -78
rect 5762 -650 6461 -622
rect 6481 -78 7180 -50
rect 6481 -622 7096 -78
rect 7160 -622 7180 -78
rect 6481 -650 7180 -622
rect -7180 -778 -6481 -750
rect -7180 -1322 -6565 -778
rect -6501 -1322 -6481 -778
rect -7180 -1350 -6481 -1322
rect -6461 -778 -5762 -750
rect -6461 -1322 -5846 -778
rect -5782 -1322 -5762 -778
rect -6461 -1350 -5762 -1322
rect -5742 -778 -5043 -750
rect -5742 -1322 -5127 -778
rect -5063 -1322 -5043 -778
rect -5742 -1350 -5043 -1322
rect -5023 -778 -4324 -750
rect -5023 -1322 -4408 -778
rect -4344 -1322 -4324 -778
rect -5023 -1350 -4324 -1322
rect -4304 -778 -3605 -750
rect -4304 -1322 -3689 -778
rect -3625 -1322 -3605 -778
rect -4304 -1350 -3605 -1322
rect -3585 -778 -2886 -750
rect -3585 -1322 -2970 -778
rect -2906 -1322 -2886 -778
rect -3585 -1350 -2886 -1322
rect -2866 -778 -2167 -750
rect -2866 -1322 -2251 -778
rect -2187 -1322 -2167 -778
rect -2866 -1350 -2167 -1322
rect -2147 -778 -1448 -750
rect -2147 -1322 -1532 -778
rect -1468 -1322 -1448 -778
rect -2147 -1350 -1448 -1322
rect -1428 -778 -729 -750
rect -1428 -1322 -813 -778
rect -749 -1322 -729 -778
rect -1428 -1350 -729 -1322
rect -709 -778 -10 -750
rect -709 -1322 -94 -778
rect -30 -1322 -10 -778
rect -709 -1350 -10 -1322
rect 10 -778 709 -750
rect 10 -1322 625 -778
rect 689 -1322 709 -778
rect 10 -1350 709 -1322
rect 729 -778 1428 -750
rect 729 -1322 1344 -778
rect 1408 -1322 1428 -778
rect 729 -1350 1428 -1322
rect 1448 -778 2147 -750
rect 1448 -1322 2063 -778
rect 2127 -1322 2147 -778
rect 1448 -1350 2147 -1322
rect 2167 -778 2866 -750
rect 2167 -1322 2782 -778
rect 2846 -1322 2866 -778
rect 2167 -1350 2866 -1322
rect 2886 -778 3585 -750
rect 2886 -1322 3501 -778
rect 3565 -1322 3585 -778
rect 2886 -1350 3585 -1322
rect 3605 -778 4304 -750
rect 3605 -1322 4220 -778
rect 4284 -1322 4304 -778
rect 3605 -1350 4304 -1322
rect 4324 -778 5023 -750
rect 4324 -1322 4939 -778
rect 5003 -1322 5023 -778
rect 4324 -1350 5023 -1322
rect 5043 -778 5742 -750
rect 5043 -1322 5658 -778
rect 5722 -1322 5742 -778
rect 5043 -1350 5742 -1322
rect 5762 -778 6461 -750
rect 5762 -1322 6377 -778
rect 6441 -1322 6461 -778
rect 5762 -1350 6461 -1322
rect 6481 -778 7180 -750
rect 6481 -1322 7096 -778
rect 7160 -1322 7180 -778
rect 6481 -1350 7180 -1322
rect -7180 -1478 -6481 -1450
rect -7180 -2022 -6565 -1478
rect -6501 -2022 -6481 -1478
rect -7180 -2050 -6481 -2022
rect -6461 -1478 -5762 -1450
rect -6461 -2022 -5846 -1478
rect -5782 -2022 -5762 -1478
rect -6461 -2050 -5762 -2022
rect -5742 -1478 -5043 -1450
rect -5742 -2022 -5127 -1478
rect -5063 -2022 -5043 -1478
rect -5742 -2050 -5043 -2022
rect -5023 -1478 -4324 -1450
rect -5023 -2022 -4408 -1478
rect -4344 -2022 -4324 -1478
rect -5023 -2050 -4324 -2022
rect -4304 -1478 -3605 -1450
rect -4304 -2022 -3689 -1478
rect -3625 -2022 -3605 -1478
rect -4304 -2050 -3605 -2022
rect -3585 -1478 -2886 -1450
rect -3585 -2022 -2970 -1478
rect -2906 -2022 -2886 -1478
rect -3585 -2050 -2886 -2022
rect -2866 -1478 -2167 -1450
rect -2866 -2022 -2251 -1478
rect -2187 -2022 -2167 -1478
rect -2866 -2050 -2167 -2022
rect -2147 -1478 -1448 -1450
rect -2147 -2022 -1532 -1478
rect -1468 -2022 -1448 -1478
rect -2147 -2050 -1448 -2022
rect -1428 -1478 -729 -1450
rect -1428 -2022 -813 -1478
rect -749 -2022 -729 -1478
rect -1428 -2050 -729 -2022
rect -709 -1478 -10 -1450
rect -709 -2022 -94 -1478
rect -30 -2022 -10 -1478
rect -709 -2050 -10 -2022
rect 10 -1478 709 -1450
rect 10 -2022 625 -1478
rect 689 -2022 709 -1478
rect 10 -2050 709 -2022
rect 729 -1478 1428 -1450
rect 729 -2022 1344 -1478
rect 1408 -2022 1428 -1478
rect 729 -2050 1428 -2022
rect 1448 -1478 2147 -1450
rect 1448 -2022 2063 -1478
rect 2127 -2022 2147 -1478
rect 1448 -2050 2147 -2022
rect 2167 -1478 2866 -1450
rect 2167 -2022 2782 -1478
rect 2846 -2022 2866 -1478
rect 2167 -2050 2866 -2022
rect 2886 -1478 3585 -1450
rect 2886 -2022 3501 -1478
rect 3565 -2022 3585 -1478
rect 2886 -2050 3585 -2022
rect 3605 -1478 4304 -1450
rect 3605 -2022 4220 -1478
rect 4284 -2022 4304 -1478
rect 3605 -2050 4304 -2022
rect 4324 -1478 5023 -1450
rect 4324 -2022 4939 -1478
rect 5003 -2022 5023 -1478
rect 4324 -2050 5023 -2022
rect 5043 -1478 5742 -1450
rect 5043 -2022 5658 -1478
rect 5722 -2022 5742 -1478
rect 5043 -2050 5742 -2022
rect 5762 -1478 6461 -1450
rect 5762 -2022 6377 -1478
rect 6441 -2022 6461 -1478
rect 5762 -2050 6461 -2022
rect 6481 -1478 7180 -1450
rect 6481 -2022 7096 -1478
rect 7160 -2022 7180 -1478
rect 6481 -2050 7180 -2022
rect -7180 -2178 -6481 -2150
rect -7180 -2722 -6565 -2178
rect -6501 -2722 -6481 -2178
rect -7180 -2750 -6481 -2722
rect -6461 -2178 -5762 -2150
rect -6461 -2722 -5846 -2178
rect -5782 -2722 -5762 -2178
rect -6461 -2750 -5762 -2722
rect -5742 -2178 -5043 -2150
rect -5742 -2722 -5127 -2178
rect -5063 -2722 -5043 -2178
rect -5742 -2750 -5043 -2722
rect -5023 -2178 -4324 -2150
rect -5023 -2722 -4408 -2178
rect -4344 -2722 -4324 -2178
rect -5023 -2750 -4324 -2722
rect -4304 -2178 -3605 -2150
rect -4304 -2722 -3689 -2178
rect -3625 -2722 -3605 -2178
rect -4304 -2750 -3605 -2722
rect -3585 -2178 -2886 -2150
rect -3585 -2722 -2970 -2178
rect -2906 -2722 -2886 -2178
rect -3585 -2750 -2886 -2722
rect -2866 -2178 -2167 -2150
rect -2866 -2722 -2251 -2178
rect -2187 -2722 -2167 -2178
rect -2866 -2750 -2167 -2722
rect -2147 -2178 -1448 -2150
rect -2147 -2722 -1532 -2178
rect -1468 -2722 -1448 -2178
rect -2147 -2750 -1448 -2722
rect -1428 -2178 -729 -2150
rect -1428 -2722 -813 -2178
rect -749 -2722 -729 -2178
rect -1428 -2750 -729 -2722
rect -709 -2178 -10 -2150
rect -709 -2722 -94 -2178
rect -30 -2722 -10 -2178
rect -709 -2750 -10 -2722
rect 10 -2178 709 -2150
rect 10 -2722 625 -2178
rect 689 -2722 709 -2178
rect 10 -2750 709 -2722
rect 729 -2178 1428 -2150
rect 729 -2722 1344 -2178
rect 1408 -2722 1428 -2178
rect 729 -2750 1428 -2722
rect 1448 -2178 2147 -2150
rect 1448 -2722 2063 -2178
rect 2127 -2722 2147 -2178
rect 1448 -2750 2147 -2722
rect 2167 -2178 2866 -2150
rect 2167 -2722 2782 -2178
rect 2846 -2722 2866 -2178
rect 2167 -2750 2866 -2722
rect 2886 -2178 3585 -2150
rect 2886 -2722 3501 -2178
rect 3565 -2722 3585 -2178
rect 2886 -2750 3585 -2722
rect 3605 -2178 4304 -2150
rect 3605 -2722 4220 -2178
rect 4284 -2722 4304 -2178
rect 3605 -2750 4304 -2722
rect 4324 -2178 5023 -2150
rect 4324 -2722 4939 -2178
rect 5003 -2722 5023 -2178
rect 4324 -2750 5023 -2722
rect 5043 -2178 5742 -2150
rect 5043 -2722 5658 -2178
rect 5722 -2722 5742 -2178
rect 5043 -2750 5742 -2722
rect 5762 -2178 6461 -2150
rect 5762 -2722 6377 -2178
rect 6441 -2722 6461 -2178
rect 5762 -2750 6461 -2722
rect 6481 -2178 7180 -2150
rect 6481 -2722 7096 -2178
rect 7160 -2722 7180 -2178
rect 6481 -2750 7180 -2722
rect -7180 -2878 -6481 -2850
rect -7180 -3422 -6565 -2878
rect -6501 -3422 -6481 -2878
rect -7180 -3450 -6481 -3422
rect -6461 -2878 -5762 -2850
rect -6461 -3422 -5846 -2878
rect -5782 -3422 -5762 -2878
rect -6461 -3450 -5762 -3422
rect -5742 -2878 -5043 -2850
rect -5742 -3422 -5127 -2878
rect -5063 -3422 -5043 -2878
rect -5742 -3450 -5043 -3422
rect -5023 -2878 -4324 -2850
rect -5023 -3422 -4408 -2878
rect -4344 -3422 -4324 -2878
rect -5023 -3450 -4324 -3422
rect -4304 -2878 -3605 -2850
rect -4304 -3422 -3689 -2878
rect -3625 -3422 -3605 -2878
rect -4304 -3450 -3605 -3422
rect -3585 -2878 -2886 -2850
rect -3585 -3422 -2970 -2878
rect -2906 -3422 -2886 -2878
rect -3585 -3450 -2886 -3422
rect -2866 -2878 -2167 -2850
rect -2866 -3422 -2251 -2878
rect -2187 -3422 -2167 -2878
rect -2866 -3450 -2167 -3422
rect -2147 -2878 -1448 -2850
rect -2147 -3422 -1532 -2878
rect -1468 -3422 -1448 -2878
rect -2147 -3450 -1448 -3422
rect -1428 -2878 -729 -2850
rect -1428 -3422 -813 -2878
rect -749 -3422 -729 -2878
rect -1428 -3450 -729 -3422
rect -709 -2878 -10 -2850
rect -709 -3422 -94 -2878
rect -30 -3422 -10 -2878
rect -709 -3450 -10 -3422
rect 10 -2878 709 -2850
rect 10 -3422 625 -2878
rect 689 -3422 709 -2878
rect 10 -3450 709 -3422
rect 729 -2878 1428 -2850
rect 729 -3422 1344 -2878
rect 1408 -3422 1428 -2878
rect 729 -3450 1428 -3422
rect 1448 -2878 2147 -2850
rect 1448 -3422 2063 -2878
rect 2127 -3422 2147 -2878
rect 1448 -3450 2147 -3422
rect 2167 -2878 2866 -2850
rect 2167 -3422 2782 -2878
rect 2846 -3422 2866 -2878
rect 2167 -3450 2866 -3422
rect 2886 -2878 3585 -2850
rect 2886 -3422 3501 -2878
rect 3565 -3422 3585 -2878
rect 2886 -3450 3585 -3422
rect 3605 -2878 4304 -2850
rect 3605 -3422 4220 -2878
rect 4284 -3422 4304 -2878
rect 3605 -3450 4304 -3422
rect 4324 -2878 5023 -2850
rect 4324 -3422 4939 -2878
rect 5003 -3422 5023 -2878
rect 4324 -3450 5023 -3422
rect 5043 -2878 5742 -2850
rect 5043 -3422 5658 -2878
rect 5722 -3422 5742 -2878
rect 5043 -3450 5742 -3422
rect 5762 -2878 6461 -2850
rect 5762 -3422 6377 -2878
rect 6441 -3422 6461 -2878
rect 5762 -3450 6461 -3422
rect 6481 -2878 7180 -2850
rect 6481 -3422 7096 -2878
rect 7160 -3422 7180 -2878
rect 6481 -3450 7180 -3422
rect -7180 -3578 -6481 -3550
rect -7180 -4122 -6565 -3578
rect -6501 -4122 -6481 -3578
rect -7180 -4150 -6481 -4122
rect -6461 -3578 -5762 -3550
rect -6461 -4122 -5846 -3578
rect -5782 -4122 -5762 -3578
rect -6461 -4150 -5762 -4122
rect -5742 -3578 -5043 -3550
rect -5742 -4122 -5127 -3578
rect -5063 -4122 -5043 -3578
rect -5742 -4150 -5043 -4122
rect -5023 -3578 -4324 -3550
rect -5023 -4122 -4408 -3578
rect -4344 -4122 -4324 -3578
rect -5023 -4150 -4324 -4122
rect -4304 -3578 -3605 -3550
rect -4304 -4122 -3689 -3578
rect -3625 -4122 -3605 -3578
rect -4304 -4150 -3605 -4122
rect -3585 -3578 -2886 -3550
rect -3585 -4122 -2970 -3578
rect -2906 -4122 -2886 -3578
rect -3585 -4150 -2886 -4122
rect -2866 -3578 -2167 -3550
rect -2866 -4122 -2251 -3578
rect -2187 -4122 -2167 -3578
rect -2866 -4150 -2167 -4122
rect -2147 -3578 -1448 -3550
rect -2147 -4122 -1532 -3578
rect -1468 -4122 -1448 -3578
rect -2147 -4150 -1448 -4122
rect -1428 -3578 -729 -3550
rect -1428 -4122 -813 -3578
rect -749 -4122 -729 -3578
rect -1428 -4150 -729 -4122
rect -709 -3578 -10 -3550
rect -709 -4122 -94 -3578
rect -30 -4122 -10 -3578
rect -709 -4150 -10 -4122
rect 10 -3578 709 -3550
rect 10 -4122 625 -3578
rect 689 -4122 709 -3578
rect 10 -4150 709 -4122
rect 729 -3578 1428 -3550
rect 729 -4122 1344 -3578
rect 1408 -4122 1428 -3578
rect 729 -4150 1428 -4122
rect 1448 -3578 2147 -3550
rect 1448 -4122 2063 -3578
rect 2127 -4122 2147 -3578
rect 1448 -4150 2147 -4122
rect 2167 -3578 2866 -3550
rect 2167 -4122 2782 -3578
rect 2846 -4122 2866 -3578
rect 2167 -4150 2866 -4122
rect 2886 -3578 3585 -3550
rect 2886 -4122 3501 -3578
rect 3565 -4122 3585 -3578
rect 2886 -4150 3585 -4122
rect 3605 -3578 4304 -3550
rect 3605 -4122 4220 -3578
rect 4284 -4122 4304 -3578
rect 3605 -4150 4304 -4122
rect 4324 -3578 5023 -3550
rect 4324 -4122 4939 -3578
rect 5003 -4122 5023 -3578
rect 4324 -4150 5023 -4122
rect 5043 -3578 5742 -3550
rect 5043 -4122 5658 -3578
rect 5722 -4122 5742 -3578
rect 5043 -4150 5742 -4122
rect 5762 -3578 6461 -3550
rect 5762 -4122 6377 -3578
rect 6441 -4122 6461 -3578
rect 5762 -4150 6461 -4122
rect 6481 -3578 7180 -3550
rect 6481 -4122 7096 -3578
rect 7160 -4122 7180 -3578
rect 6481 -4150 7180 -4122
rect -7180 -4278 -6481 -4250
rect -7180 -4822 -6565 -4278
rect -6501 -4822 -6481 -4278
rect -7180 -4850 -6481 -4822
rect -6461 -4278 -5762 -4250
rect -6461 -4822 -5846 -4278
rect -5782 -4822 -5762 -4278
rect -6461 -4850 -5762 -4822
rect -5742 -4278 -5043 -4250
rect -5742 -4822 -5127 -4278
rect -5063 -4822 -5043 -4278
rect -5742 -4850 -5043 -4822
rect -5023 -4278 -4324 -4250
rect -5023 -4822 -4408 -4278
rect -4344 -4822 -4324 -4278
rect -5023 -4850 -4324 -4822
rect -4304 -4278 -3605 -4250
rect -4304 -4822 -3689 -4278
rect -3625 -4822 -3605 -4278
rect -4304 -4850 -3605 -4822
rect -3585 -4278 -2886 -4250
rect -3585 -4822 -2970 -4278
rect -2906 -4822 -2886 -4278
rect -3585 -4850 -2886 -4822
rect -2866 -4278 -2167 -4250
rect -2866 -4822 -2251 -4278
rect -2187 -4822 -2167 -4278
rect -2866 -4850 -2167 -4822
rect -2147 -4278 -1448 -4250
rect -2147 -4822 -1532 -4278
rect -1468 -4822 -1448 -4278
rect -2147 -4850 -1448 -4822
rect -1428 -4278 -729 -4250
rect -1428 -4822 -813 -4278
rect -749 -4822 -729 -4278
rect -1428 -4850 -729 -4822
rect -709 -4278 -10 -4250
rect -709 -4822 -94 -4278
rect -30 -4822 -10 -4278
rect -709 -4850 -10 -4822
rect 10 -4278 709 -4250
rect 10 -4822 625 -4278
rect 689 -4822 709 -4278
rect 10 -4850 709 -4822
rect 729 -4278 1428 -4250
rect 729 -4822 1344 -4278
rect 1408 -4822 1428 -4278
rect 729 -4850 1428 -4822
rect 1448 -4278 2147 -4250
rect 1448 -4822 2063 -4278
rect 2127 -4822 2147 -4278
rect 1448 -4850 2147 -4822
rect 2167 -4278 2866 -4250
rect 2167 -4822 2782 -4278
rect 2846 -4822 2866 -4278
rect 2167 -4850 2866 -4822
rect 2886 -4278 3585 -4250
rect 2886 -4822 3501 -4278
rect 3565 -4822 3585 -4278
rect 2886 -4850 3585 -4822
rect 3605 -4278 4304 -4250
rect 3605 -4822 4220 -4278
rect 4284 -4822 4304 -4278
rect 3605 -4850 4304 -4822
rect 4324 -4278 5023 -4250
rect 4324 -4822 4939 -4278
rect 5003 -4822 5023 -4278
rect 4324 -4850 5023 -4822
rect 5043 -4278 5742 -4250
rect 5043 -4822 5658 -4278
rect 5722 -4822 5742 -4278
rect 5043 -4850 5742 -4822
rect 5762 -4278 6461 -4250
rect 5762 -4822 6377 -4278
rect 6441 -4822 6461 -4278
rect 5762 -4850 6461 -4822
rect 6481 -4278 7180 -4250
rect 6481 -4822 7096 -4278
rect 7160 -4822 7180 -4278
rect 6481 -4850 7180 -4822
rect -7180 -4978 -6481 -4950
rect -7180 -5522 -6565 -4978
rect -6501 -5522 -6481 -4978
rect -7180 -5550 -6481 -5522
rect -6461 -4978 -5762 -4950
rect -6461 -5522 -5846 -4978
rect -5782 -5522 -5762 -4978
rect -6461 -5550 -5762 -5522
rect -5742 -4978 -5043 -4950
rect -5742 -5522 -5127 -4978
rect -5063 -5522 -5043 -4978
rect -5742 -5550 -5043 -5522
rect -5023 -4978 -4324 -4950
rect -5023 -5522 -4408 -4978
rect -4344 -5522 -4324 -4978
rect -5023 -5550 -4324 -5522
rect -4304 -4978 -3605 -4950
rect -4304 -5522 -3689 -4978
rect -3625 -5522 -3605 -4978
rect -4304 -5550 -3605 -5522
rect -3585 -4978 -2886 -4950
rect -3585 -5522 -2970 -4978
rect -2906 -5522 -2886 -4978
rect -3585 -5550 -2886 -5522
rect -2866 -4978 -2167 -4950
rect -2866 -5522 -2251 -4978
rect -2187 -5522 -2167 -4978
rect -2866 -5550 -2167 -5522
rect -2147 -4978 -1448 -4950
rect -2147 -5522 -1532 -4978
rect -1468 -5522 -1448 -4978
rect -2147 -5550 -1448 -5522
rect -1428 -4978 -729 -4950
rect -1428 -5522 -813 -4978
rect -749 -5522 -729 -4978
rect -1428 -5550 -729 -5522
rect -709 -4978 -10 -4950
rect -709 -5522 -94 -4978
rect -30 -5522 -10 -4978
rect -709 -5550 -10 -5522
rect 10 -4978 709 -4950
rect 10 -5522 625 -4978
rect 689 -5522 709 -4978
rect 10 -5550 709 -5522
rect 729 -4978 1428 -4950
rect 729 -5522 1344 -4978
rect 1408 -5522 1428 -4978
rect 729 -5550 1428 -5522
rect 1448 -4978 2147 -4950
rect 1448 -5522 2063 -4978
rect 2127 -5522 2147 -4978
rect 1448 -5550 2147 -5522
rect 2167 -4978 2866 -4950
rect 2167 -5522 2782 -4978
rect 2846 -5522 2866 -4978
rect 2167 -5550 2866 -5522
rect 2886 -4978 3585 -4950
rect 2886 -5522 3501 -4978
rect 3565 -5522 3585 -4978
rect 2886 -5550 3585 -5522
rect 3605 -4978 4304 -4950
rect 3605 -5522 4220 -4978
rect 4284 -5522 4304 -4978
rect 3605 -5550 4304 -5522
rect 4324 -4978 5023 -4950
rect 4324 -5522 4939 -4978
rect 5003 -5522 5023 -4978
rect 4324 -5550 5023 -5522
rect 5043 -4978 5742 -4950
rect 5043 -5522 5658 -4978
rect 5722 -5522 5742 -4978
rect 5043 -5550 5742 -5522
rect 5762 -4978 6461 -4950
rect 5762 -5522 6377 -4978
rect 6441 -5522 6461 -4978
rect 5762 -5550 6461 -5522
rect 6481 -4978 7180 -4950
rect 6481 -5522 7096 -4978
rect 7160 -5522 7180 -4978
rect 6481 -5550 7180 -5522
rect -7180 -5678 -6481 -5650
rect -7180 -6222 -6565 -5678
rect -6501 -6222 -6481 -5678
rect -7180 -6250 -6481 -6222
rect -6461 -5678 -5762 -5650
rect -6461 -6222 -5846 -5678
rect -5782 -6222 -5762 -5678
rect -6461 -6250 -5762 -6222
rect -5742 -5678 -5043 -5650
rect -5742 -6222 -5127 -5678
rect -5063 -6222 -5043 -5678
rect -5742 -6250 -5043 -6222
rect -5023 -5678 -4324 -5650
rect -5023 -6222 -4408 -5678
rect -4344 -6222 -4324 -5678
rect -5023 -6250 -4324 -6222
rect -4304 -5678 -3605 -5650
rect -4304 -6222 -3689 -5678
rect -3625 -6222 -3605 -5678
rect -4304 -6250 -3605 -6222
rect -3585 -5678 -2886 -5650
rect -3585 -6222 -2970 -5678
rect -2906 -6222 -2886 -5678
rect -3585 -6250 -2886 -6222
rect -2866 -5678 -2167 -5650
rect -2866 -6222 -2251 -5678
rect -2187 -6222 -2167 -5678
rect -2866 -6250 -2167 -6222
rect -2147 -5678 -1448 -5650
rect -2147 -6222 -1532 -5678
rect -1468 -6222 -1448 -5678
rect -2147 -6250 -1448 -6222
rect -1428 -5678 -729 -5650
rect -1428 -6222 -813 -5678
rect -749 -6222 -729 -5678
rect -1428 -6250 -729 -6222
rect -709 -5678 -10 -5650
rect -709 -6222 -94 -5678
rect -30 -6222 -10 -5678
rect -709 -6250 -10 -6222
rect 10 -5678 709 -5650
rect 10 -6222 625 -5678
rect 689 -6222 709 -5678
rect 10 -6250 709 -6222
rect 729 -5678 1428 -5650
rect 729 -6222 1344 -5678
rect 1408 -6222 1428 -5678
rect 729 -6250 1428 -6222
rect 1448 -5678 2147 -5650
rect 1448 -6222 2063 -5678
rect 2127 -6222 2147 -5678
rect 1448 -6250 2147 -6222
rect 2167 -5678 2866 -5650
rect 2167 -6222 2782 -5678
rect 2846 -6222 2866 -5678
rect 2167 -6250 2866 -6222
rect 2886 -5678 3585 -5650
rect 2886 -6222 3501 -5678
rect 3565 -6222 3585 -5678
rect 2886 -6250 3585 -6222
rect 3605 -5678 4304 -5650
rect 3605 -6222 4220 -5678
rect 4284 -6222 4304 -5678
rect 3605 -6250 4304 -6222
rect 4324 -5678 5023 -5650
rect 4324 -6222 4939 -5678
rect 5003 -6222 5023 -5678
rect 4324 -6250 5023 -6222
rect 5043 -5678 5742 -5650
rect 5043 -6222 5658 -5678
rect 5722 -6222 5742 -5678
rect 5043 -6250 5742 -6222
rect 5762 -5678 6461 -5650
rect 5762 -6222 6377 -5678
rect 6441 -6222 6461 -5678
rect 5762 -6250 6461 -6222
rect 6481 -5678 7180 -5650
rect 6481 -6222 7096 -5678
rect 7160 -6222 7180 -5678
rect 6481 -6250 7180 -6222
rect -7180 -6378 -6481 -6350
rect -7180 -6922 -6565 -6378
rect -6501 -6922 -6481 -6378
rect -7180 -6950 -6481 -6922
rect -6461 -6378 -5762 -6350
rect -6461 -6922 -5846 -6378
rect -5782 -6922 -5762 -6378
rect -6461 -6950 -5762 -6922
rect -5742 -6378 -5043 -6350
rect -5742 -6922 -5127 -6378
rect -5063 -6922 -5043 -6378
rect -5742 -6950 -5043 -6922
rect -5023 -6378 -4324 -6350
rect -5023 -6922 -4408 -6378
rect -4344 -6922 -4324 -6378
rect -5023 -6950 -4324 -6922
rect -4304 -6378 -3605 -6350
rect -4304 -6922 -3689 -6378
rect -3625 -6922 -3605 -6378
rect -4304 -6950 -3605 -6922
rect -3585 -6378 -2886 -6350
rect -3585 -6922 -2970 -6378
rect -2906 -6922 -2886 -6378
rect -3585 -6950 -2886 -6922
rect -2866 -6378 -2167 -6350
rect -2866 -6922 -2251 -6378
rect -2187 -6922 -2167 -6378
rect -2866 -6950 -2167 -6922
rect -2147 -6378 -1448 -6350
rect -2147 -6922 -1532 -6378
rect -1468 -6922 -1448 -6378
rect -2147 -6950 -1448 -6922
rect -1428 -6378 -729 -6350
rect -1428 -6922 -813 -6378
rect -749 -6922 -729 -6378
rect -1428 -6950 -729 -6922
rect -709 -6378 -10 -6350
rect -709 -6922 -94 -6378
rect -30 -6922 -10 -6378
rect -709 -6950 -10 -6922
rect 10 -6378 709 -6350
rect 10 -6922 625 -6378
rect 689 -6922 709 -6378
rect 10 -6950 709 -6922
rect 729 -6378 1428 -6350
rect 729 -6922 1344 -6378
rect 1408 -6922 1428 -6378
rect 729 -6950 1428 -6922
rect 1448 -6378 2147 -6350
rect 1448 -6922 2063 -6378
rect 2127 -6922 2147 -6378
rect 1448 -6950 2147 -6922
rect 2167 -6378 2866 -6350
rect 2167 -6922 2782 -6378
rect 2846 -6922 2866 -6378
rect 2167 -6950 2866 -6922
rect 2886 -6378 3585 -6350
rect 2886 -6922 3501 -6378
rect 3565 -6922 3585 -6378
rect 2886 -6950 3585 -6922
rect 3605 -6378 4304 -6350
rect 3605 -6922 4220 -6378
rect 4284 -6922 4304 -6378
rect 3605 -6950 4304 -6922
rect 4324 -6378 5023 -6350
rect 4324 -6922 4939 -6378
rect 5003 -6922 5023 -6378
rect 4324 -6950 5023 -6922
rect 5043 -6378 5742 -6350
rect 5043 -6922 5658 -6378
rect 5722 -6922 5742 -6378
rect 5043 -6950 5742 -6922
rect 5762 -6378 6461 -6350
rect 5762 -6922 6377 -6378
rect 6441 -6922 6461 -6378
rect 5762 -6950 6461 -6922
rect 6481 -6378 7180 -6350
rect 6481 -6922 7096 -6378
rect 7160 -6922 7180 -6378
rect 6481 -6950 7180 -6922
<< via3 >>
rect -6565 6378 -6501 6922
rect -5846 6378 -5782 6922
rect -5127 6378 -5063 6922
rect -4408 6378 -4344 6922
rect -3689 6378 -3625 6922
rect -2970 6378 -2906 6922
rect -2251 6378 -2187 6922
rect -1532 6378 -1468 6922
rect -813 6378 -749 6922
rect -94 6378 -30 6922
rect 625 6378 689 6922
rect 1344 6378 1408 6922
rect 2063 6378 2127 6922
rect 2782 6378 2846 6922
rect 3501 6378 3565 6922
rect 4220 6378 4284 6922
rect 4939 6378 5003 6922
rect 5658 6378 5722 6922
rect 6377 6378 6441 6922
rect 7096 6378 7160 6922
rect -6565 5678 -6501 6222
rect -5846 5678 -5782 6222
rect -5127 5678 -5063 6222
rect -4408 5678 -4344 6222
rect -3689 5678 -3625 6222
rect -2970 5678 -2906 6222
rect -2251 5678 -2187 6222
rect -1532 5678 -1468 6222
rect -813 5678 -749 6222
rect -94 5678 -30 6222
rect 625 5678 689 6222
rect 1344 5678 1408 6222
rect 2063 5678 2127 6222
rect 2782 5678 2846 6222
rect 3501 5678 3565 6222
rect 4220 5678 4284 6222
rect 4939 5678 5003 6222
rect 5658 5678 5722 6222
rect 6377 5678 6441 6222
rect 7096 5678 7160 6222
rect -6565 4978 -6501 5522
rect -5846 4978 -5782 5522
rect -5127 4978 -5063 5522
rect -4408 4978 -4344 5522
rect -3689 4978 -3625 5522
rect -2970 4978 -2906 5522
rect -2251 4978 -2187 5522
rect -1532 4978 -1468 5522
rect -813 4978 -749 5522
rect -94 4978 -30 5522
rect 625 4978 689 5522
rect 1344 4978 1408 5522
rect 2063 4978 2127 5522
rect 2782 4978 2846 5522
rect 3501 4978 3565 5522
rect 4220 4978 4284 5522
rect 4939 4978 5003 5522
rect 5658 4978 5722 5522
rect 6377 4978 6441 5522
rect 7096 4978 7160 5522
rect -6565 4278 -6501 4822
rect -5846 4278 -5782 4822
rect -5127 4278 -5063 4822
rect -4408 4278 -4344 4822
rect -3689 4278 -3625 4822
rect -2970 4278 -2906 4822
rect -2251 4278 -2187 4822
rect -1532 4278 -1468 4822
rect -813 4278 -749 4822
rect -94 4278 -30 4822
rect 625 4278 689 4822
rect 1344 4278 1408 4822
rect 2063 4278 2127 4822
rect 2782 4278 2846 4822
rect 3501 4278 3565 4822
rect 4220 4278 4284 4822
rect 4939 4278 5003 4822
rect 5658 4278 5722 4822
rect 6377 4278 6441 4822
rect 7096 4278 7160 4822
rect -6565 3578 -6501 4122
rect -5846 3578 -5782 4122
rect -5127 3578 -5063 4122
rect -4408 3578 -4344 4122
rect -3689 3578 -3625 4122
rect -2970 3578 -2906 4122
rect -2251 3578 -2187 4122
rect -1532 3578 -1468 4122
rect -813 3578 -749 4122
rect -94 3578 -30 4122
rect 625 3578 689 4122
rect 1344 3578 1408 4122
rect 2063 3578 2127 4122
rect 2782 3578 2846 4122
rect 3501 3578 3565 4122
rect 4220 3578 4284 4122
rect 4939 3578 5003 4122
rect 5658 3578 5722 4122
rect 6377 3578 6441 4122
rect 7096 3578 7160 4122
rect -6565 2878 -6501 3422
rect -5846 2878 -5782 3422
rect -5127 2878 -5063 3422
rect -4408 2878 -4344 3422
rect -3689 2878 -3625 3422
rect -2970 2878 -2906 3422
rect -2251 2878 -2187 3422
rect -1532 2878 -1468 3422
rect -813 2878 -749 3422
rect -94 2878 -30 3422
rect 625 2878 689 3422
rect 1344 2878 1408 3422
rect 2063 2878 2127 3422
rect 2782 2878 2846 3422
rect 3501 2878 3565 3422
rect 4220 2878 4284 3422
rect 4939 2878 5003 3422
rect 5658 2878 5722 3422
rect 6377 2878 6441 3422
rect 7096 2878 7160 3422
rect -6565 2178 -6501 2722
rect -5846 2178 -5782 2722
rect -5127 2178 -5063 2722
rect -4408 2178 -4344 2722
rect -3689 2178 -3625 2722
rect -2970 2178 -2906 2722
rect -2251 2178 -2187 2722
rect -1532 2178 -1468 2722
rect -813 2178 -749 2722
rect -94 2178 -30 2722
rect 625 2178 689 2722
rect 1344 2178 1408 2722
rect 2063 2178 2127 2722
rect 2782 2178 2846 2722
rect 3501 2178 3565 2722
rect 4220 2178 4284 2722
rect 4939 2178 5003 2722
rect 5658 2178 5722 2722
rect 6377 2178 6441 2722
rect 7096 2178 7160 2722
rect -6565 1478 -6501 2022
rect -5846 1478 -5782 2022
rect -5127 1478 -5063 2022
rect -4408 1478 -4344 2022
rect -3689 1478 -3625 2022
rect -2970 1478 -2906 2022
rect -2251 1478 -2187 2022
rect -1532 1478 -1468 2022
rect -813 1478 -749 2022
rect -94 1478 -30 2022
rect 625 1478 689 2022
rect 1344 1478 1408 2022
rect 2063 1478 2127 2022
rect 2782 1478 2846 2022
rect 3501 1478 3565 2022
rect 4220 1478 4284 2022
rect 4939 1478 5003 2022
rect 5658 1478 5722 2022
rect 6377 1478 6441 2022
rect 7096 1478 7160 2022
rect -6565 778 -6501 1322
rect -5846 778 -5782 1322
rect -5127 778 -5063 1322
rect -4408 778 -4344 1322
rect -3689 778 -3625 1322
rect -2970 778 -2906 1322
rect -2251 778 -2187 1322
rect -1532 778 -1468 1322
rect -813 778 -749 1322
rect -94 778 -30 1322
rect 625 778 689 1322
rect 1344 778 1408 1322
rect 2063 778 2127 1322
rect 2782 778 2846 1322
rect 3501 778 3565 1322
rect 4220 778 4284 1322
rect 4939 778 5003 1322
rect 5658 778 5722 1322
rect 6377 778 6441 1322
rect 7096 778 7160 1322
rect -6565 78 -6501 622
rect -5846 78 -5782 622
rect -5127 78 -5063 622
rect -4408 78 -4344 622
rect -3689 78 -3625 622
rect -2970 78 -2906 622
rect -2251 78 -2187 622
rect -1532 78 -1468 622
rect -813 78 -749 622
rect -94 78 -30 622
rect 625 78 689 622
rect 1344 78 1408 622
rect 2063 78 2127 622
rect 2782 78 2846 622
rect 3501 78 3565 622
rect 4220 78 4284 622
rect 4939 78 5003 622
rect 5658 78 5722 622
rect 6377 78 6441 622
rect 7096 78 7160 622
rect -6565 -622 -6501 -78
rect -5846 -622 -5782 -78
rect -5127 -622 -5063 -78
rect -4408 -622 -4344 -78
rect -3689 -622 -3625 -78
rect -2970 -622 -2906 -78
rect -2251 -622 -2187 -78
rect -1532 -622 -1468 -78
rect -813 -622 -749 -78
rect -94 -622 -30 -78
rect 625 -622 689 -78
rect 1344 -622 1408 -78
rect 2063 -622 2127 -78
rect 2782 -622 2846 -78
rect 3501 -622 3565 -78
rect 4220 -622 4284 -78
rect 4939 -622 5003 -78
rect 5658 -622 5722 -78
rect 6377 -622 6441 -78
rect 7096 -622 7160 -78
rect -6565 -1322 -6501 -778
rect -5846 -1322 -5782 -778
rect -5127 -1322 -5063 -778
rect -4408 -1322 -4344 -778
rect -3689 -1322 -3625 -778
rect -2970 -1322 -2906 -778
rect -2251 -1322 -2187 -778
rect -1532 -1322 -1468 -778
rect -813 -1322 -749 -778
rect -94 -1322 -30 -778
rect 625 -1322 689 -778
rect 1344 -1322 1408 -778
rect 2063 -1322 2127 -778
rect 2782 -1322 2846 -778
rect 3501 -1322 3565 -778
rect 4220 -1322 4284 -778
rect 4939 -1322 5003 -778
rect 5658 -1322 5722 -778
rect 6377 -1322 6441 -778
rect 7096 -1322 7160 -778
rect -6565 -2022 -6501 -1478
rect -5846 -2022 -5782 -1478
rect -5127 -2022 -5063 -1478
rect -4408 -2022 -4344 -1478
rect -3689 -2022 -3625 -1478
rect -2970 -2022 -2906 -1478
rect -2251 -2022 -2187 -1478
rect -1532 -2022 -1468 -1478
rect -813 -2022 -749 -1478
rect -94 -2022 -30 -1478
rect 625 -2022 689 -1478
rect 1344 -2022 1408 -1478
rect 2063 -2022 2127 -1478
rect 2782 -2022 2846 -1478
rect 3501 -2022 3565 -1478
rect 4220 -2022 4284 -1478
rect 4939 -2022 5003 -1478
rect 5658 -2022 5722 -1478
rect 6377 -2022 6441 -1478
rect 7096 -2022 7160 -1478
rect -6565 -2722 -6501 -2178
rect -5846 -2722 -5782 -2178
rect -5127 -2722 -5063 -2178
rect -4408 -2722 -4344 -2178
rect -3689 -2722 -3625 -2178
rect -2970 -2722 -2906 -2178
rect -2251 -2722 -2187 -2178
rect -1532 -2722 -1468 -2178
rect -813 -2722 -749 -2178
rect -94 -2722 -30 -2178
rect 625 -2722 689 -2178
rect 1344 -2722 1408 -2178
rect 2063 -2722 2127 -2178
rect 2782 -2722 2846 -2178
rect 3501 -2722 3565 -2178
rect 4220 -2722 4284 -2178
rect 4939 -2722 5003 -2178
rect 5658 -2722 5722 -2178
rect 6377 -2722 6441 -2178
rect 7096 -2722 7160 -2178
rect -6565 -3422 -6501 -2878
rect -5846 -3422 -5782 -2878
rect -5127 -3422 -5063 -2878
rect -4408 -3422 -4344 -2878
rect -3689 -3422 -3625 -2878
rect -2970 -3422 -2906 -2878
rect -2251 -3422 -2187 -2878
rect -1532 -3422 -1468 -2878
rect -813 -3422 -749 -2878
rect -94 -3422 -30 -2878
rect 625 -3422 689 -2878
rect 1344 -3422 1408 -2878
rect 2063 -3422 2127 -2878
rect 2782 -3422 2846 -2878
rect 3501 -3422 3565 -2878
rect 4220 -3422 4284 -2878
rect 4939 -3422 5003 -2878
rect 5658 -3422 5722 -2878
rect 6377 -3422 6441 -2878
rect 7096 -3422 7160 -2878
rect -6565 -4122 -6501 -3578
rect -5846 -4122 -5782 -3578
rect -5127 -4122 -5063 -3578
rect -4408 -4122 -4344 -3578
rect -3689 -4122 -3625 -3578
rect -2970 -4122 -2906 -3578
rect -2251 -4122 -2187 -3578
rect -1532 -4122 -1468 -3578
rect -813 -4122 -749 -3578
rect -94 -4122 -30 -3578
rect 625 -4122 689 -3578
rect 1344 -4122 1408 -3578
rect 2063 -4122 2127 -3578
rect 2782 -4122 2846 -3578
rect 3501 -4122 3565 -3578
rect 4220 -4122 4284 -3578
rect 4939 -4122 5003 -3578
rect 5658 -4122 5722 -3578
rect 6377 -4122 6441 -3578
rect 7096 -4122 7160 -3578
rect -6565 -4822 -6501 -4278
rect -5846 -4822 -5782 -4278
rect -5127 -4822 -5063 -4278
rect -4408 -4822 -4344 -4278
rect -3689 -4822 -3625 -4278
rect -2970 -4822 -2906 -4278
rect -2251 -4822 -2187 -4278
rect -1532 -4822 -1468 -4278
rect -813 -4822 -749 -4278
rect -94 -4822 -30 -4278
rect 625 -4822 689 -4278
rect 1344 -4822 1408 -4278
rect 2063 -4822 2127 -4278
rect 2782 -4822 2846 -4278
rect 3501 -4822 3565 -4278
rect 4220 -4822 4284 -4278
rect 4939 -4822 5003 -4278
rect 5658 -4822 5722 -4278
rect 6377 -4822 6441 -4278
rect 7096 -4822 7160 -4278
rect -6565 -5522 -6501 -4978
rect -5846 -5522 -5782 -4978
rect -5127 -5522 -5063 -4978
rect -4408 -5522 -4344 -4978
rect -3689 -5522 -3625 -4978
rect -2970 -5522 -2906 -4978
rect -2251 -5522 -2187 -4978
rect -1532 -5522 -1468 -4978
rect -813 -5522 -749 -4978
rect -94 -5522 -30 -4978
rect 625 -5522 689 -4978
rect 1344 -5522 1408 -4978
rect 2063 -5522 2127 -4978
rect 2782 -5522 2846 -4978
rect 3501 -5522 3565 -4978
rect 4220 -5522 4284 -4978
rect 4939 -5522 5003 -4978
rect 5658 -5522 5722 -4978
rect 6377 -5522 6441 -4978
rect 7096 -5522 7160 -4978
rect -6565 -6222 -6501 -5678
rect -5846 -6222 -5782 -5678
rect -5127 -6222 -5063 -5678
rect -4408 -6222 -4344 -5678
rect -3689 -6222 -3625 -5678
rect -2970 -6222 -2906 -5678
rect -2251 -6222 -2187 -5678
rect -1532 -6222 -1468 -5678
rect -813 -6222 -749 -5678
rect -94 -6222 -30 -5678
rect 625 -6222 689 -5678
rect 1344 -6222 1408 -5678
rect 2063 -6222 2127 -5678
rect 2782 -6222 2846 -5678
rect 3501 -6222 3565 -5678
rect 4220 -6222 4284 -5678
rect 4939 -6222 5003 -5678
rect 5658 -6222 5722 -5678
rect 6377 -6222 6441 -5678
rect 7096 -6222 7160 -5678
rect -6565 -6922 -6501 -6378
rect -5846 -6922 -5782 -6378
rect -5127 -6922 -5063 -6378
rect -4408 -6922 -4344 -6378
rect -3689 -6922 -3625 -6378
rect -2970 -6922 -2906 -6378
rect -2251 -6922 -2187 -6378
rect -1532 -6922 -1468 -6378
rect -813 -6922 -749 -6378
rect -94 -6922 -30 -6378
rect 625 -6922 689 -6378
rect 1344 -6922 1408 -6378
rect 2063 -6922 2127 -6378
rect 2782 -6922 2846 -6378
rect 3501 -6922 3565 -6378
rect 4220 -6922 4284 -6378
rect 4939 -6922 5003 -6378
rect 5658 -6922 5722 -6378
rect 6377 -6922 6441 -6378
rect 7096 -6922 7160 -6378
<< mimcap >>
rect -7080 6810 -6680 6850
rect -7080 6490 -7040 6810
rect -6720 6490 -6680 6810
rect -7080 6450 -6680 6490
rect -6361 6810 -5961 6850
rect -6361 6490 -6321 6810
rect -6001 6490 -5961 6810
rect -6361 6450 -5961 6490
rect -5642 6810 -5242 6850
rect -5642 6490 -5602 6810
rect -5282 6490 -5242 6810
rect -5642 6450 -5242 6490
rect -4923 6810 -4523 6850
rect -4923 6490 -4883 6810
rect -4563 6490 -4523 6810
rect -4923 6450 -4523 6490
rect -4204 6810 -3804 6850
rect -4204 6490 -4164 6810
rect -3844 6490 -3804 6810
rect -4204 6450 -3804 6490
rect -3485 6810 -3085 6850
rect -3485 6490 -3445 6810
rect -3125 6490 -3085 6810
rect -3485 6450 -3085 6490
rect -2766 6810 -2366 6850
rect -2766 6490 -2726 6810
rect -2406 6490 -2366 6810
rect -2766 6450 -2366 6490
rect -2047 6810 -1647 6850
rect -2047 6490 -2007 6810
rect -1687 6490 -1647 6810
rect -2047 6450 -1647 6490
rect -1328 6810 -928 6850
rect -1328 6490 -1288 6810
rect -968 6490 -928 6810
rect -1328 6450 -928 6490
rect -609 6810 -209 6850
rect -609 6490 -569 6810
rect -249 6490 -209 6810
rect -609 6450 -209 6490
rect 110 6810 510 6850
rect 110 6490 150 6810
rect 470 6490 510 6810
rect 110 6450 510 6490
rect 829 6810 1229 6850
rect 829 6490 869 6810
rect 1189 6490 1229 6810
rect 829 6450 1229 6490
rect 1548 6810 1948 6850
rect 1548 6490 1588 6810
rect 1908 6490 1948 6810
rect 1548 6450 1948 6490
rect 2267 6810 2667 6850
rect 2267 6490 2307 6810
rect 2627 6490 2667 6810
rect 2267 6450 2667 6490
rect 2986 6810 3386 6850
rect 2986 6490 3026 6810
rect 3346 6490 3386 6810
rect 2986 6450 3386 6490
rect 3705 6810 4105 6850
rect 3705 6490 3745 6810
rect 4065 6490 4105 6810
rect 3705 6450 4105 6490
rect 4424 6810 4824 6850
rect 4424 6490 4464 6810
rect 4784 6490 4824 6810
rect 4424 6450 4824 6490
rect 5143 6810 5543 6850
rect 5143 6490 5183 6810
rect 5503 6490 5543 6810
rect 5143 6450 5543 6490
rect 5862 6810 6262 6850
rect 5862 6490 5902 6810
rect 6222 6490 6262 6810
rect 5862 6450 6262 6490
rect 6581 6810 6981 6850
rect 6581 6490 6621 6810
rect 6941 6490 6981 6810
rect 6581 6450 6981 6490
rect -7080 6110 -6680 6150
rect -7080 5790 -7040 6110
rect -6720 5790 -6680 6110
rect -7080 5750 -6680 5790
rect -6361 6110 -5961 6150
rect -6361 5790 -6321 6110
rect -6001 5790 -5961 6110
rect -6361 5750 -5961 5790
rect -5642 6110 -5242 6150
rect -5642 5790 -5602 6110
rect -5282 5790 -5242 6110
rect -5642 5750 -5242 5790
rect -4923 6110 -4523 6150
rect -4923 5790 -4883 6110
rect -4563 5790 -4523 6110
rect -4923 5750 -4523 5790
rect -4204 6110 -3804 6150
rect -4204 5790 -4164 6110
rect -3844 5790 -3804 6110
rect -4204 5750 -3804 5790
rect -3485 6110 -3085 6150
rect -3485 5790 -3445 6110
rect -3125 5790 -3085 6110
rect -3485 5750 -3085 5790
rect -2766 6110 -2366 6150
rect -2766 5790 -2726 6110
rect -2406 5790 -2366 6110
rect -2766 5750 -2366 5790
rect -2047 6110 -1647 6150
rect -2047 5790 -2007 6110
rect -1687 5790 -1647 6110
rect -2047 5750 -1647 5790
rect -1328 6110 -928 6150
rect -1328 5790 -1288 6110
rect -968 5790 -928 6110
rect -1328 5750 -928 5790
rect -609 6110 -209 6150
rect -609 5790 -569 6110
rect -249 5790 -209 6110
rect -609 5750 -209 5790
rect 110 6110 510 6150
rect 110 5790 150 6110
rect 470 5790 510 6110
rect 110 5750 510 5790
rect 829 6110 1229 6150
rect 829 5790 869 6110
rect 1189 5790 1229 6110
rect 829 5750 1229 5790
rect 1548 6110 1948 6150
rect 1548 5790 1588 6110
rect 1908 5790 1948 6110
rect 1548 5750 1948 5790
rect 2267 6110 2667 6150
rect 2267 5790 2307 6110
rect 2627 5790 2667 6110
rect 2267 5750 2667 5790
rect 2986 6110 3386 6150
rect 2986 5790 3026 6110
rect 3346 5790 3386 6110
rect 2986 5750 3386 5790
rect 3705 6110 4105 6150
rect 3705 5790 3745 6110
rect 4065 5790 4105 6110
rect 3705 5750 4105 5790
rect 4424 6110 4824 6150
rect 4424 5790 4464 6110
rect 4784 5790 4824 6110
rect 4424 5750 4824 5790
rect 5143 6110 5543 6150
rect 5143 5790 5183 6110
rect 5503 5790 5543 6110
rect 5143 5750 5543 5790
rect 5862 6110 6262 6150
rect 5862 5790 5902 6110
rect 6222 5790 6262 6110
rect 5862 5750 6262 5790
rect 6581 6110 6981 6150
rect 6581 5790 6621 6110
rect 6941 5790 6981 6110
rect 6581 5750 6981 5790
rect -7080 5410 -6680 5450
rect -7080 5090 -7040 5410
rect -6720 5090 -6680 5410
rect -7080 5050 -6680 5090
rect -6361 5410 -5961 5450
rect -6361 5090 -6321 5410
rect -6001 5090 -5961 5410
rect -6361 5050 -5961 5090
rect -5642 5410 -5242 5450
rect -5642 5090 -5602 5410
rect -5282 5090 -5242 5410
rect -5642 5050 -5242 5090
rect -4923 5410 -4523 5450
rect -4923 5090 -4883 5410
rect -4563 5090 -4523 5410
rect -4923 5050 -4523 5090
rect -4204 5410 -3804 5450
rect -4204 5090 -4164 5410
rect -3844 5090 -3804 5410
rect -4204 5050 -3804 5090
rect -3485 5410 -3085 5450
rect -3485 5090 -3445 5410
rect -3125 5090 -3085 5410
rect -3485 5050 -3085 5090
rect -2766 5410 -2366 5450
rect -2766 5090 -2726 5410
rect -2406 5090 -2366 5410
rect -2766 5050 -2366 5090
rect -2047 5410 -1647 5450
rect -2047 5090 -2007 5410
rect -1687 5090 -1647 5410
rect -2047 5050 -1647 5090
rect -1328 5410 -928 5450
rect -1328 5090 -1288 5410
rect -968 5090 -928 5410
rect -1328 5050 -928 5090
rect -609 5410 -209 5450
rect -609 5090 -569 5410
rect -249 5090 -209 5410
rect -609 5050 -209 5090
rect 110 5410 510 5450
rect 110 5090 150 5410
rect 470 5090 510 5410
rect 110 5050 510 5090
rect 829 5410 1229 5450
rect 829 5090 869 5410
rect 1189 5090 1229 5410
rect 829 5050 1229 5090
rect 1548 5410 1948 5450
rect 1548 5090 1588 5410
rect 1908 5090 1948 5410
rect 1548 5050 1948 5090
rect 2267 5410 2667 5450
rect 2267 5090 2307 5410
rect 2627 5090 2667 5410
rect 2267 5050 2667 5090
rect 2986 5410 3386 5450
rect 2986 5090 3026 5410
rect 3346 5090 3386 5410
rect 2986 5050 3386 5090
rect 3705 5410 4105 5450
rect 3705 5090 3745 5410
rect 4065 5090 4105 5410
rect 3705 5050 4105 5090
rect 4424 5410 4824 5450
rect 4424 5090 4464 5410
rect 4784 5090 4824 5410
rect 4424 5050 4824 5090
rect 5143 5410 5543 5450
rect 5143 5090 5183 5410
rect 5503 5090 5543 5410
rect 5143 5050 5543 5090
rect 5862 5410 6262 5450
rect 5862 5090 5902 5410
rect 6222 5090 6262 5410
rect 5862 5050 6262 5090
rect 6581 5410 6981 5450
rect 6581 5090 6621 5410
rect 6941 5090 6981 5410
rect 6581 5050 6981 5090
rect -7080 4710 -6680 4750
rect -7080 4390 -7040 4710
rect -6720 4390 -6680 4710
rect -7080 4350 -6680 4390
rect -6361 4710 -5961 4750
rect -6361 4390 -6321 4710
rect -6001 4390 -5961 4710
rect -6361 4350 -5961 4390
rect -5642 4710 -5242 4750
rect -5642 4390 -5602 4710
rect -5282 4390 -5242 4710
rect -5642 4350 -5242 4390
rect -4923 4710 -4523 4750
rect -4923 4390 -4883 4710
rect -4563 4390 -4523 4710
rect -4923 4350 -4523 4390
rect -4204 4710 -3804 4750
rect -4204 4390 -4164 4710
rect -3844 4390 -3804 4710
rect -4204 4350 -3804 4390
rect -3485 4710 -3085 4750
rect -3485 4390 -3445 4710
rect -3125 4390 -3085 4710
rect -3485 4350 -3085 4390
rect -2766 4710 -2366 4750
rect -2766 4390 -2726 4710
rect -2406 4390 -2366 4710
rect -2766 4350 -2366 4390
rect -2047 4710 -1647 4750
rect -2047 4390 -2007 4710
rect -1687 4390 -1647 4710
rect -2047 4350 -1647 4390
rect -1328 4710 -928 4750
rect -1328 4390 -1288 4710
rect -968 4390 -928 4710
rect -1328 4350 -928 4390
rect -609 4710 -209 4750
rect -609 4390 -569 4710
rect -249 4390 -209 4710
rect -609 4350 -209 4390
rect 110 4710 510 4750
rect 110 4390 150 4710
rect 470 4390 510 4710
rect 110 4350 510 4390
rect 829 4710 1229 4750
rect 829 4390 869 4710
rect 1189 4390 1229 4710
rect 829 4350 1229 4390
rect 1548 4710 1948 4750
rect 1548 4390 1588 4710
rect 1908 4390 1948 4710
rect 1548 4350 1948 4390
rect 2267 4710 2667 4750
rect 2267 4390 2307 4710
rect 2627 4390 2667 4710
rect 2267 4350 2667 4390
rect 2986 4710 3386 4750
rect 2986 4390 3026 4710
rect 3346 4390 3386 4710
rect 2986 4350 3386 4390
rect 3705 4710 4105 4750
rect 3705 4390 3745 4710
rect 4065 4390 4105 4710
rect 3705 4350 4105 4390
rect 4424 4710 4824 4750
rect 4424 4390 4464 4710
rect 4784 4390 4824 4710
rect 4424 4350 4824 4390
rect 5143 4710 5543 4750
rect 5143 4390 5183 4710
rect 5503 4390 5543 4710
rect 5143 4350 5543 4390
rect 5862 4710 6262 4750
rect 5862 4390 5902 4710
rect 6222 4390 6262 4710
rect 5862 4350 6262 4390
rect 6581 4710 6981 4750
rect 6581 4390 6621 4710
rect 6941 4390 6981 4710
rect 6581 4350 6981 4390
rect -7080 4010 -6680 4050
rect -7080 3690 -7040 4010
rect -6720 3690 -6680 4010
rect -7080 3650 -6680 3690
rect -6361 4010 -5961 4050
rect -6361 3690 -6321 4010
rect -6001 3690 -5961 4010
rect -6361 3650 -5961 3690
rect -5642 4010 -5242 4050
rect -5642 3690 -5602 4010
rect -5282 3690 -5242 4010
rect -5642 3650 -5242 3690
rect -4923 4010 -4523 4050
rect -4923 3690 -4883 4010
rect -4563 3690 -4523 4010
rect -4923 3650 -4523 3690
rect -4204 4010 -3804 4050
rect -4204 3690 -4164 4010
rect -3844 3690 -3804 4010
rect -4204 3650 -3804 3690
rect -3485 4010 -3085 4050
rect -3485 3690 -3445 4010
rect -3125 3690 -3085 4010
rect -3485 3650 -3085 3690
rect -2766 4010 -2366 4050
rect -2766 3690 -2726 4010
rect -2406 3690 -2366 4010
rect -2766 3650 -2366 3690
rect -2047 4010 -1647 4050
rect -2047 3690 -2007 4010
rect -1687 3690 -1647 4010
rect -2047 3650 -1647 3690
rect -1328 4010 -928 4050
rect -1328 3690 -1288 4010
rect -968 3690 -928 4010
rect -1328 3650 -928 3690
rect -609 4010 -209 4050
rect -609 3690 -569 4010
rect -249 3690 -209 4010
rect -609 3650 -209 3690
rect 110 4010 510 4050
rect 110 3690 150 4010
rect 470 3690 510 4010
rect 110 3650 510 3690
rect 829 4010 1229 4050
rect 829 3690 869 4010
rect 1189 3690 1229 4010
rect 829 3650 1229 3690
rect 1548 4010 1948 4050
rect 1548 3690 1588 4010
rect 1908 3690 1948 4010
rect 1548 3650 1948 3690
rect 2267 4010 2667 4050
rect 2267 3690 2307 4010
rect 2627 3690 2667 4010
rect 2267 3650 2667 3690
rect 2986 4010 3386 4050
rect 2986 3690 3026 4010
rect 3346 3690 3386 4010
rect 2986 3650 3386 3690
rect 3705 4010 4105 4050
rect 3705 3690 3745 4010
rect 4065 3690 4105 4010
rect 3705 3650 4105 3690
rect 4424 4010 4824 4050
rect 4424 3690 4464 4010
rect 4784 3690 4824 4010
rect 4424 3650 4824 3690
rect 5143 4010 5543 4050
rect 5143 3690 5183 4010
rect 5503 3690 5543 4010
rect 5143 3650 5543 3690
rect 5862 4010 6262 4050
rect 5862 3690 5902 4010
rect 6222 3690 6262 4010
rect 5862 3650 6262 3690
rect 6581 4010 6981 4050
rect 6581 3690 6621 4010
rect 6941 3690 6981 4010
rect 6581 3650 6981 3690
rect -7080 3310 -6680 3350
rect -7080 2990 -7040 3310
rect -6720 2990 -6680 3310
rect -7080 2950 -6680 2990
rect -6361 3310 -5961 3350
rect -6361 2990 -6321 3310
rect -6001 2990 -5961 3310
rect -6361 2950 -5961 2990
rect -5642 3310 -5242 3350
rect -5642 2990 -5602 3310
rect -5282 2990 -5242 3310
rect -5642 2950 -5242 2990
rect -4923 3310 -4523 3350
rect -4923 2990 -4883 3310
rect -4563 2990 -4523 3310
rect -4923 2950 -4523 2990
rect -4204 3310 -3804 3350
rect -4204 2990 -4164 3310
rect -3844 2990 -3804 3310
rect -4204 2950 -3804 2990
rect -3485 3310 -3085 3350
rect -3485 2990 -3445 3310
rect -3125 2990 -3085 3310
rect -3485 2950 -3085 2990
rect -2766 3310 -2366 3350
rect -2766 2990 -2726 3310
rect -2406 2990 -2366 3310
rect -2766 2950 -2366 2990
rect -2047 3310 -1647 3350
rect -2047 2990 -2007 3310
rect -1687 2990 -1647 3310
rect -2047 2950 -1647 2990
rect -1328 3310 -928 3350
rect -1328 2990 -1288 3310
rect -968 2990 -928 3310
rect -1328 2950 -928 2990
rect -609 3310 -209 3350
rect -609 2990 -569 3310
rect -249 2990 -209 3310
rect -609 2950 -209 2990
rect 110 3310 510 3350
rect 110 2990 150 3310
rect 470 2990 510 3310
rect 110 2950 510 2990
rect 829 3310 1229 3350
rect 829 2990 869 3310
rect 1189 2990 1229 3310
rect 829 2950 1229 2990
rect 1548 3310 1948 3350
rect 1548 2990 1588 3310
rect 1908 2990 1948 3310
rect 1548 2950 1948 2990
rect 2267 3310 2667 3350
rect 2267 2990 2307 3310
rect 2627 2990 2667 3310
rect 2267 2950 2667 2990
rect 2986 3310 3386 3350
rect 2986 2990 3026 3310
rect 3346 2990 3386 3310
rect 2986 2950 3386 2990
rect 3705 3310 4105 3350
rect 3705 2990 3745 3310
rect 4065 2990 4105 3310
rect 3705 2950 4105 2990
rect 4424 3310 4824 3350
rect 4424 2990 4464 3310
rect 4784 2990 4824 3310
rect 4424 2950 4824 2990
rect 5143 3310 5543 3350
rect 5143 2990 5183 3310
rect 5503 2990 5543 3310
rect 5143 2950 5543 2990
rect 5862 3310 6262 3350
rect 5862 2990 5902 3310
rect 6222 2990 6262 3310
rect 5862 2950 6262 2990
rect 6581 3310 6981 3350
rect 6581 2990 6621 3310
rect 6941 2990 6981 3310
rect 6581 2950 6981 2990
rect -7080 2610 -6680 2650
rect -7080 2290 -7040 2610
rect -6720 2290 -6680 2610
rect -7080 2250 -6680 2290
rect -6361 2610 -5961 2650
rect -6361 2290 -6321 2610
rect -6001 2290 -5961 2610
rect -6361 2250 -5961 2290
rect -5642 2610 -5242 2650
rect -5642 2290 -5602 2610
rect -5282 2290 -5242 2610
rect -5642 2250 -5242 2290
rect -4923 2610 -4523 2650
rect -4923 2290 -4883 2610
rect -4563 2290 -4523 2610
rect -4923 2250 -4523 2290
rect -4204 2610 -3804 2650
rect -4204 2290 -4164 2610
rect -3844 2290 -3804 2610
rect -4204 2250 -3804 2290
rect -3485 2610 -3085 2650
rect -3485 2290 -3445 2610
rect -3125 2290 -3085 2610
rect -3485 2250 -3085 2290
rect -2766 2610 -2366 2650
rect -2766 2290 -2726 2610
rect -2406 2290 -2366 2610
rect -2766 2250 -2366 2290
rect -2047 2610 -1647 2650
rect -2047 2290 -2007 2610
rect -1687 2290 -1647 2610
rect -2047 2250 -1647 2290
rect -1328 2610 -928 2650
rect -1328 2290 -1288 2610
rect -968 2290 -928 2610
rect -1328 2250 -928 2290
rect -609 2610 -209 2650
rect -609 2290 -569 2610
rect -249 2290 -209 2610
rect -609 2250 -209 2290
rect 110 2610 510 2650
rect 110 2290 150 2610
rect 470 2290 510 2610
rect 110 2250 510 2290
rect 829 2610 1229 2650
rect 829 2290 869 2610
rect 1189 2290 1229 2610
rect 829 2250 1229 2290
rect 1548 2610 1948 2650
rect 1548 2290 1588 2610
rect 1908 2290 1948 2610
rect 1548 2250 1948 2290
rect 2267 2610 2667 2650
rect 2267 2290 2307 2610
rect 2627 2290 2667 2610
rect 2267 2250 2667 2290
rect 2986 2610 3386 2650
rect 2986 2290 3026 2610
rect 3346 2290 3386 2610
rect 2986 2250 3386 2290
rect 3705 2610 4105 2650
rect 3705 2290 3745 2610
rect 4065 2290 4105 2610
rect 3705 2250 4105 2290
rect 4424 2610 4824 2650
rect 4424 2290 4464 2610
rect 4784 2290 4824 2610
rect 4424 2250 4824 2290
rect 5143 2610 5543 2650
rect 5143 2290 5183 2610
rect 5503 2290 5543 2610
rect 5143 2250 5543 2290
rect 5862 2610 6262 2650
rect 5862 2290 5902 2610
rect 6222 2290 6262 2610
rect 5862 2250 6262 2290
rect 6581 2610 6981 2650
rect 6581 2290 6621 2610
rect 6941 2290 6981 2610
rect 6581 2250 6981 2290
rect -7080 1910 -6680 1950
rect -7080 1590 -7040 1910
rect -6720 1590 -6680 1910
rect -7080 1550 -6680 1590
rect -6361 1910 -5961 1950
rect -6361 1590 -6321 1910
rect -6001 1590 -5961 1910
rect -6361 1550 -5961 1590
rect -5642 1910 -5242 1950
rect -5642 1590 -5602 1910
rect -5282 1590 -5242 1910
rect -5642 1550 -5242 1590
rect -4923 1910 -4523 1950
rect -4923 1590 -4883 1910
rect -4563 1590 -4523 1910
rect -4923 1550 -4523 1590
rect -4204 1910 -3804 1950
rect -4204 1590 -4164 1910
rect -3844 1590 -3804 1910
rect -4204 1550 -3804 1590
rect -3485 1910 -3085 1950
rect -3485 1590 -3445 1910
rect -3125 1590 -3085 1910
rect -3485 1550 -3085 1590
rect -2766 1910 -2366 1950
rect -2766 1590 -2726 1910
rect -2406 1590 -2366 1910
rect -2766 1550 -2366 1590
rect -2047 1910 -1647 1950
rect -2047 1590 -2007 1910
rect -1687 1590 -1647 1910
rect -2047 1550 -1647 1590
rect -1328 1910 -928 1950
rect -1328 1590 -1288 1910
rect -968 1590 -928 1910
rect -1328 1550 -928 1590
rect -609 1910 -209 1950
rect -609 1590 -569 1910
rect -249 1590 -209 1910
rect -609 1550 -209 1590
rect 110 1910 510 1950
rect 110 1590 150 1910
rect 470 1590 510 1910
rect 110 1550 510 1590
rect 829 1910 1229 1950
rect 829 1590 869 1910
rect 1189 1590 1229 1910
rect 829 1550 1229 1590
rect 1548 1910 1948 1950
rect 1548 1590 1588 1910
rect 1908 1590 1948 1910
rect 1548 1550 1948 1590
rect 2267 1910 2667 1950
rect 2267 1590 2307 1910
rect 2627 1590 2667 1910
rect 2267 1550 2667 1590
rect 2986 1910 3386 1950
rect 2986 1590 3026 1910
rect 3346 1590 3386 1910
rect 2986 1550 3386 1590
rect 3705 1910 4105 1950
rect 3705 1590 3745 1910
rect 4065 1590 4105 1910
rect 3705 1550 4105 1590
rect 4424 1910 4824 1950
rect 4424 1590 4464 1910
rect 4784 1590 4824 1910
rect 4424 1550 4824 1590
rect 5143 1910 5543 1950
rect 5143 1590 5183 1910
rect 5503 1590 5543 1910
rect 5143 1550 5543 1590
rect 5862 1910 6262 1950
rect 5862 1590 5902 1910
rect 6222 1590 6262 1910
rect 5862 1550 6262 1590
rect 6581 1910 6981 1950
rect 6581 1590 6621 1910
rect 6941 1590 6981 1910
rect 6581 1550 6981 1590
rect -7080 1210 -6680 1250
rect -7080 890 -7040 1210
rect -6720 890 -6680 1210
rect -7080 850 -6680 890
rect -6361 1210 -5961 1250
rect -6361 890 -6321 1210
rect -6001 890 -5961 1210
rect -6361 850 -5961 890
rect -5642 1210 -5242 1250
rect -5642 890 -5602 1210
rect -5282 890 -5242 1210
rect -5642 850 -5242 890
rect -4923 1210 -4523 1250
rect -4923 890 -4883 1210
rect -4563 890 -4523 1210
rect -4923 850 -4523 890
rect -4204 1210 -3804 1250
rect -4204 890 -4164 1210
rect -3844 890 -3804 1210
rect -4204 850 -3804 890
rect -3485 1210 -3085 1250
rect -3485 890 -3445 1210
rect -3125 890 -3085 1210
rect -3485 850 -3085 890
rect -2766 1210 -2366 1250
rect -2766 890 -2726 1210
rect -2406 890 -2366 1210
rect -2766 850 -2366 890
rect -2047 1210 -1647 1250
rect -2047 890 -2007 1210
rect -1687 890 -1647 1210
rect -2047 850 -1647 890
rect -1328 1210 -928 1250
rect -1328 890 -1288 1210
rect -968 890 -928 1210
rect -1328 850 -928 890
rect -609 1210 -209 1250
rect -609 890 -569 1210
rect -249 890 -209 1210
rect -609 850 -209 890
rect 110 1210 510 1250
rect 110 890 150 1210
rect 470 890 510 1210
rect 110 850 510 890
rect 829 1210 1229 1250
rect 829 890 869 1210
rect 1189 890 1229 1210
rect 829 850 1229 890
rect 1548 1210 1948 1250
rect 1548 890 1588 1210
rect 1908 890 1948 1210
rect 1548 850 1948 890
rect 2267 1210 2667 1250
rect 2267 890 2307 1210
rect 2627 890 2667 1210
rect 2267 850 2667 890
rect 2986 1210 3386 1250
rect 2986 890 3026 1210
rect 3346 890 3386 1210
rect 2986 850 3386 890
rect 3705 1210 4105 1250
rect 3705 890 3745 1210
rect 4065 890 4105 1210
rect 3705 850 4105 890
rect 4424 1210 4824 1250
rect 4424 890 4464 1210
rect 4784 890 4824 1210
rect 4424 850 4824 890
rect 5143 1210 5543 1250
rect 5143 890 5183 1210
rect 5503 890 5543 1210
rect 5143 850 5543 890
rect 5862 1210 6262 1250
rect 5862 890 5902 1210
rect 6222 890 6262 1210
rect 5862 850 6262 890
rect 6581 1210 6981 1250
rect 6581 890 6621 1210
rect 6941 890 6981 1210
rect 6581 850 6981 890
rect -7080 510 -6680 550
rect -7080 190 -7040 510
rect -6720 190 -6680 510
rect -7080 150 -6680 190
rect -6361 510 -5961 550
rect -6361 190 -6321 510
rect -6001 190 -5961 510
rect -6361 150 -5961 190
rect -5642 510 -5242 550
rect -5642 190 -5602 510
rect -5282 190 -5242 510
rect -5642 150 -5242 190
rect -4923 510 -4523 550
rect -4923 190 -4883 510
rect -4563 190 -4523 510
rect -4923 150 -4523 190
rect -4204 510 -3804 550
rect -4204 190 -4164 510
rect -3844 190 -3804 510
rect -4204 150 -3804 190
rect -3485 510 -3085 550
rect -3485 190 -3445 510
rect -3125 190 -3085 510
rect -3485 150 -3085 190
rect -2766 510 -2366 550
rect -2766 190 -2726 510
rect -2406 190 -2366 510
rect -2766 150 -2366 190
rect -2047 510 -1647 550
rect -2047 190 -2007 510
rect -1687 190 -1647 510
rect -2047 150 -1647 190
rect -1328 510 -928 550
rect -1328 190 -1288 510
rect -968 190 -928 510
rect -1328 150 -928 190
rect -609 510 -209 550
rect -609 190 -569 510
rect -249 190 -209 510
rect -609 150 -209 190
rect 110 510 510 550
rect 110 190 150 510
rect 470 190 510 510
rect 110 150 510 190
rect 829 510 1229 550
rect 829 190 869 510
rect 1189 190 1229 510
rect 829 150 1229 190
rect 1548 510 1948 550
rect 1548 190 1588 510
rect 1908 190 1948 510
rect 1548 150 1948 190
rect 2267 510 2667 550
rect 2267 190 2307 510
rect 2627 190 2667 510
rect 2267 150 2667 190
rect 2986 510 3386 550
rect 2986 190 3026 510
rect 3346 190 3386 510
rect 2986 150 3386 190
rect 3705 510 4105 550
rect 3705 190 3745 510
rect 4065 190 4105 510
rect 3705 150 4105 190
rect 4424 510 4824 550
rect 4424 190 4464 510
rect 4784 190 4824 510
rect 4424 150 4824 190
rect 5143 510 5543 550
rect 5143 190 5183 510
rect 5503 190 5543 510
rect 5143 150 5543 190
rect 5862 510 6262 550
rect 5862 190 5902 510
rect 6222 190 6262 510
rect 5862 150 6262 190
rect 6581 510 6981 550
rect 6581 190 6621 510
rect 6941 190 6981 510
rect 6581 150 6981 190
rect -7080 -190 -6680 -150
rect -7080 -510 -7040 -190
rect -6720 -510 -6680 -190
rect -7080 -550 -6680 -510
rect -6361 -190 -5961 -150
rect -6361 -510 -6321 -190
rect -6001 -510 -5961 -190
rect -6361 -550 -5961 -510
rect -5642 -190 -5242 -150
rect -5642 -510 -5602 -190
rect -5282 -510 -5242 -190
rect -5642 -550 -5242 -510
rect -4923 -190 -4523 -150
rect -4923 -510 -4883 -190
rect -4563 -510 -4523 -190
rect -4923 -550 -4523 -510
rect -4204 -190 -3804 -150
rect -4204 -510 -4164 -190
rect -3844 -510 -3804 -190
rect -4204 -550 -3804 -510
rect -3485 -190 -3085 -150
rect -3485 -510 -3445 -190
rect -3125 -510 -3085 -190
rect -3485 -550 -3085 -510
rect -2766 -190 -2366 -150
rect -2766 -510 -2726 -190
rect -2406 -510 -2366 -190
rect -2766 -550 -2366 -510
rect -2047 -190 -1647 -150
rect -2047 -510 -2007 -190
rect -1687 -510 -1647 -190
rect -2047 -550 -1647 -510
rect -1328 -190 -928 -150
rect -1328 -510 -1288 -190
rect -968 -510 -928 -190
rect -1328 -550 -928 -510
rect -609 -190 -209 -150
rect -609 -510 -569 -190
rect -249 -510 -209 -190
rect -609 -550 -209 -510
rect 110 -190 510 -150
rect 110 -510 150 -190
rect 470 -510 510 -190
rect 110 -550 510 -510
rect 829 -190 1229 -150
rect 829 -510 869 -190
rect 1189 -510 1229 -190
rect 829 -550 1229 -510
rect 1548 -190 1948 -150
rect 1548 -510 1588 -190
rect 1908 -510 1948 -190
rect 1548 -550 1948 -510
rect 2267 -190 2667 -150
rect 2267 -510 2307 -190
rect 2627 -510 2667 -190
rect 2267 -550 2667 -510
rect 2986 -190 3386 -150
rect 2986 -510 3026 -190
rect 3346 -510 3386 -190
rect 2986 -550 3386 -510
rect 3705 -190 4105 -150
rect 3705 -510 3745 -190
rect 4065 -510 4105 -190
rect 3705 -550 4105 -510
rect 4424 -190 4824 -150
rect 4424 -510 4464 -190
rect 4784 -510 4824 -190
rect 4424 -550 4824 -510
rect 5143 -190 5543 -150
rect 5143 -510 5183 -190
rect 5503 -510 5543 -190
rect 5143 -550 5543 -510
rect 5862 -190 6262 -150
rect 5862 -510 5902 -190
rect 6222 -510 6262 -190
rect 5862 -550 6262 -510
rect 6581 -190 6981 -150
rect 6581 -510 6621 -190
rect 6941 -510 6981 -190
rect 6581 -550 6981 -510
rect -7080 -890 -6680 -850
rect -7080 -1210 -7040 -890
rect -6720 -1210 -6680 -890
rect -7080 -1250 -6680 -1210
rect -6361 -890 -5961 -850
rect -6361 -1210 -6321 -890
rect -6001 -1210 -5961 -890
rect -6361 -1250 -5961 -1210
rect -5642 -890 -5242 -850
rect -5642 -1210 -5602 -890
rect -5282 -1210 -5242 -890
rect -5642 -1250 -5242 -1210
rect -4923 -890 -4523 -850
rect -4923 -1210 -4883 -890
rect -4563 -1210 -4523 -890
rect -4923 -1250 -4523 -1210
rect -4204 -890 -3804 -850
rect -4204 -1210 -4164 -890
rect -3844 -1210 -3804 -890
rect -4204 -1250 -3804 -1210
rect -3485 -890 -3085 -850
rect -3485 -1210 -3445 -890
rect -3125 -1210 -3085 -890
rect -3485 -1250 -3085 -1210
rect -2766 -890 -2366 -850
rect -2766 -1210 -2726 -890
rect -2406 -1210 -2366 -890
rect -2766 -1250 -2366 -1210
rect -2047 -890 -1647 -850
rect -2047 -1210 -2007 -890
rect -1687 -1210 -1647 -890
rect -2047 -1250 -1647 -1210
rect -1328 -890 -928 -850
rect -1328 -1210 -1288 -890
rect -968 -1210 -928 -890
rect -1328 -1250 -928 -1210
rect -609 -890 -209 -850
rect -609 -1210 -569 -890
rect -249 -1210 -209 -890
rect -609 -1250 -209 -1210
rect 110 -890 510 -850
rect 110 -1210 150 -890
rect 470 -1210 510 -890
rect 110 -1250 510 -1210
rect 829 -890 1229 -850
rect 829 -1210 869 -890
rect 1189 -1210 1229 -890
rect 829 -1250 1229 -1210
rect 1548 -890 1948 -850
rect 1548 -1210 1588 -890
rect 1908 -1210 1948 -890
rect 1548 -1250 1948 -1210
rect 2267 -890 2667 -850
rect 2267 -1210 2307 -890
rect 2627 -1210 2667 -890
rect 2267 -1250 2667 -1210
rect 2986 -890 3386 -850
rect 2986 -1210 3026 -890
rect 3346 -1210 3386 -890
rect 2986 -1250 3386 -1210
rect 3705 -890 4105 -850
rect 3705 -1210 3745 -890
rect 4065 -1210 4105 -890
rect 3705 -1250 4105 -1210
rect 4424 -890 4824 -850
rect 4424 -1210 4464 -890
rect 4784 -1210 4824 -890
rect 4424 -1250 4824 -1210
rect 5143 -890 5543 -850
rect 5143 -1210 5183 -890
rect 5503 -1210 5543 -890
rect 5143 -1250 5543 -1210
rect 5862 -890 6262 -850
rect 5862 -1210 5902 -890
rect 6222 -1210 6262 -890
rect 5862 -1250 6262 -1210
rect 6581 -890 6981 -850
rect 6581 -1210 6621 -890
rect 6941 -1210 6981 -890
rect 6581 -1250 6981 -1210
rect -7080 -1590 -6680 -1550
rect -7080 -1910 -7040 -1590
rect -6720 -1910 -6680 -1590
rect -7080 -1950 -6680 -1910
rect -6361 -1590 -5961 -1550
rect -6361 -1910 -6321 -1590
rect -6001 -1910 -5961 -1590
rect -6361 -1950 -5961 -1910
rect -5642 -1590 -5242 -1550
rect -5642 -1910 -5602 -1590
rect -5282 -1910 -5242 -1590
rect -5642 -1950 -5242 -1910
rect -4923 -1590 -4523 -1550
rect -4923 -1910 -4883 -1590
rect -4563 -1910 -4523 -1590
rect -4923 -1950 -4523 -1910
rect -4204 -1590 -3804 -1550
rect -4204 -1910 -4164 -1590
rect -3844 -1910 -3804 -1590
rect -4204 -1950 -3804 -1910
rect -3485 -1590 -3085 -1550
rect -3485 -1910 -3445 -1590
rect -3125 -1910 -3085 -1590
rect -3485 -1950 -3085 -1910
rect -2766 -1590 -2366 -1550
rect -2766 -1910 -2726 -1590
rect -2406 -1910 -2366 -1590
rect -2766 -1950 -2366 -1910
rect -2047 -1590 -1647 -1550
rect -2047 -1910 -2007 -1590
rect -1687 -1910 -1647 -1590
rect -2047 -1950 -1647 -1910
rect -1328 -1590 -928 -1550
rect -1328 -1910 -1288 -1590
rect -968 -1910 -928 -1590
rect -1328 -1950 -928 -1910
rect -609 -1590 -209 -1550
rect -609 -1910 -569 -1590
rect -249 -1910 -209 -1590
rect -609 -1950 -209 -1910
rect 110 -1590 510 -1550
rect 110 -1910 150 -1590
rect 470 -1910 510 -1590
rect 110 -1950 510 -1910
rect 829 -1590 1229 -1550
rect 829 -1910 869 -1590
rect 1189 -1910 1229 -1590
rect 829 -1950 1229 -1910
rect 1548 -1590 1948 -1550
rect 1548 -1910 1588 -1590
rect 1908 -1910 1948 -1590
rect 1548 -1950 1948 -1910
rect 2267 -1590 2667 -1550
rect 2267 -1910 2307 -1590
rect 2627 -1910 2667 -1590
rect 2267 -1950 2667 -1910
rect 2986 -1590 3386 -1550
rect 2986 -1910 3026 -1590
rect 3346 -1910 3386 -1590
rect 2986 -1950 3386 -1910
rect 3705 -1590 4105 -1550
rect 3705 -1910 3745 -1590
rect 4065 -1910 4105 -1590
rect 3705 -1950 4105 -1910
rect 4424 -1590 4824 -1550
rect 4424 -1910 4464 -1590
rect 4784 -1910 4824 -1590
rect 4424 -1950 4824 -1910
rect 5143 -1590 5543 -1550
rect 5143 -1910 5183 -1590
rect 5503 -1910 5543 -1590
rect 5143 -1950 5543 -1910
rect 5862 -1590 6262 -1550
rect 5862 -1910 5902 -1590
rect 6222 -1910 6262 -1590
rect 5862 -1950 6262 -1910
rect 6581 -1590 6981 -1550
rect 6581 -1910 6621 -1590
rect 6941 -1910 6981 -1590
rect 6581 -1950 6981 -1910
rect -7080 -2290 -6680 -2250
rect -7080 -2610 -7040 -2290
rect -6720 -2610 -6680 -2290
rect -7080 -2650 -6680 -2610
rect -6361 -2290 -5961 -2250
rect -6361 -2610 -6321 -2290
rect -6001 -2610 -5961 -2290
rect -6361 -2650 -5961 -2610
rect -5642 -2290 -5242 -2250
rect -5642 -2610 -5602 -2290
rect -5282 -2610 -5242 -2290
rect -5642 -2650 -5242 -2610
rect -4923 -2290 -4523 -2250
rect -4923 -2610 -4883 -2290
rect -4563 -2610 -4523 -2290
rect -4923 -2650 -4523 -2610
rect -4204 -2290 -3804 -2250
rect -4204 -2610 -4164 -2290
rect -3844 -2610 -3804 -2290
rect -4204 -2650 -3804 -2610
rect -3485 -2290 -3085 -2250
rect -3485 -2610 -3445 -2290
rect -3125 -2610 -3085 -2290
rect -3485 -2650 -3085 -2610
rect -2766 -2290 -2366 -2250
rect -2766 -2610 -2726 -2290
rect -2406 -2610 -2366 -2290
rect -2766 -2650 -2366 -2610
rect -2047 -2290 -1647 -2250
rect -2047 -2610 -2007 -2290
rect -1687 -2610 -1647 -2290
rect -2047 -2650 -1647 -2610
rect -1328 -2290 -928 -2250
rect -1328 -2610 -1288 -2290
rect -968 -2610 -928 -2290
rect -1328 -2650 -928 -2610
rect -609 -2290 -209 -2250
rect -609 -2610 -569 -2290
rect -249 -2610 -209 -2290
rect -609 -2650 -209 -2610
rect 110 -2290 510 -2250
rect 110 -2610 150 -2290
rect 470 -2610 510 -2290
rect 110 -2650 510 -2610
rect 829 -2290 1229 -2250
rect 829 -2610 869 -2290
rect 1189 -2610 1229 -2290
rect 829 -2650 1229 -2610
rect 1548 -2290 1948 -2250
rect 1548 -2610 1588 -2290
rect 1908 -2610 1948 -2290
rect 1548 -2650 1948 -2610
rect 2267 -2290 2667 -2250
rect 2267 -2610 2307 -2290
rect 2627 -2610 2667 -2290
rect 2267 -2650 2667 -2610
rect 2986 -2290 3386 -2250
rect 2986 -2610 3026 -2290
rect 3346 -2610 3386 -2290
rect 2986 -2650 3386 -2610
rect 3705 -2290 4105 -2250
rect 3705 -2610 3745 -2290
rect 4065 -2610 4105 -2290
rect 3705 -2650 4105 -2610
rect 4424 -2290 4824 -2250
rect 4424 -2610 4464 -2290
rect 4784 -2610 4824 -2290
rect 4424 -2650 4824 -2610
rect 5143 -2290 5543 -2250
rect 5143 -2610 5183 -2290
rect 5503 -2610 5543 -2290
rect 5143 -2650 5543 -2610
rect 5862 -2290 6262 -2250
rect 5862 -2610 5902 -2290
rect 6222 -2610 6262 -2290
rect 5862 -2650 6262 -2610
rect 6581 -2290 6981 -2250
rect 6581 -2610 6621 -2290
rect 6941 -2610 6981 -2290
rect 6581 -2650 6981 -2610
rect -7080 -2990 -6680 -2950
rect -7080 -3310 -7040 -2990
rect -6720 -3310 -6680 -2990
rect -7080 -3350 -6680 -3310
rect -6361 -2990 -5961 -2950
rect -6361 -3310 -6321 -2990
rect -6001 -3310 -5961 -2990
rect -6361 -3350 -5961 -3310
rect -5642 -2990 -5242 -2950
rect -5642 -3310 -5602 -2990
rect -5282 -3310 -5242 -2990
rect -5642 -3350 -5242 -3310
rect -4923 -2990 -4523 -2950
rect -4923 -3310 -4883 -2990
rect -4563 -3310 -4523 -2990
rect -4923 -3350 -4523 -3310
rect -4204 -2990 -3804 -2950
rect -4204 -3310 -4164 -2990
rect -3844 -3310 -3804 -2990
rect -4204 -3350 -3804 -3310
rect -3485 -2990 -3085 -2950
rect -3485 -3310 -3445 -2990
rect -3125 -3310 -3085 -2990
rect -3485 -3350 -3085 -3310
rect -2766 -2990 -2366 -2950
rect -2766 -3310 -2726 -2990
rect -2406 -3310 -2366 -2990
rect -2766 -3350 -2366 -3310
rect -2047 -2990 -1647 -2950
rect -2047 -3310 -2007 -2990
rect -1687 -3310 -1647 -2990
rect -2047 -3350 -1647 -3310
rect -1328 -2990 -928 -2950
rect -1328 -3310 -1288 -2990
rect -968 -3310 -928 -2990
rect -1328 -3350 -928 -3310
rect -609 -2990 -209 -2950
rect -609 -3310 -569 -2990
rect -249 -3310 -209 -2990
rect -609 -3350 -209 -3310
rect 110 -2990 510 -2950
rect 110 -3310 150 -2990
rect 470 -3310 510 -2990
rect 110 -3350 510 -3310
rect 829 -2990 1229 -2950
rect 829 -3310 869 -2990
rect 1189 -3310 1229 -2990
rect 829 -3350 1229 -3310
rect 1548 -2990 1948 -2950
rect 1548 -3310 1588 -2990
rect 1908 -3310 1948 -2990
rect 1548 -3350 1948 -3310
rect 2267 -2990 2667 -2950
rect 2267 -3310 2307 -2990
rect 2627 -3310 2667 -2990
rect 2267 -3350 2667 -3310
rect 2986 -2990 3386 -2950
rect 2986 -3310 3026 -2990
rect 3346 -3310 3386 -2990
rect 2986 -3350 3386 -3310
rect 3705 -2990 4105 -2950
rect 3705 -3310 3745 -2990
rect 4065 -3310 4105 -2990
rect 3705 -3350 4105 -3310
rect 4424 -2990 4824 -2950
rect 4424 -3310 4464 -2990
rect 4784 -3310 4824 -2990
rect 4424 -3350 4824 -3310
rect 5143 -2990 5543 -2950
rect 5143 -3310 5183 -2990
rect 5503 -3310 5543 -2990
rect 5143 -3350 5543 -3310
rect 5862 -2990 6262 -2950
rect 5862 -3310 5902 -2990
rect 6222 -3310 6262 -2990
rect 5862 -3350 6262 -3310
rect 6581 -2990 6981 -2950
rect 6581 -3310 6621 -2990
rect 6941 -3310 6981 -2990
rect 6581 -3350 6981 -3310
rect -7080 -3690 -6680 -3650
rect -7080 -4010 -7040 -3690
rect -6720 -4010 -6680 -3690
rect -7080 -4050 -6680 -4010
rect -6361 -3690 -5961 -3650
rect -6361 -4010 -6321 -3690
rect -6001 -4010 -5961 -3690
rect -6361 -4050 -5961 -4010
rect -5642 -3690 -5242 -3650
rect -5642 -4010 -5602 -3690
rect -5282 -4010 -5242 -3690
rect -5642 -4050 -5242 -4010
rect -4923 -3690 -4523 -3650
rect -4923 -4010 -4883 -3690
rect -4563 -4010 -4523 -3690
rect -4923 -4050 -4523 -4010
rect -4204 -3690 -3804 -3650
rect -4204 -4010 -4164 -3690
rect -3844 -4010 -3804 -3690
rect -4204 -4050 -3804 -4010
rect -3485 -3690 -3085 -3650
rect -3485 -4010 -3445 -3690
rect -3125 -4010 -3085 -3690
rect -3485 -4050 -3085 -4010
rect -2766 -3690 -2366 -3650
rect -2766 -4010 -2726 -3690
rect -2406 -4010 -2366 -3690
rect -2766 -4050 -2366 -4010
rect -2047 -3690 -1647 -3650
rect -2047 -4010 -2007 -3690
rect -1687 -4010 -1647 -3690
rect -2047 -4050 -1647 -4010
rect -1328 -3690 -928 -3650
rect -1328 -4010 -1288 -3690
rect -968 -4010 -928 -3690
rect -1328 -4050 -928 -4010
rect -609 -3690 -209 -3650
rect -609 -4010 -569 -3690
rect -249 -4010 -209 -3690
rect -609 -4050 -209 -4010
rect 110 -3690 510 -3650
rect 110 -4010 150 -3690
rect 470 -4010 510 -3690
rect 110 -4050 510 -4010
rect 829 -3690 1229 -3650
rect 829 -4010 869 -3690
rect 1189 -4010 1229 -3690
rect 829 -4050 1229 -4010
rect 1548 -3690 1948 -3650
rect 1548 -4010 1588 -3690
rect 1908 -4010 1948 -3690
rect 1548 -4050 1948 -4010
rect 2267 -3690 2667 -3650
rect 2267 -4010 2307 -3690
rect 2627 -4010 2667 -3690
rect 2267 -4050 2667 -4010
rect 2986 -3690 3386 -3650
rect 2986 -4010 3026 -3690
rect 3346 -4010 3386 -3690
rect 2986 -4050 3386 -4010
rect 3705 -3690 4105 -3650
rect 3705 -4010 3745 -3690
rect 4065 -4010 4105 -3690
rect 3705 -4050 4105 -4010
rect 4424 -3690 4824 -3650
rect 4424 -4010 4464 -3690
rect 4784 -4010 4824 -3690
rect 4424 -4050 4824 -4010
rect 5143 -3690 5543 -3650
rect 5143 -4010 5183 -3690
rect 5503 -4010 5543 -3690
rect 5143 -4050 5543 -4010
rect 5862 -3690 6262 -3650
rect 5862 -4010 5902 -3690
rect 6222 -4010 6262 -3690
rect 5862 -4050 6262 -4010
rect 6581 -3690 6981 -3650
rect 6581 -4010 6621 -3690
rect 6941 -4010 6981 -3690
rect 6581 -4050 6981 -4010
rect -7080 -4390 -6680 -4350
rect -7080 -4710 -7040 -4390
rect -6720 -4710 -6680 -4390
rect -7080 -4750 -6680 -4710
rect -6361 -4390 -5961 -4350
rect -6361 -4710 -6321 -4390
rect -6001 -4710 -5961 -4390
rect -6361 -4750 -5961 -4710
rect -5642 -4390 -5242 -4350
rect -5642 -4710 -5602 -4390
rect -5282 -4710 -5242 -4390
rect -5642 -4750 -5242 -4710
rect -4923 -4390 -4523 -4350
rect -4923 -4710 -4883 -4390
rect -4563 -4710 -4523 -4390
rect -4923 -4750 -4523 -4710
rect -4204 -4390 -3804 -4350
rect -4204 -4710 -4164 -4390
rect -3844 -4710 -3804 -4390
rect -4204 -4750 -3804 -4710
rect -3485 -4390 -3085 -4350
rect -3485 -4710 -3445 -4390
rect -3125 -4710 -3085 -4390
rect -3485 -4750 -3085 -4710
rect -2766 -4390 -2366 -4350
rect -2766 -4710 -2726 -4390
rect -2406 -4710 -2366 -4390
rect -2766 -4750 -2366 -4710
rect -2047 -4390 -1647 -4350
rect -2047 -4710 -2007 -4390
rect -1687 -4710 -1647 -4390
rect -2047 -4750 -1647 -4710
rect -1328 -4390 -928 -4350
rect -1328 -4710 -1288 -4390
rect -968 -4710 -928 -4390
rect -1328 -4750 -928 -4710
rect -609 -4390 -209 -4350
rect -609 -4710 -569 -4390
rect -249 -4710 -209 -4390
rect -609 -4750 -209 -4710
rect 110 -4390 510 -4350
rect 110 -4710 150 -4390
rect 470 -4710 510 -4390
rect 110 -4750 510 -4710
rect 829 -4390 1229 -4350
rect 829 -4710 869 -4390
rect 1189 -4710 1229 -4390
rect 829 -4750 1229 -4710
rect 1548 -4390 1948 -4350
rect 1548 -4710 1588 -4390
rect 1908 -4710 1948 -4390
rect 1548 -4750 1948 -4710
rect 2267 -4390 2667 -4350
rect 2267 -4710 2307 -4390
rect 2627 -4710 2667 -4390
rect 2267 -4750 2667 -4710
rect 2986 -4390 3386 -4350
rect 2986 -4710 3026 -4390
rect 3346 -4710 3386 -4390
rect 2986 -4750 3386 -4710
rect 3705 -4390 4105 -4350
rect 3705 -4710 3745 -4390
rect 4065 -4710 4105 -4390
rect 3705 -4750 4105 -4710
rect 4424 -4390 4824 -4350
rect 4424 -4710 4464 -4390
rect 4784 -4710 4824 -4390
rect 4424 -4750 4824 -4710
rect 5143 -4390 5543 -4350
rect 5143 -4710 5183 -4390
rect 5503 -4710 5543 -4390
rect 5143 -4750 5543 -4710
rect 5862 -4390 6262 -4350
rect 5862 -4710 5902 -4390
rect 6222 -4710 6262 -4390
rect 5862 -4750 6262 -4710
rect 6581 -4390 6981 -4350
rect 6581 -4710 6621 -4390
rect 6941 -4710 6981 -4390
rect 6581 -4750 6981 -4710
rect -7080 -5090 -6680 -5050
rect -7080 -5410 -7040 -5090
rect -6720 -5410 -6680 -5090
rect -7080 -5450 -6680 -5410
rect -6361 -5090 -5961 -5050
rect -6361 -5410 -6321 -5090
rect -6001 -5410 -5961 -5090
rect -6361 -5450 -5961 -5410
rect -5642 -5090 -5242 -5050
rect -5642 -5410 -5602 -5090
rect -5282 -5410 -5242 -5090
rect -5642 -5450 -5242 -5410
rect -4923 -5090 -4523 -5050
rect -4923 -5410 -4883 -5090
rect -4563 -5410 -4523 -5090
rect -4923 -5450 -4523 -5410
rect -4204 -5090 -3804 -5050
rect -4204 -5410 -4164 -5090
rect -3844 -5410 -3804 -5090
rect -4204 -5450 -3804 -5410
rect -3485 -5090 -3085 -5050
rect -3485 -5410 -3445 -5090
rect -3125 -5410 -3085 -5090
rect -3485 -5450 -3085 -5410
rect -2766 -5090 -2366 -5050
rect -2766 -5410 -2726 -5090
rect -2406 -5410 -2366 -5090
rect -2766 -5450 -2366 -5410
rect -2047 -5090 -1647 -5050
rect -2047 -5410 -2007 -5090
rect -1687 -5410 -1647 -5090
rect -2047 -5450 -1647 -5410
rect -1328 -5090 -928 -5050
rect -1328 -5410 -1288 -5090
rect -968 -5410 -928 -5090
rect -1328 -5450 -928 -5410
rect -609 -5090 -209 -5050
rect -609 -5410 -569 -5090
rect -249 -5410 -209 -5090
rect -609 -5450 -209 -5410
rect 110 -5090 510 -5050
rect 110 -5410 150 -5090
rect 470 -5410 510 -5090
rect 110 -5450 510 -5410
rect 829 -5090 1229 -5050
rect 829 -5410 869 -5090
rect 1189 -5410 1229 -5090
rect 829 -5450 1229 -5410
rect 1548 -5090 1948 -5050
rect 1548 -5410 1588 -5090
rect 1908 -5410 1948 -5090
rect 1548 -5450 1948 -5410
rect 2267 -5090 2667 -5050
rect 2267 -5410 2307 -5090
rect 2627 -5410 2667 -5090
rect 2267 -5450 2667 -5410
rect 2986 -5090 3386 -5050
rect 2986 -5410 3026 -5090
rect 3346 -5410 3386 -5090
rect 2986 -5450 3386 -5410
rect 3705 -5090 4105 -5050
rect 3705 -5410 3745 -5090
rect 4065 -5410 4105 -5090
rect 3705 -5450 4105 -5410
rect 4424 -5090 4824 -5050
rect 4424 -5410 4464 -5090
rect 4784 -5410 4824 -5090
rect 4424 -5450 4824 -5410
rect 5143 -5090 5543 -5050
rect 5143 -5410 5183 -5090
rect 5503 -5410 5543 -5090
rect 5143 -5450 5543 -5410
rect 5862 -5090 6262 -5050
rect 5862 -5410 5902 -5090
rect 6222 -5410 6262 -5090
rect 5862 -5450 6262 -5410
rect 6581 -5090 6981 -5050
rect 6581 -5410 6621 -5090
rect 6941 -5410 6981 -5090
rect 6581 -5450 6981 -5410
rect -7080 -5790 -6680 -5750
rect -7080 -6110 -7040 -5790
rect -6720 -6110 -6680 -5790
rect -7080 -6150 -6680 -6110
rect -6361 -5790 -5961 -5750
rect -6361 -6110 -6321 -5790
rect -6001 -6110 -5961 -5790
rect -6361 -6150 -5961 -6110
rect -5642 -5790 -5242 -5750
rect -5642 -6110 -5602 -5790
rect -5282 -6110 -5242 -5790
rect -5642 -6150 -5242 -6110
rect -4923 -5790 -4523 -5750
rect -4923 -6110 -4883 -5790
rect -4563 -6110 -4523 -5790
rect -4923 -6150 -4523 -6110
rect -4204 -5790 -3804 -5750
rect -4204 -6110 -4164 -5790
rect -3844 -6110 -3804 -5790
rect -4204 -6150 -3804 -6110
rect -3485 -5790 -3085 -5750
rect -3485 -6110 -3445 -5790
rect -3125 -6110 -3085 -5790
rect -3485 -6150 -3085 -6110
rect -2766 -5790 -2366 -5750
rect -2766 -6110 -2726 -5790
rect -2406 -6110 -2366 -5790
rect -2766 -6150 -2366 -6110
rect -2047 -5790 -1647 -5750
rect -2047 -6110 -2007 -5790
rect -1687 -6110 -1647 -5790
rect -2047 -6150 -1647 -6110
rect -1328 -5790 -928 -5750
rect -1328 -6110 -1288 -5790
rect -968 -6110 -928 -5790
rect -1328 -6150 -928 -6110
rect -609 -5790 -209 -5750
rect -609 -6110 -569 -5790
rect -249 -6110 -209 -5790
rect -609 -6150 -209 -6110
rect 110 -5790 510 -5750
rect 110 -6110 150 -5790
rect 470 -6110 510 -5790
rect 110 -6150 510 -6110
rect 829 -5790 1229 -5750
rect 829 -6110 869 -5790
rect 1189 -6110 1229 -5790
rect 829 -6150 1229 -6110
rect 1548 -5790 1948 -5750
rect 1548 -6110 1588 -5790
rect 1908 -6110 1948 -5790
rect 1548 -6150 1948 -6110
rect 2267 -5790 2667 -5750
rect 2267 -6110 2307 -5790
rect 2627 -6110 2667 -5790
rect 2267 -6150 2667 -6110
rect 2986 -5790 3386 -5750
rect 2986 -6110 3026 -5790
rect 3346 -6110 3386 -5790
rect 2986 -6150 3386 -6110
rect 3705 -5790 4105 -5750
rect 3705 -6110 3745 -5790
rect 4065 -6110 4105 -5790
rect 3705 -6150 4105 -6110
rect 4424 -5790 4824 -5750
rect 4424 -6110 4464 -5790
rect 4784 -6110 4824 -5790
rect 4424 -6150 4824 -6110
rect 5143 -5790 5543 -5750
rect 5143 -6110 5183 -5790
rect 5503 -6110 5543 -5790
rect 5143 -6150 5543 -6110
rect 5862 -5790 6262 -5750
rect 5862 -6110 5902 -5790
rect 6222 -6110 6262 -5790
rect 5862 -6150 6262 -6110
rect 6581 -5790 6981 -5750
rect 6581 -6110 6621 -5790
rect 6941 -6110 6981 -5790
rect 6581 -6150 6981 -6110
rect -7080 -6490 -6680 -6450
rect -7080 -6810 -7040 -6490
rect -6720 -6810 -6680 -6490
rect -7080 -6850 -6680 -6810
rect -6361 -6490 -5961 -6450
rect -6361 -6810 -6321 -6490
rect -6001 -6810 -5961 -6490
rect -6361 -6850 -5961 -6810
rect -5642 -6490 -5242 -6450
rect -5642 -6810 -5602 -6490
rect -5282 -6810 -5242 -6490
rect -5642 -6850 -5242 -6810
rect -4923 -6490 -4523 -6450
rect -4923 -6810 -4883 -6490
rect -4563 -6810 -4523 -6490
rect -4923 -6850 -4523 -6810
rect -4204 -6490 -3804 -6450
rect -4204 -6810 -4164 -6490
rect -3844 -6810 -3804 -6490
rect -4204 -6850 -3804 -6810
rect -3485 -6490 -3085 -6450
rect -3485 -6810 -3445 -6490
rect -3125 -6810 -3085 -6490
rect -3485 -6850 -3085 -6810
rect -2766 -6490 -2366 -6450
rect -2766 -6810 -2726 -6490
rect -2406 -6810 -2366 -6490
rect -2766 -6850 -2366 -6810
rect -2047 -6490 -1647 -6450
rect -2047 -6810 -2007 -6490
rect -1687 -6810 -1647 -6490
rect -2047 -6850 -1647 -6810
rect -1328 -6490 -928 -6450
rect -1328 -6810 -1288 -6490
rect -968 -6810 -928 -6490
rect -1328 -6850 -928 -6810
rect -609 -6490 -209 -6450
rect -609 -6810 -569 -6490
rect -249 -6810 -209 -6490
rect -609 -6850 -209 -6810
rect 110 -6490 510 -6450
rect 110 -6810 150 -6490
rect 470 -6810 510 -6490
rect 110 -6850 510 -6810
rect 829 -6490 1229 -6450
rect 829 -6810 869 -6490
rect 1189 -6810 1229 -6490
rect 829 -6850 1229 -6810
rect 1548 -6490 1948 -6450
rect 1548 -6810 1588 -6490
rect 1908 -6810 1948 -6490
rect 1548 -6850 1948 -6810
rect 2267 -6490 2667 -6450
rect 2267 -6810 2307 -6490
rect 2627 -6810 2667 -6490
rect 2267 -6850 2667 -6810
rect 2986 -6490 3386 -6450
rect 2986 -6810 3026 -6490
rect 3346 -6810 3386 -6490
rect 2986 -6850 3386 -6810
rect 3705 -6490 4105 -6450
rect 3705 -6810 3745 -6490
rect 4065 -6810 4105 -6490
rect 3705 -6850 4105 -6810
rect 4424 -6490 4824 -6450
rect 4424 -6810 4464 -6490
rect 4784 -6810 4824 -6490
rect 4424 -6850 4824 -6810
rect 5143 -6490 5543 -6450
rect 5143 -6810 5183 -6490
rect 5503 -6810 5543 -6490
rect 5143 -6850 5543 -6810
rect 5862 -6490 6262 -6450
rect 5862 -6810 5902 -6490
rect 6222 -6810 6262 -6490
rect 5862 -6850 6262 -6810
rect 6581 -6490 6981 -6450
rect 6581 -6810 6621 -6490
rect 6941 -6810 6981 -6490
rect 6581 -6850 6981 -6810
<< mimcapcontact >>
rect -7040 6490 -6720 6810
rect -6321 6490 -6001 6810
rect -5602 6490 -5282 6810
rect -4883 6490 -4563 6810
rect -4164 6490 -3844 6810
rect -3445 6490 -3125 6810
rect -2726 6490 -2406 6810
rect -2007 6490 -1687 6810
rect -1288 6490 -968 6810
rect -569 6490 -249 6810
rect 150 6490 470 6810
rect 869 6490 1189 6810
rect 1588 6490 1908 6810
rect 2307 6490 2627 6810
rect 3026 6490 3346 6810
rect 3745 6490 4065 6810
rect 4464 6490 4784 6810
rect 5183 6490 5503 6810
rect 5902 6490 6222 6810
rect 6621 6490 6941 6810
rect -7040 5790 -6720 6110
rect -6321 5790 -6001 6110
rect -5602 5790 -5282 6110
rect -4883 5790 -4563 6110
rect -4164 5790 -3844 6110
rect -3445 5790 -3125 6110
rect -2726 5790 -2406 6110
rect -2007 5790 -1687 6110
rect -1288 5790 -968 6110
rect -569 5790 -249 6110
rect 150 5790 470 6110
rect 869 5790 1189 6110
rect 1588 5790 1908 6110
rect 2307 5790 2627 6110
rect 3026 5790 3346 6110
rect 3745 5790 4065 6110
rect 4464 5790 4784 6110
rect 5183 5790 5503 6110
rect 5902 5790 6222 6110
rect 6621 5790 6941 6110
rect -7040 5090 -6720 5410
rect -6321 5090 -6001 5410
rect -5602 5090 -5282 5410
rect -4883 5090 -4563 5410
rect -4164 5090 -3844 5410
rect -3445 5090 -3125 5410
rect -2726 5090 -2406 5410
rect -2007 5090 -1687 5410
rect -1288 5090 -968 5410
rect -569 5090 -249 5410
rect 150 5090 470 5410
rect 869 5090 1189 5410
rect 1588 5090 1908 5410
rect 2307 5090 2627 5410
rect 3026 5090 3346 5410
rect 3745 5090 4065 5410
rect 4464 5090 4784 5410
rect 5183 5090 5503 5410
rect 5902 5090 6222 5410
rect 6621 5090 6941 5410
rect -7040 4390 -6720 4710
rect -6321 4390 -6001 4710
rect -5602 4390 -5282 4710
rect -4883 4390 -4563 4710
rect -4164 4390 -3844 4710
rect -3445 4390 -3125 4710
rect -2726 4390 -2406 4710
rect -2007 4390 -1687 4710
rect -1288 4390 -968 4710
rect -569 4390 -249 4710
rect 150 4390 470 4710
rect 869 4390 1189 4710
rect 1588 4390 1908 4710
rect 2307 4390 2627 4710
rect 3026 4390 3346 4710
rect 3745 4390 4065 4710
rect 4464 4390 4784 4710
rect 5183 4390 5503 4710
rect 5902 4390 6222 4710
rect 6621 4390 6941 4710
rect -7040 3690 -6720 4010
rect -6321 3690 -6001 4010
rect -5602 3690 -5282 4010
rect -4883 3690 -4563 4010
rect -4164 3690 -3844 4010
rect -3445 3690 -3125 4010
rect -2726 3690 -2406 4010
rect -2007 3690 -1687 4010
rect -1288 3690 -968 4010
rect -569 3690 -249 4010
rect 150 3690 470 4010
rect 869 3690 1189 4010
rect 1588 3690 1908 4010
rect 2307 3690 2627 4010
rect 3026 3690 3346 4010
rect 3745 3690 4065 4010
rect 4464 3690 4784 4010
rect 5183 3690 5503 4010
rect 5902 3690 6222 4010
rect 6621 3690 6941 4010
rect -7040 2990 -6720 3310
rect -6321 2990 -6001 3310
rect -5602 2990 -5282 3310
rect -4883 2990 -4563 3310
rect -4164 2990 -3844 3310
rect -3445 2990 -3125 3310
rect -2726 2990 -2406 3310
rect -2007 2990 -1687 3310
rect -1288 2990 -968 3310
rect -569 2990 -249 3310
rect 150 2990 470 3310
rect 869 2990 1189 3310
rect 1588 2990 1908 3310
rect 2307 2990 2627 3310
rect 3026 2990 3346 3310
rect 3745 2990 4065 3310
rect 4464 2990 4784 3310
rect 5183 2990 5503 3310
rect 5902 2990 6222 3310
rect 6621 2990 6941 3310
rect -7040 2290 -6720 2610
rect -6321 2290 -6001 2610
rect -5602 2290 -5282 2610
rect -4883 2290 -4563 2610
rect -4164 2290 -3844 2610
rect -3445 2290 -3125 2610
rect -2726 2290 -2406 2610
rect -2007 2290 -1687 2610
rect -1288 2290 -968 2610
rect -569 2290 -249 2610
rect 150 2290 470 2610
rect 869 2290 1189 2610
rect 1588 2290 1908 2610
rect 2307 2290 2627 2610
rect 3026 2290 3346 2610
rect 3745 2290 4065 2610
rect 4464 2290 4784 2610
rect 5183 2290 5503 2610
rect 5902 2290 6222 2610
rect 6621 2290 6941 2610
rect -7040 1590 -6720 1910
rect -6321 1590 -6001 1910
rect -5602 1590 -5282 1910
rect -4883 1590 -4563 1910
rect -4164 1590 -3844 1910
rect -3445 1590 -3125 1910
rect -2726 1590 -2406 1910
rect -2007 1590 -1687 1910
rect -1288 1590 -968 1910
rect -569 1590 -249 1910
rect 150 1590 470 1910
rect 869 1590 1189 1910
rect 1588 1590 1908 1910
rect 2307 1590 2627 1910
rect 3026 1590 3346 1910
rect 3745 1590 4065 1910
rect 4464 1590 4784 1910
rect 5183 1590 5503 1910
rect 5902 1590 6222 1910
rect 6621 1590 6941 1910
rect -7040 890 -6720 1210
rect -6321 890 -6001 1210
rect -5602 890 -5282 1210
rect -4883 890 -4563 1210
rect -4164 890 -3844 1210
rect -3445 890 -3125 1210
rect -2726 890 -2406 1210
rect -2007 890 -1687 1210
rect -1288 890 -968 1210
rect -569 890 -249 1210
rect 150 890 470 1210
rect 869 890 1189 1210
rect 1588 890 1908 1210
rect 2307 890 2627 1210
rect 3026 890 3346 1210
rect 3745 890 4065 1210
rect 4464 890 4784 1210
rect 5183 890 5503 1210
rect 5902 890 6222 1210
rect 6621 890 6941 1210
rect -7040 190 -6720 510
rect -6321 190 -6001 510
rect -5602 190 -5282 510
rect -4883 190 -4563 510
rect -4164 190 -3844 510
rect -3445 190 -3125 510
rect -2726 190 -2406 510
rect -2007 190 -1687 510
rect -1288 190 -968 510
rect -569 190 -249 510
rect 150 190 470 510
rect 869 190 1189 510
rect 1588 190 1908 510
rect 2307 190 2627 510
rect 3026 190 3346 510
rect 3745 190 4065 510
rect 4464 190 4784 510
rect 5183 190 5503 510
rect 5902 190 6222 510
rect 6621 190 6941 510
rect -7040 -510 -6720 -190
rect -6321 -510 -6001 -190
rect -5602 -510 -5282 -190
rect -4883 -510 -4563 -190
rect -4164 -510 -3844 -190
rect -3445 -510 -3125 -190
rect -2726 -510 -2406 -190
rect -2007 -510 -1687 -190
rect -1288 -510 -968 -190
rect -569 -510 -249 -190
rect 150 -510 470 -190
rect 869 -510 1189 -190
rect 1588 -510 1908 -190
rect 2307 -510 2627 -190
rect 3026 -510 3346 -190
rect 3745 -510 4065 -190
rect 4464 -510 4784 -190
rect 5183 -510 5503 -190
rect 5902 -510 6222 -190
rect 6621 -510 6941 -190
rect -7040 -1210 -6720 -890
rect -6321 -1210 -6001 -890
rect -5602 -1210 -5282 -890
rect -4883 -1210 -4563 -890
rect -4164 -1210 -3844 -890
rect -3445 -1210 -3125 -890
rect -2726 -1210 -2406 -890
rect -2007 -1210 -1687 -890
rect -1288 -1210 -968 -890
rect -569 -1210 -249 -890
rect 150 -1210 470 -890
rect 869 -1210 1189 -890
rect 1588 -1210 1908 -890
rect 2307 -1210 2627 -890
rect 3026 -1210 3346 -890
rect 3745 -1210 4065 -890
rect 4464 -1210 4784 -890
rect 5183 -1210 5503 -890
rect 5902 -1210 6222 -890
rect 6621 -1210 6941 -890
rect -7040 -1910 -6720 -1590
rect -6321 -1910 -6001 -1590
rect -5602 -1910 -5282 -1590
rect -4883 -1910 -4563 -1590
rect -4164 -1910 -3844 -1590
rect -3445 -1910 -3125 -1590
rect -2726 -1910 -2406 -1590
rect -2007 -1910 -1687 -1590
rect -1288 -1910 -968 -1590
rect -569 -1910 -249 -1590
rect 150 -1910 470 -1590
rect 869 -1910 1189 -1590
rect 1588 -1910 1908 -1590
rect 2307 -1910 2627 -1590
rect 3026 -1910 3346 -1590
rect 3745 -1910 4065 -1590
rect 4464 -1910 4784 -1590
rect 5183 -1910 5503 -1590
rect 5902 -1910 6222 -1590
rect 6621 -1910 6941 -1590
rect -7040 -2610 -6720 -2290
rect -6321 -2610 -6001 -2290
rect -5602 -2610 -5282 -2290
rect -4883 -2610 -4563 -2290
rect -4164 -2610 -3844 -2290
rect -3445 -2610 -3125 -2290
rect -2726 -2610 -2406 -2290
rect -2007 -2610 -1687 -2290
rect -1288 -2610 -968 -2290
rect -569 -2610 -249 -2290
rect 150 -2610 470 -2290
rect 869 -2610 1189 -2290
rect 1588 -2610 1908 -2290
rect 2307 -2610 2627 -2290
rect 3026 -2610 3346 -2290
rect 3745 -2610 4065 -2290
rect 4464 -2610 4784 -2290
rect 5183 -2610 5503 -2290
rect 5902 -2610 6222 -2290
rect 6621 -2610 6941 -2290
rect -7040 -3310 -6720 -2990
rect -6321 -3310 -6001 -2990
rect -5602 -3310 -5282 -2990
rect -4883 -3310 -4563 -2990
rect -4164 -3310 -3844 -2990
rect -3445 -3310 -3125 -2990
rect -2726 -3310 -2406 -2990
rect -2007 -3310 -1687 -2990
rect -1288 -3310 -968 -2990
rect -569 -3310 -249 -2990
rect 150 -3310 470 -2990
rect 869 -3310 1189 -2990
rect 1588 -3310 1908 -2990
rect 2307 -3310 2627 -2990
rect 3026 -3310 3346 -2990
rect 3745 -3310 4065 -2990
rect 4464 -3310 4784 -2990
rect 5183 -3310 5503 -2990
rect 5902 -3310 6222 -2990
rect 6621 -3310 6941 -2990
rect -7040 -4010 -6720 -3690
rect -6321 -4010 -6001 -3690
rect -5602 -4010 -5282 -3690
rect -4883 -4010 -4563 -3690
rect -4164 -4010 -3844 -3690
rect -3445 -4010 -3125 -3690
rect -2726 -4010 -2406 -3690
rect -2007 -4010 -1687 -3690
rect -1288 -4010 -968 -3690
rect -569 -4010 -249 -3690
rect 150 -4010 470 -3690
rect 869 -4010 1189 -3690
rect 1588 -4010 1908 -3690
rect 2307 -4010 2627 -3690
rect 3026 -4010 3346 -3690
rect 3745 -4010 4065 -3690
rect 4464 -4010 4784 -3690
rect 5183 -4010 5503 -3690
rect 5902 -4010 6222 -3690
rect 6621 -4010 6941 -3690
rect -7040 -4710 -6720 -4390
rect -6321 -4710 -6001 -4390
rect -5602 -4710 -5282 -4390
rect -4883 -4710 -4563 -4390
rect -4164 -4710 -3844 -4390
rect -3445 -4710 -3125 -4390
rect -2726 -4710 -2406 -4390
rect -2007 -4710 -1687 -4390
rect -1288 -4710 -968 -4390
rect -569 -4710 -249 -4390
rect 150 -4710 470 -4390
rect 869 -4710 1189 -4390
rect 1588 -4710 1908 -4390
rect 2307 -4710 2627 -4390
rect 3026 -4710 3346 -4390
rect 3745 -4710 4065 -4390
rect 4464 -4710 4784 -4390
rect 5183 -4710 5503 -4390
rect 5902 -4710 6222 -4390
rect 6621 -4710 6941 -4390
rect -7040 -5410 -6720 -5090
rect -6321 -5410 -6001 -5090
rect -5602 -5410 -5282 -5090
rect -4883 -5410 -4563 -5090
rect -4164 -5410 -3844 -5090
rect -3445 -5410 -3125 -5090
rect -2726 -5410 -2406 -5090
rect -2007 -5410 -1687 -5090
rect -1288 -5410 -968 -5090
rect -569 -5410 -249 -5090
rect 150 -5410 470 -5090
rect 869 -5410 1189 -5090
rect 1588 -5410 1908 -5090
rect 2307 -5410 2627 -5090
rect 3026 -5410 3346 -5090
rect 3745 -5410 4065 -5090
rect 4464 -5410 4784 -5090
rect 5183 -5410 5503 -5090
rect 5902 -5410 6222 -5090
rect 6621 -5410 6941 -5090
rect -7040 -6110 -6720 -5790
rect -6321 -6110 -6001 -5790
rect -5602 -6110 -5282 -5790
rect -4883 -6110 -4563 -5790
rect -4164 -6110 -3844 -5790
rect -3445 -6110 -3125 -5790
rect -2726 -6110 -2406 -5790
rect -2007 -6110 -1687 -5790
rect -1288 -6110 -968 -5790
rect -569 -6110 -249 -5790
rect 150 -6110 470 -5790
rect 869 -6110 1189 -5790
rect 1588 -6110 1908 -5790
rect 2307 -6110 2627 -5790
rect 3026 -6110 3346 -5790
rect 3745 -6110 4065 -5790
rect 4464 -6110 4784 -5790
rect 5183 -6110 5503 -5790
rect 5902 -6110 6222 -5790
rect 6621 -6110 6941 -5790
rect -7040 -6810 -6720 -6490
rect -6321 -6810 -6001 -6490
rect -5602 -6810 -5282 -6490
rect -4883 -6810 -4563 -6490
rect -4164 -6810 -3844 -6490
rect -3445 -6810 -3125 -6490
rect -2726 -6810 -2406 -6490
rect -2007 -6810 -1687 -6490
rect -1288 -6810 -968 -6490
rect -569 -6810 -249 -6490
rect 150 -6810 470 -6490
rect 869 -6810 1189 -6490
rect 1588 -6810 1908 -6490
rect 2307 -6810 2627 -6490
rect 3026 -6810 3346 -6490
rect 3745 -6810 4065 -6490
rect 4464 -6810 4784 -6490
rect 5183 -6810 5503 -6490
rect 5902 -6810 6222 -6490
rect 6621 -6810 6941 -6490
<< metal4 >>
rect -6932 6811 -6828 7000
rect -6612 6938 -6508 7000
rect -6612 6922 -6485 6938
rect -7041 6810 -6719 6811
rect -7041 6490 -7040 6810
rect -6720 6490 -6719 6810
rect -7041 6489 -6719 6490
rect -6932 6111 -6828 6489
rect -6612 6378 -6565 6922
rect -6501 6378 -6485 6922
rect -6213 6811 -6109 7000
rect -5893 6938 -5789 7000
rect -5893 6922 -5766 6938
rect -6322 6810 -6000 6811
rect -6322 6490 -6321 6810
rect -6001 6490 -6000 6810
rect -6322 6489 -6000 6490
rect -6612 6362 -6485 6378
rect -6612 6238 -6508 6362
rect -6612 6222 -6485 6238
rect -7041 6110 -6719 6111
rect -7041 5790 -7040 6110
rect -6720 5790 -6719 6110
rect -7041 5789 -6719 5790
rect -6932 5411 -6828 5789
rect -6612 5678 -6565 6222
rect -6501 5678 -6485 6222
rect -6213 6111 -6109 6489
rect -5893 6378 -5846 6922
rect -5782 6378 -5766 6922
rect -5494 6811 -5390 7000
rect -5174 6938 -5070 7000
rect -5174 6922 -5047 6938
rect -5603 6810 -5281 6811
rect -5603 6490 -5602 6810
rect -5282 6490 -5281 6810
rect -5603 6489 -5281 6490
rect -5893 6362 -5766 6378
rect -5893 6238 -5789 6362
rect -5893 6222 -5766 6238
rect -6322 6110 -6000 6111
rect -6322 5790 -6321 6110
rect -6001 5790 -6000 6110
rect -6322 5789 -6000 5790
rect -6612 5662 -6485 5678
rect -6612 5538 -6508 5662
rect -6612 5522 -6485 5538
rect -7041 5410 -6719 5411
rect -7041 5090 -7040 5410
rect -6720 5090 -6719 5410
rect -7041 5089 -6719 5090
rect -6932 4711 -6828 5089
rect -6612 4978 -6565 5522
rect -6501 4978 -6485 5522
rect -6213 5411 -6109 5789
rect -5893 5678 -5846 6222
rect -5782 5678 -5766 6222
rect -5494 6111 -5390 6489
rect -5174 6378 -5127 6922
rect -5063 6378 -5047 6922
rect -4775 6811 -4671 7000
rect -4455 6938 -4351 7000
rect -4455 6922 -4328 6938
rect -4884 6810 -4562 6811
rect -4884 6490 -4883 6810
rect -4563 6490 -4562 6810
rect -4884 6489 -4562 6490
rect -5174 6362 -5047 6378
rect -5174 6238 -5070 6362
rect -5174 6222 -5047 6238
rect -5603 6110 -5281 6111
rect -5603 5790 -5602 6110
rect -5282 5790 -5281 6110
rect -5603 5789 -5281 5790
rect -5893 5662 -5766 5678
rect -5893 5538 -5789 5662
rect -5893 5522 -5766 5538
rect -6322 5410 -6000 5411
rect -6322 5090 -6321 5410
rect -6001 5090 -6000 5410
rect -6322 5089 -6000 5090
rect -6612 4962 -6485 4978
rect -6612 4838 -6508 4962
rect -6612 4822 -6485 4838
rect -7041 4710 -6719 4711
rect -7041 4390 -7040 4710
rect -6720 4390 -6719 4710
rect -7041 4389 -6719 4390
rect -6932 4011 -6828 4389
rect -6612 4278 -6565 4822
rect -6501 4278 -6485 4822
rect -6213 4711 -6109 5089
rect -5893 4978 -5846 5522
rect -5782 4978 -5766 5522
rect -5494 5411 -5390 5789
rect -5174 5678 -5127 6222
rect -5063 5678 -5047 6222
rect -4775 6111 -4671 6489
rect -4455 6378 -4408 6922
rect -4344 6378 -4328 6922
rect -4056 6811 -3952 7000
rect -3736 6938 -3632 7000
rect -3736 6922 -3609 6938
rect -4165 6810 -3843 6811
rect -4165 6490 -4164 6810
rect -3844 6490 -3843 6810
rect -4165 6489 -3843 6490
rect -4455 6362 -4328 6378
rect -4455 6238 -4351 6362
rect -4455 6222 -4328 6238
rect -4884 6110 -4562 6111
rect -4884 5790 -4883 6110
rect -4563 5790 -4562 6110
rect -4884 5789 -4562 5790
rect -5174 5662 -5047 5678
rect -5174 5538 -5070 5662
rect -5174 5522 -5047 5538
rect -5603 5410 -5281 5411
rect -5603 5090 -5602 5410
rect -5282 5090 -5281 5410
rect -5603 5089 -5281 5090
rect -5893 4962 -5766 4978
rect -5893 4838 -5789 4962
rect -5893 4822 -5766 4838
rect -6322 4710 -6000 4711
rect -6322 4390 -6321 4710
rect -6001 4390 -6000 4710
rect -6322 4389 -6000 4390
rect -6612 4262 -6485 4278
rect -6612 4138 -6508 4262
rect -6612 4122 -6485 4138
rect -7041 4010 -6719 4011
rect -7041 3690 -7040 4010
rect -6720 3690 -6719 4010
rect -7041 3689 -6719 3690
rect -6932 3311 -6828 3689
rect -6612 3578 -6565 4122
rect -6501 3578 -6485 4122
rect -6213 4011 -6109 4389
rect -5893 4278 -5846 4822
rect -5782 4278 -5766 4822
rect -5494 4711 -5390 5089
rect -5174 4978 -5127 5522
rect -5063 4978 -5047 5522
rect -4775 5411 -4671 5789
rect -4455 5678 -4408 6222
rect -4344 5678 -4328 6222
rect -4056 6111 -3952 6489
rect -3736 6378 -3689 6922
rect -3625 6378 -3609 6922
rect -3337 6811 -3233 7000
rect -3017 6938 -2913 7000
rect -3017 6922 -2890 6938
rect -3446 6810 -3124 6811
rect -3446 6490 -3445 6810
rect -3125 6490 -3124 6810
rect -3446 6489 -3124 6490
rect -3736 6362 -3609 6378
rect -3736 6238 -3632 6362
rect -3736 6222 -3609 6238
rect -4165 6110 -3843 6111
rect -4165 5790 -4164 6110
rect -3844 5790 -3843 6110
rect -4165 5789 -3843 5790
rect -4455 5662 -4328 5678
rect -4455 5538 -4351 5662
rect -4455 5522 -4328 5538
rect -4884 5410 -4562 5411
rect -4884 5090 -4883 5410
rect -4563 5090 -4562 5410
rect -4884 5089 -4562 5090
rect -5174 4962 -5047 4978
rect -5174 4838 -5070 4962
rect -5174 4822 -5047 4838
rect -5603 4710 -5281 4711
rect -5603 4390 -5602 4710
rect -5282 4390 -5281 4710
rect -5603 4389 -5281 4390
rect -5893 4262 -5766 4278
rect -5893 4138 -5789 4262
rect -5893 4122 -5766 4138
rect -6322 4010 -6000 4011
rect -6322 3690 -6321 4010
rect -6001 3690 -6000 4010
rect -6322 3689 -6000 3690
rect -6612 3562 -6485 3578
rect -6612 3438 -6508 3562
rect -6612 3422 -6485 3438
rect -7041 3310 -6719 3311
rect -7041 2990 -7040 3310
rect -6720 2990 -6719 3310
rect -7041 2989 -6719 2990
rect -6932 2611 -6828 2989
rect -6612 2878 -6565 3422
rect -6501 2878 -6485 3422
rect -6213 3311 -6109 3689
rect -5893 3578 -5846 4122
rect -5782 3578 -5766 4122
rect -5494 4011 -5390 4389
rect -5174 4278 -5127 4822
rect -5063 4278 -5047 4822
rect -4775 4711 -4671 5089
rect -4455 4978 -4408 5522
rect -4344 4978 -4328 5522
rect -4056 5411 -3952 5789
rect -3736 5678 -3689 6222
rect -3625 5678 -3609 6222
rect -3337 6111 -3233 6489
rect -3017 6378 -2970 6922
rect -2906 6378 -2890 6922
rect -2618 6811 -2514 7000
rect -2298 6938 -2194 7000
rect -2298 6922 -2171 6938
rect -2727 6810 -2405 6811
rect -2727 6490 -2726 6810
rect -2406 6490 -2405 6810
rect -2727 6489 -2405 6490
rect -3017 6362 -2890 6378
rect -3017 6238 -2913 6362
rect -3017 6222 -2890 6238
rect -3446 6110 -3124 6111
rect -3446 5790 -3445 6110
rect -3125 5790 -3124 6110
rect -3446 5789 -3124 5790
rect -3736 5662 -3609 5678
rect -3736 5538 -3632 5662
rect -3736 5522 -3609 5538
rect -4165 5410 -3843 5411
rect -4165 5090 -4164 5410
rect -3844 5090 -3843 5410
rect -4165 5089 -3843 5090
rect -4455 4962 -4328 4978
rect -4455 4838 -4351 4962
rect -4455 4822 -4328 4838
rect -4884 4710 -4562 4711
rect -4884 4390 -4883 4710
rect -4563 4390 -4562 4710
rect -4884 4389 -4562 4390
rect -5174 4262 -5047 4278
rect -5174 4138 -5070 4262
rect -5174 4122 -5047 4138
rect -5603 4010 -5281 4011
rect -5603 3690 -5602 4010
rect -5282 3690 -5281 4010
rect -5603 3689 -5281 3690
rect -5893 3562 -5766 3578
rect -5893 3438 -5789 3562
rect -5893 3422 -5766 3438
rect -6322 3310 -6000 3311
rect -6322 2990 -6321 3310
rect -6001 2990 -6000 3310
rect -6322 2989 -6000 2990
rect -6612 2862 -6485 2878
rect -6612 2738 -6508 2862
rect -6612 2722 -6485 2738
rect -7041 2610 -6719 2611
rect -7041 2290 -7040 2610
rect -6720 2290 -6719 2610
rect -7041 2289 -6719 2290
rect -6932 1911 -6828 2289
rect -6612 2178 -6565 2722
rect -6501 2178 -6485 2722
rect -6213 2611 -6109 2989
rect -5893 2878 -5846 3422
rect -5782 2878 -5766 3422
rect -5494 3311 -5390 3689
rect -5174 3578 -5127 4122
rect -5063 3578 -5047 4122
rect -4775 4011 -4671 4389
rect -4455 4278 -4408 4822
rect -4344 4278 -4328 4822
rect -4056 4711 -3952 5089
rect -3736 4978 -3689 5522
rect -3625 4978 -3609 5522
rect -3337 5411 -3233 5789
rect -3017 5678 -2970 6222
rect -2906 5678 -2890 6222
rect -2618 6111 -2514 6489
rect -2298 6378 -2251 6922
rect -2187 6378 -2171 6922
rect -1899 6811 -1795 7000
rect -1579 6938 -1475 7000
rect -1579 6922 -1452 6938
rect -2008 6810 -1686 6811
rect -2008 6490 -2007 6810
rect -1687 6490 -1686 6810
rect -2008 6489 -1686 6490
rect -2298 6362 -2171 6378
rect -2298 6238 -2194 6362
rect -2298 6222 -2171 6238
rect -2727 6110 -2405 6111
rect -2727 5790 -2726 6110
rect -2406 5790 -2405 6110
rect -2727 5789 -2405 5790
rect -3017 5662 -2890 5678
rect -3017 5538 -2913 5662
rect -3017 5522 -2890 5538
rect -3446 5410 -3124 5411
rect -3446 5090 -3445 5410
rect -3125 5090 -3124 5410
rect -3446 5089 -3124 5090
rect -3736 4962 -3609 4978
rect -3736 4838 -3632 4962
rect -3736 4822 -3609 4838
rect -4165 4710 -3843 4711
rect -4165 4390 -4164 4710
rect -3844 4390 -3843 4710
rect -4165 4389 -3843 4390
rect -4455 4262 -4328 4278
rect -4455 4138 -4351 4262
rect -4455 4122 -4328 4138
rect -4884 4010 -4562 4011
rect -4884 3690 -4883 4010
rect -4563 3690 -4562 4010
rect -4884 3689 -4562 3690
rect -5174 3562 -5047 3578
rect -5174 3438 -5070 3562
rect -5174 3422 -5047 3438
rect -5603 3310 -5281 3311
rect -5603 2990 -5602 3310
rect -5282 2990 -5281 3310
rect -5603 2989 -5281 2990
rect -5893 2862 -5766 2878
rect -5893 2738 -5789 2862
rect -5893 2722 -5766 2738
rect -6322 2610 -6000 2611
rect -6322 2290 -6321 2610
rect -6001 2290 -6000 2610
rect -6322 2289 -6000 2290
rect -6612 2162 -6485 2178
rect -6612 2038 -6508 2162
rect -6612 2022 -6485 2038
rect -7041 1910 -6719 1911
rect -7041 1590 -7040 1910
rect -6720 1590 -6719 1910
rect -7041 1589 -6719 1590
rect -6932 1211 -6828 1589
rect -6612 1478 -6565 2022
rect -6501 1478 -6485 2022
rect -6213 1911 -6109 2289
rect -5893 2178 -5846 2722
rect -5782 2178 -5766 2722
rect -5494 2611 -5390 2989
rect -5174 2878 -5127 3422
rect -5063 2878 -5047 3422
rect -4775 3311 -4671 3689
rect -4455 3578 -4408 4122
rect -4344 3578 -4328 4122
rect -4056 4011 -3952 4389
rect -3736 4278 -3689 4822
rect -3625 4278 -3609 4822
rect -3337 4711 -3233 5089
rect -3017 4978 -2970 5522
rect -2906 4978 -2890 5522
rect -2618 5411 -2514 5789
rect -2298 5678 -2251 6222
rect -2187 5678 -2171 6222
rect -1899 6111 -1795 6489
rect -1579 6378 -1532 6922
rect -1468 6378 -1452 6922
rect -1180 6811 -1076 7000
rect -860 6938 -756 7000
rect -860 6922 -733 6938
rect -1289 6810 -967 6811
rect -1289 6490 -1288 6810
rect -968 6490 -967 6810
rect -1289 6489 -967 6490
rect -1579 6362 -1452 6378
rect -1579 6238 -1475 6362
rect -1579 6222 -1452 6238
rect -2008 6110 -1686 6111
rect -2008 5790 -2007 6110
rect -1687 5790 -1686 6110
rect -2008 5789 -1686 5790
rect -2298 5662 -2171 5678
rect -2298 5538 -2194 5662
rect -2298 5522 -2171 5538
rect -2727 5410 -2405 5411
rect -2727 5090 -2726 5410
rect -2406 5090 -2405 5410
rect -2727 5089 -2405 5090
rect -3017 4962 -2890 4978
rect -3017 4838 -2913 4962
rect -3017 4822 -2890 4838
rect -3446 4710 -3124 4711
rect -3446 4390 -3445 4710
rect -3125 4390 -3124 4710
rect -3446 4389 -3124 4390
rect -3736 4262 -3609 4278
rect -3736 4138 -3632 4262
rect -3736 4122 -3609 4138
rect -4165 4010 -3843 4011
rect -4165 3690 -4164 4010
rect -3844 3690 -3843 4010
rect -4165 3689 -3843 3690
rect -4455 3562 -4328 3578
rect -4455 3438 -4351 3562
rect -4455 3422 -4328 3438
rect -4884 3310 -4562 3311
rect -4884 2990 -4883 3310
rect -4563 2990 -4562 3310
rect -4884 2989 -4562 2990
rect -5174 2862 -5047 2878
rect -5174 2738 -5070 2862
rect -5174 2722 -5047 2738
rect -5603 2610 -5281 2611
rect -5603 2290 -5602 2610
rect -5282 2290 -5281 2610
rect -5603 2289 -5281 2290
rect -5893 2162 -5766 2178
rect -5893 2038 -5789 2162
rect -5893 2022 -5766 2038
rect -6322 1910 -6000 1911
rect -6322 1590 -6321 1910
rect -6001 1590 -6000 1910
rect -6322 1589 -6000 1590
rect -6612 1462 -6485 1478
rect -6612 1338 -6508 1462
rect -6612 1322 -6485 1338
rect -7041 1210 -6719 1211
rect -7041 890 -7040 1210
rect -6720 890 -6719 1210
rect -7041 889 -6719 890
rect -6932 511 -6828 889
rect -6612 778 -6565 1322
rect -6501 778 -6485 1322
rect -6213 1211 -6109 1589
rect -5893 1478 -5846 2022
rect -5782 1478 -5766 2022
rect -5494 1911 -5390 2289
rect -5174 2178 -5127 2722
rect -5063 2178 -5047 2722
rect -4775 2611 -4671 2989
rect -4455 2878 -4408 3422
rect -4344 2878 -4328 3422
rect -4056 3311 -3952 3689
rect -3736 3578 -3689 4122
rect -3625 3578 -3609 4122
rect -3337 4011 -3233 4389
rect -3017 4278 -2970 4822
rect -2906 4278 -2890 4822
rect -2618 4711 -2514 5089
rect -2298 4978 -2251 5522
rect -2187 4978 -2171 5522
rect -1899 5411 -1795 5789
rect -1579 5678 -1532 6222
rect -1468 5678 -1452 6222
rect -1180 6111 -1076 6489
rect -860 6378 -813 6922
rect -749 6378 -733 6922
rect -461 6811 -357 7000
rect -141 6938 -37 7000
rect -141 6922 -14 6938
rect -570 6810 -248 6811
rect -570 6490 -569 6810
rect -249 6490 -248 6810
rect -570 6489 -248 6490
rect -860 6362 -733 6378
rect -860 6238 -756 6362
rect -860 6222 -733 6238
rect -1289 6110 -967 6111
rect -1289 5790 -1288 6110
rect -968 5790 -967 6110
rect -1289 5789 -967 5790
rect -1579 5662 -1452 5678
rect -1579 5538 -1475 5662
rect -1579 5522 -1452 5538
rect -2008 5410 -1686 5411
rect -2008 5090 -2007 5410
rect -1687 5090 -1686 5410
rect -2008 5089 -1686 5090
rect -2298 4962 -2171 4978
rect -2298 4838 -2194 4962
rect -2298 4822 -2171 4838
rect -2727 4710 -2405 4711
rect -2727 4390 -2726 4710
rect -2406 4390 -2405 4710
rect -2727 4389 -2405 4390
rect -3017 4262 -2890 4278
rect -3017 4138 -2913 4262
rect -3017 4122 -2890 4138
rect -3446 4010 -3124 4011
rect -3446 3690 -3445 4010
rect -3125 3690 -3124 4010
rect -3446 3689 -3124 3690
rect -3736 3562 -3609 3578
rect -3736 3438 -3632 3562
rect -3736 3422 -3609 3438
rect -4165 3310 -3843 3311
rect -4165 2990 -4164 3310
rect -3844 2990 -3843 3310
rect -4165 2989 -3843 2990
rect -4455 2862 -4328 2878
rect -4455 2738 -4351 2862
rect -4455 2722 -4328 2738
rect -4884 2610 -4562 2611
rect -4884 2290 -4883 2610
rect -4563 2290 -4562 2610
rect -4884 2289 -4562 2290
rect -5174 2162 -5047 2178
rect -5174 2038 -5070 2162
rect -5174 2022 -5047 2038
rect -5603 1910 -5281 1911
rect -5603 1590 -5602 1910
rect -5282 1590 -5281 1910
rect -5603 1589 -5281 1590
rect -5893 1462 -5766 1478
rect -5893 1338 -5789 1462
rect -5893 1322 -5766 1338
rect -6322 1210 -6000 1211
rect -6322 890 -6321 1210
rect -6001 890 -6000 1210
rect -6322 889 -6000 890
rect -6612 762 -6485 778
rect -6612 638 -6508 762
rect -6612 622 -6485 638
rect -7041 510 -6719 511
rect -7041 190 -7040 510
rect -6720 190 -6719 510
rect -7041 189 -6719 190
rect -6932 -189 -6828 189
rect -6612 78 -6565 622
rect -6501 78 -6485 622
rect -6213 511 -6109 889
rect -5893 778 -5846 1322
rect -5782 778 -5766 1322
rect -5494 1211 -5390 1589
rect -5174 1478 -5127 2022
rect -5063 1478 -5047 2022
rect -4775 1911 -4671 2289
rect -4455 2178 -4408 2722
rect -4344 2178 -4328 2722
rect -4056 2611 -3952 2989
rect -3736 2878 -3689 3422
rect -3625 2878 -3609 3422
rect -3337 3311 -3233 3689
rect -3017 3578 -2970 4122
rect -2906 3578 -2890 4122
rect -2618 4011 -2514 4389
rect -2298 4278 -2251 4822
rect -2187 4278 -2171 4822
rect -1899 4711 -1795 5089
rect -1579 4978 -1532 5522
rect -1468 4978 -1452 5522
rect -1180 5411 -1076 5789
rect -860 5678 -813 6222
rect -749 5678 -733 6222
rect -461 6111 -357 6489
rect -141 6378 -94 6922
rect -30 6378 -14 6922
rect 258 6811 362 7000
rect 578 6938 682 7000
rect 578 6922 705 6938
rect 149 6810 471 6811
rect 149 6490 150 6810
rect 470 6490 471 6810
rect 149 6489 471 6490
rect -141 6362 -14 6378
rect -141 6238 -37 6362
rect -141 6222 -14 6238
rect -570 6110 -248 6111
rect -570 5790 -569 6110
rect -249 5790 -248 6110
rect -570 5789 -248 5790
rect -860 5662 -733 5678
rect -860 5538 -756 5662
rect -860 5522 -733 5538
rect -1289 5410 -967 5411
rect -1289 5090 -1288 5410
rect -968 5090 -967 5410
rect -1289 5089 -967 5090
rect -1579 4962 -1452 4978
rect -1579 4838 -1475 4962
rect -1579 4822 -1452 4838
rect -2008 4710 -1686 4711
rect -2008 4390 -2007 4710
rect -1687 4390 -1686 4710
rect -2008 4389 -1686 4390
rect -2298 4262 -2171 4278
rect -2298 4138 -2194 4262
rect -2298 4122 -2171 4138
rect -2727 4010 -2405 4011
rect -2727 3690 -2726 4010
rect -2406 3690 -2405 4010
rect -2727 3689 -2405 3690
rect -3017 3562 -2890 3578
rect -3017 3438 -2913 3562
rect -3017 3422 -2890 3438
rect -3446 3310 -3124 3311
rect -3446 2990 -3445 3310
rect -3125 2990 -3124 3310
rect -3446 2989 -3124 2990
rect -3736 2862 -3609 2878
rect -3736 2738 -3632 2862
rect -3736 2722 -3609 2738
rect -4165 2610 -3843 2611
rect -4165 2290 -4164 2610
rect -3844 2290 -3843 2610
rect -4165 2289 -3843 2290
rect -4455 2162 -4328 2178
rect -4455 2038 -4351 2162
rect -4455 2022 -4328 2038
rect -4884 1910 -4562 1911
rect -4884 1590 -4883 1910
rect -4563 1590 -4562 1910
rect -4884 1589 -4562 1590
rect -5174 1462 -5047 1478
rect -5174 1338 -5070 1462
rect -5174 1322 -5047 1338
rect -5603 1210 -5281 1211
rect -5603 890 -5602 1210
rect -5282 890 -5281 1210
rect -5603 889 -5281 890
rect -5893 762 -5766 778
rect -5893 638 -5789 762
rect -5893 622 -5766 638
rect -6322 510 -6000 511
rect -6322 190 -6321 510
rect -6001 190 -6000 510
rect -6322 189 -6000 190
rect -6612 62 -6485 78
rect -6612 -62 -6508 62
rect -6612 -78 -6485 -62
rect -7041 -190 -6719 -189
rect -7041 -510 -7040 -190
rect -6720 -510 -6719 -190
rect -7041 -511 -6719 -510
rect -6932 -889 -6828 -511
rect -6612 -622 -6565 -78
rect -6501 -622 -6485 -78
rect -6213 -189 -6109 189
rect -5893 78 -5846 622
rect -5782 78 -5766 622
rect -5494 511 -5390 889
rect -5174 778 -5127 1322
rect -5063 778 -5047 1322
rect -4775 1211 -4671 1589
rect -4455 1478 -4408 2022
rect -4344 1478 -4328 2022
rect -4056 1911 -3952 2289
rect -3736 2178 -3689 2722
rect -3625 2178 -3609 2722
rect -3337 2611 -3233 2989
rect -3017 2878 -2970 3422
rect -2906 2878 -2890 3422
rect -2618 3311 -2514 3689
rect -2298 3578 -2251 4122
rect -2187 3578 -2171 4122
rect -1899 4011 -1795 4389
rect -1579 4278 -1532 4822
rect -1468 4278 -1452 4822
rect -1180 4711 -1076 5089
rect -860 4978 -813 5522
rect -749 4978 -733 5522
rect -461 5411 -357 5789
rect -141 5678 -94 6222
rect -30 5678 -14 6222
rect 258 6111 362 6489
rect 578 6378 625 6922
rect 689 6378 705 6922
rect 977 6811 1081 7000
rect 1297 6938 1401 7000
rect 1297 6922 1424 6938
rect 868 6810 1190 6811
rect 868 6490 869 6810
rect 1189 6490 1190 6810
rect 868 6489 1190 6490
rect 578 6362 705 6378
rect 578 6238 682 6362
rect 578 6222 705 6238
rect 149 6110 471 6111
rect 149 5790 150 6110
rect 470 5790 471 6110
rect 149 5789 471 5790
rect -141 5662 -14 5678
rect -141 5538 -37 5662
rect -141 5522 -14 5538
rect -570 5410 -248 5411
rect -570 5090 -569 5410
rect -249 5090 -248 5410
rect -570 5089 -248 5090
rect -860 4962 -733 4978
rect -860 4838 -756 4962
rect -860 4822 -733 4838
rect -1289 4710 -967 4711
rect -1289 4390 -1288 4710
rect -968 4390 -967 4710
rect -1289 4389 -967 4390
rect -1579 4262 -1452 4278
rect -1579 4138 -1475 4262
rect -1579 4122 -1452 4138
rect -2008 4010 -1686 4011
rect -2008 3690 -2007 4010
rect -1687 3690 -1686 4010
rect -2008 3689 -1686 3690
rect -2298 3562 -2171 3578
rect -2298 3438 -2194 3562
rect -2298 3422 -2171 3438
rect -2727 3310 -2405 3311
rect -2727 2990 -2726 3310
rect -2406 2990 -2405 3310
rect -2727 2989 -2405 2990
rect -3017 2862 -2890 2878
rect -3017 2738 -2913 2862
rect -3017 2722 -2890 2738
rect -3446 2610 -3124 2611
rect -3446 2290 -3445 2610
rect -3125 2290 -3124 2610
rect -3446 2289 -3124 2290
rect -3736 2162 -3609 2178
rect -3736 2038 -3632 2162
rect -3736 2022 -3609 2038
rect -4165 1910 -3843 1911
rect -4165 1590 -4164 1910
rect -3844 1590 -3843 1910
rect -4165 1589 -3843 1590
rect -4455 1462 -4328 1478
rect -4455 1338 -4351 1462
rect -4455 1322 -4328 1338
rect -4884 1210 -4562 1211
rect -4884 890 -4883 1210
rect -4563 890 -4562 1210
rect -4884 889 -4562 890
rect -5174 762 -5047 778
rect -5174 638 -5070 762
rect -5174 622 -5047 638
rect -5603 510 -5281 511
rect -5603 190 -5602 510
rect -5282 190 -5281 510
rect -5603 189 -5281 190
rect -5893 62 -5766 78
rect -5893 -62 -5789 62
rect -5893 -78 -5766 -62
rect -6322 -190 -6000 -189
rect -6322 -510 -6321 -190
rect -6001 -510 -6000 -190
rect -6322 -511 -6000 -510
rect -6612 -638 -6485 -622
rect -6612 -762 -6508 -638
rect -6612 -778 -6485 -762
rect -7041 -890 -6719 -889
rect -7041 -1210 -7040 -890
rect -6720 -1210 -6719 -890
rect -7041 -1211 -6719 -1210
rect -6932 -1589 -6828 -1211
rect -6612 -1322 -6565 -778
rect -6501 -1322 -6485 -778
rect -6213 -889 -6109 -511
rect -5893 -622 -5846 -78
rect -5782 -622 -5766 -78
rect -5494 -189 -5390 189
rect -5174 78 -5127 622
rect -5063 78 -5047 622
rect -4775 511 -4671 889
rect -4455 778 -4408 1322
rect -4344 778 -4328 1322
rect -4056 1211 -3952 1589
rect -3736 1478 -3689 2022
rect -3625 1478 -3609 2022
rect -3337 1911 -3233 2289
rect -3017 2178 -2970 2722
rect -2906 2178 -2890 2722
rect -2618 2611 -2514 2989
rect -2298 2878 -2251 3422
rect -2187 2878 -2171 3422
rect -1899 3311 -1795 3689
rect -1579 3578 -1532 4122
rect -1468 3578 -1452 4122
rect -1180 4011 -1076 4389
rect -860 4278 -813 4822
rect -749 4278 -733 4822
rect -461 4711 -357 5089
rect -141 4978 -94 5522
rect -30 4978 -14 5522
rect 258 5411 362 5789
rect 578 5678 625 6222
rect 689 5678 705 6222
rect 977 6111 1081 6489
rect 1297 6378 1344 6922
rect 1408 6378 1424 6922
rect 1696 6811 1800 7000
rect 2016 6938 2120 7000
rect 2016 6922 2143 6938
rect 1587 6810 1909 6811
rect 1587 6490 1588 6810
rect 1908 6490 1909 6810
rect 1587 6489 1909 6490
rect 1297 6362 1424 6378
rect 1297 6238 1401 6362
rect 1297 6222 1424 6238
rect 868 6110 1190 6111
rect 868 5790 869 6110
rect 1189 5790 1190 6110
rect 868 5789 1190 5790
rect 578 5662 705 5678
rect 578 5538 682 5662
rect 578 5522 705 5538
rect 149 5410 471 5411
rect 149 5090 150 5410
rect 470 5090 471 5410
rect 149 5089 471 5090
rect -141 4962 -14 4978
rect -141 4838 -37 4962
rect -141 4822 -14 4838
rect -570 4710 -248 4711
rect -570 4390 -569 4710
rect -249 4390 -248 4710
rect -570 4389 -248 4390
rect -860 4262 -733 4278
rect -860 4138 -756 4262
rect -860 4122 -733 4138
rect -1289 4010 -967 4011
rect -1289 3690 -1288 4010
rect -968 3690 -967 4010
rect -1289 3689 -967 3690
rect -1579 3562 -1452 3578
rect -1579 3438 -1475 3562
rect -1579 3422 -1452 3438
rect -2008 3310 -1686 3311
rect -2008 2990 -2007 3310
rect -1687 2990 -1686 3310
rect -2008 2989 -1686 2990
rect -2298 2862 -2171 2878
rect -2298 2738 -2194 2862
rect -2298 2722 -2171 2738
rect -2727 2610 -2405 2611
rect -2727 2290 -2726 2610
rect -2406 2290 -2405 2610
rect -2727 2289 -2405 2290
rect -3017 2162 -2890 2178
rect -3017 2038 -2913 2162
rect -3017 2022 -2890 2038
rect -3446 1910 -3124 1911
rect -3446 1590 -3445 1910
rect -3125 1590 -3124 1910
rect -3446 1589 -3124 1590
rect -3736 1462 -3609 1478
rect -3736 1338 -3632 1462
rect -3736 1322 -3609 1338
rect -4165 1210 -3843 1211
rect -4165 890 -4164 1210
rect -3844 890 -3843 1210
rect -4165 889 -3843 890
rect -4455 762 -4328 778
rect -4455 638 -4351 762
rect -4455 622 -4328 638
rect -4884 510 -4562 511
rect -4884 190 -4883 510
rect -4563 190 -4562 510
rect -4884 189 -4562 190
rect -5174 62 -5047 78
rect -5174 -62 -5070 62
rect -5174 -78 -5047 -62
rect -5603 -190 -5281 -189
rect -5603 -510 -5602 -190
rect -5282 -510 -5281 -190
rect -5603 -511 -5281 -510
rect -5893 -638 -5766 -622
rect -5893 -762 -5789 -638
rect -5893 -778 -5766 -762
rect -6322 -890 -6000 -889
rect -6322 -1210 -6321 -890
rect -6001 -1210 -6000 -890
rect -6322 -1211 -6000 -1210
rect -6612 -1338 -6485 -1322
rect -6612 -1462 -6508 -1338
rect -6612 -1478 -6485 -1462
rect -7041 -1590 -6719 -1589
rect -7041 -1910 -7040 -1590
rect -6720 -1910 -6719 -1590
rect -7041 -1911 -6719 -1910
rect -6932 -2289 -6828 -1911
rect -6612 -2022 -6565 -1478
rect -6501 -2022 -6485 -1478
rect -6213 -1589 -6109 -1211
rect -5893 -1322 -5846 -778
rect -5782 -1322 -5766 -778
rect -5494 -889 -5390 -511
rect -5174 -622 -5127 -78
rect -5063 -622 -5047 -78
rect -4775 -189 -4671 189
rect -4455 78 -4408 622
rect -4344 78 -4328 622
rect -4056 511 -3952 889
rect -3736 778 -3689 1322
rect -3625 778 -3609 1322
rect -3337 1211 -3233 1589
rect -3017 1478 -2970 2022
rect -2906 1478 -2890 2022
rect -2618 1911 -2514 2289
rect -2298 2178 -2251 2722
rect -2187 2178 -2171 2722
rect -1899 2611 -1795 2989
rect -1579 2878 -1532 3422
rect -1468 2878 -1452 3422
rect -1180 3311 -1076 3689
rect -860 3578 -813 4122
rect -749 3578 -733 4122
rect -461 4011 -357 4389
rect -141 4278 -94 4822
rect -30 4278 -14 4822
rect 258 4711 362 5089
rect 578 4978 625 5522
rect 689 4978 705 5522
rect 977 5411 1081 5789
rect 1297 5678 1344 6222
rect 1408 5678 1424 6222
rect 1696 6111 1800 6489
rect 2016 6378 2063 6922
rect 2127 6378 2143 6922
rect 2415 6811 2519 7000
rect 2735 6938 2839 7000
rect 2735 6922 2862 6938
rect 2306 6810 2628 6811
rect 2306 6490 2307 6810
rect 2627 6490 2628 6810
rect 2306 6489 2628 6490
rect 2016 6362 2143 6378
rect 2016 6238 2120 6362
rect 2016 6222 2143 6238
rect 1587 6110 1909 6111
rect 1587 5790 1588 6110
rect 1908 5790 1909 6110
rect 1587 5789 1909 5790
rect 1297 5662 1424 5678
rect 1297 5538 1401 5662
rect 1297 5522 1424 5538
rect 868 5410 1190 5411
rect 868 5090 869 5410
rect 1189 5090 1190 5410
rect 868 5089 1190 5090
rect 578 4962 705 4978
rect 578 4838 682 4962
rect 578 4822 705 4838
rect 149 4710 471 4711
rect 149 4390 150 4710
rect 470 4390 471 4710
rect 149 4389 471 4390
rect -141 4262 -14 4278
rect -141 4138 -37 4262
rect -141 4122 -14 4138
rect -570 4010 -248 4011
rect -570 3690 -569 4010
rect -249 3690 -248 4010
rect -570 3689 -248 3690
rect -860 3562 -733 3578
rect -860 3438 -756 3562
rect -860 3422 -733 3438
rect -1289 3310 -967 3311
rect -1289 2990 -1288 3310
rect -968 2990 -967 3310
rect -1289 2989 -967 2990
rect -1579 2862 -1452 2878
rect -1579 2738 -1475 2862
rect -1579 2722 -1452 2738
rect -2008 2610 -1686 2611
rect -2008 2290 -2007 2610
rect -1687 2290 -1686 2610
rect -2008 2289 -1686 2290
rect -2298 2162 -2171 2178
rect -2298 2038 -2194 2162
rect -2298 2022 -2171 2038
rect -2727 1910 -2405 1911
rect -2727 1590 -2726 1910
rect -2406 1590 -2405 1910
rect -2727 1589 -2405 1590
rect -3017 1462 -2890 1478
rect -3017 1338 -2913 1462
rect -3017 1322 -2890 1338
rect -3446 1210 -3124 1211
rect -3446 890 -3445 1210
rect -3125 890 -3124 1210
rect -3446 889 -3124 890
rect -3736 762 -3609 778
rect -3736 638 -3632 762
rect -3736 622 -3609 638
rect -4165 510 -3843 511
rect -4165 190 -4164 510
rect -3844 190 -3843 510
rect -4165 189 -3843 190
rect -4455 62 -4328 78
rect -4455 -62 -4351 62
rect -4455 -78 -4328 -62
rect -4884 -190 -4562 -189
rect -4884 -510 -4883 -190
rect -4563 -510 -4562 -190
rect -4884 -511 -4562 -510
rect -5174 -638 -5047 -622
rect -5174 -762 -5070 -638
rect -5174 -778 -5047 -762
rect -5603 -890 -5281 -889
rect -5603 -1210 -5602 -890
rect -5282 -1210 -5281 -890
rect -5603 -1211 -5281 -1210
rect -5893 -1338 -5766 -1322
rect -5893 -1462 -5789 -1338
rect -5893 -1478 -5766 -1462
rect -6322 -1590 -6000 -1589
rect -6322 -1910 -6321 -1590
rect -6001 -1910 -6000 -1590
rect -6322 -1911 -6000 -1910
rect -6612 -2038 -6485 -2022
rect -6612 -2162 -6508 -2038
rect -6612 -2178 -6485 -2162
rect -7041 -2290 -6719 -2289
rect -7041 -2610 -7040 -2290
rect -6720 -2610 -6719 -2290
rect -7041 -2611 -6719 -2610
rect -6932 -2989 -6828 -2611
rect -6612 -2722 -6565 -2178
rect -6501 -2722 -6485 -2178
rect -6213 -2289 -6109 -1911
rect -5893 -2022 -5846 -1478
rect -5782 -2022 -5766 -1478
rect -5494 -1589 -5390 -1211
rect -5174 -1322 -5127 -778
rect -5063 -1322 -5047 -778
rect -4775 -889 -4671 -511
rect -4455 -622 -4408 -78
rect -4344 -622 -4328 -78
rect -4056 -189 -3952 189
rect -3736 78 -3689 622
rect -3625 78 -3609 622
rect -3337 511 -3233 889
rect -3017 778 -2970 1322
rect -2906 778 -2890 1322
rect -2618 1211 -2514 1589
rect -2298 1478 -2251 2022
rect -2187 1478 -2171 2022
rect -1899 1911 -1795 2289
rect -1579 2178 -1532 2722
rect -1468 2178 -1452 2722
rect -1180 2611 -1076 2989
rect -860 2878 -813 3422
rect -749 2878 -733 3422
rect -461 3311 -357 3689
rect -141 3578 -94 4122
rect -30 3578 -14 4122
rect 258 4011 362 4389
rect 578 4278 625 4822
rect 689 4278 705 4822
rect 977 4711 1081 5089
rect 1297 4978 1344 5522
rect 1408 4978 1424 5522
rect 1696 5411 1800 5789
rect 2016 5678 2063 6222
rect 2127 5678 2143 6222
rect 2415 6111 2519 6489
rect 2735 6378 2782 6922
rect 2846 6378 2862 6922
rect 3134 6811 3238 7000
rect 3454 6938 3558 7000
rect 3454 6922 3581 6938
rect 3025 6810 3347 6811
rect 3025 6490 3026 6810
rect 3346 6490 3347 6810
rect 3025 6489 3347 6490
rect 2735 6362 2862 6378
rect 2735 6238 2839 6362
rect 2735 6222 2862 6238
rect 2306 6110 2628 6111
rect 2306 5790 2307 6110
rect 2627 5790 2628 6110
rect 2306 5789 2628 5790
rect 2016 5662 2143 5678
rect 2016 5538 2120 5662
rect 2016 5522 2143 5538
rect 1587 5410 1909 5411
rect 1587 5090 1588 5410
rect 1908 5090 1909 5410
rect 1587 5089 1909 5090
rect 1297 4962 1424 4978
rect 1297 4838 1401 4962
rect 1297 4822 1424 4838
rect 868 4710 1190 4711
rect 868 4390 869 4710
rect 1189 4390 1190 4710
rect 868 4389 1190 4390
rect 578 4262 705 4278
rect 578 4138 682 4262
rect 578 4122 705 4138
rect 149 4010 471 4011
rect 149 3690 150 4010
rect 470 3690 471 4010
rect 149 3689 471 3690
rect -141 3562 -14 3578
rect -141 3438 -37 3562
rect -141 3422 -14 3438
rect -570 3310 -248 3311
rect -570 2990 -569 3310
rect -249 2990 -248 3310
rect -570 2989 -248 2990
rect -860 2862 -733 2878
rect -860 2738 -756 2862
rect -860 2722 -733 2738
rect -1289 2610 -967 2611
rect -1289 2290 -1288 2610
rect -968 2290 -967 2610
rect -1289 2289 -967 2290
rect -1579 2162 -1452 2178
rect -1579 2038 -1475 2162
rect -1579 2022 -1452 2038
rect -2008 1910 -1686 1911
rect -2008 1590 -2007 1910
rect -1687 1590 -1686 1910
rect -2008 1589 -1686 1590
rect -2298 1462 -2171 1478
rect -2298 1338 -2194 1462
rect -2298 1322 -2171 1338
rect -2727 1210 -2405 1211
rect -2727 890 -2726 1210
rect -2406 890 -2405 1210
rect -2727 889 -2405 890
rect -3017 762 -2890 778
rect -3017 638 -2913 762
rect -3017 622 -2890 638
rect -3446 510 -3124 511
rect -3446 190 -3445 510
rect -3125 190 -3124 510
rect -3446 189 -3124 190
rect -3736 62 -3609 78
rect -3736 -62 -3632 62
rect -3736 -78 -3609 -62
rect -4165 -190 -3843 -189
rect -4165 -510 -4164 -190
rect -3844 -510 -3843 -190
rect -4165 -511 -3843 -510
rect -4455 -638 -4328 -622
rect -4455 -762 -4351 -638
rect -4455 -778 -4328 -762
rect -4884 -890 -4562 -889
rect -4884 -1210 -4883 -890
rect -4563 -1210 -4562 -890
rect -4884 -1211 -4562 -1210
rect -5174 -1338 -5047 -1322
rect -5174 -1462 -5070 -1338
rect -5174 -1478 -5047 -1462
rect -5603 -1590 -5281 -1589
rect -5603 -1910 -5602 -1590
rect -5282 -1910 -5281 -1590
rect -5603 -1911 -5281 -1910
rect -5893 -2038 -5766 -2022
rect -5893 -2162 -5789 -2038
rect -5893 -2178 -5766 -2162
rect -6322 -2290 -6000 -2289
rect -6322 -2610 -6321 -2290
rect -6001 -2610 -6000 -2290
rect -6322 -2611 -6000 -2610
rect -6612 -2738 -6485 -2722
rect -6612 -2862 -6508 -2738
rect -6612 -2878 -6485 -2862
rect -7041 -2990 -6719 -2989
rect -7041 -3310 -7040 -2990
rect -6720 -3310 -6719 -2990
rect -7041 -3311 -6719 -3310
rect -6932 -3689 -6828 -3311
rect -6612 -3422 -6565 -2878
rect -6501 -3422 -6485 -2878
rect -6213 -2989 -6109 -2611
rect -5893 -2722 -5846 -2178
rect -5782 -2722 -5766 -2178
rect -5494 -2289 -5390 -1911
rect -5174 -2022 -5127 -1478
rect -5063 -2022 -5047 -1478
rect -4775 -1589 -4671 -1211
rect -4455 -1322 -4408 -778
rect -4344 -1322 -4328 -778
rect -4056 -889 -3952 -511
rect -3736 -622 -3689 -78
rect -3625 -622 -3609 -78
rect -3337 -189 -3233 189
rect -3017 78 -2970 622
rect -2906 78 -2890 622
rect -2618 511 -2514 889
rect -2298 778 -2251 1322
rect -2187 778 -2171 1322
rect -1899 1211 -1795 1589
rect -1579 1478 -1532 2022
rect -1468 1478 -1452 2022
rect -1180 1911 -1076 2289
rect -860 2178 -813 2722
rect -749 2178 -733 2722
rect -461 2611 -357 2989
rect -141 2878 -94 3422
rect -30 2878 -14 3422
rect 258 3311 362 3689
rect 578 3578 625 4122
rect 689 3578 705 4122
rect 977 4011 1081 4389
rect 1297 4278 1344 4822
rect 1408 4278 1424 4822
rect 1696 4711 1800 5089
rect 2016 4978 2063 5522
rect 2127 4978 2143 5522
rect 2415 5411 2519 5789
rect 2735 5678 2782 6222
rect 2846 5678 2862 6222
rect 3134 6111 3238 6489
rect 3454 6378 3501 6922
rect 3565 6378 3581 6922
rect 3853 6811 3957 7000
rect 4173 6938 4277 7000
rect 4173 6922 4300 6938
rect 3744 6810 4066 6811
rect 3744 6490 3745 6810
rect 4065 6490 4066 6810
rect 3744 6489 4066 6490
rect 3454 6362 3581 6378
rect 3454 6238 3558 6362
rect 3454 6222 3581 6238
rect 3025 6110 3347 6111
rect 3025 5790 3026 6110
rect 3346 5790 3347 6110
rect 3025 5789 3347 5790
rect 2735 5662 2862 5678
rect 2735 5538 2839 5662
rect 2735 5522 2862 5538
rect 2306 5410 2628 5411
rect 2306 5090 2307 5410
rect 2627 5090 2628 5410
rect 2306 5089 2628 5090
rect 2016 4962 2143 4978
rect 2016 4838 2120 4962
rect 2016 4822 2143 4838
rect 1587 4710 1909 4711
rect 1587 4390 1588 4710
rect 1908 4390 1909 4710
rect 1587 4389 1909 4390
rect 1297 4262 1424 4278
rect 1297 4138 1401 4262
rect 1297 4122 1424 4138
rect 868 4010 1190 4011
rect 868 3690 869 4010
rect 1189 3690 1190 4010
rect 868 3689 1190 3690
rect 578 3562 705 3578
rect 578 3438 682 3562
rect 578 3422 705 3438
rect 149 3310 471 3311
rect 149 2990 150 3310
rect 470 2990 471 3310
rect 149 2989 471 2990
rect -141 2862 -14 2878
rect -141 2738 -37 2862
rect -141 2722 -14 2738
rect -570 2610 -248 2611
rect -570 2290 -569 2610
rect -249 2290 -248 2610
rect -570 2289 -248 2290
rect -860 2162 -733 2178
rect -860 2038 -756 2162
rect -860 2022 -733 2038
rect -1289 1910 -967 1911
rect -1289 1590 -1288 1910
rect -968 1590 -967 1910
rect -1289 1589 -967 1590
rect -1579 1462 -1452 1478
rect -1579 1338 -1475 1462
rect -1579 1322 -1452 1338
rect -2008 1210 -1686 1211
rect -2008 890 -2007 1210
rect -1687 890 -1686 1210
rect -2008 889 -1686 890
rect -2298 762 -2171 778
rect -2298 638 -2194 762
rect -2298 622 -2171 638
rect -2727 510 -2405 511
rect -2727 190 -2726 510
rect -2406 190 -2405 510
rect -2727 189 -2405 190
rect -3017 62 -2890 78
rect -3017 -62 -2913 62
rect -3017 -78 -2890 -62
rect -3446 -190 -3124 -189
rect -3446 -510 -3445 -190
rect -3125 -510 -3124 -190
rect -3446 -511 -3124 -510
rect -3736 -638 -3609 -622
rect -3736 -762 -3632 -638
rect -3736 -778 -3609 -762
rect -4165 -890 -3843 -889
rect -4165 -1210 -4164 -890
rect -3844 -1210 -3843 -890
rect -4165 -1211 -3843 -1210
rect -4455 -1338 -4328 -1322
rect -4455 -1462 -4351 -1338
rect -4455 -1478 -4328 -1462
rect -4884 -1590 -4562 -1589
rect -4884 -1910 -4883 -1590
rect -4563 -1910 -4562 -1590
rect -4884 -1911 -4562 -1910
rect -5174 -2038 -5047 -2022
rect -5174 -2162 -5070 -2038
rect -5174 -2178 -5047 -2162
rect -5603 -2290 -5281 -2289
rect -5603 -2610 -5602 -2290
rect -5282 -2610 -5281 -2290
rect -5603 -2611 -5281 -2610
rect -5893 -2738 -5766 -2722
rect -5893 -2862 -5789 -2738
rect -5893 -2878 -5766 -2862
rect -6322 -2990 -6000 -2989
rect -6322 -3310 -6321 -2990
rect -6001 -3310 -6000 -2990
rect -6322 -3311 -6000 -3310
rect -6612 -3438 -6485 -3422
rect -6612 -3562 -6508 -3438
rect -6612 -3578 -6485 -3562
rect -7041 -3690 -6719 -3689
rect -7041 -4010 -7040 -3690
rect -6720 -4010 -6719 -3690
rect -7041 -4011 -6719 -4010
rect -6932 -4389 -6828 -4011
rect -6612 -4122 -6565 -3578
rect -6501 -4122 -6485 -3578
rect -6213 -3689 -6109 -3311
rect -5893 -3422 -5846 -2878
rect -5782 -3422 -5766 -2878
rect -5494 -2989 -5390 -2611
rect -5174 -2722 -5127 -2178
rect -5063 -2722 -5047 -2178
rect -4775 -2289 -4671 -1911
rect -4455 -2022 -4408 -1478
rect -4344 -2022 -4328 -1478
rect -4056 -1589 -3952 -1211
rect -3736 -1322 -3689 -778
rect -3625 -1322 -3609 -778
rect -3337 -889 -3233 -511
rect -3017 -622 -2970 -78
rect -2906 -622 -2890 -78
rect -2618 -189 -2514 189
rect -2298 78 -2251 622
rect -2187 78 -2171 622
rect -1899 511 -1795 889
rect -1579 778 -1532 1322
rect -1468 778 -1452 1322
rect -1180 1211 -1076 1589
rect -860 1478 -813 2022
rect -749 1478 -733 2022
rect -461 1911 -357 2289
rect -141 2178 -94 2722
rect -30 2178 -14 2722
rect 258 2611 362 2989
rect 578 2878 625 3422
rect 689 2878 705 3422
rect 977 3311 1081 3689
rect 1297 3578 1344 4122
rect 1408 3578 1424 4122
rect 1696 4011 1800 4389
rect 2016 4278 2063 4822
rect 2127 4278 2143 4822
rect 2415 4711 2519 5089
rect 2735 4978 2782 5522
rect 2846 4978 2862 5522
rect 3134 5411 3238 5789
rect 3454 5678 3501 6222
rect 3565 5678 3581 6222
rect 3853 6111 3957 6489
rect 4173 6378 4220 6922
rect 4284 6378 4300 6922
rect 4572 6811 4676 7000
rect 4892 6938 4996 7000
rect 4892 6922 5019 6938
rect 4463 6810 4785 6811
rect 4463 6490 4464 6810
rect 4784 6490 4785 6810
rect 4463 6489 4785 6490
rect 4173 6362 4300 6378
rect 4173 6238 4277 6362
rect 4173 6222 4300 6238
rect 3744 6110 4066 6111
rect 3744 5790 3745 6110
rect 4065 5790 4066 6110
rect 3744 5789 4066 5790
rect 3454 5662 3581 5678
rect 3454 5538 3558 5662
rect 3454 5522 3581 5538
rect 3025 5410 3347 5411
rect 3025 5090 3026 5410
rect 3346 5090 3347 5410
rect 3025 5089 3347 5090
rect 2735 4962 2862 4978
rect 2735 4838 2839 4962
rect 2735 4822 2862 4838
rect 2306 4710 2628 4711
rect 2306 4390 2307 4710
rect 2627 4390 2628 4710
rect 2306 4389 2628 4390
rect 2016 4262 2143 4278
rect 2016 4138 2120 4262
rect 2016 4122 2143 4138
rect 1587 4010 1909 4011
rect 1587 3690 1588 4010
rect 1908 3690 1909 4010
rect 1587 3689 1909 3690
rect 1297 3562 1424 3578
rect 1297 3438 1401 3562
rect 1297 3422 1424 3438
rect 868 3310 1190 3311
rect 868 2990 869 3310
rect 1189 2990 1190 3310
rect 868 2989 1190 2990
rect 578 2862 705 2878
rect 578 2738 682 2862
rect 578 2722 705 2738
rect 149 2610 471 2611
rect 149 2290 150 2610
rect 470 2290 471 2610
rect 149 2289 471 2290
rect -141 2162 -14 2178
rect -141 2038 -37 2162
rect -141 2022 -14 2038
rect -570 1910 -248 1911
rect -570 1590 -569 1910
rect -249 1590 -248 1910
rect -570 1589 -248 1590
rect -860 1462 -733 1478
rect -860 1338 -756 1462
rect -860 1322 -733 1338
rect -1289 1210 -967 1211
rect -1289 890 -1288 1210
rect -968 890 -967 1210
rect -1289 889 -967 890
rect -1579 762 -1452 778
rect -1579 638 -1475 762
rect -1579 622 -1452 638
rect -2008 510 -1686 511
rect -2008 190 -2007 510
rect -1687 190 -1686 510
rect -2008 189 -1686 190
rect -2298 62 -2171 78
rect -2298 -62 -2194 62
rect -2298 -78 -2171 -62
rect -2727 -190 -2405 -189
rect -2727 -510 -2726 -190
rect -2406 -510 -2405 -190
rect -2727 -511 -2405 -510
rect -3017 -638 -2890 -622
rect -3017 -762 -2913 -638
rect -3017 -778 -2890 -762
rect -3446 -890 -3124 -889
rect -3446 -1210 -3445 -890
rect -3125 -1210 -3124 -890
rect -3446 -1211 -3124 -1210
rect -3736 -1338 -3609 -1322
rect -3736 -1462 -3632 -1338
rect -3736 -1478 -3609 -1462
rect -4165 -1590 -3843 -1589
rect -4165 -1910 -4164 -1590
rect -3844 -1910 -3843 -1590
rect -4165 -1911 -3843 -1910
rect -4455 -2038 -4328 -2022
rect -4455 -2162 -4351 -2038
rect -4455 -2178 -4328 -2162
rect -4884 -2290 -4562 -2289
rect -4884 -2610 -4883 -2290
rect -4563 -2610 -4562 -2290
rect -4884 -2611 -4562 -2610
rect -5174 -2738 -5047 -2722
rect -5174 -2862 -5070 -2738
rect -5174 -2878 -5047 -2862
rect -5603 -2990 -5281 -2989
rect -5603 -3310 -5602 -2990
rect -5282 -3310 -5281 -2990
rect -5603 -3311 -5281 -3310
rect -5893 -3438 -5766 -3422
rect -5893 -3562 -5789 -3438
rect -5893 -3578 -5766 -3562
rect -6322 -3690 -6000 -3689
rect -6322 -4010 -6321 -3690
rect -6001 -4010 -6000 -3690
rect -6322 -4011 -6000 -4010
rect -6612 -4138 -6485 -4122
rect -6612 -4262 -6508 -4138
rect -6612 -4278 -6485 -4262
rect -7041 -4390 -6719 -4389
rect -7041 -4710 -7040 -4390
rect -6720 -4710 -6719 -4390
rect -7041 -4711 -6719 -4710
rect -6932 -5089 -6828 -4711
rect -6612 -4822 -6565 -4278
rect -6501 -4822 -6485 -4278
rect -6213 -4389 -6109 -4011
rect -5893 -4122 -5846 -3578
rect -5782 -4122 -5766 -3578
rect -5494 -3689 -5390 -3311
rect -5174 -3422 -5127 -2878
rect -5063 -3422 -5047 -2878
rect -4775 -2989 -4671 -2611
rect -4455 -2722 -4408 -2178
rect -4344 -2722 -4328 -2178
rect -4056 -2289 -3952 -1911
rect -3736 -2022 -3689 -1478
rect -3625 -2022 -3609 -1478
rect -3337 -1589 -3233 -1211
rect -3017 -1322 -2970 -778
rect -2906 -1322 -2890 -778
rect -2618 -889 -2514 -511
rect -2298 -622 -2251 -78
rect -2187 -622 -2171 -78
rect -1899 -189 -1795 189
rect -1579 78 -1532 622
rect -1468 78 -1452 622
rect -1180 511 -1076 889
rect -860 778 -813 1322
rect -749 778 -733 1322
rect -461 1211 -357 1589
rect -141 1478 -94 2022
rect -30 1478 -14 2022
rect 258 1911 362 2289
rect 578 2178 625 2722
rect 689 2178 705 2722
rect 977 2611 1081 2989
rect 1297 2878 1344 3422
rect 1408 2878 1424 3422
rect 1696 3311 1800 3689
rect 2016 3578 2063 4122
rect 2127 3578 2143 4122
rect 2415 4011 2519 4389
rect 2735 4278 2782 4822
rect 2846 4278 2862 4822
rect 3134 4711 3238 5089
rect 3454 4978 3501 5522
rect 3565 4978 3581 5522
rect 3853 5411 3957 5789
rect 4173 5678 4220 6222
rect 4284 5678 4300 6222
rect 4572 6111 4676 6489
rect 4892 6378 4939 6922
rect 5003 6378 5019 6922
rect 5291 6811 5395 7000
rect 5611 6938 5715 7000
rect 5611 6922 5738 6938
rect 5182 6810 5504 6811
rect 5182 6490 5183 6810
rect 5503 6490 5504 6810
rect 5182 6489 5504 6490
rect 4892 6362 5019 6378
rect 4892 6238 4996 6362
rect 4892 6222 5019 6238
rect 4463 6110 4785 6111
rect 4463 5790 4464 6110
rect 4784 5790 4785 6110
rect 4463 5789 4785 5790
rect 4173 5662 4300 5678
rect 4173 5538 4277 5662
rect 4173 5522 4300 5538
rect 3744 5410 4066 5411
rect 3744 5090 3745 5410
rect 4065 5090 4066 5410
rect 3744 5089 4066 5090
rect 3454 4962 3581 4978
rect 3454 4838 3558 4962
rect 3454 4822 3581 4838
rect 3025 4710 3347 4711
rect 3025 4390 3026 4710
rect 3346 4390 3347 4710
rect 3025 4389 3347 4390
rect 2735 4262 2862 4278
rect 2735 4138 2839 4262
rect 2735 4122 2862 4138
rect 2306 4010 2628 4011
rect 2306 3690 2307 4010
rect 2627 3690 2628 4010
rect 2306 3689 2628 3690
rect 2016 3562 2143 3578
rect 2016 3438 2120 3562
rect 2016 3422 2143 3438
rect 1587 3310 1909 3311
rect 1587 2990 1588 3310
rect 1908 2990 1909 3310
rect 1587 2989 1909 2990
rect 1297 2862 1424 2878
rect 1297 2738 1401 2862
rect 1297 2722 1424 2738
rect 868 2610 1190 2611
rect 868 2290 869 2610
rect 1189 2290 1190 2610
rect 868 2289 1190 2290
rect 578 2162 705 2178
rect 578 2038 682 2162
rect 578 2022 705 2038
rect 149 1910 471 1911
rect 149 1590 150 1910
rect 470 1590 471 1910
rect 149 1589 471 1590
rect -141 1462 -14 1478
rect -141 1338 -37 1462
rect -141 1322 -14 1338
rect -570 1210 -248 1211
rect -570 890 -569 1210
rect -249 890 -248 1210
rect -570 889 -248 890
rect -860 762 -733 778
rect -860 638 -756 762
rect -860 622 -733 638
rect -1289 510 -967 511
rect -1289 190 -1288 510
rect -968 190 -967 510
rect -1289 189 -967 190
rect -1579 62 -1452 78
rect -1579 -62 -1475 62
rect -1579 -78 -1452 -62
rect -2008 -190 -1686 -189
rect -2008 -510 -2007 -190
rect -1687 -510 -1686 -190
rect -2008 -511 -1686 -510
rect -2298 -638 -2171 -622
rect -2298 -762 -2194 -638
rect -2298 -778 -2171 -762
rect -2727 -890 -2405 -889
rect -2727 -1210 -2726 -890
rect -2406 -1210 -2405 -890
rect -2727 -1211 -2405 -1210
rect -3017 -1338 -2890 -1322
rect -3017 -1462 -2913 -1338
rect -3017 -1478 -2890 -1462
rect -3446 -1590 -3124 -1589
rect -3446 -1910 -3445 -1590
rect -3125 -1910 -3124 -1590
rect -3446 -1911 -3124 -1910
rect -3736 -2038 -3609 -2022
rect -3736 -2162 -3632 -2038
rect -3736 -2178 -3609 -2162
rect -4165 -2290 -3843 -2289
rect -4165 -2610 -4164 -2290
rect -3844 -2610 -3843 -2290
rect -4165 -2611 -3843 -2610
rect -4455 -2738 -4328 -2722
rect -4455 -2862 -4351 -2738
rect -4455 -2878 -4328 -2862
rect -4884 -2990 -4562 -2989
rect -4884 -3310 -4883 -2990
rect -4563 -3310 -4562 -2990
rect -4884 -3311 -4562 -3310
rect -5174 -3438 -5047 -3422
rect -5174 -3562 -5070 -3438
rect -5174 -3578 -5047 -3562
rect -5603 -3690 -5281 -3689
rect -5603 -4010 -5602 -3690
rect -5282 -4010 -5281 -3690
rect -5603 -4011 -5281 -4010
rect -5893 -4138 -5766 -4122
rect -5893 -4262 -5789 -4138
rect -5893 -4278 -5766 -4262
rect -6322 -4390 -6000 -4389
rect -6322 -4710 -6321 -4390
rect -6001 -4710 -6000 -4390
rect -6322 -4711 -6000 -4710
rect -6612 -4838 -6485 -4822
rect -6612 -4962 -6508 -4838
rect -6612 -4978 -6485 -4962
rect -7041 -5090 -6719 -5089
rect -7041 -5410 -7040 -5090
rect -6720 -5410 -6719 -5090
rect -7041 -5411 -6719 -5410
rect -6932 -5789 -6828 -5411
rect -6612 -5522 -6565 -4978
rect -6501 -5522 -6485 -4978
rect -6213 -5089 -6109 -4711
rect -5893 -4822 -5846 -4278
rect -5782 -4822 -5766 -4278
rect -5494 -4389 -5390 -4011
rect -5174 -4122 -5127 -3578
rect -5063 -4122 -5047 -3578
rect -4775 -3689 -4671 -3311
rect -4455 -3422 -4408 -2878
rect -4344 -3422 -4328 -2878
rect -4056 -2989 -3952 -2611
rect -3736 -2722 -3689 -2178
rect -3625 -2722 -3609 -2178
rect -3337 -2289 -3233 -1911
rect -3017 -2022 -2970 -1478
rect -2906 -2022 -2890 -1478
rect -2618 -1589 -2514 -1211
rect -2298 -1322 -2251 -778
rect -2187 -1322 -2171 -778
rect -1899 -889 -1795 -511
rect -1579 -622 -1532 -78
rect -1468 -622 -1452 -78
rect -1180 -189 -1076 189
rect -860 78 -813 622
rect -749 78 -733 622
rect -461 511 -357 889
rect -141 778 -94 1322
rect -30 778 -14 1322
rect 258 1211 362 1589
rect 578 1478 625 2022
rect 689 1478 705 2022
rect 977 1911 1081 2289
rect 1297 2178 1344 2722
rect 1408 2178 1424 2722
rect 1696 2611 1800 2989
rect 2016 2878 2063 3422
rect 2127 2878 2143 3422
rect 2415 3311 2519 3689
rect 2735 3578 2782 4122
rect 2846 3578 2862 4122
rect 3134 4011 3238 4389
rect 3454 4278 3501 4822
rect 3565 4278 3581 4822
rect 3853 4711 3957 5089
rect 4173 4978 4220 5522
rect 4284 4978 4300 5522
rect 4572 5411 4676 5789
rect 4892 5678 4939 6222
rect 5003 5678 5019 6222
rect 5291 6111 5395 6489
rect 5611 6378 5658 6922
rect 5722 6378 5738 6922
rect 6010 6811 6114 7000
rect 6330 6938 6434 7000
rect 6330 6922 6457 6938
rect 5901 6810 6223 6811
rect 5901 6490 5902 6810
rect 6222 6490 6223 6810
rect 5901 6489 6223 6490
rect 5611 6362 5738 6378
rect 5611 6238 5715 6362
rect 5611 6222 5738 6238
rect 5182 6110 5504 6111
rect 5182 5790 5183 6110
rect 5503 5790 5504 6110
rect 5182 5789 5504 5790
rect 4892 5662 5019 5678
rect 4892 5538 4996 5662
rect 4892 5522 5019 5538
rect 4463 5410 4785 5411
rect 4463 5090 4464 5410
rect 4784 5090 4785 5410
rect 4463 5089 4785 5090
rect 4173 4962 4300 4978
rect 4173 4838 4277 4962
rect 4173 4822 4300 4838
rect 3744 4710 4066 4711
rect 3744 4390 3745 4710
rect 4065 4390 4066 4710
rect 3744 4389 4066 4390
rect 3454 4262 3581 4278
rect 3454 4138 3558 4262
rect 3454 4122 3581 4138
rect 3025 4010 3347 4011
rect 3025 3690 3026 4010
rect 3346 3690 3347 4010
rect 3025 3689 3347 3690
rect 2735 3562 2862 3578
rect 2735 3438 2839 3562
rect 2735 3422 2862 3438
rect 2306 3310 2628 3311
rect 2306 2990 2307 3310
rect 2627 2990 2628 3310
rect 2306 2989 2628 2990
rect 2016 2862 2143 2878
rect 2016 2738 2120 2862
rect 2016 2722 2143 2738
rect 1587 2610 1909 2611
rect 1587 2290 1588 2610
rect 1908 2290 1909 2610
rect 1587 2289 1909 2290
rect 1297 2162 1424 2178
rect 1297 2038 1401 2162
rect 1297 2022 1424 2038
rect 868 1910 1190 1911
rect 868 1590 869 1910
rect 1189 1590 1190 1910
rect 868 1589 1190 1590
rect 578 1462 705 1478
rect 578 1338 682 1462
rect 578 1322 705 1338
rect 149 1210 471 1211
rect 149 890 150 1210
rect 470 890 471 1210
rect 149 889 471 890
rect -141 762 -14 778
rect -141 638 -37 762
rect -141 622 -14 638
rect -570 510 -248 511
rect -570 190 -569 510
rect -249 190 -248 510
rect -570 189 -248 190
rect -860 62 -733 78
rect -860 -62 -756 62
rect -860 -78 -733 -62
rect -1289 -190 -967 -189
rect -1289 -510 -1288 -190
rect -968 -510 -967 -190
rect -1289 -511 -967 -510
rect -1579 -638 -1452 -622
rect -1579 -762 -1475 -638
rect -1579 -778 -1452 -762
rect -2008 -890 -1686 -889
rect -2008 -1210 -2007 -890
rect -1687 -1210 -1686 -890
rect -2008 -1211 -1686 -1210
rect -2298 -1338 -2171 -1322
rect -2298 -1462 -2194 -1338
rect -2298 -1478 -2171 -1462
rect -2727 -1590 -2405 -1589
rect -2727 -1910 -2726 -1590
rect -2406 -1910 -2405 -1590
rect -2727 -1911 -2405 -1910
rect -3017 -2038 -2890 -2022
rect -3017 -2162 -2913 -2038
rect -3017 -2178 -2890 -2162
rect -3446 -2290 -3124 -2289
rect -3446 -2610 -3445 -2290
rect -3125 -2610 -3124 -2290
rect -3446 -2611 -3124 -2610
rect -3736 -2738 -3609 -2722
rect -3736 -2862 -3632 -2738
rect -3736 -2878 -3609 -2862
rect -4165 -2990 -3843 -2989
rect -4165 -3310 -4164 -2990
rect -3844 -3310 -3843 -2990
rect -4165 -3311 -3843 -3310
rect -4455 -3438 -4328 -3422
rect -4455 -3562 -4351 -3438
rect -4455 -3578 -4328 -3562
rect -4884 -3690 -4562 -3689
rect -4884 -4010 -4883 -3690
rect -4563 -4010 -4562 -3690
rect -4884 -4011 -4562 -4010
rect -5174 -4138 -5047 -4122
rect -5174 -4262 -5070 -4138
rect -5174 -4278 -5047 -4262
rect -5603 -4390 -5281 -4389
rect -5603 -4710 -5602 -4390
rect -5282 -4710 -5281 -4390
rect -5603 -4711 -5281 -4710
rect -5893 -4838 -5766 -4822
rect -5893 -4962 -5789 -4838
rect -5893 -4978 -5766 -4962
rect -6322 -5090 -6000 -5089
rect -6322 -5410 -6321 -5090
rect -6001 -5410 -6000 -5090
rect -6322 -5411 -6000 -5410
rect -6612 -5538 -6485 -5522
rect -6612 -5662 -6508 -5538
rect -6612 -5678 -6485 -5662
rect -7041 -5790 -6719 -5789
rect -7041 -6110 -7040 -5790
rect -6720 -6110 -6719 -5790
rect -7041 -6111 -6719 -6110
rect -6932 -6489 -6828 -6111
rect -6612 -6222 -6565 -5678
rect -6501 -6222 -6485 -5678
rect -6213 -5789 -6109 -5411
rect -5893 -5522 -5846 -4978
rect -5782 -5522 -5766 -4978
rect -5494 -5089 -5390 -4711
rect -5174 -4822 -5127 -4278
rect -5063 -4822 -5047 -4278
rect -4775 -4389 -4671 -4011
rect -4455 -4122 -4408 -3578
rect -4344 -4122 -4328 -3578
rect -4056 -3689 -3952 -3311
rect -3736 -3422 -3689 -2878
rect -3625 -3422 -3609 -2878
rect -3337 -2989 -3233 -2611
rect -3017 -2722 -2970 -2178
rect -2906 -2722 -2890 -2178
rect -2618 -2289 -2514 -1911
rect -2298 -2022 -2251 -1478
rect -2187 -2022 -2171 -1478
rect -1899 -1589 -1795 -1211
rect -1579 -1322 -1532 -778
rect -1468 -1322 -1452 -778
rect -1180 -889 -1076 -511
rect -860 -622 -813 -78
rect -749 -622 -733 -78
rect -461 -189 -357 189
rect -141 78 -94 622
rect -30 78 -14 622
rect 258 511 362 889
rect 578 778 625 1322
rect 689 778 705 1322
rect 977 1211 1081 1589
rect 1297 1478 1344 2022
rect 1408 1478 1424 2022
rect 1696 1911 1800 2289
rect 2016 2178 2063 2722
rect 2127 2178 2143 2722
rect 2415 2611 2519 2989
rect 2735 2878 2782 3422
rect 2846 2878 2862 3422
rect 3134 3311 3238 3689
rect 3454 3578 3501 4122
rect 3565 3578 3581 4122
rect 3853 4011 3957 4389
rect 4173 4278 4220 4822
rect 4284 4278 4300 4822
rect 4572 4711 4676 5089
rect 4892 4978 4939 5522
rect 5003 4978 5019 5522
rect 5291 5411 5395 5789
rect 5611 5678 5658 6222
rect 5722 5678 5738 6222
rect 6010 6111 6114 6489
rect 6330 6378 6377 6922
rect 6441 6378 6457 6922
rect 6729 6811 6833 7000
rect 7049 6938 7153 7000
rect 7049 6922 7176 6938
rect 6620 6810 6942 6811
rect 6620 6490 6621 6810
rect 6941 6490 6942 6810
rect 6620 6489 6942 6490
rect 6330 6362 6457 6378
rect 6330 6238 6434 6362
rect 6330 6222 6457 6238
rect 5901 6110 6223 6111
rect 5901 5790 5902 6110
rect 6222 5790 6223 6110
rect 5901 5789 6223 5790
rect 5611 5662 5738 5678
rect 5611 5538 5715 5662
rect 5611 5522 5738 5538
rect 5182 5410 5504 5411
rect 5182 5090 5183 5410
rect 5503 5090 5504 5410
rect 5182 5089 5504 5090
rect 4892 4962 5019 4978
rect 4892 4838 4996 4962
rect 4892 4822 5019 4838
rect 4463 4710 4785 4711
rect 4463 4390 4464 4710
rect 4784 4390 4785 4710
rect 4463 4389 4785 4390
rect 4173 4262 4300 4278
rect 4173 4138 4277 4262
rect 4173 4122 4300 4138
rect 3744 4010 4066 4011
rect 3744 3690 3745 4010
rect 4065 3690 4066 4010
rect 3744 3689 4066 3690
rect 3454 3562 3581 3578
rect 3454 3438 3558 3562
rect 3454 3422 3581 3438
rect 3025 3310 3347 3311
rect 3025 2990 3026 3310
rect 3346 2990 3347 3310
rect 3025 2989 3347 2990
rect 2735 2862 2862 2878
rect 2735 2738 2839 2862
rect 2735 2722 2862 2738
rect 2306 2610 2628 2611
rect 2306 2290 2307 2610
rect 2627 2290 2628 2610
rect 2306 2289 2628 2290
rect 2016 2162 2143 2178
rect 2016 2038 2120 2162
rect 2016 2022 2143 2038
rect 1587 1910 1909 1911
rect 1587 1590 1588 1910
rect 1908 1590 1909 1910
rect 1587 1589 1909 1590
rect 1297 1462 1424 1478
rect 1297 1338 1401 1462
rect 1297 1322 1424 1338
rect 868 1210 1190 1211
rect 868 890 869 1210
rect 1189 890 1190 1210
rect 868 889 1190 890
rect 578 762 705 778
rect 578 638 682 762
rect 578 622 705 638
rect 149 510 471 511
rect 149 190 150 510
rect 470 190 471 510
rect 149 189 471 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -570 -190 -248 -189
rect -570 -510 -569 -190
rect -249 -510 -248 -190
rect -570 -511 -248 -510
rect -860 -638 -733 -622
rect -860 -762 -756 -638
rect -860 -778 -733 -762
rect -1289 -890 -967 -889
rect -1289 -1210 -1288 -890
rect -968 -1210 -967 -890
rect -1289 -1211 -967 -1210
rect -1579 -1338 -1452 -1322
rect -1579 -1462 -1475 -1338
rect -1579 -1478 -1452 -1462
rect -2008 -1590 -1686 -1589
rect -2008 -1910 -2007 -1590
rect -1687 -1910 -1686 -1590
rect -2008 -1911 -1686 -1910
rect -2298 -2038 -2171 -2022
rect -2298 -2162 -2194 -2038
rect -2298 -2178 -2171 -2162
rect -2727 -2290 -2405 -2289
rect -2727 -2610 -2726 -2290
rect -2406 -2610 -2405 -2290
rect -2727 -2611 -2405 -2610
rect -3017 -2738 -2890 -2722
rect -3017 -2862 -2913 -2738
rect -3017 -2878 -2890 -2862
rect -3446 -2990 -3124 -2989
rect -3446 -3310 -3445 -2990
rect -3125 -3310 -3124 -2990
rect -3446 -3311 -3124 -3310
rect -3736 -3438 -3609 -3422
rect -3736 -3562 -3632 -3438
rect -3736 -3578 -3609 -3562
rect -4165 -3690 -3843 -3689
rect -4165 -4010 -4164 -3690
rect -3844 -4010 -3843 -3690
rect -4165 -4011 -3843 -4010
rect -4455 -4138 -4328 -4122
rect -4455 -4262 -4351 -4138
rect -4455 -4278 -4328 -4262
rect -4884 -4390 -4562 -4389
rect -4884 -4710 -4883 -4390
rect -4563 -4710 -4562 -4390
rect -4884 -4711 -4562 -4710
rect -5174 -4838 -5047 -4822
rect -5174 -4962 -5070 -4838
rect -5174 -4978 -5047 -4962
rect -5603 -5090 -5281 -5089
rect -5603 -5410 -5602 -5090
rect -5282 -5410 -5281 -5090
rect -5603 -5411 -5281 -5410
rect -5893 -5538 -5766 -5522
rect -5893 -5662 -5789 -5538
rect -5893 -5678 -5766 -5662
rect -6322 -5790 -6000 -5789
rect -6322 -6110 -6321 -5790
rect -6001 -6110 -6000 -5790
rect -6322 -6111 -6000 -6110
rect -6612 -6238 -6485 -6222
rect -6612 -6362 -6508 -6238
rect -6612 -6378 -6485 -6362
rect -7041 -6490 -6719 -6489
rect -7041 -6810 -7040 -6490
rect -6720 -6810 -6719 -6490
rect -7041 -6811 -6719 -6810
rect -6932 -7000 -6828 -6811
rect -6612 -6922 -6565 -6378
rect -6501 -6922 -6485 -6378
rect -6213 -6489 -6109 -6111
rect -5893 -6222 -5846 -5678
rect -5782 -6222 -5766 -5678
rect -5494 -5789 -5390 -5411
rect -5174 -5522 -5127 -4978
rect -5063 -5522 -5047 -4978
rect -4775 -5089 -4671 -4711
rect -4455 -4822 -4408 -4278
rect -4344 -4822 -4328 -4278
rect -4056 -4389 -3952 -4011
rect -3736 -4122 -3689 -3578
rect -3625 -4122 -3609 -3578
rect -3337 -3689 -3233 -3311
rect -3017 -3422 -2970 -2878
rect -2906 -3422 -2890 -2878
rect -2618 -2989 -2514 -2611
rect -2298 -2722 -2251 -2178
rect -2187 -2722 -2171 -2178
rect -1899 -2289 -1795 -1911
rect -1579 -2022 -1532 -1478
rect -1468 -2022 -1452 -1478
rect -1180 -1589 -1076 -1211
rect -860 -1322 -813 -778
rect -749 -1322 -733 -778
rect -461 -889 -357 -511
rect -141 -622 -94 -78
rect -30 -622 -14 -78
rect 258 -189 362 189
rect 578 78 625 622
rect 689 78 705 622
rect 977 511 1081 889
rect 1297 778 1344 1322
rect 1408 778 1424 1322
rect 1696 1211 1800 1589
rect 2016 1478 2063 2022
rect 2127 1478 2143 2022
rect 2415 1911 2519 2289
rect 2735 2178 2782 2722
rect 2846 2178 2862 2722
rect 3134 2611 3238 2989
rect 3454 2878 3501 3422
rect 3565 2878 3581 3422
rect 3853 3311 3957 3689
rect 4173 3578 4220 4122
rect 4284 3578 4300 4122
rect 4572 4011 4676 4389
rect 4892 4278 4939 4822
rect 5003 4278 5019 4822
rect 5291 4711 5395 5089
rect 5611 4978 5658 5522
rect 5722 4978 5738 5522
rect 6010 5411 6114 5789
rect 6330 5678 6377 6222
rect 6441 5678 6457 6222
rect 6729 6111 6833 6489
rect 7049 6378 7096 6922
rect 7160 6378 7176 6922
rect 7049 6362 7176 6378
rect 7049 6238 7153 6362
rect 7049 6222 7176 6238
rect 6620 6110 6942 6111
rect 6620 5790 6621 6110
rect 6941 5790 6942 6110
rect 6620 5789 6942 5790
rect 6330 5662 6457 5678
rect 6330 5538 6434 5662
rect 6330 5522 6457 5538
rect 5901 5410 6223 5411
rect 5901 5090 5902 5410
rect 6222 5090 6223 5410
rect 5901 5089 6223 5090
rect 5611 4962 5738 4978
rect 5611 4838 5715 4962
rect 5611 4822 5738 4838
rect 5182 4710 5504 4711
rect 5182 4390 5183 4710
rect 5503 4390 5504 4710
rect 5182 4389 5504 4390
rect 4892 4262 5019 4278
rect 4892 4138 4996 4262
rect 4892 4122 5019 4138
rect 4463 4010 4785 4011
rect 4463 3690 4464 4010
rect 4784 3690 4785 4010
rect 4463 3689 4785 3690
rect 4173 3562 4300 3578
rect 4173 3438 4277 3562
rect 4173 3422 4300 3438
rect 3744 3310 4066 3311
rect 3744 2990 3745 3310
rect 4065 2990 4066 3310
rect 3744 2989 4066 2990
rect 3454 2862 3581 2878
rect 3454 2738 3558 2862
rect 3454 2722 3581 2738
rect 3025 2610 3347 2611
rect 3025 2290 3026 2610
rect 3346 2290 3347 2610
rect 3025 2289 3347 2290
rect 2735 2162 2862 2178
rect 2735 2038 2839 2162
rect 2735 2022 2862 2038
rect 2306 1910 2628 1911
rect 2306 1590 2307 1910
rect 2627 1590 2628 1910
rect 2306 1589 2628 1590
rect 2016 1462 2143 1478
rect 2016 1338 2120 1462
rect 2016 1322 2143 1338
rect 1587 1210 1909 1211
rect 1587 890 1588 1210
rect 1908 890 1909 1210
rect 1587 889 1909 890
rect 1297 762 1424 778
rect 1297 638 1401 762
rect 1297 622 1424 638
rect 868 510 1190 511
rect 868 190 869 510
rect 1189 190 1190 510
rect 868 189 1190 190
rect 578 62 705 78
rect 578 -62 682 62
rect 578 -78 705 -62
rect 149 -190 471 -189
rect 149 -510 150 -190
rect 470 -510 471 -190
rect 149 -511 471 -510
rect -141 -638 -14 -622
rect -141 -762 -37 -638
rect -141 -778 -14 -762
rect -570 -890 -248 -889
rect -570 -1210 -569 -890
rect -249 -1210 -248 -890
rect -570 -1211 -248 -1210
rect -860 -1338 -733 -1322
rect -860 -1462 -756 -1338
rect -860 -1478 -733 -1462
rect -1289 -1590 -967 -1589
rect -1289 -1910 -1288 -1590
rect -968 -1910 -967 -1590
rect -1289 -1911 -967 -1910
rect -1579 -2038 -1452 -2022
rect -1579 -2162 -1475 -2038
rect -1579 -2178 -1452 -2162
rect -2008 -2290 -1686 -2289
rect -2008 -2610 -2007 -2290
rect -1687 -2610 -1686 -2290
rect -2008 -2611 -1686 -2610
rect -2298 -2738 -2171 -2722
rect -2298 -2862 -2194 -2738
rect -2298 -2878 -2171 -2862
rect -2727 -2990 -2405 -2989
rect -2727 -3310 -2726 -2990
rect -2406 -3310 -2405 -2990
rect -2727 -3311 -2405 -3310
rect -3017 -3438 -2890 -3422
rect -3017 -3562 -2913 -3438
rect -3017 -3578 -2890 -3562
rect -3446 -3690 -3124 -3689
rect -3446 -4010 -3445 -3690
rect -3125 -4010 -3124 -3690
rect -3446 -4011 -3124 -4010
rect -3736 -4138 -3609 -4122
rect -3736 -4262 -3632 -4138
rect -3736 -4278 -3609 -4262
rect -4165 -4390 -3843 -4389
rect -4165 -4710 -4164 -4390
rect -3844 -4710 -3843 -4390
rect -4165 -4711 -3843 -4710
rect -4455 -4838 -4328 -4822
rect -4455 -4962 -4351 -4838
rect -4455 -4978 -4328 -4962
rect -4884 -5090 -4562 -5089
rect -4884 -5410 -4883 -5090
rect -4563 -5410 -4562 -5090
rect -4884 -5411 -4562 -5410
rect -5174 -5538 -5047 -5522
rect -5174 -5662 -5070 -5538
rect -5174 -5678 -5047 -5662
rect -5603 -5790 -5281 -5789
rect -5603 -6110 -5602 -5790
rect -5282 -6110 -5281 -5790
rect -5603 -6111 -5281 -6110
rect -5893 -6238 -5766 -6222
rect -5893 -6362 -5789 -6238
rect -5893 -6378 -5766 -6362
rect -6322 -6490 -6000 -6489
rect -6322 -6810 -6321 -6490
rect -6001 -6810 -6000 -6490
rect -6322 -6811 -6000 -6810
rect -6612 -6938 -6485 -6922
rect -6612 -7000 -6508 -6938
rect -6213 -7000 -6109 -6811
rect -5893 -6922 -5846 -6378
rect -5782 -6922 -5766 -6378
rect -5494 -6489 -5390 -6111
rect -5174 -6222 -5127 -5678
rect -5063 -6222 -5047 -5678
rect -4775 -5789 -4671 -5411
rect -4455 -5522 -4408 -4978
rect -4344 -5522 -4328 -4978
rect -4056 -5089 -3952 -4711
rect -3736 -4822 -3689 -4278
rect -3625 -4822 -3609 -4278
rect -3337 -4389 -3233 -4011
rect -3017 -4122 -2970 -3578
rect -2906 -4122 -2890 -3578
rect -2618 -3689 -2514 -3311
rect -2298 -3422 -2251 -2878
rect -2187 -3422 -2171 -2878
rect -1899 -2989 -1795 -2611
rect -1579 -2722 -1532 -2178
rect -1468 -2722 -1452 -2178
rect -1180 -2289 -1076 -1911
rect -860 -2022 -813 -1478
rect -749 -2022 -733 -1478
rect -461 -1589 -357 -1211
rect -141 -1322 -94 -778
rect -30 -1322 -14 -778
rect 258 -889 362 -511
rect 578 -622 625 -78
rect 689 -622 705 -78
rect 977 -189 1081 189
rect 1297 78 1344 622
rect 1408 78 1424 622
rect 1696 511 1800 889
rect 2016 778 2063 1322
rect 2127 778 2143 1322
rect 2415 1211 2519 1589
rect 2735 1478 2782 2022
rect 2846 1478 2862 2022
rect 3134 1911 3238 2289
rect 3454 2178 3501 2722
rect 3565 2178 3581 2722
rect 3853 2611 3957 2989
rect 4173 2878 4220 3422
rect 4284 2878 4300 3422
rect 4572 3311 4676 3689
rect 4892 3578 4939 4122
rect 5003 3578 5019 4122
rect 5291 4011 5395 4389
rect 5611 4278 5658 4822
rect 5722 4278 5738 4822
rect 6010 4711 6114 5089
rect 6330 4978 6377 5522
rect 6441 4978 6457 5522
rect 6729 5411 6833 5789
rect 7049 5678 7096 6222
rect 7160 5678 7176 6222
rect 7049 5662 7176 5678
rect 7049 5538 7153 5662
rect 7049 5522 7176 5538
rect 6620 5410 6942 5411
rect 6620 5090 6621 5410
rect 6941 5090 6942 5410
rect 6620 5089 6942 5090
rect 6330 4962 6457 4978
rect 6330 4838 6434 4962
rect 6330 4822 6457 4838
rect 5901 4710 6223 4711
rect 5901 4390 5902 4710
rect 6222 4390 6223 4710
rect 5901 4389 6223 4390
rect 5611 4262 5738 4278
rect 5611 4138 5715 4262
rect 5611 4122 5738 4138
rect 5182 4010 5504 4011
rect 5182 3690 5183 4010
rect 5503 3690 5504 4010
rect 5182 3689 5504 3690
rect 4892 3562 5019 3578
rect 4892 3438 4996 3562
rect 4892 3422 5019 3438
rect 4463 3310 4785 3311
rect 4463 2990 4464 3310
rect 4784 2990 4785 3310
rect 4463 2989 4785 2990
rect 4173 2862 4300 2878
rect 4173 2738 4277 2862
rect 4173 2722 4300 2738
rect 3744 2610 4066 2611
rect 3744 2290 3745 2610
rect 4065 2290 4066 2610
rect 3744 2289 4066 2290
rect 3454 2162 3581 2178
rect 3454 2038 3558 2162
rect 3454 2022 3581 2038
rect 3025 1910 3347 1911
rect 3025 1590 3026 1910
rect 3346 1590 3347 1910
rect 3025 1589 3347 1590
rect 2735 1462 2862 1478
rect 2735 1338 2839 1462
rect 2735 1322 2862 1338
rect 2306 1210 2628 1211
rect 2306 890 2307 1210
rect 2627 890 2628 1210
rect 2306 889 2628 890
rect 2016 762 2143 778
rect 2016 638 2120 762
rect 2016 622 2143 638
rect 1587 510 1909 511
rect 1587 190 1588 510
rect 1908 190 1909 510
rect 1587 189 1909 190
rect 1297 62 1424 78
rect 1297 -62 1401 62
rect 1297 -78 1424 -62
rect 868 -190 1190 -189
rect 868 -510 869 -190
rect 1189 -510 1190 -190
rect 868 -511 1190 -510
rect 578 -638 705 -622
rect 578 -762 682 -638
rect 578 -778 705 -762
rect 149 -890 471 -889
rect 149 -1210 150 -890
rect 470 -1210 471 -890
rect 149 -1211 471 -1210
rect -141 -1338 -14 -1322
rect -141 -1462 -37 -1338
rect -141 -1478 -14 -1462
rect -570 -1590 -248 -1589
rect -570 -1910 -569 -1590
rect -249 -1910 -248 -1590
rect -570 -1911 -248 -1910
rect -860 -2038 -733 -2022
rect -860 -2162 -756 -2038
rect -860 -2178 -733 -2162
rect -1289 -2290 -967 -2289
rect -1289 -2610 -1288 -2290
rect -968 -2610 -967 -2290
rect -1289 -2611 -967 -2610
rect -1579 -2738 -1452 -2722
rect -1579 -2862 -1475 -2738
rect -1579 -2878 -1452 -2862
rect -2008 -2990 -1686 -2989
rect -2008 -3310 -2007 -2990
rect -1687 -3310 -1686 -2990
rect -2008 -3311 -1686 -3310
rect -2298 -3438 -2171 -3422
rect -2298 -3562 -2194 -3438
rect -2298 -3578 -2171 -3562
rect -2727 -3690 -2405 -3689
rect -2727 -4010 -2726 -3690
rect -2406 -4010 -2405 -3690
rect -2727 -4011 -2405 -4010
rect -3017 -4138 -2890 -4122
rect -3017 -4262 -2913 -4138
rect -3017 -4278 -2890 -4262
rect -3446 -4390 -3124 -4389
rect -3446 -4710 -3445 -4390
rect -3125 -4710 -3124 -4390
rect -3446 -4711 -3124 -4710
rect -3736 -4838 -3609 -4822
rect -3736 -4962 -3632 -4838
rect -3736 -4978 -3609 -4962
rect -4165 -5090 -3843 -5089
rect -4165 -5410 -4164 -5090
rect -3844 -5410 -3843 -5090
rect -4165 -5411 -3843 -5410
rect -4455 -5538 -4328 -5522
rect -4455 -5662 -4351 -5538
rect -4455 -5678 -4328 -5662
rect -4884 -5790 -4562 -5789
rect -4884 -6110 -4883 -5790
rect -4563 -6110 -4562 -5790
rect -4884 -6111 -4562 -6110
rect -5174 -6238 -5047 -6222
rect -5174 -6362 -5070 -6238
rect -5174 -6378 -5047 -6362
rect -5603 -6490 -5281 -6489
rect -5603 -6810 -5602 -6490
rect -5282 -6810 -5281 -6490
rect -5603 -6811 -5281 -6810
rect -5893 -6938 -5766 -6922
rect -5893 -7000 -5789 -6938
rect -5494 -7000 -5390 -6811
rect -5174 -6922 -5127 -6378
rect -5063 -6922 -5047 -6378
rect -4775 -6489 -4671 -6111
rect -4455 -6222 -4408 -5678
rect -4344 -6222 -4328 -5678
rect -4056 -5789 -3952 -5411
rect -3736 -5522 -3689 -4978
rect -3625 -5522 -3609 -4978
rect -3337 -5089 -3233 -4711
rect -3017 -4822 -2970 -4278
rect -2906 -4822 -2890 -4278
rect -2618 -4389 -2514 -4011
rect -2298 -4122 -2251 -3578
rect -2187 -4122 -2171 -3578
rect -1899 -3689 -1795 -3311
rect -1579 -3422 -1532 -2878
rect -1468 -3422 -1452 -2878
rect -1180 -2989 -1076 -2611
rect -860 -2722 -813 -2178
rect -749 -2722 -733 -2178
rect -461 -2289 -357 -1911
rect -141 -2022 -94 -1478
rect -30 -2022 -14 -1478
rect 258 -1589 362 -1211
rect 578 -1322 625 -778
rect 689 -1322 705 -778
rect 977 -889 1081 -511
rect 1297 -622 1344 -78
rect 1408 -622 1424 -78
rect 1696 -189 1800 189
rect 2016 78 2063 622
rect 2127 78 2143 622
rect 2415 511 2519 889
rect 2735 778 2782 1322
rect 2846 778 2862 1322
rect 3134 1211 3238 1589
rect 3454 1478 3501 2022
rect 3565 1478 3581 2022
rect 3853 1911 3957 2289
rect 4173 2178 4220 2722
rect 4284 2178 4300 2722
rect 4572 2611 4676 2989
rect 4892 2878 4939 3422
rect 5003 2878 5019 3422
rect 5291 3311 5395 3689
rect 5611 3578 5658 4122
rect 5722 3578 5738 4122
rect 6010 4011 6114 4389
rect 6330 4278 6377 4822
rect 6441 4278 6457 4822
rect 6729 4711 6833 5089
rect 7049 4978 7096 5522
rect 7160 4978 7176 5522
rect 7049 4962 7176 4978
rect 7049 4838 7153 4962
rect 7049 4822 7176 4838
rect 6620 4710 6942 4711
rect 6620 4390 6621 4710
rect 6941 4390 6942 4710
rect 6620 4389 6942 4390
rect 6330 4262 6457 4278
rect 6330 4138 6434 4262
rect 6330 4122 6457 4138
rect 5901 4010 6223 4011
rect 5901 3690 5902 4010
rect 6222 3690 6223 4010
rect 5901 3689 6223 3690
rect 5611 3562 5738 3578
rect 5611 3438 5715 3562
rect 5611 3422 5738 3438
rect 5182 3310 5504 3311
rect 5182 2990 5183 3310
rect 5503 2990 5504 3310
rect 5182 2989 5504 2990
rect 4892 2862 5019 2878
rect 4892 2738 4996 2862
rect 4892 2722 5019 2738
rect 4463 2610 4785 2611
rect 4463 2290 4464 2610
rect 4784 2290 4785 2610
rect 4463 2289 4785 2290
rect 4173 2162 4300 2178
rect 4173 2038 4277 2162
rect 4173 2022 4300 2038
rect 3744 1910 4066 1911
rect 3744 1590 3745 1910
rect 4065 1590 4066 1910
rect 3744 1589 4066 1590
rect 3454 1462 3581 1478
rect 3454 1338 3558 1462
rect 3454 1322 3581 1338
rect 3025 1210 3347 1211
rect 3025 890 3026 1210
rect 3346 890 3347 1210
rect 3025 889 3347 890
rect 2735 762 2862 778
rect 2735 638 2839 762
rect 2735 622 2862 638
rect 2306 510 2628 511
rect 2306 190 2307 510
rect 2627 190 2628 510
rect 2306 189 2628 190
rect 2016 62 2143 78
rect 2016 -62 2120 62
rect 2016 -78 2143 -62
rect 1587 -190 1909 -189
rect 1587 -510 1588 -190
rect 1908 -510 1909 -190
rect 1587 -511 1909 -510
rect 1297 -638 1424 -622
rect 1297 -762 1401 -638
rect 1297 -778 1424 -762
rect 868 -890 1190 -889
rect 868 -1210 869 -890
rect 1189 -1210 1190 -890
rect 868 -1211 1190 -1210
rect 578 -1338 705 -1322
rect 578 -1462 682 -1338
rect 578 -1478 705 -1462
rect 149 -1590 471 -1589
rect 149 -1910 150 -1590
rect 470 -1910 471 -1590
rect 149 -1911 471 -1910
rect -141 -2038 -14 -2022
rect -141 -2162 -37 -2038
rect -141 -2178 -14 -2162
rect -570 -2290 -248 -2289
rect -570 -2610 -569 -2290
rect -249 -2610 -248 -2290
rect -570 -2611 -248 -2610
rect -860 -2738 -733 -2722
rect -860 -2862 -756 -2738
rect -860 -2878 -733 -2862
rect -1289 -2990 -967 -2989
rect -1289 -3310 -1288 -2990
rect -968 -3310 -967 -2990
rect -1289 -3311 -967 -3310
rect -1579 -3438 -1452 -3422
rect -1579 -3562 -1475 -3438
rect -1579 -3578 -1452 -3562
rect -2008 -3690 -1686 -3689
rect -2008 -4010 -2007 -3690
rect -1687 -4010 -1686 -3690
rect -2008 -4011 -1686 -4010
rect -2298 -4138 -2171 -4122
rect -2298 -4262 -2194 -4138
rect -2298 -4278 -2171 -4262
rect -2727 -4390 -2405 -4389
rect -2727 -4710 -2726 -4390
rect -2406 -4710 -2405 -4390
rect -2727 -4711 -2405 -4710
rect -3017 -4838 -2890 -4822
rect -3017 -4962 -2913 -4838
rect -3017 -4978 -2890 -4962
rect -3446 -5090 -3124 -5089
rect -3446 -5410 -3445 -5090
rect -3125 -5410 -3124 -5090
rect -3446 -5411 -3124 -5410
rect -3736 -5538 -3609 -5522
rect -3736 -5662 -3632 -5538
rect -3736 -5678 -3609 -5662
rect -4165 -5790 -3843 -5789
rect -4165 -6110 -4164 -5790
rect -3844 -6110 -3843 -5790
rect -4165 -6111 -3843 -6110
rect -4455 -6238 -4328 -6222
rect -4455 -6362 -4351 -6238
rect -4455 -6378 -4328 -6362
rect -4884 -6490 -4562 -6489
rect -4884 -6810 -4883 -6490
rect -4563 -6810 -4562 -6490
rect -4884 -6811 -4562 -6810
rect -5174 -6938 -5047 -6922
rect -5174 -7000 -5070 -6938
rect -4775 -7000 -4671 -6811
rect -4455 -6922 -4408 -6378
rect -4344 -6922 -4328 -6378
rect -4056 -6489 -3952 -6111
rect -3736 -6222 -3689 -5678
rect -3625 -6222 -3609 -5678
rect -3337 -5789 -3233 -5411
rect -3017 -5522 -2970 -4978
rect -2906 -5522 -2890 -4978
rect -2618 -5089 -2514 -4711
rect -2298 -4822 -2251 -4278
rect -2187 -4822 -2171 -4278
rect -1899 -4389 -1795 -4011
rect -1579 -4122 -1532 -3578
rect -1468 -4122 -1452 -3578
rect -1180 -3689 -1076 -3311
rect -860 -3422 -813 -2878
rect -749 -3422 -733 -2878
rect -461 -2989 -357 -2611
rect -141 -2722 -94 -2178
rect -30 -2722 -14 -2178
rect 258 -2289 362 -1911
rect 578 -2022 625 -1478
rect 689 -2022 705 -1478
rect 977 -1589 1081 -1211
rect 1297 -1322 1344 -778
rect 1408 -1322 1424 -778
rect 1696 -889 1800 -511
rect 2016 -622 2063 -78
rect 2127 -622 2143 -78
rect 2415 -189 2519 189
rect 2735 78 2782 622
rect 2846 78 2862 622
rect 3134 511 3238 889
rect 3454 778 3501 1322
rect 3565 778 3581 1322
rect 3853 1211 3957 1589
rect 4173 1478 4220 2022
rect 4284 1478 4300 2022
rect 4572 1911 4676 2289
rect 4892 2178 4939 2722
rect 5003 2178 5019 2722
rect 5291 2611 5395 2989
rect 5611 2878 5658 3422
rect 5722 2878 5738 3422
rect 6010 3311 6114 3689
rect 6330 3578 6377 4122
rect 6441 3578 6457 4122
rect 6729 4011 6833 4389
rect 7049 4278 7096 4822
rect 7160 4278 7176 4822
rect 7049 4262 7176 4278
rect 7049 4138 7153 4262
rect 7049 4122 7176 4138
rect 6620 4010 6942 4011
rect 6620 3690 6621 4010
rect 6941 3690 6942 4010
rect 6620 3689 6942 3690
rect 6330 3562 6457 3578
rect 6330 3438 6434 3562
rect 6330 3422 6457 3438
rect 5901 3310 6223 3311
rect 5901 2990 5902 3310
rect 6222 2990 6223 3310
rect 5901 2989 6223 2990
rect 5611 2862 5738 2878
rect 5611 2738 5715 2862
rect 5611 2722 5738 2738
rect 5182 2610 5504 2611
rect 5182 2290 5183 2610
rect 5503 2290 5504 2610
rect 5182 2289 5504 2290
rect 4892 2162 5019 2178
rect 4892 2038 4996 2162
rect 4892 2022 5019 2038
rect 4463 1910 4785 1911
rect 4463 1590 4464 1910
rect 4784 1590 4785 1910
rect 4463 1589 4785 1590
rect 4173 1462 4300 1478
rect 4173 1338 4277 1462
rect 4173 1322 4300 1338
rect 3744 1210 4066 1211
rect 3744 890 3745 1210
rect 4065 890 4066 1210
rect 3744 889 4066 890
rect 3454 762 3581 778
rect 3454 638 3558 762
rect 3454 622 3581 638
rect 3025 510 3347 511
rect 3025 190 3026 510
rect 3346 190 3347 510
rect 3025 189 3347 190
rect 2735 62 2862 78
rect 2735 -62 2839 62
rect 2735 -78 2862 -62
rect 2306 -190 2628 -189
rect 2306 -510 2307 -190
rect 2627 -510 2628 -190
rect 2306 -511 2628 -510
rect 2016 -638 2143 -622
rect 2016 -762 2120 -638
rect 2016 -778 2143 -762
rect 1587 -890 1909 -889
rect 1587 -1210 1588 -890
rect 1908 -1210 1909 -890
rect 1587 -1211 1909 -1210
rect 1297 -1338 1424 -1322
rect 1297 -1462 1401 -1338
rect 1297 -1478 1424 -1462
rect 868 -1590 1190 -1589
rect 868 -1910 869 -1590
rect 1189 -1910 1190 -1590
rect 868 -1911 1190 -1910
rect 578 -2038 705 -2022
rect 578 -2162 682 -2038
rect 578 -2178 705 -2162
rect 149 -2290 471 -2289
rect 149 -2610 150 -2290
rect 470 -2610 471 -2290
rect 149 -2611 471 -2610
rect -141 -2738 -14 -2722
rect -141 -2862 -37 -2738
rect -141 -2878 -14 -2862
rect -570 -2990 -248 -2989
rect -570 -3310 -569 -2990
rect -249 -3310 -248 -2990
rect -570 -3311 -248 -3310
rect -860 -3438 -733 -3422
rect -860 -3562 -756 -3438
rect -860 -3578 -733 -3562
rect -1289 -3690 -967 -3689
rect -1289 -4010 -1288 -3690
rect -968 -4010 -967 -3690
rect -1289 -4011 -967 -4010
rect -1579 -4138 -1452 -4122
rect -1579 -4262 -1475 -4138
rect -1579 -4278 -1452 -4262
rect -2008 -4390 -1686 -4389
rect -2008 -4710 -2007 -4390
rect -1687 -4710 -1686 -4390
rect -2008 -4711 -1686 -4710
rect -2298 -4838 -2171 -4822
rect -2298 -4962 -2194 -4838
rect -2298 -4978 -2171 -4962
rect -2727 -5090 -2405 -5089
rect -2727 -5410 -2726 -5090
rect -2406 -5410 -2405 -5090
rect -2727 -5411 -2405 -5410
rect -3017 -5538 -2890 -5522
rect -3017 -5662 -2913 -5538
rect -3017 -5678 -2890 -5662
rect -3446 -5790 -3124 -5789
rect -3446 -6110 -3445 -5790
rect -3125 -6110 -3124 -5790
rect -3446 -6111 -3124 -6110
rect -3736 -6238 -3609 -6222
rect -3736 -6362 -3632 -6238
rect -3736 -6378 -3609 -6362
rect -4165 -6490 -3843 -6489
rect -4165 -6810 -4164 -6490
rect -3844 -6810 -3843 -6490
rect -4165 -6811 -3843 -6810
rect -4455 -6938 -4328 -6922
rect -4455 -7000 -4351 -6938
rect -4056 -7000 -3952 -6811
rect -3736 -6922 -3689 -6378
rect -3625 -6922 -3609 -6378
rect -3337 -6489 -3233 -6111
rect -3017 -6222 -2970 -5678
rect -2906 -6222 -2890 -5678
rect -2618 -5789 -2514 -5411
rect -2298 -5522 -2251 -4978
rect -2187 -5522 -2171 -4978
rect -1899 -5089 -1795 -4711
rect -1579 -4822 -1532 -4278
rect -1468 -4822 -1452 -4278
rect -1180 -4389 -1076 -4011
rect -860 -4122 -813 -3578
rect -749 -4122 -733 -3578
rect -461 -3689 -357 -3311
rect -141 -3422 -94 -2878
rect -30 -3422 -14 -2878
rect 258 -2989 362 -2611
rect 578 -2722 625 -2178
rect 689 -2722 705 -2178
rect 977 -2289 1081 -1911
rect 1297 -2022 1344 -1478
rect 1408 -2022 1424 -1478
rect 1696 -1589 1800 -1211
rect 2016 -1322 2063 -778
rect 2127 -1322 2143 -778
rect 2415 -889 2519 -511
rect 2735 -622 2782 -78
rect 2846 -622 2862 -78
rect 3134 -189 3238 189
rect 3454 78 3501 622
rect 3565 78 3581 622
rect 3853 511 3957 889
rect 4173 778 4220 1322
rect 4284 778 4300 1322
rect 4572 1211 4676 1589
rect 4892 1478 4939 2022
rect 5003 1478 5019 2022
rect 5291 1911 5395 2289
rect 5611 2178 5658 2722
rect 5722 2178 5738 2722
rect 6010 2611 6114 2989
rect 6330 2878 6377 3422
rect 6441 2878 6457 3422
rect 6729 3311 6833 3689
rect 7049 3578 7096 4122
rect 7160 3578 7176 4122
rect 7049 3562 7176 3578
rect 7049 3438 7153 3562
rect 7049 3422 7176 3438
rect 6620 3310 6942 3311
rect 6620 2990 6621 3310
rect 6941 2990 6942 3310
rect 6620 2989 6942 2990
rect 6330 2862 6457 2878
rect 6330 2738 6434 2862
rect 6330 2722 6457 2738
rect 5901 2610 6223 2611
rect 5901 2290 5902 2610
rect 6222 2290 6223 2610
rect 5901 2289 6223 2290
rect 5611 2162 5738 2178
rect 5611 2038 5715 2162
rect 5611 2022 5738 2038
rect 5182 1910 5504 1911
rect 5182 1590 5183 1910
rect 5503 1590 5504 1910
rect 5182 1589 5504 1590
rect 4892 1462 5019 1478
rect 4892 1338 4996 1462
rect 4892 1322 5019 1338
rect 4463 1210 4785 1211
rect 4463 890 4464 1210
rect 4784 890 4785 1210
rect 4463 889 4785 890
rect 4173 762 4300 778
rect 4173 638 4277 762
rect 4173 622 4300 638
rect 3744 510 4066 511
rect 3744 190 3745 510
rect 4065 190 4066 510
rect 3744 189 4066 190
rect 3454 62 3581 78
rect 3454 -62 3558 62
rect 3454 -78 3581 -62
rect 3025 -190 3347 -189
rect 3025 -510 3026 -190
rect 3346 -510 3347 -190
rect 3025 -511 3347 -510
rect 2735 -638 2862 -622
rect 2735 -762 2839 -638
rect 2735 -778 2862 -762
rect 2306 -890 2628 -889
rect 2306 -1210 2307 -890
rect 2627 -1210 2628 -890
rect 2306 -1211 2628 -1210
rect 2016 -1338 2143 -1322
rect 2016 -1462 2120 -1338
rect 2016 -1478 2143 -1462
rect 1587 -1590 1909 -1589
rect 1587 -1910 1588 -1590
rect 1908 -1910 1909 -1590
rect 1587 -1911 1909 -1910
rect 1297 -2038 1424 -2022
rect 1297 -2162 1401 -2038
rect 1297 -2178 1424 -2162
rect 868 -2290 1190 -2289
rect 868 -2610 869 -2290
rect 1189 -2610 1190 -2290
rect 868 -2611 1190 -2610
rect 578 -2738 705 -2722
rect 578 -2862 682 -2738
rect 578 -2878 705 -2862
rect 149 -2990 471 -2989
rect 149 -3310 150 -2990
rect 470 -3310 471 -2990
rect 149 -3311 471 -3310
rect -141 -3438 -14 -3422
rect -141 -3562 -37 -3438
rect -141 -3578 -14 -3562
rect -570 -3690 -248 -3689
rect -570 -4010 -569 -3690
rect -249 -4010 -248 -3690
rect -570 -4011 -248 -4010
rect -860 -4138 -733 -4122
rect -860 -4262 -756 -4138
rect -860 -4278 -733 -4262
rect -1289 -4390 -967 -4389
rect -1289 -4710 -1288 -4390
rect -968 -4710 -967 -4390
rect -1289 -4711 -967 -4710
rect -1579 -4838 -1452 -4822
rect -1579 -4962 -1475 -4838
rect -1579 -4978 -1452 -4962
rect -2008 -5090 -1686 -5089
rect -2008 -5410 -2007 -5090
rect -1687 -5410 -1686 -5090
rect -2008 -5411 -1686 -5410
rect -2298 -5538 -2171 -5522
rect -2298 -5662 -2194 -5538
rect -2298 -5678 -2171 -5662
rect -2727 -5790 -2405 -5789
rect -2727 -6110 -2726 -5790
rect -2406 -6110 -2405 -5790
rect -2727 -6111 -2405 -6110
rect -3017 -6238 -2890 -6222
rect -3017 -6362 -2913 -6238
rect -3017 -6378 -2890 -6362
rect -3446 -6490 -3124 -6489
rect -3446 -6810 -3445 -6490
rect -3125 -6810 -3124 -6490
rect -3446 -6811 -3124 -6810
rect -3736 -6938 -3609 -6922
rect -3736 -7000 -3632 -6938
rect -3337 -7000 -3233 -6811
rect -3017 -6922 -2970 -6378
rect -2906 -6922 -2890 -6378
rect -2618 -6489 -2514 -6111
rect -2298 -6222 -2251 -5678
rect -2187 -6222 -2171 -5678
rect -1899 -5789 -1795 -5411
rect -1579 -5522 -1532 -4978
rect -1468 -5522 -1452 -4978
rect -1180 -5089 -1076 -4711
rect -860 -4822 -813 -4278
rect -749 -4822 -733 -4278
rect -461 -4389 -357 -4011
rect -141 -4122 -94 -3578
rect -30 -4122 -14 -3578
rect 258 -3689 362 -3311
rect 578 -3422 625 -2878
rect 689 -3422 705 -2878
rect 977 -2989 1081 -2611
rect 1297 -2722 1344 -2178
rect 1408 -2722 1424 -2178
rect 1696 -2289 1800 -1911
rect 2016 -2022 2063 -1478
rect 2127 -2022 2143 -1478
rect 2415 -1589 2519 -1211
rect 2735 -1322 2782 -778
rect 2846 -1322 2862 -778
rect 3134 -889 3238 -511
rect 3454 -622 3501 -78
rect 3565 -622 3581 -78
rect 3853 -189 3957 189
rect 4173 78 4220 622
rect 4284 78 4300 622
rect 4572 511 4676 889
rect 4892 778 4939 1322
rect 5003 778 5019 1322
rect 5291 1211 5395 1589
rect 5611 1478 5658 2022
rect 5722 1478 5738 2022
rect 6010 1911 6114 2289
rect 6330 2178 6377 2722
rect 6441 2178 6457 2722
rect 6729 2611 6833 2989
rect 7049 2878 7096 3422
rect 7160 2878 7176 3422
rect 7049 2862 7176 2878
rect 7049 2738 7153 2862
rect 7049 2722 7176 2738
rect 6620 2610 6942 2611
rect 6620 2290 6621 2610
rect 6941 2290 6942 2610
rect 6620 2289 6942 2290
rect 6330 2162 6457 2178
rect 6330 2038 6434 2162
rect 6330 2022 6457 2038
rect 5901 1910 6223 1911
rect 5901 1590 5902 1910
rect 6222 1590 6223 1910
rect 5901 1589 6223 1590
rect 5611 1462 5738 1478
rect 5611 1338 5715 1462
rect 5611 1322 5738 1338
rect 5182 1210 5504 1211
rect 5182 890 5183 1210
rect 5503 890 5504 1210
rect 5182 889 5504 890
rect 4892 762 5019 778
rect 4892 638 4996 762
rect 4892 622 5019 638
rect 4463 510 4785 511
rect 4463 190 4464 510
rect 4784 190 4785 510
rect 4463 189 4785 190
rect 4173 62 4300 78
rect 4173 -62 4277 62
rect 4173 -78 4300 -62
rect 3744 -190 4066 -189
rect 3744 -510 3745 -190
rect 4065 -510 4066 -190
rect 3744 -511 4066 -510
rect 3454 -638 3581 -622
rect 3454 -762 3558 -638
rect 3454 -778 3581 -762
rect 3025 -890 3347 -889
rect 3025 -1210 3026 -890
rect 3346 -1210 3347 -890
rect 3025 -1211 3347 -1210
rect 2735 -1338 2862 -1322
rect 2735 -1462 2839 -1338
rect 2735 -1478 2862 -1462
rect 2306 -1590 2628 -1589
rect 2306 -1910 2307 -1590
rect 2627 -1910 2628 -1590
rect 2306 -1911 2628 -1910
rect 2016 -2038 2143 -2022
rect 2016 -2162 2120 -2038
rect 2016 -2178 2143 -2162
rect 1587 -2290 1909 -2289
rect 1587 -2610 1588 -2290
rect 1908 -2610 1909 -2290
rect 1587 -2611 1909 -2610
rect 1297 -2738 1424 -2722
rect 1297 -2862 1401 -2738
rect 1297 -2878 1424 -2862
rect 868 -2990 1190 -2989
rect 868 -3310 869 -2990
rect 1189 -3310 1190 -2990
rect 868 -3311 1190 -3310
rect 578 -3438 705 -3422
rect 578 -3562 682 -3438
rect 578 -3578 705 -3562
rect 149 -3690 471 -3689
rect 149 -4010 150 -3690
rect 470 -4010 471 -3690
rect 149 -4011 471 -4010
rect -141 -4138 -14 -4122
rect -141 -4262 -37 -4138
rect -141 -4278 -14 -4262
rect -570 -4390 -248 -4389
rect -570 -4710 -569 -4390
rect -249 -4710 -248 -4390
rect -570 -4711 -248 -4710
rect -860 -4838 -733 -4822
rect -860 -4962 -756 -4838
rect -860 -4978 -733 -4962
rect -1289 -5090 -967 -5089
rect -1289 -5410 -1288 -5090
rect -968 -5410 -967 -5090
rect -1289 -5411 -967 -5410
rect -1579 -5538 -1452 -5522
rect -1579 -5662 -1475 -5538
rect -1579 -5678 -1452 -5662
rect -2008 -5790 -1686 -5789
rect -2008 -6110 -2007 -5790
rect -1687 -6110 -1686 -5790
rect -2008 -6111 -1686 -6110
rect -2298 -6238 -2171 -6222
rect -2298 -6362 -2194 -6238
rect -2298 -6378 -2171 -6362
rect -2727 -6490 -2405 -6489
rect -2727 -6810 -2726 -6490
rect -2406 -6810 -2405 -6490
rect -2727 -6811 -2405 -6810
rect -3017 -6938 -2890 -6922
rect -3017 -7000 -2913 -6938
rect -2618 -7000 -2514 -6811
rect -2298 -6922 -2251 -6378
rect -2187 -6922 -2171 -6378
rect -1899 -6489 -1795 -6111
rect -1579 -6222 -1532 -5678
rect -1468 -6222 -1452 -5678
rect -1180 -5789 -1076 -5411
rect -860 -5522 -813 -4978
rect -749 -5522 -733 -4978
rect -461 -5089 -357 -4711
rect -141 -4822 -94 -4278
rect -30 -4822 -14 -4278
rect 258 -4389 362 -4011
rect 578 -4122 625 -3578
rect 689 -4122 705 -3578
rect 977 -3689 1081 -3311
rect 1297 -3422 1344 -2878
rect 1408 -3422 1424 -2878
rect 1696 -2989 1800 -2611
rect 2016 -2722 2063 -2178
rect 2127 -2722 2143 -2178
rect 2415 -2289 2519 -1911
rect 2735 -2022 2782 -1478
rect 2846 -2022 2862 -1478
rect 3134 -1589 3238 -1211
rect 3454 -1322 3501 -778
rect 3565 -1322 3581 -778
rect 3853 -889 3957 -511
rect 4173 -622 4220 -78
rect 4284 -622 4300 -78
rect 4572 -189 4676 189
rect 4892 78 4939 622
rect 5003 78 5019 622
rect 5291 511 5395 889
rect 5611 778 5658 1322
rect 5722 778 5738 1322
rect 6010 1211 6114 1589
rect 6330 1478 6377 2022
rect 6441 1478 6457 2022
rect 6729 1911 6833 2289
rect 7049 2178 7096 2722
rect 7160 2178 7176 2722
rect 7049 2162 7176 2178
rect 7049 2038 7153 2162
rect 7049 2022 7176 2038
rect 6620 1910 6942 1911
rect 6620 1590 6621 1910
rect 6941 1590 6942 1910
rect 6620 1589 6942 1590
rect 6330 1462 6457 1478
rect 6330 1338 6434 1462
rect 6330 1322 6457 1338
rect 5901 1210 6223 1211
rect 5901 890 5902 1210
rect 6222 890 6223 1210
rect 5901 889 6223 890
rect 5611 762 5738 778
rect 5611 638 5715 762
rect 5611 622 5738 638
rect 5182 510 5504 511
rect 5182 190 5183 510
rect 5503 190 5504 510
rect 5182 189 5504 190
rect 4892 62 5019 78
rect 4892 -62 4996 62
rect 4892 -78 5019 -62
rect 4463 -190 4785 -189
rect 4463 -510 4464 -190
rect 4784 -510 4785 -190
rect 4463 -511 4785 -510
rect 4173 -638 4300 -622
rect 4173 -762 4277 -638
rect 4173 -778 4300 -762
rect 3744 -890 4066 -889
rect 3744 -1210 3745 -890
rect 4065 -1210 4066 -890
rect 3744 -1211 4066 -1210
rect 3454 -1338 3581 -1322
rect 3454 -1462 3558 -1338
rect 3454 -1478 3581 -1462
rect 3025 -1590 3347 -1589
rect 3025 -1910 3026 -1590
rect 3346 -1910 3347 -1590
rect 3025 -1911 3347 -1910
rect 2735 -2038 2862 -2022
rect 2735 -2162 2839 -2038
rect 2735 -2178 2862 -2162
rect 2306 -2290 2628 -2289
rect 2306 -2610 2307 -2290
rect 2627 -2610 2628 -2290
rect 2306 -2611 2628 -2610
rect 2016 -2738 2143 -2722
rect 2016 -2862 2120 -2738
rect 2016 -2878 2143 -2862
rect 1587 -2990 1909 -2989
rect 1587 -3310 1588 -2990
rect 1908 -3310 1909 -2990
rect 1587 -3311 1909 -3310
rect 1297 -3438 1424 -3422
rect 1297 -3562 1401 -3438
rect 1297 -3578 1424 -3562
rect 868 -3690 1190 -3689
rect 868 -4010 869 -3690
rect 1189 -4010 1190 -3690
rect 868 -4011 1190 -4010
rect 578 -4138 705 -4122
rect 578 -4262 682 -4138
rect 578 -4278 705 -4262
rect 149 -4390 471 -4389
rect 149 -4710 150 -4390
rect 470 -4710 471 -4390
rect 149 -4711 471 -4710
rect -141 -4838 -14 -4822
rect -141 -4962 -37 -4838
rect -141 -4978 -14 -4962
rect -570 -5090 -248 -5089
rect -570 -5410 -569 -5090
rect -249 -5410 -248 -5090
rect -570 -5411 -248 -5410
rect -860 -5538 -733 -5522
rect -860 -5662 -756 -5538
rect -860 -5678 -733 -5662
rect -1289 -5790 -967 -5789
rect -1289 -6110 -1288 -5790
rect -968 -6110 -967 -5790
rect -1289 -6111 -967 -6110
rect -1579 -6238 -1452 -6222
rect -1579 -6362 -1475 -6238
rect -1579 -6378 -1452 -6362
rect -2008 -6490 -1686 -6489
rect -2008 -6810 -2007 -6490
rect -1687 -6810 -1686 -6490
rect -2008 -6811 -1686 -6810
rect -2298 -6938 -2171 -6922
rect -2298 -7000 -2194 -6938
rect -1899 -7000 -1795 -6811
rect -1579 -6922 -1532 -6378
rect -1468 -6922 -1452 -6378
rect -1180 -6489 -1076 -6111
rect -860 -6222 -813 -5678
rect -749 -6222 -733 -5678
rect -461 -5789 -357 -5411
rect -141 -5522 -94 -4978
rect -30 -5522 -14 -4978
rect 258 -5089 362 -4711
rect 578 -4822 625 -4278
rect 689 -4822 705 -4278
rect 977 -4389 1081 -4011
rect 1297 -4122 1344 -3578
rect 1408 -4122 1424 -3578
rect 1696 -3689 1800 -3311
rect 2016 -3422 2063 -2878
rect 2127 -3422 2143 -2878
rect 2415 -2989 2519 -2611
rect 2735 -2722 2782 -2178
rect 2846 -2722 2862 -2178
rect 3134 -2289 3238 -1911
rect 3454 -2022 3501 -1478
rect 3565 -2022 3581 -1478
rect 3853 -1589 3957 -1211
rect 4173 -1322 4220 -778
rect 4284 -1322 4300 -778
rect 4572 -889 4676 -511
rect 4892 -622 4939 -78
rect 5003 -622 5019 -78
rect 5291 -189 5395 189
rect 5611 78 5658 622
rect 5722 78 5738 622
rect 6010 511 6114 889
rect 6330 778 6377 1322
rect 6441 778 6457 1322
rect 6729 1211 6833 1589
rect 7049 1478 7096 2022
rect 7160 1478 7176 2022
rect 7049 1462 7176 1478
rect 7049 1338 7153 1462
rect 7049 1322 7176 1338
rect 6620 1210 6942 1211
rect 6620 890 6621 1210
rect 6941 890 6942 1210
rect 6620 889 6942 890
rect 6330 762 6457 778
rect 6330 638 6434 762
rect 6330 622 6457 638
rect 5901 510 6223 511
rect 5901 190 5902 510
rect 6222 190 6223 510
rect 5901 189 6223 190
rect 5611 62 5738 78
rect 5611 -62 5715 62
rect 5611 -78 5738 -62
rect 5182 -190 5504 -189
rect 5182 -510 5183 -190
rect 5503 -510 5504 -190
rect 5182 -511 5504 -510
rect 4892 -638 5019 -622
rect 4892 -762 4996 -638
rect 4892 -778 5019 -762
rect 4463 -890 4785 -889
rect 4463 -1210 4464 -890
rect 4784 -1210 4785 -890
rect 4463 -1211 4785 -1210
rect 4173 -1338 4300 -1322
rect 4173 -1462 4277 -1338
rect 4173 -1478 4300 -1462
rect 3744 -1590 4066 -1589
rect 3744 -1910 3745 -1590
rect 4065 -1910 4066 -1590
rect 3744 -1911 4066 -1910
rect 3454 -2038 3581 -2022
rect 3454 -2162 3558 -2038
rect 3454 -2178 3581 -2162
rect 3025 -2290 3347 -2289
rect 3025 -2610 3026 -2290
rect 3346 -2610 3347 -2290
rect 3025 -2611 3347 -2610
rect 2735 -2738 2862 -2722
rect 2735 -2862 2839 -2738
rect 2735 -2878 2862 -2862
rect 2306 -2990 2628 -2989
rect 2306 -3310 2307 -2990
rect 2627 -3310 2628 -2990
rect 2306 -3311 2628 -3310
rect 2016 -3438 2143 -3422
rect 2016 -3562 2120 -3438
rect 2016 -3578 2143 -3562
rect 1587 -3690 1909 -3689
rect 1587 -4010 1588 -3690
rect 1908 -4010 1909 -3690
rect 1587 -4011 1909 -4010
rect 1297 -4138 1424 -4122
rect 1297 -4262 1401 -4138
rect 1297 -4278 1424 -4262
rect 868 -4390 1190 -4389
rect 868 -4710 869 -4390
rect 1189 -4710 1190 -4390
rect 868 -4711 1190 -4710
rect 578 -4838 705 -4822
rect 578 -4962 682 -4838
rect 578 -4978 705 -4962
rect 149 -5090 471 -5089
rect 149 -5410 150 -5090
rect 470 -5410 471 -5090
rect 149 -5411 471 -5410
rect -141 -5538 -14 -5522
rect -141 -5662 -37 -5538
rect -141 -5678 -14 -5662
rect -570 -5790 -248 -5789
rect -570 -6110 -569 -5790
rect -249 -6110 -248 -5790
rect -570 -6111 -248 -6110
rect -860 -6238 -733 -6222
rect -860 -6362 -756 -6238
rect -860 -6378 -733 -6362
rect -1289 -6490 -967 -6489
rect -1289 -6810 -1288 -6490
rect -968 -6810 -967 -6490
rect -1289 -6811 -967 -6810
rect -1579 -6938 -1452 -6922
rect -1579 -7000 -1475 -6938
rect -1180 -7000 -1076 -6811
rect -860 -6922 -813 -6378
rect -749 -6922 -733 -6378
rect -461 -6489 -357 -6111
rect -141 -6222 -94 -5678
rect -30 -6222 -14 -5678
rect 258 -5789 362 -5411
rect 578 -5522 625 -4978
rect 689 -5522 705 -4978
rect 977 -5089 1081 -4711
rect 1297 -4822 1344 -4278
rect 1408 -4822 1424 -4278
rect 1696 -4389 1800 -4011
rect 2016 -4122 2063 -3578
rect 2127 -4122 2143 -3578
rect 2415 -3689 2519 -3311
rect 2735 -3422 2782 -2878
rect 2846 -3422 2862 -2878
rect 3134 -2989 3238 -2611
rect 3454 -2722 3501 -2178
rect 3565 -2722 3581 -2178
rect 3853 -2289 3957 -1911
rect 4173 -2022 4220 -1478
rect 4284 -2022 4300 -1478
rect 4572 -1589 4676 -1211
rect 4892 -1322 4939 -778
rect 5003 -1322 5019 -778
rect 5291 -889 5395 -511
rect 5611 -622 5658 -78
rect 5722 -622 5738 -78
rect 6010 -189 6114 189
rect 6330 78 6377 622
rect 6441 78 6457 622
rect 6729 511 6833 889
rect 7049 778 7096 1322
rect 7160 778 7176 1322
rect 7049 762 7176 778
rect 7049 638 7153 762
rect 7049 622 7176 638
rect 6620 510 6942 511
rect 6620 190 6621 510
rect 6941 190 6942 510
rect 6620 189 6942 190
rect 6330 62 6457 78
rect 6330 -62 6434 62
rect 6330 -78 6457 -62
rect 5901 -190 6223 -189
rect 5901 -510 5902 -190
rect 6222 -510 6223 -190
rect 5901 -511 6223 -510
rect 5611 -638 5738 -622
rect 5611 -762 5715 -638
rect 5611 -778 5738 -762
rect 5182 -890 5504 -889
rect 5182 -1210 5183 -890
rect 5503 -1210 5504 -890
rect 5182 -1211 5504 -1210
rect 4892 -1338 5019 -1322
rect 4892 -1462 4996 -1338
rect 4892 -1478 5019 -1462
rect 4463 -1590 4785 -1589
rect 4463 -1910 4464 -1590
rect 4784 -1910 4785 -1590
rect 4463 -1911 4785 -1910
rect 4173 -2038 4300 -2022
rect 4173 -2162 4277 -2038
rect 4173 -2178 4300 -2162
rect 3744 -2290 4066 -2289
rect 3744 -2610 3745 -2290
rect 4065 -2610 4066 -2290
rect 3744 -2611 4066 -2610
rect 3454 -2738 3581 -2722
rect 3454 -2862 3558 -2738
rect 3454 -2878 3581 -2862
rect 3025 -2990 3347 -2989
rect 3025 -3310 3026 -2990
rect 3346 -3310 3347 -2990
rect 3025 -3311 3347 -3310
rect 2735 -3438 2862 -3422
rect 2735 -3562 2839 -3438
rect 2735 -3578 2862 -3562
rect 2306 -3690 2628 -3689
rect 2306 -4010 2307 -3690
rect 2627 -4010 2628 -3690
rect 2306 -4011 2628 -4010
rect 2016 -4138 2143 -4122
rect 2016 -4262 2120 -4138
rect 2016 -4278 2143 -4262
rect 1587 -4390 1909 -4389
rect 1587 -4710 1588 -4390
rect 1908 -4710 1909 -4390
rect 1587 -4711 1909 -4710
rect 1297 -4838 1424 -4822
rect 1297 -4962 1401 -4838
rect 1297 -4978 1424 -4962
rect 868 -5090 1190 -5089
rect 868 -5410 869 -5090
rect 1189 -5410 1190 -5090
rect 868 -5411 1190 -5410
rect 578 -5538 705 -5522
rect 578 -5662 682 -5538
rect 578 -5678 705 -5662
rect 149 -5790 471 -5789
rect 149 -6110 150 -5790
rect 470 -6110 471 -5790
rect 149 -6111 471 -6110
rect -141 -6238 -14 -6222
rect -141 -6362 -37 -6238
rect -141 -6378 -14 -6362
rect -570 -6490 -248 -6489
rect -570 -6810 -569 -6490
rect -249 -6810 -248 -6490
rect -570 -6811 -248 -6810
rect -860 -6938 -733 -6922
rect -860 -7000 -756 -6938
rect -461 -7000 -357 -6811
rect -141 -6922 -94 -6378
rect -30 -6922 -14 -6378
rect 258 -6489 362 -6111
rect 578 -6222 625 -5678
rect 689 -6222 705 -5678
rect 977 -5789 1081 -5411
rect 1297 -5522 1344 -4978
rect 1408 -5522 1424 -4978
rect 1696 -5089 1800 -4711
rect 2016 -4822 2063 -4278
rect 2127 -4822 2143 -4278
rect 2415 -4389 2519 -4011
rect 2735 -4122 2782 -3578
rect 2846 -4122 2862 -3578
rect 3134 -3689 3238 -3311
rect 3454 -3422 3501 -2878
rect 3565 -3422 3581 -2878
rect 3853 -2989 3957 -2611
rect 4173 -2722 4220 -2178
rect 4284 -2722 4300 -2178
rect 4572 -2289 4676 -1911
rect 4892 -2022 4939 -1478
rect 5003 -2022 5019 -1478
rect 5291 -1589 5395 -1211
rect 5611 -1322 5658 -778
rect 5722 -1322 5738 -778
rect 6010 -889 6114 -511
rect 6330 -622 6377 -78
rect 6441 -622 6457 -78
rect 6729 -189 6833 189
rect 7049 78 7096 622
rect 7160 78 7176 622
rect 7049 62 7176 78
rect 7049 -62 7153 62
rect 7049 -78 7176 -62
rect 6620 -190 6942 -189
rect 6620 -510 6621 -190
rect 6941 -510 6942 -190
rect 6620 -511 6942 -510
rect 6330 -638 6457 -622
rect 6330 -762 6434 -638
rect 6330 -778 6457 -762
rect 5901 -890 6223 -889
rect 5901 -1210 5902 -890
rect 6222 -1210 6223 -890
rect 5901 -1211 6223 -1210
rect 5611 -1338 5738 -1322
rect 5611 -1462 5715 -1338
rect 5611 -1478 5738 -1462
rect 5182 -1590 5504 -1589
rect 5182 -1910 5183 -1590
rect 5503 -1910 5504 -1590
rect 5182 -1911 5504 -1910
rect 4892 -2038 5019 -2022
rect 4892 -2162 4996 -2038
rect 4892 -2178 5019 -2162
rect 4463 -2290 4785 -2289
rect 4463 -2610 4464 -2290
rect 4784 -2610 4785 -2290
rect 4463 -2611 4785 -2610
rect 4173 -2738 4300 -2722
rect 4173 -2862 4277 -2738
rect 4173 -2878 4300 -2862
rect 3744 -2990 4066 -2989
rect 3744 -3310 3745 -2990
rect 4065 -3310 4066 -2990
rect 3744 -3311 4066 -3310
rect 3454 -3438 3581 -3422
rect 3454 -3562 3558 -3438
rect 3454 -3578 3581 -3562
rect 3025 -3690 3347 -3689
rect 3025 -4010 3026 -3690
rect 3346 -4010 3347 -3690
rect 3025 -4011 3347 -4010
rect 2735 -4138 2862 -4122
rect 2735 -4262 2839 -4138
rect 2735 -4278 2862 -4262
rect 2306 -4390 2628 -4389
rect 2306 -4710 2307 -4390
rect 2627 -4710 2628 -4390
rect 2306 -4711 2628 -4710
rect 2016 -4838 2143 -4822
rect 2016 -4962 2120 -4838
rect 2016 -4978 2143 -4962
rect 1587 -5090 1909 -5089
rect 1587 -5410 1588 -5090
rect 1908 -5410 1909 -5090
rect 1587 -5411 1909 -5410
rect 1297 -5538 1424 -5522
rect 1297 -5662 1401 -5538
rect 1297 -5678 1424 -5662
rect 868 -5790 1190 -5789
rect 868 -6110 869 -5790
rect 1189 -6110 1190 -5790
rect 868 -6111 1190 -6110
rect 578 -6238 705 -6222
rect 578 -6362 682 -6238
rect 578 -6378 705 -6362
rect 149 -6490 471 -6489
rect 149 -6810 150 -6490
rect 470 -6810 471 -6490
rect 149 -6811 471 -6810
rect -141 -6938 -14 -6922
rect -141 -7000 -37 -6938
rect 258 -7000 362 -6811
rect 578 -6922 625 -6378
rect 689 -6922 705 -6378
rect 977 -6489 1081 -6111
rect 1297 -6222 1344 -5678
rect 1408 -6222 1424 -5678
rect 1696 -5789 1800 -5411
rect 2016 -5522 2063 -4978
rect 2127 -5522 2143 -4978
rect 2415 -5089 2519 -4711
rect 2735 -4822 2782 -4278
rect 2846 -4822 2862 -4278
rect 3134 -4389 3238 -4011
rect 3454 -4122 3501 -3578
rect 3565 -4122 3581 -3578
rect 3853 -3689 3957 -3311
rect 4173 -3422 4220 -2878
rect 4284 -3422 4300 -2878
rect 4572 -2989 4676 -2611
rect 4892 -2722 4939 -2178
rect 5003 -2722 5019 -2178
rect 5291 -2289 5395 -1911
rect 5611 -2022 5658 -1478
rect 5722 -2022 5738 -1478
rect 6010 -1589 6114 -1211
rect 6330 -1322 6377 -778
rect 6441 -1322 6457 -778
rect 6729 -889 6833 -511
rect 7049 -622 7096 -78
rect 7160 -622 7176 -78
rect 7049 -638 7176 -622
rect 7049 -762 7153 -638
rect 7049 -778 7176 -762
rect 6620 -890 6942 -889
rect 6620 -1210 6621 -890
rect 6941 -1210 6942 -890
rect 6620 -1211 6942 -1210
rect 6330 -1338 6457 -1322
rect 6330 -1462 6434 -1338
rect 6330 -1478 6457 -1462
rect 5901 -1590 6223 -1589
rect 5901 -1910 5902 -1590
rect 6222 -1910 6223 -1590
rect 5901 -1911 6223 -1910
rect 5611 -2038 5738 -2022
rect 5611 -2162 5715 -2038
rect 5611 -2178 5738 -2162
rect 5182 -2290 5504 -2289
rect 5182 -2610 5183 -2290
rect 5503 -2610 5504 -2290
rect 5182 -2611 5504 -2610
rect 4892 -2738 5019 -2722
rect 4892 -2862 4996 -2738
rect 4892 -2878 5019 -2862
rect 4463 -2990 4785 -2989
rect 4463 -3310 4464 -2990
rect 4784 -3310 4785 -2990
rect 4463 -3311 4785 -3310
rect 4173 -3438 4300 -3422
rect 4173 -3562 4277 -3438
rect 4173 -3578 4300 -3562
rect 3744 -3690 4066 -3689
rect 3744 -4010 3745 -3690
rect 4065 -4010 4066 -3690
rect 3744 -4011 4066 -4010
rect 3454 -4138 3581 -4122
rect 3454 -4262 3558 -4138
rect 3454 -4278 3581 -4262
rect 3025 -4390 3347 -4389
rect 3025 -4710 3026 -4390
rect 3346 -4710 3347 -4390
rect 3025 -4711 3347 -4710
rect 2735 -4838 2862 -4822
rect 2735 -4962 2839 -4838
rect 2735 -4978 2862 -4962
rect 2306 -5090 2628 -5089
rect 2306 -5410 2307 -5090
rect 2627 -5410 2628 -5090
rect 2306 -5411 2628 -5410
rect 2016 -5538 2143 -5522
rect 2016 -5662 2120 -5538
rect 2016 -5678 2143 -5662
rect 1587 -5790 1909 -5789
rect 1587 -6110 1588 -5790
rect 1908 -6110 1909 -5790
rect 1587 -6111 1909 -6110
rect 1297 -6238 1424 -6222
rect 1297 -6362 1401 -6238
rect 1297 -6378 1424 -6362
rect 868 -6490 1190 -6489
rect 868 -6810 869 -6490
rect 1189 -6810 1190 -6490
rect 868 -6811 1190 -6810
rect 578 -6938 705 -6922
rect 578 -7000 682 -6938
rect 977 -7000 1081 -6811
rect 1297 -6922 1344 -6378
rect 1408 -6922 1424 -6378
rect 1696 -6489 1800 -6111
rect 2016 -6222 2063 -5678
rect 2127 -6222 2143 -5678
rect 2415 -5789 2519 -5411
rect 2735 -5522 2782 -4978
rect 2846 -5522 2862 -4978
rect 3134 -5089 3238 -4711
rect 3454 -4822 3501 -4278
rect 3565 -4822 3581 -4278
rect 3853 -4389 3957 -4011
rect 4173 -4122 4220 -3578
rect 4284 -4122 4300 -3578
rect 4572 -3689 4676 -3311
rect 4892 -3422 4939 -2878
rect 5003 -3422 5019 -2878
rect 5291 -2989 5395 -2611
rect 5611 -2722 5658 -2178
rect 5722 -2722 5738 -2178
rect 6010 -2289 6114 -1911
rect 6330 -2022 6377 -1478
rect 6441 -2022 6457 -1478
rect 6729 -1589 6833 -1211
rect 7049 -1322 7096 -778
rect 7160 -1322 7176 -778
rect 7049 -1338 7176 -1322
rect 7049 -1462 7153 -1338
rect 7049 -1478 7176 -1462
rect 6620 -1590 6942 -1589
rect 6620 -1910 6621 -1590
rect 6941 -1910 6942 -1590
rect 6620 -1911 6942 -1910
rect 6330 -2038 6457 -2022
rect 6330 -2162 6434 -2038
rect 6330 -2178 6457 -2162
rect 5901 -2290 6223 -2289
rect 5901 -2610 5902 -2290
rect 6222 -2610 6223 -2290
rect 5901 -2611 6223 -2610
rect 5611 -2738 5738 -2722
rect 5611 -2862 5715 -2738
rect 5611 -2878 5738 -2862
rect 5182 -2990 5504 -2989
rect 5182 -3310 5183 -2990
rect 5503 -3310 5504 -2990
rect 5182 -3311 5504 -3310
rect 4892 -3438 5019 -3422
rect 4892 -3562 4996 -3438
rect 4892 -3578 5019 -3562
rect 4463 -3690 4785 -3689
rect 4463 -4010 4464 -3690
rect 4784 -4010 4785 -3690
rect 4463 -4011 4785 -4010
rect 4173 -4138 4300 -4122
rect 4173 -4262 4277 -4138
rect 4173 -4278 4300 -4262
rect 3744 -4390 4066 -4389
rect 3744 -4710 3745 -4390
rect 4065 -4710 4066 -4390
rect 3744 -4711 4066 -4710
rect 3454 -4838 3581 -4822
rect 3454 -4962 3558 -4838
rect 3454 -4978 3581 -4962
rect 3025 -5090 3347 -5089
rect 3025 -5410 3026 -5090
rect 3346 -5410 3347 -5090
rect 3025 -5411 3347 -5410
rect 2735 -5538 2862 -5522
rect 2735 -5662 2839 -5538
rect 2735 -5678 2862 -5662
rect 2306 -5790 2628 -5789
rect 2306 -6110 2307 -5790
rect 2627 -6110 2628 -5790
rect 2306 -6111 2628 -6110
rect 2016 -6238 2143 -6222
rect 2016 -6362 2120 -6238
rect 2016 -6378 2143 -6362
rect 1587 -6490 1909 -6489
rect 1587 -6810 1588 -6490
rect 1908 -6810 1909 -6490
rect 1587 -6811 1909 -6810
rect 1297 -6938 1424 -6922
rect 1297 -7000 1401 -6938
rect 1696 -7000 1800 -6811
rect 2016 -6922 2063 -6378
rect 2127 -6922 2143 -6378
rect 2415 -6489 2519 -6111
rect 2735 -6222 2782 -5678
rect 2846 -6222 2862 -5678
rect 3134 -5789 3238 -5411
rect 3454 -5522 3501 -4978
rect 3565 -5522 3581 -4978
rect 3853 -5089 3957 -4711
rect 4173 -4822 4220 -4278
rect 4284 -4822 4300 -4278
rect 4572 -4389 4676 -4011
rect 4892 -4122 4939 -3578
rect 5003 -4122 5019 -3578
rect 5291 -3689 5395 -3311
rect 5611 -3422 5658 -2878
rect 5722 -3422 5738 -2878
rect 6010 -2989 6114 -2611
rect 6330 -2722 6377 -2178
rect 6441 -2722 6457 -2178
rect 6729 -2289 6833 -1911
rect 7049 -2022 7096 -1478
rect 7160 -2022 7176 -1478
rect 7049 -2038 7176 -2022
rect 7049 -2162 7153 -2038
rect 7049 -2178 7176 -2162
rect 6620 -2290 6942 -2289
rect 6620 -2610 6621 -2290
rect 6941 -2610 6942 -2290
rect 6620 -2611 6942 -2610
rect 6330 -2738 6457 -2722
rect 6330 -2862 6434 -2738
rect 6330 -2878 6457 -2862
rect 5901 -2990 6223 -2989
rect 5901 -3310 5902 -2990
rect 6222 -3310 6223 -2990
rect 5901 -3311 6223 -3310
rect 5611 -3438 5738 -3422
rect 5611 -3562 5715 -3438
rect 5611 -3578 5738 -3562
rect 5182 -3690 5504 -3689
rect 5182 -4010 5183 -3690
rect 5503 -4010 5504 -3690
rect 5182 -4011 5504 -4010
rect 4892 -4138 5019 -4122
rect 4892 -4262 4996 -4138
rect 4892 -4278 5019 -4262
rect 4463 -4390 4785 -4389
rect 4463 -4710 4464 -4390
rect 4784 -4710 4785 -4390
rect 4463 -4711 4785 -4710
rect 4173 -4838 4300 -4822
rect 4173 -4962 4277 -4838
rect 4173 -4978 4300 -4962
rect 3744 -5090 4066 -5089
rect 3744 -5410 3745 -5090
rect 4065 -5410 4066 -5090
rect 3744 -5411 4066 -5410
rect 3454 -5538 3581 -5522
rect 3454 -5662 3558 -5538
rect 3454 -5678 3581 -5662
rect 3025 -5790 3347 -5789
rect 3025 -6110 3026 -5790
rect 3346 -6110 3347 -5790
rect 3025 -6111 3347 -6110
rect 2735 -6238 2862 -6222
rect 2735 -6362 2839 -6238
rect 2735 -6378 2862 -6362
rect 2306 -6490 2628 -6489
rect 2306 -6810 2307 -6490
rect 2627 -6810 2628 -6490
rect 2306 -6811 2628 -6810
rect 2016 -6938 2143 -6922
rect 2016 -7000 2120 -6938
rect 2415 -7000 2519 -6811
rect 2735 -6922 2782 -6378
rect 2846 -6922 2862 -6378
rect 3134 -6489 3238 -6111
rect 3454 -6222 3501 -5678
rect 3565 -6222 3581 -5678
rect 3853 -5789 3957 -5411
rect 4173 -5522 4220 -4978
rect 4284 -5522 4300 -4978
rect 4572 -5089 4676 -4711
rect 4892 -4822 4939 -4278
rect 5003 -4822 5019 -4278
rect 5291 -4389 5395 -4011
rect 5611 -4122 5658 -3578
rect 5722 -4122 5738 -3578
rect 6010 -3689 6114 -3311
rect 6330 -3422 6377 -2878
rect 6441 -3422 6457 -2878
rect 6729 -2989 6833 -2611
rect 7049 -2722 7096 -2178
rect 7160 -2722 7176 -2178
rect 7049 -2738 7176 -2722
rect 7049 -2862 7153 -2738
rect 7049 -2878 7176 -2862
rect 6620 -2990 6942 -2989
rect 6620 -3310 6621 -2990
rect 6941 -3310 6942 -2990
rect 6620 -3311 6942 -3310
rect 6330 -3438 6457 -3422
rect 6330 -3562 6434 -3438
rect 6330 -3578 6457 -3562
rect 5901 -3690 6223 -3689
rect 5901 -4010 5902 -3690
rect 6222 -4010 6223 -3690
rect 5901 -4011 6223 -4010
rect 5611 -4138 5738 -4122
rect 5611 -4262 5715 -4138
rect 5611 -4278 5738 -4262
rect 5182 -4390 5504 -4389
rect 5182 -4710 5183 -4390
rect 5503 -4710 5504 -4390
rect 5182 -4711 5504 -4710
rect 4892 -4838 5019 -4822
rect 4892 -4962 4996 -4838
rect 4892 -4978 5019 -4962
rect 4463 -5090 4785 -5089
rect 4463 -5410 4464 -5090
rect 4784 -5410 4785 -5090
rect 4463 -5411 4785 -5410
rect 4173 -5538 4300 -5522
rect 4173 -5662 4277 -5538
rect 4173 -5678 4300 -5662
rect 3744 -5790 4066 -5789
rect 3744 -6110 3745 -5790
rect 4065 -6110 4066 -5790
rect 3744 -6111 4066 -6110
rect 3454 -6238 3581 -6222
rect 3454 -6362 3558 -6238
rect 3454 -6378 3581 -6362
rect 3025 -6490 3347 -6489
rect 3025 -6810 3026 -6490
rect 3346 -6810 3347 -6490
rect 3025 -6811 3347 -6810
rect 2735 -6938 2862 -6922
rect 2735 -7000 2839 -6938
rect 3134 -7000 3238 -6811
rect 3454 -6922 3501 -6378
rect 3565 -6922 3581 -6378
rect 3853 -6489 3957 -6111
rect 4173 -6222 4220 -5678
rect 4284 -6222 4300 -5678
rect 4572 -5789 4676 -5411
rect 4892 -5522 4939 -4978
rect 5003 -5522 5019 -4978
rect 5291 -5089 5395 -4711
rect 5611 -4822 5658 -4278
rect 5722 -4822 5738 -4278
rect 6010 -4389 6114 -4011
rect 6330 -4122 6377 -3578
rect 6441 -4122 6457 -3578
rect 6729 -3689 6833 -3311
rect 7049 -3422 7096 -2878
rect 7160 -3422 7176 -2878
rect 7049 -3438 7176 -3422
rect 7049 -3562 7153 -3438
rect 7049 -3578 7176 -3562
rect 6620 -3690 6942 -3689
rect 6620 -4010 6621 -3690
rect 6941 -4010 6942 -3690
rect 6620 -4011 6942 -4010
rect 6330 -4138 6457 -4122
rect 6330 -4262 6434 -4138
rect 6330 -4278 6457 -4262
rect 5901 -4390 6223 -4389
rect 5901 -4710 5902 -4390
rect 6222 -4710 6223 -4390
rect 5901 -4711 6223 -4710
rect 5611 -4838 5738 -4822
rect 5611 -4962 5715 -4838
rect 5611 -4978 5738 -4962
rect 5182 -5090 5504 -5089
rect 5182 -5410 5183 -5090
rect 5503 -5410 5504 -5090
rect 5182 -5411 5504 -5410
rect 4892 -5538 5019 -5522
rect 4892 -5662 4996 -5538
rect 4892 -5678 5019 -5662
rect 4463 -5790 4785 -5789
rect 4463 -6110 4464 -5790
rect 4784 -6110 4785 -5790
rect 4463 -6111 4785 -6110
rect 4173 -6238 4300 -6222
rect 4173 -6362 4277 -6238
rect 4173 -6378 4300 -6362
rect 3744 -6490 4066 -6489
rect 3744 -6810 3745 -6490
rect 4065 -6810 4066 -6490
rect 3744 -6811 4066 -6810
rect 3454 -6938 3581 -6922
rect 3454 -7000 3558 -6938
rect 3853 -7000 3957 -6811
rect 4173 -6922 4220 -6378
rect 4284 -6922 4300 -6378
rect 4572 -6489 4676 -6111
rect 4892 -6222 4939 -5678
rect 5003 -6222 5019 -5678
rect 5291 -5789 5395 -5411
rect 5611 -5522 5658 -4978
rect 5722 -5522 5738 -4978
rect 6010 -5089 6114 -4711
rect 6330 -4822 6377 -4278
rect 6441 -4822 6457 -4278
rect 6729 -4389 6833 -4011
rect 7049 -4122 7096 -3578
rect 7160 -4122 7176 -3578
rect 7049 -4138 7176 -4122
rect 7049 -4262 7153 -4138
rect 7049 -4278 7176 -4262
rect 6620 -4390 6942 -4389
rect 6620 -4710 6621 -4390
rect 6941 -4710 6942 -4390
rect 6620 -4711 6942 -4710
rect 6330 -4838 6457 -4822
rect 6330 -4962 6434 -4838
rect 6330 -4978 6457 -4962
rect 5901 -5090 6223 -5089
rect 5901 -5410 5902 -5090
rect 6222 -5410 6223 -5090
rect 5901 -5411 6223 -5410
rect 5611 -5538 5738 -5522
rect 5611 -5662 5715 -5538
rect 5611 -5678 5738 -5662
rect 5182 -5790 5504 -5789
rect 5182 -6110 5183 -5790
rect 5503 -6110 5504 -5790
rect 5182 -6111 5504 -6110
rect 4892 -6238 5019 -6222
rect 4892 -6362 4996 -6238
rect 4892 -6378 5019 -6362
rect 4463 -6490 4785 -6489
rect 4463 -6810 4464 -6490
rect 4784 -6810 4785 -6490
rect 4463 -6811 4785 -6810
rect 4173 -6938 4300 -6922
rect 4173 -7000 4277 -6938
rect 4572 -7000 4676 -6811
rect 4892 -6922 4939 -6378
rect 5003 -6922 5019 -6378
rect 5291 -6489 5395 -6111
rect 5611 -6222 5658 -5678
rect 5722 -6222 5738 -5678
rect 6010 -5789 6114 -5411
rect 6330 -5522 6377 -4978
rect 6441 -5522 6457 -4978
rect 6729 -5089 6833 -4711
rect 7049 -4822 7096 -4278
rect 7160 -4822 7176 -4278
rect 7049 -4838 7176 -4822
rect 7049 -4962 7153 -4838
rect 7049 -4978 7176 -4962
rect 6620 -5090 6942 -5089
rect 6620 -5410 6621 -5090
rect 6941 -5410 6942 -5090
rect 6620 -5411 6942 -5410
rect 6330 -5538 6457 -5522
rect 6330 -5662 6434 -5538
rect 6330 -5678 6457 -5662
rect 5901 -5790 6223 -5789
rect 5901 -6110 5902 -5790
rect 6222 -6110 6223 -5790
rect 5901 -6111 6223 -6110
rect 5611 -6238 5738 -6222
rect 5611 -6362 5715 -6238
rect 5611 -6378 5738 -6362
rect 5182 -6490 5504 -6489
rect 5182 -6810 5183 -6490
rect 5503 -6810 5504 -6490
rect 5182 -6811 5504 -6810
rect 4892 -6938 5019 -6922
rect 4892 -7000 4996 -6938
rect 5291 -7000 5395 -6811
rect 5611 -6922 5658 -6378
rect 5722 -6922 5738 -6378
rect 6010 -6489 6114 -6111
rect 6330 -6222 6377 -5678
rect 6441 -6222 6457 -5678
rect 6729 -5789 6833 -5411
rect 7049 -5522 7096 -4978
rect 7160 -5522 7176 -4978
rect 7049 -5538 7176 -5522
rect 7049 -5662 7153 -5538
rect 7049 -5678 7176 -5662
rect 6620 -5790 6942 -5789
rect 6620 -6110 6621 -5790
rect 6941 -6110 6942 -5790
rect 6620 -6111 6942 -6110
rect 6330 -6238 6457 -6222
rect 6330 -6362 6434 -6238
rect 6330 -6378 6457 -6362
rect 5901 -6490 6223 -6489
rect 5901 -6810 5902 -6490
rect 6222 -6810 6223 -6490
rect 5901 -6811 6223 -6810
rect 5611 -6938 5738 -6922
rect 5611 -7000 5715 -6938
rect 6010 -7000 6114 -6811
rect 6330 -6922 6377 -6378
rect 6441 -6922 6457 -6378
rect 6729 -6489 6833 -6111
rect 7049 -6222 7096 -5678
rect 7160 -6222 7176 -5678
rect 7049 -6238 7176 -6222
rect 7049 -6362 7153 -6238
rect 7049 -6378 7176 -6362
rect 6620 -6490 6942 -6489
rect 6620 -6810 6621 -6490
rect 6941 -6810 6942 -6490
rect 6620 -6811 6942 -6810
rect 6330 -6938 6457 -6922
rect 6330 -7000 6434 -6938
rect 6729 -7000 6833 -6811
rect 7049 -6922 7096 -6378
rect 7160 -6922 7176 -6378
rect 7049 -6938 7176 -6922
rect 7049 -7000 7153 -6938
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 6481 6350 7081 6950
string parameters w 2.00 l 2.00 val 5.36 carea 1.00 cperi 0.17 nx 20 ny 20 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
