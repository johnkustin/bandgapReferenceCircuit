magic
tech sky130A
magscale 1 2
timestamp 1620836830
<< error_p >>
rect -1688 -931 -1630 869
rect -1230 -931 -1172 869
rect -1116 -931 -1058 869
rect -658 -931 -600 869
rect -544 -931 -486 869
rect -86 -931 -28 869
rect 28 -931 86 869
rect 486 -931 544 869
rect 600 -931 658 869
rect 1058 -931 1116 869
rect 1172 -931 1230 869
rect 1630 -931 1688 869
<< nmoslvt >>
rect -1630 -931 -1230 869
rect -1058 -931 -658 869
rect -486 -931 -86 869
rect 86 -931 486 869
rect 658 -931 1058 869
rect 1230 -931 1630 869
<< ndiff >>
rect -1688 857 -1630 869
rect -1688 -919 -1676 857
rect -1642 -919 -1630 857
rect -1688 -931 -1630 -919
rect -1230 857 -1172 869
rect -1230 -919 -1218 857
rect -1184 -919 -1172 857
rect -1230 -931 -1172 -919
rect -1116 857 -1058 869
rect -1116 -919 -1104 857
rect -1070 -919 -1058 857
rect -1116 -931 -1058 -919
rect -658 857 -600 869
rect -658 -919 -646 857
rect -612 -919 -600 857
rect -658 -931 -600 -919
rect -544 857 -486 869
rect -544 -919 -532 857
rect -498 -919 -486 857
rect -544 -931 -486 -919
rect -86 857 -28 869
rect -86 -919 -74 857
rect -40 -919 -28 857
rect -86 -931 -28 -919
rect 28 857 86 869
rect 28 -919 40 857
rect 74 -919 86 857
rect 28 -931 86 -919
rect 486 857 544 869
rect 486 -919 498 857
rect 532 -919 544 857
rect 486 -931 544 -919
rect 600 857 658 869
rect 600 -919 612 857
rect 646 -919 658 857
rect 600 -931 658 -919
rect 1058 857 1116 869
rect 1058 -919 1070 857
rect 1104 -919 1116 857
rect 1058 -931 1116 -919
rect 1172 857 1230 869
rect 1172 -919 1184 857
rect 1218 -919 1230 857
rect 1172 -931 1230 -919
rect 1630 857 1688 869
rect 1630 -919 1642 857
rect 1676 -919 1688 857
rect 1630 -931 1688 -919
<< ndiffc >>
rect -1676 -919 -1642 857
rect -1218 -919 -1184 857
rect -1104 -919 -1070 857
rect -646 -919 -612 857
rect -532 -919 -498 857
rect -74 -919 -40 857
rect 40 -919 74 857
rect 498 -919 532 857
rect 612 -919 646 857
rect 1070 -919 1104 857
rect 1184 -919 1218 857
rect 1642 -919 1676 857
<< poly >>
rect -1630 941 -1230 957
rect -1630 907 -1614 941
rect -1246 907 -1230 941
rect -1630 869 -1230 907
rect -1058 941 -658 957
rect -1058 907 -1042 941
rect -674 907 -658 941
rect -1058 869 -658 907
rect -486 941 -86 957
rect -486 907 -470 941
rect -102 907 -86 941
rect -486 869 -86 907
rect 86 941 486 957
rect 86 907 102 941
rect 470 907 486 941
rect 86 869 486 907
rect 658 941 1058 957
rect 658 907 674 941
rect 1042 907 1058 941
rect 658 869 1058 907
rect 1230 941 1630 957
rect 1230 907 1246 941
rect 1614 907 1630 941
rect 1230 869 1630 907
rect -1630 -957 -1230 -931
rect -1058 -957 -658 -931
rect -486 -957 -86 -931
rect 86 -957 486 -931
rect 658 -957 1058 -931
rect 1230 -957 1630 -931
<< polycont >>
rect -1614 907 -1246 941
rect -1042 907 -674 941
rect -470 907 -102 941
rect 102 907 470 941
rect 674 907 1042 941
rect 1246 907 1614 941
<< locali >>
rect -1630 907 -1614 941
rect -1246 907 -1230 941
rect -1058 907 -1042 941
rect -674 907 -658 941
rect -486 907 -470 941
rect -102 907 -86 941
rect 86 907 102 941
rect 470 907 486 941
rect 658 907 674 941
rect 1042 907 1058 941
rect 1230 907 1246 941
rect 1614 907 1630 941
rect -1676 857 -1642 873
rect -1676 -935 -1642 -919
rect -1218 857 -1184 873
rect -1218 -935 -1184 -919
rect -1104 857 -1070 873
rect -1104 -935 -1070 -919
rect -646 857 -612 873
rect -646 -935 -612 -919
rect -532 857 -498 873
rect -532 -935 -498 -919
rect -74 857 -40 873
rect -74 -935 -40 -919
rect 40 857 74 873
rect 40 -935 74 -919
rect 498 857 532 873
rect 498 -935 532 -919
rect 612 857 646 873
rect 612 -935 646 -919
rect 1070 857 1104 873
rect 1070 -935 1104 -919
rect 1184 857 1218 873
rect 1184 -935 1218 -919
rect 1642 857 1676 873
rect 1642 -935 1676 -919
<< viali >>
rect -1522 907 -1338 941
rect -950 907 -766 941
rect -378 907 -194 941
rect 194 907 378 941
rect 766 907 950 941
rect 1338 907 1522 941
rect -1676 -919 -1642 857
rect -1218 -919 -1184 857
rect -1104 -919 -1070 857
rect -646 -919 -612 857
rect -532 -919 -498 857
rect -74 -919 -40 857
rect 40 -919 74 857
rect 498 -919 532 857
rect 612 -919 646 857
rect 1070 -919 1104 857
rect 1184 -919 1218 857
rect 1642 -919 1676 857
<< metal1 >>
rect -1534 941 -1326 947
rect -1534 907 -1522 941
rect -1338 907 -1326 941
rect -1534 901 -1326 907
rect -962 941 -754 947
rect -962 907 -950 941
rect -766 907 -754 941
rect -962 901 -754 907
rect -390 941 -182 947
rect -390 907 -378 941
rect -194 907 -182 941
rect -390 901 -182 907
rect 182 941 390 947
rect 182 907 194 941
rect 378 907 390 941
rect 182 901 390 907
rect 754 941 962 947
rect 754 907 766 941
rect 950 907 962 941
rect 754 901 962 907
rect 1326 941 1534 947
rect 1326 907 1338 941
rect 1522 907 1534 941
rect 1326 901 1534 907
rect -1682 857 -1636 869
rect -1682 -919 -1676 857
rect -1642 -919 -1636 857
rect -1682 -931 -1636 -919
rect -1224 857 -1178 869
rect -1224 -919 -1218 857
rect -1184 -919 -1178 857
rect -1224 -931 -1178 -919
rect -1110 857 -1064 869
rect -1110 -919 -1104 857
rect -1070 -919 -1064 857
rect -1110 -931 -1064 -919
rect -652 857 -606 869
rect -652 -919 -646 857
rect -612 -919 -606 857
rect -652 -931 -606 -919
rect -538 857 -492 869
rect -538 -919 -532 857
rect -498 -919 -492 857
rect -538 -931 -492 -919
rect -80 857 -34 869
rect -80 -919 -74 857
rect -40 -919 -34 857
rect -80 -931 -34 -919
rect 34 857 80 869
rect 34 -919 40 857
rect 74 -919 80 857
rect 34 -931 80 -919
rect 492 857 538 869
rect 492 -919 498 857
rect 532 -919 538 857
rect 492 -931 538 -919
rect 606 857 652 869
rect 606 -919 612 857
rect 646 -919 652 857
rect 606 -931 652 -919
rect 1064 857 1110 869
rect 1064 -919 1070 857
rect 1104 -919 1110 857
rect 1064 -931 1110 -919
rect 1178 857 1224 869
rect 1178 -919 1184 857
rect 1218 -919 1224 857
rect 1178 -931 1224 -919
rect 1636 857 1682 869
rect 1636 -919 1642 857
rect 1676 -919 1682 857
rect 1636 -931 1682 -919
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 9 l 2 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
