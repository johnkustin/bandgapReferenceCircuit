magic
tech sky130A
magscale 1 2
timestamp 1620793367
<< xpolycontact >>
rect 10102 6600 10172 7032
rect 10902 6600 10972 7032
rect 12102 6600 12172 7032
<< locali >>
rect 8400 -5000 8600 5300
rect 9500 -5000 9900 5200
rect 10800 -5000 11200 5200
rect 12100 -5000 12500 5200
rect 13300 -5000 13800 5300
rect 14600 5100 14800 5300
rect 14600 4300 14700 5100
rect 14600 -5000 14800 4300
<< viali >>
rect 10118 6618 10156 7015
rect 10918 6618 10956 7015
rect 12118 6618 12156 7015
rect 14700 4300 14800 5100
<< metal1 >>
rect 8102 8196 8172 8216
rect 8102 8144 8108 8196
rect 8160 8144 8172 8196
rect 8102 7784 8172 8144
rect 8502 7864 8572 8216
rect 8502 7812 8508 7864
rect 8560 7812 8572 7864
rect 8502 7784 8572 7812
rect 8902 8196 8972 8216
rect 8902 8144 8908 8196
rect 8960 8144 8972 8196
rect 8902 7784 8972 8144
rect 9302 7864 9372 8216
rect 9302 7812 9308 7864
rect 9360 7812 9372 7864
rect 9302 7784 9372 7812
rect 9702 8196 9772 8216
rect 9702 8144 9708 8196
rect 9760 8144 9772 8196
rect 9702 7784 9772 8144
rect 10102 7864 10172 8216
rect 10102 7812 10108 7864
rect 10160 7812 10172 7864
rect 10102 7784 10172 7812
rect 10502 8196 10572 8216
rect 10502 8144 10508 8196
rect 10560 8144 10572 8196
rect 10502 7784 10572 8144
rect 10902 7864 10972 8216
rect 10902 7812 10908 7864
rect 10960 7812 10972 7864
rect 10902 7784 10972 7812
rect 8502 7448 8572 7468
rect 8502 7396 8510 7448
rect 8562 7396 8572 7448
rect 8102 5900 8172 7032
rect 8502 6492 8572 7396
rect 11302 7448 11372 8216
rect 11702 8196 11772 8216
rect 11702 8144 11708 8196
rect 11760 8144 11772 8196
rect 11702 7784 11772 8144
rect 12102 7864 12172 8216
rect 12102 7812 12108 7864
rect 12160 7812 12172 7864
rect 12102 7784 12172 7812
rect 12502 8196 12572 8202
rect 12502 8144 12508 8196
rect 12560 8144 12572 8196
rect 12502 7754 12572 8144
rect 12902 7864 12972 8186
rect 12902 7812 12908 7864
rect 12960 7812 12972 7864
rect 12902 7754 12972 7812
rect 11302 7396 11308 7448
rect 11360 7396 11372 7448
rect 11302 7368 11372 7396
rect 8902 6680 8972 7032
rect 8902 6628 8908 6680
rect 8960 6628 8972 6680
rect 8902 6600 8972 6628
rect 9302 7012 9372 7032
rect 9302 6960 9308 7012
rect 9360 6960 9372 7012
rect 9302 6600 9372 6960
rect 9702 6680 9772 7032
rect 9702 6628 9708 6680
rect 9760 6628 9772 6680
rect 9702 6600 9772 6628
rect 10102 7015 10172 7032
rect 10102 7012 10118 7015
rect 10156 7012 10172 7015
rect 10102 6960 10108 7012
rect 10160 6960 10172 7012
rect 10102 6618 10118 6960
rect 10156 6618 10172 6960
rect 10102 6600 10172 6618
rect 10502 6680 10572 7032
rect 10502 6628 10508 6680
rect 10560 6628 10572 6680
rect 10502 6600 10572 6628
rect 10902 7015 10972 7032
rect 10902 7012 10918 7015
rect 10956 7012 10972 7015
rect 10902 6960 10908 7012
rect 10960 6960 10972 7012
rect 10902 6618 10918 6960
rect 10956 6618 10972 6960
rect 10902 6600 10972 6618
rect 11302 6500 11372 7032
rect 11702 6680 11772 7032
rect 11702 6628 11708 6680
rect 11760 6628 11772 6680
rect 11702 6600 11772 6628
rect 12102 7015 12172 7032
rect 12102 7012 12118 7015
rect 12156 7012 12172 7015
rect 12102 6960 12108 7012
rect 12160 6960 12172 7012
rect 12102 6618 12118 6960
rect 12156 6618 12172 6960
rect 12502 6886 12572 7248
rect 12502 6834 12508 6886
rect 12560 6834 12572 6886
rect 12502 6816 12572 6834
rect 12902 7228 12972 7248
rect 12902 7176 12908 7228
rect 12960 7176 12972 7228
rect 12902 6816 12972 7176
rect 12102 6600 12172 6618
rect 8444 6486 8630 6492
rect 8444 6300 8450 6486
rect 8624 6300 8630 6486
rect 8444 6294 8630 6300
rect 8102 5686 9400 5900
rect 8102 5500 8450 5686
rect 8624 5500 9400 5686
rect 8102 4300 9400 5500
rect 11000 5000 11700 6500
rect 14800 5200 15400 5300
rect 14600 5100 15400 5200
rect 10000 3900 14500 5000
rect 14600 4300 14700 5100
rect 14800 4300 15000 5100
rect 14600 4100 15000 4300
rect 15300 4100 15400 5100
rect 14800 3900 15400 4100
rect 10000 3700 14600 3900
rect 8700 -4700 14600 3700
<< via1 >>
rect 8108 8144 8160 8196
rect 8508 7812 8560 7864
rect 8908 8144 8960 8196
rect 9308 7812 9360 7864
rect 9708 8144 9760 8196
rect 10108 7812 10160 7864
rect 10508 8144 10560 8196
rect 10908 7812 10960 7864
rect 8510 7396 8562 7448
rect 11708 8144 11760 8196
rect 12108 7812 12160 7864
rect 12508 8144 12560 8196
rect 12908 7812 12960 7864
rect 11308 7396 11360 7448
rect 8908 6628 8960 6680
rect 9308 6960 9360 7012
rect 9708 6628 9760 6680
rect 10108 6960 10118 7012
rect 10118 6960 10156 7012
rect 10156 6960 10160 7012
rect 10508 6628 10560 6680
rect 10908 6960 10918 7012
rect 10918 6960 10956 7012
rect 10956 6960 10960 7012
rect 11708 6628 11760 6680
rect 12108 6960 12118 7012
rect 12118 6960 12156 7012
rect 12156 6960 12160 7012
rect 12508 6834 12560 6886
rect 12908 7176 12960 7228
rect 8450 6300 8624 6486
rect 8450 5500 8624 5686
rect 15000 4100 15300 5100
<< metal2 >>
rect 8090 8196 8990 8216
rect 8090 8144 8108 8196
rect 8160 8144 8908 8196
rect 8960 8144 8990 8196
rect 8090 8116 8990 8144
rect 9690 8196 10590 8216
rect 9690 8144 9708 8196
rect 9760 8144 10508 8196
rect 10560 8144 10590 8196
rect 9690 8116 10590 8144
rect 11690 8196 12572 8216
rect 11690 8144 11708 8196
rect 11760 8144 12508 8196
rect 12560 8144 12572 8196
rect 11690 8116 12572 8144
rect 8490 7864 9390 7884
rect 8490 7812 8508 7864
rect 8560 7812 9308 7864
rect 9360 7812 9390 7864
rect 8490 7784 9390 7812
rect 10090 7864 10990 7884
rect 10090 7812 10108 7864
rect 10160 7812 10908 7864
rect 10960 7812 10990 7864
rect 10090 7784 10990 7812
rect 12090 7864 12972 7884
rect 12090 7812 12108 7864
rect 12160 7812 12908 7864
rect 12960 7812 12972 7864
rect 12090 7784 12972 7812
rect 8500 7448 11390 7468
rect 8500 7396 8510 7448
rect 8562 7396 11308 7448
rect 11360 7396 11390 7448
rect 8500 7368 11390 7396
rect 14900 7248 15400 8790
rect 12902 7228 15400 7248
rect 12902 7176 12908 7228
rect 12960 7176 15400 7228
rect 12902 7148 12972 7176
rect 9290 7012 10190 7032
rect 9290 6960 9308 7012
rect 9360 6960 10108 7012
rect 10160 6960 10190 7012
rect 9290 6932 10190 6960
rect 10890 7012 12190 7032
rect 10890 6960 10908 7012
rect 10960 6960 12108 7012
rect 12160 6960 12190 7012
rect 10890 6932 12190 6960
rect 12502 6886 12572 6906
rect 14900 6886 15400 7176
rect 12502 6834 12508 6886
rect 12560 6834 15400 6886
rect 12502 6806 15400 6834
rect 8890 6680 9790 6700
rect 8890 6628 8908 6680
rect 8960 6628 9708 6680
rect 9760 6628 9790 6680
rect 8890 6600 9790 6628
rect 10490 6680 11790 6700
rect 10490 6628 10508 6680
rect 10560 6628 11708 6680
rect 11760 6628 11790 6680
rect 10490 6600 11790 6628
rect 8444 6486 8630 6492
rect 8444 6300 8450 6486
rect 8624 6300 8630 6486
rect 8444 6294 8630 6300
rect 8444 5686 8630 5692
rect 8444 5500 8450 5686
rect 8624 5500 8630 5686
rect 8444 5494 8630 5500
rect 14900 5100 15400 6806
rect 14900 4100 15000 5100
rect 15300 4100 15400 5100
rect 14900 4000 15400 4100
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_2
timestamp 1620683974
transform 1 0 8937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_3
timestamp 1620683974
transform 1 0 9337 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_4
timestamp 1620683974
transform 1 0 9737 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_1
timestamp 1620683974
transform 1 0 8537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_0
timestamp 1620683974
transform 1 0 8137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_8
timestamp 1620683974
transform 1 0 11337 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_5
timestamp 1620683974
transform 1 0 10137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_6
timestamp 1620683974
transform 1 0 10537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_7
timestamp 1620683974
transform 1 0 10937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_8LEWSR  sky130_fd_pr__res_xhigh_po_0p35_8LEWSR_1
timestamp 1620793367
transform 1 0 12937 0 1 7501
box -37 -685 37 685
use sky130_fd_pr__res_xhigh_po_0p35_8LEWSR  sky130_fd_pr__res_xhigh_po_0p35_8LEWSR_0
timestamp 1620793367
transform 1 0 12537 0 1 7501
box -37 -685 37 685
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_9
timestamp 1620683974
transform 1 0 11737 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_10
timestamp 1620683974
transform 1 0 12137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 7 1288
timestamp 1620596431
transform 1 0 8374 0 1 -5042
box 26 26 1314 1314
<< labels >>
flabel metal2 14900 6100 15400 6400 1 FreeSans 1600 0 0 0 GND!
port 2 n
flabel metal1 11240 5360 11440 5580 1 FreeSans 800 0 0 0 Vbneg
flabel metal1 8700 5500 9000 5800 1 FreeSans 1600 0 0 0 Va
port 1 n
flabel via1 8458 6304 8606 6468 1 FreeSans 1600 0 0 0 Vb
port 0 n
<< end >>
