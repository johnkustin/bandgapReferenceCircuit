magic
tech sky130A
magscale 1 2
timestamp 1621270775
<< xpolycontact >>
rect -6829 3152 -6259 3584
rect -6829 -3584 -6259 -3152
rect -6011 3152 -5441 3584
rect -6011 -3584 -5441 -3152
rect -5193 3152 -4623 3584
rect -5193 -3584 -4623 -3152
rect -4375 3152 -3805 3584
rect -4375 -3584 -3805 -3152
rect -3557 3152 -2987 3584
rect -3557 -3584 -2987 -3152
rect -2739 3152 -2169 3584
rect -2739 -3584 -2169 -3152
rect -1921 3152 -1351 3584
rect -1921 -3584 -1351 -3152
rect -1103 3152 -533 3584
rect -1103 -3584 -533 -3152
rect -285 3152 285 3584
rect -285 -3584 285 -3152
rect 533 3152 1103 3584
rect 533 -3584 1103 -3152
rect 1351 3152 1921 3584
rect 1351 -3584 1921 -3152
rect 2169 3152 2739 3584
rect 2169 -3584 2739 -3152
rect 2987 3152 3557 3584
rect 2987 -3584 3557 -3152
rect 3805 3152 4375 3584
rect 3805 -3584 4375 -3152
rect 4623 3152 5193 3584
rect 4623 -3584 5193 -3152
rect 5441 3152 6011 3584
rect 5441 -3584 6011 -3152
rect 6259 3152 6829 3584
rect 6259 -3584 6829 -3152
<< xpolyres >>
rect -6829 -3152 -6259 3152
rect -6011 -3152 -5441 3152
rect -5193 -3152 -4623 3152
rect -4375 -3152 -3805 3152
rect -3557 -3152 -2987 3152
rect -2739 -3152 -2169 3152
rect -1921 -3152 -1351 3152
rect -1103 -3152 -533 3152
rect -285 -3152 285 3152
rect 533 -3152 1103 3152
rect 1351 -3152 1921 3152
rect 2169 -3152 2739 3152
rect 2987 -3152 3557 3152
rect 3805 -3152 4375 3152
rect 4623 -3152 5193 3152
rect 5441 -3152 6011 3152
rect 6259 -3152 6829 3152
<< viali >>
rect -6813 3169 -6275 3566
rect -5995 3169 -5457 3566
rect -5177 3169 -4639 3566
rect -4359 3169 -3821 3566
rect -3541 3169 -3003 3566
rect -2723 3169 -2185 3566
rect -1905 3169 -1367 3566
rect -1087 3169 -549 3566
rect -269 3169 269 3566
rect 549 3169 1087 3566
rect 1367 3169 1905 3566
rect 2185 3169 2723 3566
rect 3003 3169 3541 3566
rect 3821 3169 4359 3566
rect 4639 3169 5177 3566
rect 5457 3169 5995 3566
rect 6275 3169 6813 3566
rect -6813 -3566 -6275 -3169
rect -5995 -3566 -5457 -3169
rect -5177 -3566 -4639 -3169
rect -4359 -3566 -3821 -3169
rect -3541 -3566 -3003 -3169
rect -2723 -3566 -2185 -3169
rect -1905 -3566 -1367 -3169
rect -1087 -3566 -549 -3169
rect -269 -3566 269 -3169
rect 549 -3566 1087 -3169
rect 1367 -3566 1905 -3169
rect 2185 -3566 2723 -3169
rect 3003 -3566 3541 -3169
rect 3821 -3566 4359 -3169
rect 4639 -3566 5177 -3169
rect 5457 -3566 5995 -3169
rect 6275 -3566 6813 -3169
<< metal1 >>
rect -6825 3566 -6263 3572
rect -6825 3169 -6813 3566
rect -6275 3169 -6263 3566
rect -6825 3163 -6263 3169
rect -6007 3566 -5445 3572
rect -6007 3169 -5995 3566
rect -5457 3169 -5445 3566
rect -6007 3163 -5445 3169
rect -5189 3566 -4627 3572
rect -5189 3169 -5177 3566
rect -4639 3169 -4627 3566
rect -5189 3163 -4627 3169
rect -4371 3566 -3809 3572
rect -4371 3169 -4359 3566
rect -3821 3169 -3809 3566
rect -4371 3163 -3809 3169
rect -3553 3566 -2991 3572
rect -3553 3169 -3541 3566
rect -3003 3169 -2991 3566
rect -3553 3163 -2991 3169
rect -2735 3566 -2173 3572
rect -2735 3169 -2723 3566
rect -2185 3169 -2173 3566
rect -2735 3163 -2173 3169
rect -1917 3566 -1355 3572
rect -1917 3169 -1905 3566
rect -1367 3169 -1355 3566
rect -1917 3163 -1355 3169
rect -1099 3566 -537 3572
rect -1099 3169 -1087 3566
rect -549 3169 -537 3566
rect -1099 3163 -537 3169
rect -281 3566 281 3572
rect -281 3169 -269 3566
rect 269 3169 281 3566
rect -281 3163 281 3169
rect 537 3566 1099 3572
rect 537 3169 549 3566
rect 1087 3169 1099 3566
rect 537 3163 1099 3169
rect 1355 3566 1917 3572
rect 1355 3169 1367 3566
rect 1905 3169 1917 3566
rect 1355 3163 1917 3169
rect 2173 3566 2735 3572
rect 2173 3169 2185 3566
rect 2723 3169 2735 3566
rect 2173 3163 2735 3169
rect 2991 3566 3553 3572
rect 2991 3169 3003 3566
rect 3541 3169 3553 3566
rect 2991 3163 3553 3169
rect 3809 3566 4371 3572
rect 3809 3169 3821 3566
rect 4359 3169 4371 3566
rect 3809 3163 4371 3169
rect 4627 3566 5189 3572
rect 4627 3169 4639 3566
rect 5177 3169 5189 3566
rect 4627 3163 5189 3169
rect 5445 3566 6007 3572
rect 5445 3169 5457 3566
rect 5995 3169 6007 3566
rect 5445 3163 6007 3169
rect 6263 3566 6825 3572
rect 6263 3169 6275 3566
rect 6813 3169 6825 3566
rect 6263 3163 6825 3169
rect -6825 -3169 -6263 -3163
rect -6825 -3566 -6813 -3169
rect -6275 -3566 -6263 -3169
rect -6825 -3572 -6263 -3566
rect -6007 -3169 -5445 -3163
rect -6007 -3566 -5995 -3169
rect -5457 -3566 -5445 -3169
rect -6007 -3572 -5445 -3566
rect -5189 -3169 -4627 -3163
rect -5189 -3566 -5177 -3169
rect -4639 -3566 -4627 -3169
rect -5189 -3572 -4627 -3566
rect -4371 -3169 -3809 -3163
rect -4371 -3566 -4359 -3169
rect -3821 -3566 -3809 -3169
rect -4371 -3572 -3809 -3566
rect -3553 -3169 -2991 -3163
rect -3553 -3566 -3541 -3169
rect -3003 -3566 -2991 -3169
rect -3553 -3572 -2991 -3566
rect -2735 -3169 -2173 -3163
rect -2735 -3566 -2723 -3169
rect -2185 -3566 -2173 -3169
rect -2735 -3572 -2173 -3566
rect -1917 -3169 -1355 -3163
rect -1917 -3566 -1905 -3169
rect -1367 -3566 -1355 -3169
rect -1917 -3572 -1355 -3566
rect -1099 -3169 -537 -3163
rect -1099 -3566 -1087 -3169
rect -549 -3566 -537 -3169
rect -1099 -3572 -537 -3566
rect -281 -3169 281 -3163
rect -281 -3566 -269 -3169
rect 269 -3566 281 -3169
rect -281 -3572 281 -3566
rect 537 -3169 1099 -3163
rect 537 -3566 549 -3169
rect 1087 -3566 1099 -3169
rect 537 -3572 1099 -3566
rect 1355 -3169 1917 -3163
rect 1355 -3566 1367 -3169
rect 1905 -3566 1917 -3169
rect 1355 -3572 1917 -3566
rect 2173 -3169 2735 -3163
rect 2173 -3566 2185 -3169
rect 2723 -3566 2735 -3169
rect 2173 -3572 2735 -3566
rect 2991 -3169 3553 -3163
rect 2991 -3566 3003 -3169
rect 3541 -3566 3553 -3169
rect 2991 -3572 3553 -3566
rect 3809 -3169 4371 -3163
rect 3809 -3566 3821 -3169
rect 4359 -3566 4371 -3169
rect 3809 -3572 4371 -3566
rect 4627 -3169 5189 -3163
rect 4627 -3566 4639 -3169
rect 5177 -3566 5189 -3169
rect 4627 -3572 5189 -3566
rect 5445 -3169 6007 -3163
rect 5445 -3566 5457 -3169
rect 5995 -3566 6007 -3169
rect 5445 -3572 6007 -3566
rect 6263 -3169 6825 -3163
rect 6263 -3566 6275 -3169
rect 6813 -3566 6825 -3169
rect 6263 -3572 6825 -3566
<< res2p85 >>
rect -6831 -3154 -6257 3154
rect -6013 -3154 -5439 3154
rect -5195 -3154 -4621 3154
rect -4377 -3154 -3803 3154
rect -3559 -3154 -2985 3154
rect -2741 -3154 -2167 3154
rect -1923 -3154 -1349 3154
rect -1105 -3154 -531 3154
rect -287 -3154 287 3154
rect 531 -3154 1105 3154
rect 1349 -3154 1923 3154
rect 2167 -3154 2741 3154
rect 2985 -3154 3559 3154
rect 3803 -3154 4377 3154
rect 4621 -3154 5195 3154
rect 5439 -3154 6013 3154
rect 6257 -3154 6831 3154
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_2p85
string parameters w 2.850 l 31.52 m 1 nx 17 wmin 2.850 lmin 0.50 rho 2000 val 22.132k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 2.850 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
