magic
tech sky130A
magscale 1 2
timestamp 1620244706
<< nwell >>
rect -396 -84467 396 84467
<< pmoslvt >>
rect -200 84048 200 84248
rect -200 83612 200 83812
rect -200 83176 200 83376
rect -200 82740 200 82940
rect -200 82304 200 82504
rect -200 81868 200 82068
rect -200 81432 200 81632
rect -200 80996 200 81196
rect -200 80560 200 80760
rect -200 80124 200 80324
rect -200 79688 200 79888
rect -200 79252 200 79452
rect -200 78816 200 79016
rect -200 78380 200 78580
rect -200 77944 200 78144
rect -200 77508 200 77708
rect -200 77072 200 77272
rect -200 76636 200 76836
rect -200 76200 200 76400
rect -200 75764 200 75964
rect -200 75328 200 75528
rect -200 74892 200 75092
rect -200 74456 200 74656
rect -200 74020 200 74220
rect -200 73584 200 73784
rect -200 73148 200 73348
rect -200 72712 200 72912
rect -200 72276 200 72476
rect -200 71840 200 72040
rect -200 71404 200 71604
rect -200 70968 200 71168
rect -200 70532 200 70732
rect -200 70096 200 70296
rect -200 69660 200 69860
rect -200 69224 200 69424
rect -200 68788 200 68988
rect -200 68352 200 68552
rect -200 67916 200 68116
rect -200 67480 200 67680
rect -200 67044 200 67244
rect -200 66608 200 66808
rect -200 66172 200 66372
rect -200 65736 200 65936
rect -200 65300 200 65500
rect -200 64864 200 65064
rect -200 64428 200 64628
rect -200 63992 200 64192
rect -200 63556 200 63756
rect -200 63120 200 63320
rect -200 62684 200 62884
rect -200 62248 200 62448
rect -200 61812 200 62012
rect -200 61376 200 61576
rect -200 60940 200 61140
rect -200 60504 200 60704
rect -200 60068 200 60268
rect -200 59632 200 59832
rect -200 59196 200 59396
rect -200 58760 200 58960
rect -200 58324 200 58524
rect -200 57888 200 58088
rect -200 57452 200 57652
rect -200 57016 200 57216
rect -200 56580 200 56780
rect -200 56144 200 56344
rect -200 55708 200 55908
rect -200 55272 200 55472
rect -200 54836 200 55036
rect -200 54400 200 54600
rect -200 53964 200 54164
rect -200 53528 200 53728
rect -200 53092 200 53292
rect -200 52656 200 52856
rect -200 52220 200 52420
rect -200 51784 200 51984
rect -200 51348 200 51548
rect -200 50912 200 51112
rect -200 50476 200 50676
rect -200 50040 200 50240
rect -200 49604 200 49804
rect -200 49168 200 49368
rect -200 48732 200 48932
rect -200 48296 200 48496
rect -200 47860 200 48060
rect -200 47424 200 47624
rect -200 46988 200 47188
rect -200 46552 200 46752
rect -200 46116 200 46316
rect -200 45680 200 45880
rect -200 45244 200 45444
rect -200 44808 200 45008
rect -200 44372 200 44572
rect -200 43936 200 44136
rect -200 43500 200 43700
rect -200 43064 200 43264
rect -200 42628 200 42828
rect -200 42192 200 42392
rect -200 41756 200 41956
rect -200 41320 200 41520
rect -200 40884 200 41084
rect -200 40448 200 40648
rect -200 40012 200 40212
rect -200 39576 200 39776
rect -200 39140 200 39340
rect -200 38704 200 38904
rect -200 38268 200 38468
rect -200 37832 200 38032
rect -200 37396 200 37596
rect -200 36960 200 37160
rect -200 36524 200 36724
rect -200 36088 200 36288
rect -200 35652 200 35852
rect -200 35216 200 35416
rect -200 34780 200 34980
rect -200 34344 200 34544
rect -200 33908 200 34108
rect -200 33472 200 33672
rect -200 33036 200 33236
rect -200 32600 200 32800
rect -200 32164 200 32364
rect -200 31728 200 31928
rect -200 31292 200 31492
rect -200 30856 200 31056
rect -200 30420 200 30620
rect -200 29984 200 30184
rect -200 29548 200 29748
rect -200 29112 200 29312
rect -200 28676 200 28876
rect -200 28240 200 28440
rect -200 27804 200 28004
rect -200 27368 200 27568
rect -200 26932 200 27132
rect -200 26496 200 26696
rect -200 26060 200 26260
rect -200 25624 200 25824
rect -200 25188 200 25388
rect -200 24752 200 24952
rect -200 24316 200 24516
rect -200 23880 200 24080
rect -200 23444 200 23644
rect -200 23008 200 23208
rect -200 22572 200 22772
rect -200 22136 200 22336
rect -200 21700 200 21900
rect -200 21264 200 21464
rect -200 20828 200 21028
rect -200 20392 200 20592
rect -200 19956 200 20156
rect -200 19520 200 19720
rect -200 19084 200 19284
rect -200 18648 200 18848
rect -200 18212 200 18412
rect -200 17776 200 17976
rect -200 17340 200 17540
rect -200 16904 200 17104
rect -200 16468 200 16668
rect -200 16032 200 16232
rect -200 15596 200 15796
rect -200 15160 200 15360
rect -200 14724 200 14924
rect -200 14288 200 14488
rect -200 13852 200 14052
rect -200 13416 200 13616
rect -200 12980 200 13180
rect -200 12544 200 12744
rect -200 12108 200 12308
rect -200 11672 200 11872
rect -200 11236 200 11436
rect -200 10800 200 11000
rect -200 10364 200 10564
rect -200 9928 200 10128
rect -200 9492 200 9692
rect -200 9056 200 9256
rect -200 8620 200 8820
rect -200 8184 200 8384
rect -200 7748 200 7948
rect -200 7312 200 7512
rect -200 6876 200 7076
rect -200 6440 200 6640
rect -200 6004 200 6204
rect -200 5568 200 5768
rect -200 5132 200 5332
rect -200 4696 200 4896
rect -200 4260 200 4460
rect -200 3824 200 4024
rect -200 3388 200 3588
rect -200 2952 200 3152
rect -200 2516 200 2716
rect -200 2080 200 2280
rect -200 1644 200 1844
rect -200 1208 200 1408
rect -200 772 200 972
rect -200 336 200 536
rect -200 -100 200 100
rect -200 -536 200 -336
rect -200 -972 200 -772
rect -200 -1408 200 -1208
rect -200 -1844 200 -1644
rect -200 -2280 200 -2080
rect -200 -2716 200 -2516
rect -200 -3152 200 -2952
rect -200 -3588 200 -3388
rect -200 -4024 200 -3824
rect -200 -4460 200 -4260
rect -200 -4896 200 -4696
rect -200 -5332 200 -5132
rect -200 -5768 200 -5568
rect -200 -6204 200 -6004
rect -200 -6640 200 -6440
rect -200 -7076 200 -6876
rect -200 -7512 200 -7312
rect -200 -7948 200 -7748
rect -200 -8384 200 -8184
rect -200 -8820 200 -8620
rect -200 -9256 200 -9056
rect -200 -9692 200 -9492
rect -200 -10128 200 -9928
rect -200 -10564 200 -10364
rect -200 -11000 200 -10800
rect -200 -11436 200 -11236
rect -200 -11872 200 -11672
rect -200 -12308 200 -12108
rect -200 -12744 200 -12544
rect -200 -13180 200 -12980
rect -200 -13616 200 -13416
rect -200 -14052 200 -13852
rect -200 -14488 200 -14288
rect -200 -14924 200 -14724
rect -200 -15360 200 -15160
rect -200 -15796 200 -15596
rect -200 -16232 200 -16032
rect -200 -16668 200 -16468
rect -200 -17104 200 -16904
rect -200 -17540 200 -17340
rect -200 -17976 200 -17776
rect -200 -18412 200 -18212
rect -200 -18848 200 -18648
rect -200 -19284 200 -19084
rect -200 -19720 200 -19520
rect -200 -20156 200 -19956
rect -200 -20592 200 -20392
rect -200 -21028 200 -20828
rect -200 -21464 200 -21264
rect -200 -21900 200 -21700
rect -200 -22336 200 -22136
rect -200 -22772 200 -22572
rect -200 -23208 200 -23008
rect -200 -23644 200 -23444
rect -200 -24080 200 -23880
rect -200 -24516 200 -24316
rect -200 -24952 200 -24752
rect -200 -25388 200 -25188
rect -200 -25824 200 -25624
rect -200 -26260 200 -26060
rect -200 -26696 200 -26496
rect -200 -27132 200 -26932
rect -200 -27568 200 -27368
rect -200 -28004 200 -27804
rect -200 -28440 200 -28240
rect -200 -28876 200 -28676
rect -200 -29312 200 -29112
rect -200 -29748 200 -29548
rect -200 -30184 200 -29984
rect -200 -30620 200 -30420
rect -200 -31056 200 -30856
rect -200 -31492 200 -31292
rect -200 -31928 200 -31728
rect -200 -32364 200 -32164
rect -200 -32800 200 -32600
rect -200 -33236 200 -33036
rect -200 -33672 200 -33472
rect -200 -34108 200 -33908
rect -200 -34544 200 -34344
rect -200 -34980 200 -34780
rect -200 -35416 200 -35216
rect -200 -35852 200 -35652
rect -200 -36288 200 -36088
rect -200 -36724 200 -36524
rect -200 -37160 200 -36960
rect -200 -37596 200 -37396
rect -200 -38032 200 -37832
rect -200 -38468 200 -38268
rect -200 -38904 200 -38704
rect -200 -39340 200 -39140
rect -200 -39776 200 -39576
rect -200 -40212 200 -40012
rect -200 -40648 200 -40448
rect -200 -41084 200 -40884
rect -200 -41520 200 -41320
rect -200 -41956 200 -41756
rect -200 -42392 200 -42192
rect -200 -42828 200 -42628
rect -200 -43264 200 -43064
rect -200 -43700 200 -43500
rect -200 -44136 200 -43936
rect -200 -44572 200 -44372
rect -200 -45008 200 -44808
rect -200 -45444 200 -45244
rect -200 -45880 200 -45680
rect -200 -46316 200 -46116
rect -200 -46752 200 -46552
rect -200 -47188 200 -46988
rect -200 -47624 200 -47424
rect -200 -48060 200 -47860
rect -200 -48496 200 -48296
rect -200 -48932 200 -48732
rect -200 -49368 200 -49168
rect -200 -49804 200 -49604
rect -200 -50240 200 -50040
rect -200 -50676 200 -50476
rect -200 -51112 200 -50912
rect -200 -51548 200 -51348
rect -200 -51984 200 -51784
rect -200 -52420 200 -52220
rect -200 -52856 200 -52656
rect -200 -53292 200 -53092
rect -200 -53728 200 -53528
rect -200 -54164 200 -53964
rect -200 -54600 200 -54400
rect -200 -55036 200 -54836
rect -200 -55472 200 -55272
rect -200 -55908 200 -55708
rect -200 -56344 200 -56144
rect -200 -56780 200 -56580
rect -200 -57216 200 -57016
rect -200 -57652 200 -57452
rect -200 -58088 200 -57888
rect -200 -58524 200 -58324
rect -200 -58960 200 -58760
rect -200 -59396 200 -59196
rect -200 -59832 200 -59632
rect -200 -60268 200 -60068
rect -200 -60704 200 -60504
rect -200 -61140 200 -60940
rect -200 -61576 200 -61376
rect -200 -62012 200 -61812
rect -200 -62448 200 -62248
rect -200 -62884 200 -62684
rect -200 -63320 200 -63120
rect -200 -63756 200 -63556
rect -200 -64192 200 -63992
rect -200 -64628 200 -64428
rect -200 -65064 200 -64864
rect -200 -65500 200 -65300
rect -200 -65936 200 -65736
rect -200 -66372 200 -66172
rect -200 -66808 200 -66608
rect -200 -67244 200 -67044
rect -200 -67680 200 -67480
rect -200 -68116 200 -67916
rect -200 -68552 200 -68352
rect -200 -68988 200 -68788
rect -200 -69424 200 -69224
rect -200 -69860 200 -69660
rect -200 -70296 200 -70096
rect -200 -70732 200 -70532
rect -200 -71168 200 -70968
rect -200 -71604 200 -71404
rect -200 -72040 200 -71840
rect -200 -72476 200 -72276
rect -200 -72912 200 -72712
rect -200 -73348 200 -73148
rect -200 -73784 200 -73584
rect -200 -74220 200 -74020
rect -200 -74656 200 -74456
rect -200 -75092 200 -74892
rect -200 -75528 200 -75328
rect -200 -75964 200 -75764
rect -200 -76400 200 -76200
rect -200 -76836 200 -76636
rect -200 -77272 200 -77072
rect -200 -77708 200 -77508
rect -200 -78144 200 -77944
rect -200 -78580 200 -78380
rect -200 -79016 200 -78816
rect -200 -79452 200 -79252
rect -200 -79888 200 -79688
rect -200 -80324 200 -80124
rect -200 -80760 200 -80560
rect -200 -81196 200 -80996
rect -200 -81632 200 -81432
rect -200 -82068 200 -81868
rect -200 -82504 200 -82304
rect -200 -82940 200 -82740
rect -200 -83376 200 -83176
rect -200 -83812 200 -83612
rect -200 -84248 200 -84048
<< pdiff >>
rect -258 84236 -200 84248
rect -258 84060 -246 84236
rect -212 84060 -200 84236
rect -258 84048 -200 84060
rect 200 84236 258 84248
rect 200 84060 212 84236
rect 246 84060 258 84236
rect 200 84048 258 84060
rect -258 83800 -200 83812
rect -258 83624 -246 83800
rect -212 83624 -200 83800
rect -258 83612 -200 83624
rect 200 83800 258 83812
rect 200 83624 212 83800
rect 246 83624 258 83800
rect 200 83612 258 83624
rect -258 83364 -200 83376
rect -258 83188 -246 83364
rect -212 83188 -200 83364
rect -258 83176 -200 83188
rect 200 83364 258 83376
rect 200 83188 212 83364
rect 246 83188 258 83364
rect 200 83176 258 83188
rect -258 82928 -200 82940
rect -258 82752 -246 82928
rect -212 82752 -200 82928
rect -258 82740 -200 82752
rect 200 82928 258 82940
rect 200 82752 212 82928
rect 246 82752 258 82928
rect 200 82740 258 82752
rect -258 82492 -200 82504
rect -258 82316 -246 82492
rect -212 82316 -200 82492
rect -258 82304 -200 82316
rect 200 82492 258 82504
rect 200 82316 212 82492
rect 246 82316 258 82492
rect 200 82304 258 82316
rect -258 82056 -200 82068
rect -258 81880 -246 82056
rect -212 81880 -200 82056
rect -258 81868 -200 81880
rect 200 82056 258 82068
rect 200 81880 212 82056
rect 246 81880 258 82056
rect 200 81868 258 81880
rect -258 81620 -200 81632
rect -258 81444 -246 81620
rect -212 81444 -200 81620
rect -258 81432 -200 81444
rect 200 81620 258 81632
rect 200 81444 212 81620
rect 246 81444 258 81620
rect 200 81432 258 81444
rect -258 81184 -200 81196
rect -258 81008 -246 81184
rect -212 81008 -200 81184
rect -258 80996 -200 81008
rect 200 81184 258 81196
rect 200 81008 212 81184
rect 246 81008 258 81184
rect 200 80996 258 81008
rect -258 80748 -200 80760
rect -258 80572 -246 80748
rect -212 80572 -200 80748
rect -258 80560 -200 80572
rect 200 80748 258 80760
rect 200 80572 212 80748
rect 246 80572 258 80748
rect 200 80560 258 80572
rect -258 80312 -200 80324
rect -258 80136 -246 80312
rect -212 80136 -200 80312
rect -258 80124 -200 80136
rect 200 80312 258 80324
rect 200 80136 212 80312
rect 246 80136 258 80312
rect 200 80124 258 80136
rect -258 79876 -200 79888
rect -258 79700 -246 79876
rect -212 79700 -200 79876
rect -258 79688 -200 79700
rect 200 79876 258 79888
rect 200 79700 212 79876
rect 246 79700 258 79876
rect 200 79688 258 79700
rect -258 79440 -200 79452
rect -258 79264 -246 79440
rect -212 79264 -200 79440
rect -258 79252 -200 79264
rect 200 79440 258 79452
rect 200 79264 212 79440
rect 246 79264 258 79440
rect 200 79252 258 79264
rect -258 79004 -200 79016
rect -258 78828 -246 79004
rect -212 78828 -200 79004
rect -258 78816 -200 78828
rect 200 79004 258 79016
rect 200 78828 212 79004
rect 246 78828 258 79004
rect 200 78816 258 78828
rect -258 78568 -200 78580
rect -258 78392 -246 78568
rect -212 78392 -200 78568
rect -258 78380 -200 78392
rect 200 78568 258 78580
rect 200 78392 212 78568
rect 246 78392 258 78568
rect 200 78380 258 78392
rect -258 78132 -200 78144
rect -258 77956 -246 78132
rect -212 77956 -200 78132
rect -258 77944 -200 77956
rect 200 78132 258 78144
rect 200 77956 212 78132
rect 246 77956 258 78132
rect 200 77944 258 77956
rect -258 77696 -200 77708
rect -258 77520 -246 77696
rect -212 77520 -200 77696
rect -258 77508 -200 77520
rect 200 77696 258 77708
rect 200 77520 212 77696
rect 246 77520 258 77696
rect 200 77508 258 77520
rect -258 77260 -200 77272
rect -258 77084 -246 77260
rect -212 77084 -200 77260
rect -258 77072 -200 77084
rect 200 77260 258 77272
rect 200 77084 212 77260
rect 246 77084 258 77260
rect 200 77072 258 77084
rect -258 76824 -200 76836
rect -258 76648 -246 76824
rect -212 76648 -200 76824
rect -258 76636 -200 76648
rect 200 76824 258 76836
rect 200 76648 212 76824
rect 246 76648 258 76824
rect 200 76636 258 76648
rect -258 76388 -200 76400
rect -258 76212 -246 76388
rect -212 76212 -200 76388
rect -258 76200 -200 76212
rect 200 76388 258 76400
rect 200 76212 212 76388
rect 246 76212 258 76388
rect 200 76200 258 76212
rect -258 75952 -200 75964
rect -258 75776 -246 75952
rect -212 75776 -200 75952
rect -258 75764 -200 75776
rect 200 75952 258 75964
rect 200 75776 212 75952
rect 246 75776 258 75952
rect 200 75764 258 75776
rect -258 75516 -200 75528
rect -258 75340 -246 75516
rect -212 75340 -200 75516
rect -258 75328 -200 75340
rect 200 75516 258 75528
rect 200 75340 212 75516
rect 246 75340 258 75516
rect 200 75328 258 75340
rect -258 75080 -200 75092
rect -258 74904 -246 75080
rect -212 74904 -200 75080
rect -258 74892 -200 74904
rect 200 75080 258 75092
rect 200 74904 212 75080
rect 246 74904 258 75080
rect 200 74892 258 74904
rect -258 74644 -200 74656
rect -258 74468 -246 74644
rect -212 74468 -200 74644
rect -258 74456 -200 74468
rect 200 74644 258 74656
rect 200 74468 212 74644
rect 246 74468 258 74644
rect 200 74456 258 74468
rect -258 74208 -200 74220
rect -258 74032 -246 74208
rect -212 74032 -200 74208
rect -258 74020 -200 74032
rect 200 74208 258 74220
rect 200 74032 212 74208
rect 246 74032 258 74208
rect 200 74020 258 74032
rect -258 73772 -200 73784
rect -258 73596 -246 73772
rect -212 73596 -200 73772
rect -258 73584 -200 73596
rect 200 73772 258 73784
rect 200 73596 212 73772
rect 246 73596 258 73772
rect 200 73584 258 73596
rect -258 73336 -200 73348
rect -258 73160 -246 73336
rect -212 73160 -200 73336
rect -258 73148 -200 73160
rect 200 73336 258 73348
rect 200 73160 212 73336
rect 246 73160 258 73336
rect 200 73148 258 73160
rect -258 72900 -200 72912
rect -258 72724 -246 72900
rect -212 72724 -200 72900
rect -258 72712 -200 72724
rect 200 72900 258 72912
rect 200 72724 212 72900
rect 246 72724 258 72900
rect 200 72712 258 72724
rect -258 72464 -200 72476
rect -258 72288 -246 72464
rect -212 72288 -200 72464
rect -258 72276 -200 72288
rect 200 72464 258 72476
rect 200 72288 212 72464
rect 246 72288 258 72464
rect 200 72276 258 72288
rect -258 72028 -200 72040
rect -258 71852 -246 72028
rect -212 71852 -200 72028
rect -258 71840 -200 71852
rect 200 72028 258 72040
rect 200 71852 212 72028
rect 246 71852 258 72028
rect 200 71840 258 71852
rect -258 71592 -200 71604
rect -258 71416 -246 71592
rect -212 71416 -200 71592
rect -258 71404 -200 71416
rect 200 71592 258 71604
rect 200 71416 212 71592
rect 246 71416 258 71592
rect 200 71404 258 71416
rect -258 71156 -200 71168
rect -258 70980 -246 71156
rect -212 70980 -200 71156
rect -258 70968 -200 70980
rect 200 71156 258 71168
rect 200 70980 212 71156
rect 246 70980 258 71156
rect 200 70968 258 70980
rect -258 70720 -200 70732
rect -258 70544 -246 70720
rect -212 70544 -200 70720
rect -258 70532 -200 70544
rect 200 70720 258 70732
rect 200 70544 212 70720
rect 246 70544 258 70720
rect 200 70532 258 70544
rect -258 70284 -200 70296
rect -258 70108 -246 70284
rect -212 70108 -200 70284
rect -258 70096 -200 70108
rect 200 70284 258 70296
rect 200 70108 212 70284
rect 246 70108 258 70284
rect 200 70096 258 70108
rect -258 69848 -200 69860
rect -258 69672 -246 69848
rect -212 69672 -200 69848
rect -258 69660 -200 69672
rect 200 69848 258 69860
rect 200 69672 212 69848
rect 246 69672 258 69848
rect 200 69660 258 69672
rect -258 69412 -200 69424
rect -258 69236 -246 69412
rect -212 69236 -200 69412
rect -258 69224 -200 69236
rect 200 69412 258 69424
rect 200 69236 212 69412
rect 246 69236 258 69412
rect 200 69224 258 69236
rect -258 68976 -200 68988
rect -258 68800 -246 68976
rect -212 68800 -200 68976
rect -258 68788 -200 68800
rect 200 68976 258 68988
rect 200 68800 212 68976
rect 246 68800 258 68976
rect 200 68788 258 68800
rect -258 68540 -200 68552
rect -258 68364 -246 68540
rect -212 68364 -200 68540
rect -258 68352 -200 68364
rect 200 68540 258 68552
rect 200 68364 212 68540
rect 246 68364 258 68540
rect 200 68352 258 68364
rect -258 68104 -200 68116
rect -258 67928 -246 68104
rect -212 67928 -200 68104
rect -258 67916 -200 67928
rect 200 68104 258 68116
rect 200 67928 212 68104
rect 246 67928 258 68104
rect 200 67916 258 67928
rect -258 67668 -200 67680
rect -258 67492 -246 67668
rect -212 67492 -200 67668
rect -258 67480 -200 67492
rect 200 67668 258 67680
rect 200 67492 212 67668
rect 246 67492 258 67668
rect 200 67480 258 67492
rect -258 67232 -200 67244
rect -258 67056 -246 67232
rect -212 67056 -200 67232
rect -258 67044 -200 67056
rect 200 67232 258 67244
rect 200 67056 212 67232
rect 246 67056 258 67232
rect 200 67044 258 67056
rect -258 66796 -200 66808
rect -258 66620 -246 66796
rect -212 66620 -200 66796
rect -258 66608 -200 66620
rect 200 66796 258 66808
rect 200 66620 212 66796
rect 246 66620 258 66796
rect 200 66608 258 66620
rect -258 66360 -200 66372
rect -258 66184 -246 66360
rect -212 66184 -200 66360
rect -258 66172 -200 66184
rect 200 66360 258 66372
rect 200 66184 212 66360
rect 246 66184 258 66360
rect 200 66172 258 66184
rect -258 65924 -200 65936
rect -258 65748 -246 65924
rect -212 65748 -200 65924
rect -258 65736 -200 65748
rect 200 65924 258 65936
rect 200 65748 212 65924
rect 246 65748 258 65924
rect 200 65736 258 65748
rect -258 65488 -200 65500
rect -258 65312 -246 65488
rect -212 65312 -200 65488
rect -258 65300 -200 65312
rect 200 65488 258 65500
rect 200 65312 212 65488
rect 246 65312 258 65488
rect 200 65300 258 65312
rect -258 65052 -200 65064
rect -258 64876 -246 65052
rect -212 64876 -200 65052
rect -258 64864 -200 64876
rect 200 65052 258 65064
rect 200 64876 212 65052
rect 246 64876 258 65052
rect 200 64864 258 64876
rect -258 64616 -200 64628
rect -258 64440 -246 64616
rect -212 64440 -200 64616
rect -258 64428 -200 64440
rect 200 64616 258 64628
rect 200 64440 212 64616
rect 246 64440 258 64616
rect 200 64428 258 64440
rect -258 64180 -200 64192
rect -258 64004 -246 64180
rect -212 64004 -200 64180
rect -258 63992 -200 64004
rect 200 64180 258 64192
rect 200 64004 212 64180
rect 246 64004 258 64180
rect 200 63992 258 64004
rect -258 63744 -200 63756
rect -258 63568 -246 63744
rect -212 63568 -200 63744
rect -258 63556 -200 63568
rect 200 63744 258 63756
rect 200 63568 212 63744
rect 246 63568 258 63744
rect 200 63556 258 63568
rect -258 63308 -200 63320
rect -258 63132 -246 63308
rect -212 63132 -200 63308
rect -258 63120 -200 63132
rect 200 63308 258 63320
rect 200 63132 212 63308
rect 246 63132 258 63308
rect 200 63120 258 63132
rect -258 62872 -200 62884
rect -258 62696 -246 62872
rect -212 62696 -200 62872
rect -258 62684 -200 62696
rect 200 62872 258 62884
rect 200 62696 212 62872
rect 246 62696 258 62872
rect 200 62684 258 62696
rect -258 62436 -200 62448
rect -258 62260 -246 62436
rect -212 62260 -200 62436
rect -258 62248 -200 62260
rect 200 62436 258 62448
rect 200 62260 212 62436
rect 246 62260 258 62436
rect 200 62248 258 62260
rect -258 62000 -200 62012
rect -258 61824 -246 62000
rect -212 61824 -200 62000
rect -258 61812 -200 61824
rect 200 62000 258 62012
rect 200 61824 212 62000
rect 246 61824 258 62000
rect 200 61812 258 61824
rect -258 61564 -200 61576
rect -258 61388 -246 61564
rect -212 61388 -200 61564
rect -258 61376 -200 61388
rect 200 61564 258 61576
rect 200 61388 212 61564
rect 246 61388 258 61564
rect 200 61376 258 61388
rect -258 61128 -200 61140
rect -258 60952 -246 61128
rect -212 60952 -200 61128
rect -258 60940 -200 60952
rect 200 61128 258 61140
rect 200 60952 212 61128
rect 246 60952 258 61128
rect 200 60940 258 60952
rect -258 60692 -200 60704
rect -258 60516 -246 60692
rect -212 60516 -200 60692
rect -258 60504 -200 60516
rect 200 60692 258 60704
rect 200 60516 212 60692
rect 246 60516 258 60692
rect 200 60504 258 60516
rect -258 60256 -200 60268
rect -258 60080 -246 60256
rect -212 60080 -200 60256
rect -258 60068 -200 60080
rect 200 60256 258 60268
rect 200 60080 212 60256
rect 246 60080 258 60256
rect 200 60068 258 60080
rect -258 59820 -200 59832
rect -258 59644 -246 59820
rect -212 59644 -200 59820
rect -258 59632 -200 59644
rect 200 59820 258 59832
rect 200 59644 212 59820
rect 246 59644 258 59820
rect 200 59632 258 59644
rect -258 59384 -200 59396
rect -258 59208 -246 59384
rect -212 59208 -200 59384
rect -258 59196 -200 59208
rect 200 59384 258 59396
rect 200 59208 212 59384
rect 246 59208 258 59384
rect 200 59196 258 59208
rect -258 58948 -200 58960
rect -258 58772 -246 58948
rect -212 58772 -200 58948
rect -258 58760 -200 58772
rect 200 58948 258 58960
rect 200 58772 212 58948
rect 246 58772 258 58948
rect 200 58760 258 58772
rect -258 58512 -200 58524
rect -258 58336 -246 58512
rect -212 58336 -200 58512
rect -258 58324 -200 58336
rect 200 58512 258 58524
rect 200 58336 212 58512
rect 246 58336 258 58512
rect 200 58324 258 58336
rect -258 58076 -200 58088
rect -258 57900 -246 58076
rect -212 57900 -200 58076
rect -258 57888 -200 57900
rect 200 58076 258 58088
rect 200 57900 212 58076
rect 246 57900 258 58076
rect 200 57888 258 57900
rect -258 57640 -200 57652
rect -258 57464 -246 57640
rect -212 57464 -200 57640
rect -258 57452 -200 57464
rect 200 57640 258 57652
rect 200 57464 212 57640
rect 246 57464 258 57640
rect 200 57452 258 57464
rect -258 57204 -200 57216
rect -258 57028 -246 57204
rect -212 57028 -200 57204
rect -258 57016 -200 57028
rect 200 57204 258 57216
rect 200 57028 212 57204
rect 246 57028 258 57204
rect 200 57016 258 57028
rect -258 56768 -200 56780
rect -258 56592 -246 56768
rect -212 56592 -200 56768
rect -258 56580 -200 56592
rect 200 56768 258 56780
rect 200 56592 212 56768
rect 246 56592 258 56768
rect 200 56580 258 56592
rect -258 56332 -200 56344
rect -258 56156 -246 56332
rect -212 56156 -200 56332
rect -258 56144 -200 56156
rect 200 56332 258 56344
rect 200 56156 212 56332
rect 246 56156 258 56332
rect 200 56144 258 56156
rect -258 55896 -200 55908
rect -258 55720 -246 55896
rect -212 55720 -200 55896
rect -258 55708 -200 55720
rect 200 55896 258 55908
rect 200 55720 212 55896
rect 246 55720 258 55896
rect 200 55708 258 55720
rect -258 55460 -200 55472
rect -258 55284 -246 55460
rect -212 55284 -200 55460
rect -258 55272 -200 55284
rect 200 55460 258 55472
rect 200 55284 212 55460
rect 246 55284 258 55460
rect 200 55272 258 55284
rect -258 55024 -200 55036
rect -258 54848 -246 55024
rect -212 54848 -200 55024
rect -258 54836 -200 54848
rect 200 55024 258 55036
rect 200 54848 212 55024
rect 246 54848 258 55024
rect 200 54836 258 54848
rect -258 54588 -200 54600
rect -258 54412 -246 54588
rect -212 54412 -200 54588
rect -258 54400 -200 54412
rect 200 54588 258 54600
rect 200 54412 212 54588
rect 246 54412 258 54588
rect 200 54400 258 54412
rect -258 54152 -200 54164
rect -258 53976 -246 54152
rect -212 53976 -200 54152
rect -258 53964 -200 53976
rect 200 54152 258 54164
rect 200 53976 212 54152
rect 246 53976 258 54152
rect 200 53964 258 53976
rect -258 53716 -200 53728
rect -258 53540 -246 53716
rect -212 53540 -200 53716
rect -258 53528 -200 53540
rect 200 53716 258 53728
rect 200 53540 212 53716
rect 246 53540 258 53716
rect 200 53528 258 53540
rect -258 53280 -200 53292
rect -258 53104 -246 53280
rect -212 53104 -200 53280
rect -258 53092 -200 53104
rect 200 53280 258 53292
rect 200 53104 212 53280
rect 246 53104 258 53280
rect 200 53092 258 53104
rect -258 52844 -200 52856
rect -258 52668 -246 52844
rect -212 52668 -200 52844
rect -258 52656 -200 52668
rect 200 52844 258 52856
rect 200 52668 212 52844
rect 246 52668 258 52844
rect 200 52656 258 52668
rect -258 52408 -200 52420
rect -258 52232 -246 52408
rect -212 52232 -200 52408
rect -258 52220 -200 52232
rect 200 52408 258 52420
rect 200 52232 212 52408
rect 246 52232 258 52408
rect 200 52220 258 52232
rect -258 51972 -200 51984
rect -258 51796 -246 51972
rect -212 51796 -200 51972
rect -258 51784 -200 51796
rect 200 51972 258 51984
rect 200 51796 212 51972
rect 246 51796 258 51972
rect 200 51784 258 51796
rect -258 51536 -200 51548
rect -258 51360 -246 51536
rect -212 51360 -200 51536
rect -258 51348 -200 51360
rect 200 51536 258 51548
rect 200 51360 212 51536
rect 246 51360 258 51536
rect 200 51348 258 51360
rect -258 51100 -200 51112
rect -258 50924 -246 51100
rect -212 50924 -200 51100
rect -258 50912 -200 50924
rect 200 51100 258 51112
rect 200 50924 212 51100
rect 246 50924 258 51100
rect 200 50912 258 50924
rect -258 50664 -200 50676
rect -258 50488 -246 50664
rect -212 50488 -200 50664
rect -258 50476 -200 50488
rect 200 50664 258 50676
rect 200 50488 212 50664
rect 246 50488 258 50664
rect 200 50476 258 50488
rect -258 50228 -200 50240
rect -258 50052 -246 50228
rect -212 50052 -200 50228
rect -258 50040 -200 50052
rect 200 50228 258 50240
rect 200 50052 212 50228
rect 246 50052 258 50228
rect 200 50040 258 50052
rect -258 49792 -200 49804
rect -258 49616 -246 49792
rect -212 49616 -200 49792
rect -258 49604 -200 49616
rect 200 49792 258 49804
rect 200 49616 212 49792
rect 246 49616 258 49792
rect 200 49604 258 49616
rect -258 49356 -200 49368
rect -258 49180 -246 49356
rect -212 49180 -200 49356
rect -258 49168 -200 49180
rect 200 49356 258 49368
rect 200 49180 212 49356
rect 246 49180 258 49356
rect 200 49168 258 49180
rect -258 48920 -200 48932
rect -258 48744 -246 48920
rect -212 48744 -200 48920
rect -258 48732 -200 48744
rect 200 48920 258 48932
rect 200 48744 212 48920
rect 246 48744 258 48920
rect 200 48732 258 48744
rect -258 48484 -200 48496
rect -258 48308 -246 48484
rect -212 48308 -200 48484
rect -258 48296 -200 48308
rect 200 48484 258 48496
rect 200 48308 212 48484
rect 246 48308 258 48484
rect 200 48296 258 48308
rect -258 48048 -200 48060
rect -258 47872 -246 48048
rect -212 47872 -200 48048
rect -258 47860 -200 47872
rect 200 48048 258 48060
rect 200 47872 212 48048
rect 246 47872 258 48048
rect 200 47860 258 47872
rect -258 47612 -200 47624
rect -258 47436 -246 47612
rect -212 47436 -200 47612
rect -258 47424 -200 47436
rect 200 47612 258 47624
rect 200 47436 212 47612
rect 246 47436 258 47612
rect 200 47424 258 47436
rect -258 47176 -200 47188
rect -258 47000 -246 47176
rect -212 47000 -200 47176
rect -258 46988 -200 47000
rect 200 47176 258 47188
rect 200 47000 212 47176
rect 246 47000 258 47176
rect 200 46988 258 47000
rect -258 46740 -200 46752
rect -258 46564 -246 46740
rect -212 46564 -200 46740
rect -258 46552 -200 46564
rect 200 46740 258 46752
rect 200 46564 212 46740
rect 246 46564 258 46740
rect 200 46552 258 46564
rect -258 46304 -200 46316
rect -258 46128 -246 46304
rect -212 46128 -200 46304
rect -258 46116 -200 46128
rect 200 46304 258 46316
rect 200 46128 212 46304
rect 246 46128 258 46304
rect 200 46116 258 46128
rect -258 45868 -200 45880
rect -258 45692 -246 45868
rect -212 45692 -200 45868
rect -258 45680 -200 45692
rect 200 45868 258 45880
rect 200 45692 212 45868
rect 246 45692 258 45868
rect 200 45680 258 45692
rect -258 45432 -200 45444
rect -258 45256 -246 45432
rect -212 45256 -200 45432
rect -258 45244 -200 45256
rect 200 45432 258 45444
rect 200 45256 212 45432
rect 246 45256 258 45432
rect 200 45244 258 45256
rect -258 44996 -200 45008
rect -258 44820 -246 44996
rect -212 44820 -200 44996
rect -258 44808 -200 44820
rect 200 44996 258 45008
rect 200 44820 212 44996
rect 246 44820 258 44996
rect 200 44808 258 44820
rect -258 44560 -200 44572
rect -258 44384 -246 44560
rect -212 44384 -200 44560
rect -258 44372 -200 44384
rect 200 44560 258 44572
rect 200 44384 212 44560
rect 246 44384 258 44560
rect 200 44372 258 44384
rect -258 44124 -200 44136
rect -258 43948 -246 44124
rect -212 43948 -200 44124
rect -258 43936 -200 43948
rect 200 44124 258 44136
rect 200 43948 212 44124
rect 246 43948 258 44124
rect 200 43936 258 43948
rect -258 43688 -200 43700
rect -258 43512 -246 43688
rect -212 43512 -200 43688
rect -258 43500 -200 43512
rect 200 43688 258 43700
rect 200 43512 212 43688
rect 246 43512 258 43688
rect 200 43500 258 43512
rect -258 43252 -200 43264
rect -258 43076 -246 43252
rect -212 43076 -200 43252
rect -258 43064 -200 43076
rect 200 43252 258 43264
rect 200 43076 212 43252
rect 246 43076 258 43252
rect 200 43064 258 43076
rect -258 42816 -200 42828
rect -258 42640 -246 42816
rect -212 42640 -200 42816
rect -258 42628 -200 42640
rect 200 42816 258 42828
rect 200 42640 212 42816
rect 246 42640 258 42816
rect 200 42628 258 42640
rect -258 42380 -200 42392
rect -258 42204 -246 42380
rect -212 42204 -200 42380
rect -258 42192 -200 42204
rect 200 42380 258 42392
rect 200 42204 212 42380
rect 246 42204 258 42380
rect 200 42192 258 42204
rect -258 41944 -200 41956
rect -258 41768 -246 41944
rect -212 41768 -200 41944
rect -258 41756 -200 41768
rect 200 41944 258 41956
rect 200 41768 212 41944
rect 246 41768 258 41944
rect 200 41756 258 41768
rect -258 41508 -200 41520
rect -258 41332 -246 41508
rect -212 41332 -200 41508
rect -258 41320 -200 41332
rect 200 41508 258 41520
rect 200 41332 212 41508
rect 246 41332 258 41508
rect 200 41320 258 41332
rect -258 41072 -200 41084
rect -258 40896 -246 41072
rect -212 40896 -200 41072
rect -258 40884 -200 40896
rect 200 41072 258 41084
rect 200 40896 212 41072
rect 246 40896 258 41072
rect 200 40884 258 40896
rect -258 40636 -200 40648
rect -258 40460 -246 40636
rect -212 40460 -200 40636
rect -258 40448 -200 40460
rect 200 40636 258 40648
rect 200 40460 212 40636
rect 246 40460 258 40636
rect 200 40448 258 40460
rect -258 40200 -200 40212
rect -258 40024 -246 40200
rect -212 40024 -200 40200
rect -258 40012 -200 40024
rect 200 40200 258 40212
rect 200 40024 212 40200
rect 246 40024 258 40200
rect 200 40012 258 40024
rect -258 39764 -200 39776
rect -258 39588 -246 39764
rect -212 39588 -200 39764
rect -258 39576 -200 39588
rect 200 39764 258 39776
rect 200 39588 212 39764
rect 246 39588 258 39764
rect 200 39576 258 39588
rect -258 39328 -200 39340
rect -258 39152 -246 39328
rect -212 39152 -200 39328
rect -258 39140 -200 39152
rect 200 39328 258 39340
rect 200 39152 212 39328
rect 246 39152 258 39328
rect 200 39140 258 39152
rect -258 38892 -200 38904
rect -258 38716 -246 38892
rect -212 38716 -200 38892
rect -258 38704 -200 38716
rect 200 38892 258 38904
rect 200 38716 212 38892
rect 246 38716 258 38892
rect 200 38704 258 38716
rect -258 38456 -200 38468
rect -258 38280 -246 38456
rect -212 38280 -200 38456
rect -258 38268 -200 38280
rect 200 38456 258 38468
rect 200 38280 212 38456
rect 246 38280 258 38456
rect 200 38268 258 38280
rect -258 38020 -200 38032
rect -258 37844 -246 38020
rect -212 37844 -200 38020
rect -258 37832 -200 37844
rect 200 38020 258 38032
rect 200 37844 212 38020
rect 246 37844 258 38020
rect 200 37832 258 37844
rect -258 37584 -200 37596
rect -258 37408 -246 37584
rect -212 37408 -200 37584
rect -258 37396 -200 37408
rect 200 37584 258 37596
rect 200 37408 212 37584
rect 246 37408 258 37584
rect 200 37396 258 37408
rect -258 37148 -200 37160
rect -258 36972 -246 37148
rect -212 36972 -200 37148
rect -258 36960 -200 36972
rect 200 37148 258 37160
rect 200 36972 212 37148
rect 246 36972 258 37148
rect 200 36960 258 36972
rect -258 36712 -200 36724
rect -258 36536 -246 36712
rect -212 36536 -200 36712
rect -258 36524 -200 36536
rect 200 36712 258 36724
rect 200 36536 212 36712
rect 246 36536 258 36712
rect 200 36524 258 36536
rect -258 36276 -200 36288
rect -258 36100 -246 36276
rect -212 36100 -200 36276
rect -258 36088 -200 36100
rect 200 36276 258 36288
rect 200 36100 212 36276
rect 246 36100 258 36276
rect 200 36088 258 36100
rect -258 35840 -200 35852
rect -258 35664 -246 35840
rect -212 35664 -200 35840
rect -258 35652 -200 35664
rect 200 35840 258 35852
rect 200 35664 212 35840
rect 246 35664 258 35840
rect 200 35652 258 35664
rect -258 35404 -200 35416
rect -258 35228 -246 35404
rect -212 35228 -200 35404
rect -258 35216 -200 35228
rect 200 35404 258 35416
rect 200 35228 212 35404
rect 246 35228 258 35404
rect 200 35216 258 35228
rect -258 34968 -200 34980
rect -258 34792 -246 34968
rect -212 34792 -200 34968
rect -258 34780 -200 34792
rect 200 34968 258 34980
rect 200 34792 212 34968
rect 246 34792 258 34968
rect 200 34780 258 34792
rect -258 34532 -200 34544
rect -258 34356 -246 34532
rect -212 34356 -200 34532
rect -258 34344 -200 34356
rect 200 34532 258 34544
rect 200 34356 212 34532
rect 246 34356 258 34532
rect 200 34344 258 34356
rect -258 34096 -200 34108
rect -258 33920 -246 34096
rect -212 33920 -200 34096
rect -258 33908 -200 33920
rect 200 34096 258 34108
rect 200 33920 212 34096
rect 246 33920 258 34096
rect 200 33908 258 33920
rect -258 33660 -200 33672
rect -258 33484 -246 33660
rect -212 33484 -200 33660
rect -258 33472 -200 33484
rect 200 33660 258 33672
rect 200 33484 212 33660
rect 246 33484 258 33660
rect 200 33472 258 33484
rect -258 33224 -200 33236
rect -258 33048 -246 33224
rect -212 33048 -200 33224
rect -258 33036 -200 33048
rect 200 33224 258 33236
rect 200 33048 212 33224
rect 246 33048 258 33224
rect 200 33036 258 33048
rect -258 32788 -200 32800
rect -258 32612 -246 32788
rect -212 32612 -200 32788
rect -258 32600 -200 32612
rect 200 32788 258 32800
rect 200 32612 212 32788
rect 246 32612 258 32788
rect 200 32600 258 32612
rect -258 32352 -200 32364
rect -258 32176 -246 32352
rect -212 32176 -200 32352
rect -258 32164 -200 32176
rect 200 32352 258 32364
rect 200 32176 212 32352
rect 246 32176 258 32352
rect 200 32164 258 32176
rect -258 31916 -200 31928
rect -258 31740 -246 31916
rect -212 31740 -200 31916
rect -258 31728 -200 31740
rect 200 31916 258 31928
rect 200 31740 212 31916
rect 246 31740 258 31916
rect 200 31728 258 31740
rect -258 31480 -200 31492
rect -258 31304 -246 31480
rect -212 31304 -200 31480
rect -258 31292 -200 31304
rect 200 31480 258 31492
rect 200 31304 212 31480
rect 246 31304 258 31480
rect 200 31292 258 31304
rect -258 31044 -200 31056
rect -258 30868 -246 31044
rect -212 30868 -200 31044
rect -258 30856 -200 30868
rect 200 31044 258 31056
rect 200 30868 212 31044
rect 246 30868 258 31044
rect 200 30856 258 30868
rect -258 30608 -200 30620
rect -258 30432 -246 30608
rect -212 30432 -200 30608
rect -258 30420 -200 30432
rect 200 30608 258 30620
rect 200 30432 212 30608
rect 246 30432 258 30608
rect 200 30420 258 30432
rect -258 30172 -200 30184
rect -258 29996 -246 30172
rect -212 29996 -200 30172
rect -258 29984 -200 29996
rect 200 30172 258 30184
rect 200 29996 212 30172
rect 246 29996 258 30172
rect 200 29984 258 29996
rect -258 29736 -200 29748
rect -258 29560 -246 29736
rect -212 29560 -200 29736
rect -258 29548 -200 29560
rect 200 29736 258 29748
rect 200 29560 212 29736
rect 246 29560 258 29736
rect 200 29548 258 29560
rect -258 29300 -200 29312
rect -258 29124 -246 29300
rect -212 29124 -200 29300
rect -258 29112 -200 29124
rect 200 29300 258 29312
rect 200 29124 212 29300
rect 246 29124 258 29300
rect 200 29112 258 29124
rect -258 28864 -200 28876
rect -258 28688 -246 28864
rect -212 28688 -200 28864
rect -258 28676 -200 28688
rect 200 28864 258 28876
rect 200 28688 212 28864
rect 246 28688 258 28864
rect 200 28676 258 28688
rect -258 28428 -200 28440
rect -258 28252 -246 28428
rect -212 28252 -200 28428
rect -258 28240 -200 28252
rect 200 28428 258 28440
rect 200 28252 212 28428
rect 246 28252 258 28428
rect 200 28240 258 28252
rect -258 27992 -200 28004
rect -258 27816 -246 27992
rect -212 27816 -200 27992
rect -258 27804 -200 27816
rect 200 27992 258 28004
rect 200 27816 212 27992
rect 246 27816 258 27992
rect 200 27804 258 27816
rect -258 27556 -200 27568
rect -258 27380 -246 27556
rect -212 27380 -200 27556
rect -258 27368 -200 27380
rect 200 27556 258 27568
rect 200 27380 212 27556
rect 246 27380 258 27556
rect 200 27368 258 27380
rect -258 27120 -200 27132
rect -258 26944 -246 27120
rect -212 26944 -200 27120
rect -258 26932 -200 26944
rect 200 27120 258 27132
rect 200 26944 212 27120
rect 246 26944 258 27120
rect 200 26932 258 26944
rect -258 26684 -200 26696
rect -258 26508 -246 26684
rect -212 26508 -200 26684
rect -258 26496 -200 26508
rect 200 26684 258 26696
rect 200 26508 212 26684
rect 246 26508 258 26684
rect 200 26496 258 26508
rect -258 26248 -200 26260
rect -258 26072 -246 26248
rect -212 26072 -200 26248
rect -258 26060 -200 26072
rect 200 26248 258 26260
rect 200 26072 212 26248
rect 246 26072 258 26248
rect 200 26060 258 26072
rect -258 25812 -200 25824
rect -258 25636 -246 25812
rect -212 25636 -200 25812
rect -258 25624 -200 25636
rect 200 25812 258 25824
rect 200 25636 212 25812
rect 246 25636 258 25812
rect 200 25624 258 25636
rect -258 25376 -200 25388
rect -258 25200 -246 25376
rect -212 25200 -200 25376
rect -258 25188 -200 25200
rect 200 25376 258 25388
rect 200 25200 212 25376
rect 246 25200 258 25376
rect 200 25188 258 25200
rect -258 24940 -200 24952
rect -258 24764 -246 24940
rect -212 24764 -200 24940
rect -258 24752 -200 24764
rect 200 24940 258 24952
rect 200 24764 212 24940
rect 246 24764 258 24940
rect 200 24752 258 24764
rect -258 24504 -200 24516
rect -258 24328 -246 24504
rect -212 24328 -200 24504
rect -258 24316 -200 24328
rect 200 24504 258 24516
rect 200 24328 212 24504
rect 246 24328 258 24504
rect 200 24316 258 24328
rect -258 24068 -200 24080
rect -258 23892 -246 24068
rect -212 23892 -200 24068
rect -258 23880 -200 23892
rect 200 24068 258 24080
rect 200 23892 212 24068
rect 246 23892 258 24068
rect 200 23880 258 23892
rect -258 23632 -200 23644
rect -258 23456 -246 23632
rect -212 23456 -200 23632
rect -258 23444 -200 23456
rect 200 23632 258 23644
rect 200 23456 212 23632
rect 246 23456 258 23632
rect 200 23444 258 23456
rect -258 23196 -200 23208
rect -258 23020 -246 23196
rect -212 23020 -200 23196
rect -258 23008 -200 23020
rect 200 23196 258 23208
rect 200 23020 212 23196
rect 246 23020 258 23196
rect 200 23008 258 23020
rect -258 22760 -200 22772
rect -258 22584 -246 22760
rect -212 22584 -200 22760
rect -258 22572 -200 22584
rect 200 22760 258 22772
rect 200 22584 212 22760
rect 246 22584 258 22760
rect 200 22572 258 22584
rect -258 22324 -200 22336
rect -258 22148 -246 22324
rect -212 22148 -200 22324
rect -258 22136 -200 22148
rect 200 22324 258 22336
rect 200 22148 212 22324
rect 246 22148 258 22324
rect 200 22136 258 22148
rect -258 21888 -200 21900
rect -258 21712 -246 21888
rect -212 21712 -200 21888
rect -258 21700 -200 21712
rect 200 21888 258 21900
rect 200 21712 212 21888
rect 246 21712 258 21888
rect 200 21700 258 21712
rect -258 21452 -200 21464
rect -258 21276 -246 21452
rect -212 21276 -200 21452
rect -258 21264 -200 21276
rect 200 21452 258 21464
rect 200 21276 212 21452
rect 246 21276 258 21452
rect 200 21264 258 21276
rect -258 21016 -200 21028
rect -258 20840 -246 21016
rect -212 20840 -200 21016
rect -258 20828 -200 20840
rect 200 21016 258 21028
rect 200 20840 212 21016
rect 246 20840 258 21016
rect 200 20828 258 20840
rect -258 20580 -200 20592
rect -258 20404 -246 20580
rect -212 20404 -200 20580
rect -258 20392 -200 20404
rect 200 20580 258 20592
rect 200 20404 212 20580
rect 246 20404 258 20580
rect 200 20392 258 20404
rect -258 20144 -200 20156
rect -258 19968 -246 20144
rect -212 19968 -200 20144
rect -258 19956 -200 19968
rect 200 20144 258 20156
rect 200 19968 212 20144
rect 246 19968 258 20144
rect 200 19956 258 19968
rect -258 19708 -200 19720
rect -258 19532 -246 19708
rect -212 19532 -200 19708
rect -258 19520 -200 19532
rect 200 19708 258 19720
rect 200 19532 212 19708
rect 246 19532 258 19708
rect 200 19520 258 19532
rect -258 19272 -200 19284
rect -258 19096 -246 19272
rect -212 19096 -200 19272
rect -258 19084 -200 19096
rect 200 19272 258 19284
rect 200 19096 212 19272
rect 246 19096 258 19272
rect 200 19084 258 19096
rect -258 18836 -200 18848
rect -258 18660 -246 18836
rect -212 18660 -200 18836
rect -258 18648 -200 18660
rect 200 18836 258 18848
rect 200 18660 212 18836
rect 246 18660 258 18836
rect 200 18648 258 18660
rect -258 18400 -200 18412
rect -258 18224 -246 18400
rect -212 18224 -200 18400
rect -258 18212 -200 18224
rect 200 18400 258 18412
rect 200 18224 212 18400
rect 246 18224 258 18400
rect 200 18212 258 18224
rect -258 17964 -200 17976
rect -258 17788 -246 17964
rect -212 17788 -200 17964
rect -258 17776 -200 17788
rect 200 17964 258 17976
rect 200 17788 212 17964
rect 246 17788 258 17964
rect 200 17776 258 17788
rect -258 17528 -200 17540
rect -258 17352 -246 17528
rect -212 17352 -200 17528
rect -258 17340 -200 17352
rect 200 17528 258 17540
rect 200 17352 212 17528
rect 246 17352 258 17528
rect 200 17340 258 17352
rect -258 17092 -200 17104
rect -258 16916 -246 17092
rect -212 16916 -200 17092
rect -258 16904 -200 16916
rect 200 17092 258 17104
rect 200 16916 212 17092
rect 246 16916 258 17092
rect 200 16904 258 16916
rect -258 16656 -200 16668
rect -258 16480 -246 16656
rect -212 16480 -200 16656
rect -258 16468 -200 16480
rect 200 16656 258 16668
rect 200 16480 212 16656
rect 246 16480 258 16656
rect 200 16468 258 16480
rect -258 16220 -200 16232
rect -258 16044 -246 16220
rect -212 16044 -200 16220
rect -258 16032 -200 16044
rect 200 16220 258 16232
rect 200 16044 212 16220
rect 246 16044 258 16220
rect 200 16032 258 16044
rect -258 15784 -200 15796
rect -258 15608 -246 15784
rect -212 15608 -200 15784
rect -258 15596 -200 15608
rect 200 15784 258 15796
rect 200 15608 212 15784
rect 246 15608 258 15784
rect 200 15596 258 15608
rect -258 15348 -200 15360
rect -258 15172 -246 15348
rect -212 15172 -200 15348
rect -258 15160 -200 15172
rect 200 15348 258 15360
rect 200 15172 212 15348
rect 246 15172 258 15348
rect 200 15160 258 15172
rect -258 14912 -200 14924
rect -258 14736 -246 14912
rect -212 14736 -200 14912
rect -258 14724 -200 14736
rect 200 14912 258 14924
rect 200 14736 212 14912
rect 246 14736 258 14912
rect 200 14724 258 14736
rect -258 14476 -200 14488
rect -258 14300 -246 14476
rect -212 14300 -200 14476
rect -258 14288 -200 14300
rect 200 14476 258 14488
rect 200 14300 212 14476
rect 246 14300 258 14476
rect 200 14288 258 14300
rect -258 14040 -200 14052
rect -258 13864 -246 14040
rect -212 13864 -200 14040
rect -258 13852 -200 13864
rect 200 14040 258 14052
rect 200 13864 212 14040
rect 246 13864 258 14040
rect 200 13852 258 13864
rect -258 13604 -200 13616
rect -258 13428 -246 13604
rect -212 13428 -200 13604
rect -258 13416 -200 13428
rect 200 13604 258 13616
rect 200 13428 212 13604
rect 246 13428 258 13604
rect 200 13416 258 13428
rect -258 13168 -200 13180
rect -258 12992 -246 13168
rect -212 12992 -200 13168
rect -258 12980 -200 12992
rect 200 13168 258 13180
rect 200 12992 212 13168
rect 246 12992 258 13168
rect 200 12980 258 12992
rect -258 12732 -200 12744
rect -258 12556 -246 12732
rect -212 12556 -200 12732
rect -258 12544 -200 12556
rect 200 12732 258 12744
rect 200 12556 212 12732
rect 246 12556 258 12732
rect 200 12544 258 12556
rect -258 12296 -200 12308
rect -258 12120 -246 12296
rect -212 12120 -200 12296
rect -258 12108 -200 12120
rect 200 12296 258 12308
rect 200 12120 212 12296
rect 246 12120 258 12296
rect 200 12108 258 12120
rect -258 11860 -200 11872
rect -258 11684 -246 11860
rect -212 11684 -200 11860
rect -258 11672 -200 11684
rect 200 11860 258 11872
rect 200 11684 212 11860
rect 246 11684 258 11860
rect 200 11672 258 11684
rect -258 11424 -200 11436
rect -258 11248 -246 11424
rect -212 11248 -200 11424
rect -258 11236 -200 11248
rect 200 11424 258 11436
rect 200 11248 212 11424
rect 246 11248 258 11424
rect 200 11236 258 11248
rect -258 10988 -200 11000
rect -258 10812 -246 10988
rect -212 10812 -200 10988
rect -258 10800 -200 10812
rect 200 10988 258 11000
rect 200 10812 212 10988
rect 246 10812 258 10988
rect 200 10800 258 10812
rect -258 10552 -200 10564
rect -258 10376 -246 10552
rect -212 10376 -200 10552
rect -258 10364 -200 10376
rect 200 10552 258 10564
rect 200 10376 212 10552
rect 246 10376 258 10552
rect 200 10364 258 10376
rect -258 10116 -200 10128
rect -258 9940 -246 10116
rect -212 9940 -200 10116
rect -258 9928 -200 9940
rect 200 10116 258 10128
rect 200 9940 212 10116
rect 246 9940 258 10116
rect 200 9928 258 9940
rect -258 9680 -200 9692
rect -258 9504 -246 9680
rect -212 9504 -200 9680
rect -258 9492 -200 9504
rect 200 9680 258 9692
rect 200 9504 212 9680
rect 246 9504 258 9680
rect 200 9492 258 9504
rect -258 9244 -200 9256
rect -258 9068 -246 9244
rect -212 9068 -200 9244
rect -258 9056 -200 9068
rect 200 9244 258 9256
rect 200 9068 212 9244
rect 246 9068 258 9244
rect 200 9056 258 9068
rect -258 8808 -200 8820
rect -258 8632 -246 8808
rect -212 8632 -200 8808
rect -258 8620 -200 8632
rect 200 8808 258 8820
rect 200 8632 212 8808
rect 246 8632 258 8808
rect 200 8620 258 8632
rect -258 8372 -200 8384
rect -258 8196 -246 8372
rect -212 8196 -200 8372
rect -258 8184 -200 8196
rect 200 8372 258 8384
rect 200 8196 212 8372
rect 246 8196 258 8372
rect 200 8184 258 8196
rect -258 7936 -200 7948
rect -258 7760 -246 7936
rect -212 7760 -200 7936
rect -258 7748 -200 7760
rect 200 7936 258 7948
rect 200 7760 212 7936
rect 246 7760 258 7936
rect 200 7748 258 7760
rect -258 7500 -200 7512
rect -258 7324 -246 7500
rect -212 7324 -200 7500
rect -258 7312 -200 7324
rect 200 7500 258 7512
rect 200 7324 212 7500
rect 246 7324 258 7500
rect 200 7312 258 7324
rect -258 7064 -200 7076
rect -258 6888 -246 7064
rect -212 6888 -200 7064
rect -258 6876 -200 6888
rect 200 7064 258 7076
rect 200 6888 212 7064
rect 246 6888 258 7064
rect 200 6876 258 6888
rect -258 6628 -200 6640
rect -258 6452 -246 6628
rect -212 6452 -200 6628
rect -258 6440 -200 6452
rect 200 6628 258 6640
rect 200 6452 212 6628
rect 246 6452 258 6628
rect 200 6440 258 6452
rect -258 6192 -200 6204
rect -258 6016 -246 6192
rect -212 6016 -200 6192
rect -258 6004 -200 6016
rect 200 6192 258 6204
rect 200 6016 212 6192
rect 246 6016 258 6192
rect 200 6004 258 6016
rect -258 5756 -200 5768
rect -258 5580 -246 5756
rect -212 5580 -200 5756
rect -258 5568 -200 5580
rect 200 5756 258 5768
rect 200 5580 212 5756
rect 246 5580 258 5756
rect 200 5568 258 5580
rect -258 5320 -200 5332
rect -258 5144 -246 5320
rect -212 5144 -200 5320
rect -258 5132 -200 5144
rect 200 5320 258 5332
rect 200 5144 212 5320
rect 246 5144 258 5320
rect 200 5132 258 5144
rect -258 4884 -200 4896
rect -258 4708 -246 4884
rect -212 4708 -200 4884
rect -258 4696 -200 4708
rect 200 4884 258 4896
rect 200 4708 212 4884
rect 246 4708 258 4884
rect 200 4696 258 4708
rect -258 4448 -200 4460
rect -258 4272 -246 4448
rect -212 4272 -200 4448
rect -258 4260 -200 4272
rect 200 4448 258 4460
rect 200 4272 212 4448
rect 246 4272 258 4448
rect 200 4260 258 4272
rect -258 4012 -200 4024
rect -258 3836 -246 4012
rect -212 3836 -200 4012
rect -258 3824 -200 3836
rect 200 4012 258 4024
rect 200 3836 212 4012
rect 246 3836 258 4012
rect 200 3824 258 3836
rect -258 3576 -200 3588
rect -258 3400 -246 3576
rect -212 3400 -200 3576
rect -258 3388 -200 3400
rect 200 3576 258 3588
rect 200 3400 212 3576
rect 246 3400 258 3576
rect 200 3388 258 3400
rect -258 3140 -200 3152
rect -258 2964 -246 3140
rect -212 2964 -200 3140
rect -258 2952 -200 2964
rect 200 3140 258 3152
rect 200 2964 212 3140
rect 246 2964 258 3140
rect 200 2952 258 2964
rect -258 2704 -200 2716
rect -258 2528 -246 2704
rect -212 2528 -200 2704
rect -258 2516 -200 2528
rect 200 2704 258 2716
rect 200 2528 212 2704
rect 246 2528 258 2704
rect 200 2516 258 2528
rect -258 2268 -200 2280
rect -258 2092 -246 2268
rect -212 2092 -200 2268
rect -258 2080 -200 2092
rect 200 2268 258 2280
rect 200 2092 212 2268
rect 246 2092 258 2268
rect 200 2080 258 2092
rect -258 1832 -200 1844
rect -258 1656 -246 1832
rect -212 1656 -200 1832
rect -258 1644 -200 1656
rect 200 1832 258 1844
rect 200 1656 212 1832
rect 246 1656 258 1832
rect 200 1644 258 1656
rect -258 1396 -200 1408
rect -258 1220 -246 1396
rect -212 1220 -200 1396
rect -258 1208 -200 1220
rect 200 1396 258 1408
rect 200 1220 212 1396
rect 246 1220 258 1396
rect 200 1208 258 1220
rect -258 960 -200 972
rect -258 784 -246 960
rect -212 784 -200 960
rect -258 772 -200 784
rect 200 960 258 972
rect 200 784 212 960
rect 246 784 258 960
rect 200 772 258 784
rect -258 524 -200 536
rect -258 348 -246 524
rect -212 348 -200 524
rect -258 336 -200 348
rect 200 524 258 536
rect 200 348 212 524
rect 246 348 258 524
rect 200 336 258 348
rect -258 88 -200 100
rect -258 -88 -246 88
rect -212 -88 -200 88
rect -258 -100 -200 -88
rect 200 88 258 100
rect 200 -88 212 88
rect 246 -88 258 88
rect 200 -100 258 -88
rect -258 -348 -200 -336
rect -258 -524 -246 -348
rect -212 -524 -200 -348
rect -258 -536 -200 -524
rect 200 -348 258 -336
rect 200 -524 212 -348
rect 246 -524 258 -348
rect 200 -536 258 -524
rect -258 -784 -200 -772
rect -258 -960 -246 -784
rect -212 -960 -200 -784
rect -258 -972 -200 -960
rect 200 -784 258 -772
rect 200 -960 212 -784
rect 246 -960 258 -784
rect 200 -972 258 -960
rect -258 -1220 -200 -1208
rect -258 -1396 -246 -1220
rect -212 -1396 -200 -1220
rect -258 -1408 -200 -1396
rect 200 -1220 258 -1208
rect 200 -1396 212 -1220
rect 246 -1396 258 -1220
rect 200 -1408 258 -1396
rect -258 -1656 -200 -1644
rect -258 -1832 -246 -1656
rect -212 -1832 -200 -1656
rect -258 -1844 -200 -1832
rect 200 -1656 258 -1644
rect 200 -1832 212 -1656
rect 246 -1832 258 -1656
rect 200 -1844 258 -1832
rect -258 -2092 -200 -2080
rect -258 -2268 -246 -2092
rect -212 -2268 -200 -2092
rect -258 -2280 -200 -2268
rect 200 -2092 258 -2080
rect 200 -2268 212 -2092
rect 246 -2268 258 -2092
rect 200 -2280 258 -2268
rect -258 -2528 -200 -2516
rect -258 -2704 -246 -2528
rect -212 -2704 -200 -2528
rect -258 -2716 -200 -2704
rect 200 -2528 258 -2516
rect 200 -2704 212 -2528
rect 246 -2704 258 -2528
rect 200 -2716 258 -2704
rect -258 -2964 -200 -2952
rect -258 -3140 -246 -2964
rect -212 -3140 -200 -2964
rect -258 -3152 -200 -3140
rect 200 -2964 258 -2952
rect 200 -3140 212 -2964
rect 246 -3140 258 -2964
rect 200 -3152 258 -3140
rect -258 -3400 -200 -3388
rect -258 -3576 -246 -3400
rect -212 -3576 -200 -3400
rect -258 -3588 -200 -3576
rect 200 -3400 258 -3388
rect 200 -3576 212 -3400
rect 246 -3576 258 -3400
rect 200 -3588 258 -3576
rect -258 -3836 -200 -3824
rect -258 -4012 -246 -3836
rect -212 -4012 -200 -3836
rect -258 -4024 -200 -4012
rect 200 -3836 258 -3824
rect 200 -4012 212 -3836
rect 246 -4012 258 -3836
rect 200 -4024 258 -4012
rect -258 -4272 -200 -4260
rect -258 -4448 -246 -4272
rect -212 -4448 -200 -4272
rect -258 -4460 -200 -4448
rect 200 -4272 258 -4260
rect 200 -4448 212 -4272
rect 246 -4448 258 -4272
rect 200 -4460 258 -4448
rect -258 -4708 -200 -4696
rect -258 -4884 -246 -4708
rect -212 -4884 -200 -4708
rect -258 -4896 -200 -4884
rect 200 -4708 258 -4696
rect 200 -4884 212 -4708
rect 246 -4884 258 -4708
rect 200 -4896 258 -4884
rect -258 -5144 -200 -5132
rect -258 -5320 -246 -5144
rect -212 -5320 -200 -5144
rect -258 -5332 -200 -5320
rect 200 -5144 258 -5132
rect 200 -5320 212 -5144
rect 246 -5320 258 -5144
rect 200 -5332 258 -5320
rect -258 -5580 -200 -5568
rect -258 -5756 -246 -5580
rect -212 -5756 -200 -5580
rect -258 -5768 -200 -5756
rect 200 -5580 258 -5568
rect 200 -5756 212 -5580
rect 246 -5756 258 -5580
rect 200 -5768 258 -5756
rect -258 -6016 -200 -6004
rect -258 -6192 -246 -6016
rect -212 -6192 -200 -6016
rect -258 -6204 -200 -6192
rect 200 -6016 258 -6004
rect 200 -6192 212 -6016
rect 246 -6192 258 -6016
rect 200 -6204 258 -6192
rect -258 -6452 -200 -6440
rect -258 -6628 -246 -6452
rect -212 -6628 -200 -6452
rect -258 -6640 -200 -6628
rect 200 -6452 258 -6440
rect 200 -6628 212 -6452
rect 246 -6628 258 -6452
rect 200 -6640 258 -6628
rect -258 -6888 -200 -6876
rect -258 -7064 -246 -6888
rect -212 -7064 -200 -6888
rect -258 -7076 -200 -7064
rect 200 -6888 258 -6876
rect 200 -7064 212 -6888
rect 246 -7064 258 -6888
rect 200 -7076 258 -7064
rect -258 -7324 -200 -7312
rect -258 -7500 -246 -7324
rect -212 -7500 -200 -7324
rect -258 -7512 -200 -7500
rect 200 -7324 258 -7312
rect 200 -7500 212 -7324
rect 246 -7500 258 -7324
rect 200 -7512 258 -7500
rect -258 -7760 -200 -7748
rect -258 -7936 -246 -7760
rect -212 -7936 -200 -7760
rect -258 -7948 -200 -7936
rect 200 -7760 258 -7748
rect 200 -7936 212 -7760
rect 246 -7936 258 -7760
rect 200 -7948 258 -7936
rect -258 -8196 -200 -8184
rect -258 -8372 -246 -8196
rect -212 -8372 -200 -8196
rect -258 -8384 -200 -8372
rect 200 -8196 258 -8184
rect 200 -8372 212 -8196
rect 246 -8372 258 -8196
rect 200 -8384 258 -8372
rect -258 -8632 -200 -8620
rect -258 -8808 -246 -8632
rect -212 -8808 -200 -8632
rect -258 -8820 -200 -8808
rect 200 -8632 258 -8620
rect 200 -8808 212 -8632
rect 246 -8808 258 -8632
rect 200 -8820 258 -8808
rect -258 -9068 -200 -9056
rect -258 -9244 -246 -9068
rect -212 -9244 -200 -9068
rect -258 -9256 -200 -9244
rect 200 -9068 258 -9056
rect 200 -9244 212 -9068
rect 246 -9244 258 -9068
rect 200 -9256 258 -9244
rect -258 -9504 -200 -9492
rect -258 -9680 -246 -9504
rect -212 -9680 -200 -9504
rect -258 -9692 -200 -9680
rect 200 -9504 258 -9492
rect 200 -9680 212 -9504
rect 246 -9680 258 -9504
rect 200 -9692 258 -9680
rect -258 -9940 -200 -9928
rect -258 -10116 -246 -9940
rect -212 -10116 -200 -9940
rect -258 -10128 -200 -10116
rect 200 -9940 258 -9928
rect 200 -10116 212 -9940
rect 246 -10116 258 -9940
rect 200 -10128 258 -10116
rect -258 -10376 -200 -10364
rect -258 -10552 -246 -10376
rect -212 -10552 -200 -10376
rect -258 -10564 -200 -10552
rect 200 -10376 258 -10364
rect 200 -10552 212 -10376
rect 246 -10552 258 -10376
rect 200 -10564 258 -10552
rect -258 -10812 -200 -10800
rect -258 -10988 -246 -10812
rect -212 -10988 -200 -10812
rect -258 -11000 -200 -10988
rect 200 -10812 258 -10800
rect 200 -10988 212 -10812
rect 246 -10988 258 -10812
rect 200 -11000 258 -10988
rect -258 -11248 -200 -11236
rect -258 -11424 -246 -11248
rect -212 -11424 -200 -11248
rect -258 -11436 -200 -11424
rect 200 -11248 258 -11236
rect 200 -11424 212 -11248
rect 246 -11424 258 -11248
rect 200 -11436 258 -11424
rect -258 -11684 -200 -11672
rect -258 -11860 -246 -11684
rect -212 -11860 -200 -11684
rect -258 -11872 -200 -11860
rect 200 -11684 258 -11672
rect 200 -11860 212 -11684
rect 246 -11860 258 -11684
rect 200 -11872 258 -11860
rect -258 -12120 -200 -12108
rect -258 -12296 -246 -12120
rect -212 -12296 -200 -12120
rect -258 -12308 -200 -12296
rect 200 -12120 258 -12108
rect 200 -12296 212 -12120
rect 246 -12296 258 -12120
rect 200 -12308 258 -12296
rect -258 -12556 -200 -12544
rect -258 -12732 -246 -12556
rect -212 -12732 -200 -12556
rect -258 -12744 -200 -12732
rect 200 -12556 258 -12544
rect 200 -12732 212 -12556
rect 246 -12732 258 -12556
rect 200 -12744 258 -12732
rect -258 -12992 -200 -12980
rect -258 -13168 -246 -12992
rect -212 -13168 -200 -12992
rect -258 -13180 -200 -13168
rect 200 -12992 258 -12980
rect 200 -13168 212 -12992
rect 246 -13168 258 -12992
rect 200 -13180 258 -13168
rect -258 -13428 -200 -13416
rect -258 -13604 -246 -13428
rect -212 -13604 -200 -13428
rect -258 -13616 -200 -13604
rect 200 -13428 258 -13416
rect 200 -13604 212 -13428
rect 246 -13604 258 -13428
rect 200 -13616 258 -13604
rect -258 -13864 -200 -13852
rect -258 -14040 -246 -13864
rect -212 -14040 -200 -13864
rect -258 -14052 -200 -14040
rect 200 -13864 258 -13852
rect 200 -14040 212 -13864
rect 246 -14040 258 -13864
rect 200 -14052 258 -14040
rect -258 -14300 -200 -14288
rect -258 -14476 -246 -14300
rect -212 -14476 -200 -14300
rect -258 -14488 -200 -14476
rect 200 -14300 258 -14288
rect 200 -14476 212 -14300
rect 246 -14476 258 -14300
rect 200 -14488 258 -14476
rect -258 -14736 -200 -14724
rect -258 -14912 -246 -14736
rect -212 -14912 -200 -14736
rect -258 -14924 -200 -14912
rect 200 -14736 258 -14724
rect 200 -14912 212 -14736
rect 246 -14912 258 -14736
rect 200 -14924 258 -14912
rect -258 -15172 -200 -15160
rect -258 -15348 -246 -15172
rect -212 -15348 -200 -15172
rect -258 -15360 -200 -15348
rect 200 -15172 258 -15160
rect 200 -15348 212 -15172
rect 246 -15348 258 -15172
rect 200 -15360 258 -15348
rect -258 -15608 -200 -15596
rect -258 -15784 -246 -15608
rect -212 -15784 -200 -15608
rect -258 -15796 -200 -15784
rect 200 -15608 258 -15596
rect 200 -15784 212 -15608
rect 246 -15784 258 -15608
rect 200 -15796 258 -15784
rect -258 -16044 -200 -16032
rect -258 -16220 -246 -16044
rect -212 -16220 -200 -16044
rect -258 -16232 -200 -16220
rect 200 -16044 258 -16032
rect 200 -16220 212 -16044
rect 246 -16220 258 -16044
rect 200 -16232 258 -16220
rect -258 -16480 -200 -16468
rect -258 -16656 -246 -16480
rect -212 -16656 -200 -16480
rect -258 -16668 -200 -16656
rect 200 -16480 258 -16468
rect 200 -16656 212 -16480
rect 246 -16656 258 -16480
rect 200 -16668 258 -16656
rect -258 -16916 -200 -16904
rect -258 -17092 -246 -16916
rect -212 -17092 -200 -16916
rect -258 -17104 -200 -17092
rect 200 -16916 258 -16904
rect 200 -17092 212 -16916
rect 246 -17092 258 -16916
rect 200 -17104 258 -17092
rect -258 -17352 -200 -17340
rect -258 -17528 -246 -17352
rect -212 -17528 -200 -17352
rect -258 -17540 -200 -17528
rect 200 -17352 258 -17340
rect 200 -17528 212 -17352
rect 246 -17528 258 -17352
rect 200 -17540 258 -17528
rect -258 -17788 -200 -17776
rect -258 -17964 -246 -17788
rect -212 -17964 -200 -17788
rect -258 -17976 -200 -17964
rect 200 -17788 258 -17776
rect 200 -17964 212 -17788
rect 246 -17964 258 -17788
rect 200 -17976 258 -17964
rect -258 -18224 -200 -18212
rect -258 -18400 -246 -18224
rect -212 -18400 -200 -18224
rect -258 -18412 -200 -18400
rect 200 -18224 258 -18212
rect 200 -18400 212 -18224
rect 246 -18400 258 -18224
rect 200 -18412 258 -18400
rect -258 -18660 -200 -18648
rect -258 -18836 -246 -18660
rect -212 -18836 -200 -18660
rect -258 -18848 -200 -18836
rect 200 -18660 258 -18648
rect 200 -18836 212 -18660
rect 246 -18836 258 -18660
rect 200 -18848 258 -18836
rect -258 -19096 -200 -19084
rect -258 -19272 -246 -19096
rect -212 -19272 -200 -19096
rect -258 -19284 -200 -19272
rect 200 -19096 258 -19084
rect 200 -19272 212 -19096
rect 246 -19272 258 -19096
rect 200 -19284 258 -19272
rect -258 -19532 -200 -19520
rect -258 -19708 -246 -19532
rect -212 -19708 -200 -19532
rect -258 -19720 -200 -19708
rect 200 -19532 258 -19520
rect 200 -19708 212 -19532
rect 246 -19708 258 -19532
rect 200 -19720 258 -19708
rect -258 -19968 -200 -19956
rect -258 -20144 -246 -19968
rect -212 -20144 -200 -19968
rect -258 -20156 -200 -20144
rect 200 -19968 258 -19956
rect 200 -20144 212 -19968
rect 246 -20144 258 -19968
rect 200 -20156 258 -20144
rect -258 -20404 -200 -20392
rect -258 -20580 -246 -20404
rect -212 -20580 -200 -20404
rect -258 -20592 -200 -20580
rect 200 -20404 258 -20392
rect 200 -20580 212 -20404
rect 246 -20580 258 -20404
rect 200 -20592 258 -20580
rect -258 -20840 -200 -20828
rect -258 -21016 -246 -20840
rect -212 -21016 -200 -20840
rect -258 -21028 -200 -21016
rect 200 -20840 258 -20828
rect 200 -21016 212 -20840
rect 246 -21016 258 -20840
rect 200 -21028 258 -21016
rect -258 -21276 -200 -21264
rect -258 -21452 -246 -21276
rect -212 -21452 -200 -21276
rect -258 -21464 -200 -21452
rect 200 -21276 258 -21264
rect 200 -21452 212 -21276
rect 246 -21452 258 -21276
rect 200 -21464 258 -21452
rect -258 -21712 -200 -21700
rect -258 -21888 -246 -21712
rect -212 -21888 -200 -21712
rect -258 -21900 -200 -21888
rect 200 -21712 258 -21700
rect 200 -21888 212 -21712
rect 246 -21888 258 -21712
rect 200 -21900 258 -21888
rect -258 -22148 -200 -22136
rect -258 -22324 -246 -22148
rect -212 -22324 -200 -22148
rect -258 -22336 -200 -22324
rect 200 -22148 258 -22136
rect 200 -22324 212 -22148
rect 246 -22324 258 -22148
rect 200 -22336 258 -22324
rect -258 -22584 -200 -22572
rect -258 -22760 -246 -22584
rect -212 -22760 -200 -22584
rect -258 -22772 -200 -22760
rect 200 -22584 258 -22572
rect 200 -22760 212 -22584
rect 246 -22760 258 -22584
rect 200 -22772 258 -22760
rect -258 -23020 -200 -23008
rect -258 -23196 -246 -23020
rect -212 -23196 -200 -23020
rect -258 -23208 -200 -23196
rect 200 -23020 258 -23008
rect 200 -23196 212 -23020
rect 246 -23196 258 -23020
rect 200 -23208 258 -23196
rect -258 -23456 -200 -23444
rect -258 -23632 -246 -23456
rect -212 -23632 -200 -23456
rect -258 -23644 -200 -23632
rect 200 -23456 258 -23444
rect 200 -23632 212 -23456
rect 246 -23632 258 -23456
rect 200 -23644 258 -23632
rect -258 -23892 -200 -23880
rect -258 -24068 -246 -23892
rect -212 -24068 -200 -23892
rect -258 -24080 -200 -24068
rect 200 -23892 258 -23880
rect 200 -24068 212 -23892
rect 246 -24068 258 -23892
rect 200 -24080 258 -24068
rect -258 -24328 -200 -24316
rect -258 -24504 -246 -24328
rect -212 -24504 -200 -24328
rect -258 -24516 -200 -24504
rect 200 -24328 258 -24316
rect 200 -24504 212 -24328
rect 246 -24504 258 -24328
rect 200 -24516 258 -24504
rect -258 -24764 -200 -24752
rect -258 -24940 -246 -24764
rect -212 -24940 -200 -24764
rect -258 -24952 -200 -24940
rect 200 -24764 258 -24752
rect 200 -24940 212 -24764
rect 246 -24940 258 -24764
rect 200 -24952 258 -24940
rect -258 -25200 -200 -25188
rect -258 -25376 -246 -25200
rect -212 -25376 -200 -25200
rect -258 -25388 -200 -25376
rect 200 -25200 258 -25188
rect 200 -25376 212 -25200
rect 246 -25376 258 -25200
rect 200 -25388 258 -25376
rect -258 -25636 -200 -25624
rect -258 -25812 -246 -25636
rect -212 -25812 -200 -25636
rect -258 -25824 -200 -25812
rect 200 -25636 258 -25624
rect 200 -25812 212 -25636
rect 246 -25812 258 -25636
rect 200 -25824 258 -25812
rect -258 -26072 -200 -26060
rect -258 -26248 -246 -26072
rect -212 -26248 -200 -26072
rect -258 -26260 -200 -26248
rect 200 -26072 258 -26060
rect 200 -26248 212 -26072
rect 246 -26248 258 -26072
rect 200 -26260 258 -26248
rect -258 -26508 -200 -26496
rect -258 -26684 -246 -26508
rect -212 -26684 -200 -26508
rect -258 -26696 -200 -26684
rect 200 -26508 258 -26496
rect 200 -26684 212 -26508
rect 246 -26684 258 -26508
rect 200 -26696 258 -26684
rect -258 -26944 -200 -26932
rect -258 -27120 -246 -26944
rect -212 -27120 -200 -26944
rect -258 -27132 -200 -27120
rect 200 -26944 258 -26932
rect 200 -27120 212 -26944
rect 246 -27120 258 -26944
rect 200 -27132 258 -27120
rect -258 -27380 -200 -27368
rect -258 -27556 -246 -27380
rect -212 -27556 -200 -27380
rect -258 -27568 -200 -27556
rect 200 -27380 258 -27368
rect 200 -27556 212 -27380
rect 246 -27556 258 -27380
rect 200 -27568 258 -27556
rect -258 -27816 -200 -27804
rect -258 -27992 -246 -27816
rect -212 -27992 -200 -27816
rect -258 -28004 -200 -27992
rect 200 -27816 258 -27804
rect 200 -27992 212 -27816
rect 246 -27992 258 -27816
rect 200 -28004 258 -27992
rect -258 -28252 -200 -28240
rect -258 -28428 -246 -28252
rect -212 -28428 -200 -28252
rect -258 -28440 -200 -28428
rect 200 -28252 258 -28240
rect 200 -28428 212 -28252
rect 246 -28428 258 -28252
rect 200 -28440 258 -28428
rect -258 -28688 -200 -28676
rect -258 -28864 -246 -28688
rect -212 -28864 -200 -28688
rect -258 -28876 -200 -28864
rect 200 -28688 258 -28676
rect 200 -28864 212 -28688
rect 246 -28864 258 -28688
rect 200 -28876 258 -28864
rect -258 -29124 -200 -29112
rect -258 -29300 -246 -29124
rect -212 -29300 -200 -29124
rect -258 -29312 -200 -29300
rect 200 -29124 258 -29112
rect 200 -29300 212 -29124
rect 246 -29300 258 -29124
rect 200 -29312 258 -29300
rect -258 -29560 -200 -29548
rect -258 -29736 -246 -29560
rect -212 -29736 -200 -29560
rect -258 -29748 -200 -29736
rect 200 -29560 258 -29548
rect 200 -29736 212 -29560
rect 246 -29736 258 -29560
rect 200 -29748 258 -29736
rect -258 -29996 -200 -29984
rect -258 -30172 -246 -29996
rect -212 -30172 -200 -29996
rect -258 -30184 -200 -30172
rect 200 -29996 258 -29984
rect 200 -30172 212 -29996
rect 246 -30172 258 -29996
rect 200 -30184 258 -30172
rect -258 -30432 -200 -30420
rect -258 -30608 -246 -30432
rect -212 -30608 -200 -30432
rect -258 -30620 -200 -30608
rect 200 -30432 258 -30420
rect 200 -30608 212 -30432
rect 246 -30608 258 -30432
rect 200 -30620 258 -30608
rect -258 -30868 -200 -30856
rect -258 -31044 -246 -30868
rect -212 -31044 -200 -30868
rect -258 -31056 -200 -31044
rect 200 -30868 258 -30856
rect 200 -31044 212 -30868
rect 246 -31044 258 -30868
rect 200 -31056 258 -31044
rect -258 -31304 -200 -31292
rect -258 -31480 -246 -31304
rect -212 -31480 -200 -31304
rect -258 -31492 -200 -31480
rect 200 -31304 258 -31292
rect 200 -31480 212 -31304
rect 246 -31480 258 -31304
rect 200 -31492 258 -31480
rect -258 -31740 -200 -31728
rect -258 -31916 -246 -31740
rect -212 -31916 -200 -31740
rect -258 -31928 -200 -31916
rect 200 -31740 258 -31728
rect 200 -31916 212 -31740
rect 246 -31916 258 -31740
rect 200 -31928 258 -31916
rect -258 -32176 -200 -32164
rect -258 -32352 -246 -32176
rect -212 -32352 -200 -32176
rect -258 -32364 -200 -32352
rect 200 -32176 258 -32164
rect 200 -32352 212 -32176
rect 246 -32352 258 -32176
rect 200 -32364 258 -32352
rect -258 -32612 -200 -32600
rect -258 -32788 -246 -32612
rect -212 -32788 -200 -32612
rect -258 -32800 -200 -32788
rect 200 -32612 258 -32600
rect 200 -32788 212 -32612
rect 246 -32788 258 -32612
rect 200 -32800 258 -32788
rect -258 -33048 -200 -33036
rect -258 -33224 -246 -33048
rect -212 -33224 -200 -33048
rect -258 -33236 -200 -33224
rect 200 -33048 258 -33036
rect 200 -33224 212 -33048
rect 246 -33224 258 -33048
rect 200 -33236 258 -33224
rect -258 -33484 -200 -33472
rect -258 -33660 -246 -33484
rect -212 -33660 -200 -33484
rect -258 -33672 -200 -33660
rect 200 -33484 258 -33472
rect 200 -33660 212 -33484
rect 246 -33660 258 -33484
rect 200 -33672 258 -33660
rect -258 -33920 -200 -33908
rect -258 -34096 -246 -33920
rect -212 -34096 -200 -33920
rect -258 -34108 -200 -34096
rect 200 -33920 258 -33908
rect 200 -34096 212 -33920
rect 246 -34096 258 -33920
rect 200 -34108 258 -34096
rect -258 -34356 -200 -34344
rect -258 -34532 -246 -34356
rect -212 -34532 -200 -34356
rect -258 -34544 -200 -34532
rect 200 -34356 258 -34344
rect 200 -34532 212 -34356
rect 246 -34532 258 -34356
rect 200 -34544 258 -34532
rect -258 -34792 -200 -34780
rect -258 -34968 -246 -34792
rect -212 -34968 -200 -34792
rect -258 -34980 -200 -34968
rect 200 -34792 258 -34780
rect 200 -34968 212 -34792
rect 246 -34968 258 -34792
rect 200 -34980 258 -34968
rect -258 -35228 -200 -35216
rect -258 -35404 -246 -35228
rect -212 -35404 -200 -35228
rect -258 -35416 -200 -35404
rect 200 -35228 258 -35216
rect 200 -35404 212 -35228
rect 246 -35404 258 -35228
rect 200 -35416 258 -35404
rect -258 -35664 -200 -35652
rect -258 -35840 -246 -35664
rect -212 -35840 -200 -35664
rect -258 -35852 -200 -35840
rect 200 -35664 258 -35652
rect 200 -35840 212 -35664
rect 246 -35840 258 -35664
rect 200 -35852 258 -35840
rect -258 -36100 -200 -36088
rect -258 -36276 -246 -36100
rect -212 -36276 -200 -36100
rect -258 -36288 -200 -36276
rect 200 -36100 258 -36088
rect 200 -36276 212 -36100
rect 246 -36276 258 -36100
rect 200 -36288 258 -36276
rect -258 -36536 -200 -36524
rect -258 -36712 -246 -36536
rect -212 -36712 -200 -36536
rect -258 -36724 -200 -36712
rect 200 -36536 258 -36524
rect 200 -36712 212 -36536
rect 246 -36712 258 -36536
rect 200 -36724 258 -36712
rect -258 -36972 -200 -36960
rect -258 -37148 -246 -36972
rect -212 -37148 -200 -36972
rect -258 -37160 -200 -37148
rect 200 -36972 258 -36960
rect 200 -37148 212 -36972
rect 246 -37148 258 -36972
rect 200 -37160 258 -37148
rect -258 -37408 -200 -37396
rect -258 -37584 -246 -37408
rect -212 -37584 -200 -37408
rect -258 -37596 -200 -37584
rect 200 -37408 258 -37396
rect 200 -37584 212 -37408
rect 246 -37584 258 -37408
rect 200 -37596 258 -37584
rect -258 -37844 -200 -37832
rect -258 -38020 -246 -37844
rect -212 -38020 -200 -37844
rect -258 -38032 -200 -38020
rect 200 -37844 258 -37832
rect 200 -38020 212 -37844
rect 246 -38020 258 -37844
rect 200 -38032 258 -38020
rect -258 -38280 -200 -38268
rect -258 -38456 -246 -38280
rect -212 -38456 -200 -38280
rect -258 -38468 -200 -38456
rect 200 -38280 258 -38268
rect 200 -38456 212 -38280
rect 246 -38456 258 -38280
rect 200 -38468 258 -38456
rect -258 -38716 -200 -38704
rect -258 -38892 -246 -38716
rect -212 -38892 -200 -38716
rect -258 -38904 -200 -38892
rect 200 -38716 258 -38704
rect 200 -38892 212 -38716
rect 246 -38892 258 -38716
rect 200 -38904 258 -38892
rect -258 -39152 -200 -39140
rect -258 -39328 -246 -39152
rect -212 -39328 -200 -39152
rect -258 -39340 -200 -39328
rect 200 -39152 258 -39140
rect 200 -39328 212 -39152
rect 246 -39328 258 -39152
rect 200 -39340 258 -39328
rect -258 -39588 -200 -39576
rect -258 -39764 -246 -39588
rect -212 -39764 -200 -39588
rect -258 -39776 -200 -39764
rect 200 -39588 258 -39576
rect 200 -39764 212 -39588
rect 246 -39764 258 -39588
rect 200 -39776 258 -39764
rect -258 -40024 -200 -40012
rect -258 -40200 -246 -40024
rect -212 -40200 -200 -40024
rect -258 -40212 -200 -40200
rect 200 -40024 258 -40012
rect 200 -40200 212 -40024
rect 246 -40200 258 -40024
rect 200 -40212 258 -40200
rect -258 -40460 -200 -40448
rect -258 -40636 -246 -40460
rect -212 -40636 -200 -40460
rect -258 -40648 -200 -40636
rect 200 -40460 258 -40448
rect 200 -40636 212 -40460
rect 246 -40636 258 -40460
rect 200 -40648 258 -40636
rect -258 -40896 -200 -40884
rect -258 -41072 -246 -40896
rect -212 -41072 -200 -40896
rect -258 -41084 -200 -41072
rect 200 -40896 258 -40884
rect 200 -41072 212 -40896
rect 246 -41072 258 -40896
rect 200 -41084 258 -41072
rect -258 -41332 -200 -41320
rect -258 -41508 -246 -41332
rect -212 -41508 -200 -41332
rect -258 -41520 -200 -41508
rect 200 -41332 258 -41320
rect 200 -41508 212 -41332
rect 246 -41508 258 -41332
rect 200 -41520 258 -41508
rect -258 -41768 -200 -41756
rect -258 -41944 -246 -41768
rect -212 -41944 -200 -41768
rect -258 -41956 -200 -41944
rect 200 -41768 258 -41756
rect 200 -41944 212 -41768
rect 246 -41944 258 -41768
rect 200 -41956 258 -41944
rect -258 -42204 -200 -42192
rect -258 -42380 -246 -42204
rect -212 -42380 -200 -42204
rect -258 -42392 -200 -42380
rect 200 -42204 258 -42192
rect 200 -42380 212 -42204
rect 246 -42380 258 -42204
rect 200 -42392 258 -42380
rect -258 -42640 -200 -42628
rect -258 -42816 -246 -42640
rect -212 -42816 -200 -42640
rect -258 -42828 -200 -42816
rect 200 -42640 258 -42628
rect 200 -42816 212 -42640
rect 246 -42816 258 -42640
rect 200 -42828 258 -42816
rect -258 -43076 -200 -43064
rect -258 -43252 -246 -43076
rect -212 -43252 -200 -43076
rect -258 -43264 -200 -43252
rect 200 -43076 258 -43064
rect 200 -43252 212 -43076
rect 246 -43252 258 -43076
rect 200 -43264 258 -43252
rect -258 -43512 -200 -43500
rect -258 -43688 -246 -43512
rect -212 -43688 -200 -43512
rect -258 -43700 -200 -43688
rect 200 -43512 258 -43500
rect 200 -43688 212 -43512
rect 246 -43688 258 -43512
rect 200 -43700 258 -43688
rect -258 -43948 -200 -43936
rect -258 -44124 -246 -43948
rect -212 -44124 -200 -43948
rect -258 -44136 -200 -44124
rect 200 -43948 258 -43936
rect 200 -44124 212 -43948
rect 246 -44124 258 -43948
rect 200 -44136 258 -44124
rect -258 -44384 -200 -44372
rect -258 -44560 -246 -44384
rect -212 -44560 -200 -44384
rect -258 -44572 -200 -44560
rect 200 -44384 258 -44372
rect 200 -44560 212 -44384
rect 246 -44560 258 -44384
rect 200 -44572 258 -44560
rect -258 -44820 -200 -44808
rect -258 -44996 -246 -44820
rect -212 -44996 -200 -44820
rect -258 -45008 -200 -44996
rect 200 -44820 258 -44808
rect 200 -44996 212 -44820
rect 246 -44996 258 -44820
rect 200 -45008 258 -44996
rect -258 -45256 -200 -45244
rect -258 -45432 -246 -45256
rect -212 -45432 -200 -45256
rect -258 -45444 -200 -45432
rect 200 -45256 258 -45244
rect 200 -45432 212 -45256
rect 246 -45432 258 -45256
rect 200 -45444 258 -45432
rect -258 -45692 -200 -45680
rect -258 -45868 -246 -45692
rect -212 -45868 -200 -45692
rect -258 -45880 -200 -45868
rect 200 -45692 258 -45680
rect 200 -45868 212 -45692
rect 246 -45868 258 -45692
rect 200 -45880 258 -45868
rect -258 -46128 -200 -46116
rect -258 -46304 -246 -46128
rect -212 -46304 -200 -46128
rect -258 -46316 -200 -46304
rect 200 -46128 258 -46116
rect 200 -46304 212 -46128
rect 246 -46304 258 -46128
rect 200 -46316 258 -46304
rect -258 -46564 -200 -46552
rect -258 -46740 -246 -46564
rect -212 -46740 -200 -46564
rect -258 -46752 -200 -46740
rect 200 -46564 258 -46552
rect 200 -46740 212 -46564
rect 246 -46740 258 -46564
rect 200 -46752 258 -46740
rect -258 -47000 -200 -46988
rect -258 -47176 -246 -47000
rect -212 -47176 -200 -47000
rect -258 -47188 -200 -47176
rect 200 -47000 258 -46988
rect 200 -47176 212 -47000
rect 246 -47176 258 -47000
rect 200 -47188 258 -47176
rect -258 -47436 -200 -47424
rect -258 -47612 -246 -47436
rect -212 -47612 -200 -47436
rect -258 -47624 -200 -47612
rect 200 -47436 258 -47424
rect 200 -47612 212 -47436
rect 246 -47612 258 -47436
rect 200 -47624 258 -47612
rect -258 -47872 -200 -47860
rect -258 -48048 -246 -47872
rect -212 -48048 -200 -47872
rect -258 -48060 -200 -48048
rect 200 -47872 258 -47860
rect 200 -48048 212 -47872
rect 246 -48048 258 -47872
rect 200 -48060 258 -48048
rect -258 -48308 -200 -48296
rect -258 -48484 -246 -48308
rect -212 -48484 -200 -48308
rect -258 -48496 -200 -48484
rect 200 -48308 258 -48296
rect 200 -48484 212 -48308
rect 246 -48484 258 -48308
rect 200 -48496 258 -48484
rect -258 -48744 -200 -48732
rect -258 -48920 -246 -48744
rect -212 -48920 -200 -48744
rect -258 -48932 -200 -48920
rect 200 -48744 258 -48732
rect 200 -48920 212 -48744
rect 246 -48920 258 -48744
rect 200 -48932 258 -48920
rect -258 -49180 -200 -49168
rect -258 -49356 -246 -49180
rect -212 -49356 -200 -49180
rect -258 -49368 -200 -49356
rect 200 -49180 258 -49168
rect 200 -49356 212 -49180
rect 246 -49356 258 -49180
rect 200 -49368 258 -49356
rect -258 -49616 -200 -49604
rect -258 -49792 -246 -49616
rect -212 -49792 -200 -49616
rect -258 -49804 -200 -49792
rect 200 -49616 258 -49604
rect 200 -49792 212 -49616
rect 246 -49792 258 -49616
rect 200 -49804 258 -49792
rect -258 -50052 -200 -50040
rect -258 -50228 -246 -50052
rect -212 -50228 -200 -50052
rect -258 -50240 -200 -50228
rect 200 -50052 258 -50040
rect 200 -50228 212 -50052
rect 246 -50228 258 -50052
rect 200 -50240 258 -50228
rect -258 -50488 -200 -50476
rect -258 -50664 -246 -50488
rect -212 -50664 -200 -50488
rect -258 -50676 -200 -50664
rect 200 -50488 258 -50476
rect 200 -50664 212 -50488
rect 246 -50664 258 -50488
rect 200 -50676 258 -50664
rect -258 -50924 -200 -50912
rect -258 -51100 -246 -50924
rect -212 -51100 -200 -50924
rect -258 -51112 -200 -51100
rect 200 -50924 258 -50912
rect 200 -51100 212 -50924
rect 246 -51100 258 -50924
rect 200 -51112 258 -51100
rect -258 -51360 -200 -51348
rect -258 -51536 -246 -51360
rect -212 -51536 -200 -51360
rect -258 -51548 -200 -51536
rect 200 -51360 258 -51348
rect 200 -51536 212 -51360
rect 246 -51536 258 -51360
rect 200 -51548 258 -51536
rect -258 -51796 -200 -51784
rect -258 -51972 -246 -51796
rect -212 -51972 -200 -51796
rect -258 -51984 -200 -51972
rect 200 -51796 258 -51784
rect 200 -51972 212 -51796
rect 246 -51972 258 -51796
rect 200 -51984 258 -51972
rect -258 -52232 -200 -52220
rect -258 -52408 -246 -52232
rect -212 -52408 -200 -52232
rect -258 -52420 -200 -52408
rect 200 -52232 258 -52220
rect 200 -52408 212 -52232
rect 246 -52408 258 -52232
rect 200 -52420 258 -52408
rect -258 -52668 -200 -52656
rect -258 -52844 -246 -52668
rect -212 -52844 -200 -52668
rect -258 -52856 -200 -52844
rect 200 -52668 258 -52656
rect 200 -52844 212 -52668
rect 246 -52844 258 -52668
rect 200 -52856 258 -52844
rect -258 -53104 -200 -53092
rect -258 -53280 -246 -53104
rect -212 -53280 -200 -53104
rect -258 -53292 -200 -53280
rect 200 -53104 258 -53092
rect 200 -53280 212 -53104
rect 246 -53280 258 -53104
rect 200 -53292 258 -53280
rect -258 -53540 -200 -53528
rect -258 -53716 -246 -53540
rect -212 -53716 -200 -53540
rect -258 -53728 -200 -53716
rect 200 -53540 258 -53528
rect 200 -53716 212 -53540
rect 246 -53716 258 -53540
rect 200 -53728 258 -53716
rect -258 -53976 -200 -53964
rect -258 -54152 -246 -53976
rect -212 -54152 -200 -53976
rect -258 -54164 -200 -54152
rect 200 -53976 258 -53964
rect 200 -54152 212 -53976
rect 246 -54152 258 -53976
rect 200 -54164 258 -54152
rect -258 -54412 -200 -54400
rect -258 -54588 -246 -54412
rect -212 -54588 -200 -54412
rect -258 -54600 -200 -54588
rect 200 -54412 258 -54400
rect 200 -54588 212 -54412
rect 246 -54588 258 -54412
rect 200 -54600 258 -54588
rect -258 -54848 -200 -54836
rect -258 -55024 -246 -54848
rect -212 -55024 -200 -54848
rect -258 -55036 -200 -55024
rect 200 -54848 258 -54836
rect 200 -55024 212 -54848
rect 246 -55024 258 -54848
rect 200 -55036 258 -55024
rect -258 -55284 -200 -55272
rect -258 -55460 -246 -55284
rect -212 -55460 -200 -55284
rect -258 -55472 -200 -55460
rect 200 -55284 258 -55272
rect 200 -55460 212 -55284
rect 246 -55460 258 -55284
rect 200 -55472 258 -55460
rect -258 -55720 -200 -55708
rect -258 -55896 -246 -55720
rect -212 -55896 -200 -55720
rect -258 -55908 -200 -55896
rect 200 -55720 258 -55708
rect 200 -55896 212 -55720
rect 246 -55896 258 -55720
rect 200 -55908 258 -55896
rect -258 -56156 -200 -56144
rect -258 -56332 -246 -56156
rect -212 -56332 -200 -56156
rect -258 -56344 -200 -56332
rect 200 -56156 258 -56144
rect 200 -56332 212 -56156
rect 246 -56332 258 -56156
rect 200 -56344 258 -56332
rect -258 -56592 -200 -56580
rect -258 -56768 -246 -56592
rect -212 -56768 -200 -56592
rect -258 -56780 -200 -56768
rect 200 -56592 258 -56580
rect 200 -56768 212 -56592
rect 246 -56768 258 -56592
rect 200 -56780 258 -56768
rect -258 -57028 -200 -57016
rect -258 -57204 -246 -57028
rect -212 -57204 -200 -57028
rect -258 -57216 -200 -57204
rect 200 -57028 258 -57016
rect 200 -57204 212 -57028
rect 246 -57204 258 -57028
rect 200 -57216 258 -57204
rect -258 -57464 -200 -57452
rect -258 -57640 -246 -57464
rect -212 -57640 -200 -57464
rect -258 -57652 -200 -57640
rect 200 -57464 258 -57452
rect 200 -57640 212 -57464
rect 246 -57640 258 -57464
rect 200 -57652 258 -57640
rect -258 -57900 -200 -57888
rect -258 -58076 -246 -57900
rect -212 -58076 -200 -57900
rect -258 -58088 -200 -58076
rect 200 -57900 258 -57888
rect 200 -58076 212 -57900
rect 246 -58076 258 -57900
rect 200 -58088 258 -58076
rect -258 -58336 -200 -58324
rect -258 -58512 -246 -58336
rect -212 -58512 -200 -58336
rect -258 -58524 -200 -58512
rect 200 -58336 258 -58324
rect 200 -58512 212 -58336
rect 246 -58512 258 -58336
rect 200 -58524 258 -58512
rect -258 -58772 -200 -58760
rect -258 -58948 -246 -58772
rect -212 -58948 -200 -58772
rect -258 -58960 -200 -58948
rect 200 -58772 258 -58760
rect 200 -58948 212 -58772
rect 246 -58948 258 -58772
rect 200 -58960 258 -58948
rect -258 -59208 -200 -59196
rect -258 -59384 -246 -59208
rect -212 -59384 -200 -59208
rect -258 -59396 -200 -59384
rect 200 -59208 258 -59196
rect 200 -59384 212 -59208
rect 246 -59384 258 -59208
rect 200 -59396 258 -59384
rect -258 -59644 -200 -59632
rect -258 -59820 -246 -59644
rect -212 -59820 -200 -59644
rect -258 -59832 -200 -59820
rect 200 -59644 258 -59632
rect 200 -59820 212 -59644
rect 246 -59820 258 -59644
rect 200 -59832 258 -59820
rect -258 -60080 -200 -60068
rect -258 -60256 -246 -60080
rect -212 -60256 -200 -60080
rect -258 -60268 -200 -60256
rect 200 -60080 258 -60068
rect 200 -60256 212 -60080
rect 246 -60256 258 -60080
rect 200 -60268 258 -60256
rect -258 -60516 -200 -60504
rect -258 -60692 -246 -60516
rect -212 -60692 -200 -60516
rect -258 -60704 -200 -60692
rect 200 -60516 258 -60504
rect 200 -60692 212 -60516
rect 246 -60692 258 -60516
rect 200 -60704 258 -60692
rect -258 -60952 -200 -60940
rect -258 -61128 -246 -60952
rect -212 -61128 -200 -60952
rect -258 -61140 -200 -61128
rect 200 -60952 258 -60940
rect 200 -61128 212 -60952
rect 246 -61128 258 -60952
rect 200 -61140 258 -61128
rect -258 -61388 -200 -61376
rect -258 -61564 -246 -61388
rect -212 -61564 -200 -61388
rect -258 -61576 -200 -61564
rect 200 -61388 258 -61376
rect 200 -61564 212 -61388
rect 246 -61564 258 -61388
rect 200 -61576 258 -61564
rect -258 -61824 -200 -61812
rect -258 -62000 -246 -61824
rect -212 -62000 -200 -61824
rect -258 -62012 -200 -62000
rect 200 -61824 258 -61812
rect 200 -62000 212 -61824
rect 246 -62000 258 -61824
rect 200 -62012 258 -62000
rect -258 -62260 -200 -62248
rect -258 -62436 -246 -62260
rect -212 -62436 -200 -62260
rect -258 -62448 -200 -62436
rect 200 -62260 258 -62248
rect 200 -62436 212 -62260
rect 246 -62436 258 -62260
rect 200 -62448 258 -62436
rect -258 -62696 -200 -62684
rect -258 -62872 -246 -62696
rect -212 -62872 -200 -62696
rect -258 -62884 -200 -62872
rect 200 -62696 258 -62684
rect 200 -62872 212 -62696
rect 246 -62872 258 -62696
rect 200 -62884 258 -62872
rect -258 -63132 -200 -63120
rect -258 -63308 -246 -63132
rect -212 -63308 -200 -63132
rect -258 -63320 -200 -63308
rect 200 -63132 258 -63120
rect 200 -63308 212 -63132
rect 246 -63308 258 -63132
rect 200 -63320 258 -63308
rect -258 -63568 -200 -63556
rect -258 -63744 -246 -63568
rect -212 -63744 -200 -63568
rect -258 -63756 -200 -63744
rect 200 -63568 258 -63556
rect 200 -63744 212 -63568
rect 246 -63744 258 -63568
rect 200 -63756 258 -63744
rect -258 -64004 -200 -63992
rect -258 -64180 -246 -64004
rect -212 -64180 -200 -64004
rect -258 -64192 -200 -64180
rect 200 -64004 258 -63992
rect 200 -64180 212 -64004
rect 246 -64180 258 -64004
rect 200 -64192 258 -64180
rect -258 -64440 -200 -64428
rect -258 -64616 -246 -64440
rect -212 -64616 -200 -64440
rect -258 -64628 -200 -64616
rect 200 -64440 258 -64428
rect 200 -64616 212 -64440
rect 246 -64616 258 -64440
rect 200 -64628 258 -64616
rect -258 -64876 -200 -64864
rect -258 -65052 -246 -64876
rect -212 -65052 -200 -64876
rect -258 -65064 -200 -65052
rect 200 -64876 258 -64864
rect 200 -65052 212 -64876
rect 246 -65052 258 -64876
rect 200 -65064 258 -65052
rect -258 -65312 -200 -65300
rect -258 -65488 -246 -65312
rect -212 -65488 -200 -65312
rect -258 -65500 -200 -65488
rect 200 -65312 258 -65300
rect 200 -65488 212 -65312
rect 246 -65488 258 -65312
rect 200 -65500 258 -65488
rect -258 -65748 -200 -65736
rect -258 -65924 -246 -65748
rect -212 -65924 -200 -65748
rect -258 -65936 -200 -65924
rect 200 -65748 258 -65736
rect 200 -65924 212 -65748
rect 246 -65924 258 -65748
rect 200 -65936 258 -65924
rect -258 -66184 -200 -66172
rect -258 -66360 -246 -66184
rect -212 -66360 -200 -66184
rect -258 -66372 -200 -66360
rect 200 -66184 258 -66172
rect 200 -66360 212 -66184
rect 246 -66360 258 -66184
rect 200 -66372 258 -66360
rect -258 -66620 -200 -66608
rect -258 -66796 -246 -66620
rect -212 -66796 -200 -66620
rect -258 -66808 -200 -66796
rect 200 -66620 258 -66608
rect 200 -66796 212 -66620
rect 246 -66796 258 -66620
rect 200 -66808 258 -66796
rect -258 -67056 -200 -67044
rect -258 -67232 -246 -67056
rect -212 -67232 -200 -67056
rect -258 -67244 -200 -67232
rect 200 -67056 258 -67044
rect 200 -67232 212 -67056
rect 246 -67232 258 -67056
rect 200 -67244 258 -67232
rect -258 -67492 -200 -67480
rect -258 -67668 -246 -67492
rect -212 -67668 -200 -67492
rect -258 -67680 -200 -67668
rect 200 -67492 258 -67480
rect 200 -67668 212 -67492
rect 246 -67668 258 -67492
rect 200 -67680 258 -67668
rect -258 -67928 -200 -67916
rect -258 -68104 -246 -67928
rect -212 -68104 -200 -67928
rect -258 -68116 -200 -68104
rect 200 -67928 258 -67916
rect 200 -68104 212 -67928
rect 246 -68104 258 -67928
rect 200 -68116 258 -68104
rect -258 -68364 -200 -68352
rect -258 -68540 -246 -68364
rect -212 -68540 -200 -68364
rect -258 -68552 -200 -68540
rect 200 -68364 258 -68352
rect 200 -68540 212 -68364
rect 246 -68540 258 -68364
rect 200 -68552 258 -68540
rect -258 -68800 -200 -68788
rect -258 -68976 -246 -68800
rect -212 -68976 -200 -68800
rect -258 -68988 -200 -68976
rect 200 -68800 258 -68788
rect 200 -68976 212 -68800
rect 246 -68976 258 -68800
rect 200 -68988 258 -68976
rect -258 -69236 -200 -69224
rect -258 -69412 -246 -69236
rect -212 -69412 -200 -69236
rect -258 -69424 -200 -69412
rect 200 -69236 258 -69224
rect 200 -69412 212 -69236
rect 246 -69412 258 -69236
rect 200 -69424 258 -69412
rect -258 -69672 -200 -69660
rect -258 -69848 -246 -69672
rect -212 -69848 -200 -69672
rect -258 -69860 -200 -69848
rect 200 -69672 258 -69660
rect 200 -69848 212 -69672
rect 246 -69848 258 -69672
rect 200 -69860 258 -69848
rect -258 -70108 -200 -70096
rect -258 -70284 -246 -70108
rect -212 -70284 -200 -70108
rect -258 -70296 -200 -70284
rect 200 -70108 258 -70096
rect 200 -70284 212 -70108
rect 246 -70284 258 -70108
rect 200 -70296 258 -70284
rect -258 -70544 -200 -70532
rect -258 -70720 -246 -70544
rect -212 -70720 -200 -70544
rect -258 -70732 -200 -70720
rect 200 -70544 258 -70532
rect 200 -70720 212 -70544
rect 246 -70720 258 -70544
rect 200 -70732 258 -70720
rect -258 -70980 -200 -70968
rect -258 -71156 -246 -70980
rect -212 -71156 -200 -70980
rect -258 -71168 -200 -71156
rect 200 -70980 258 -70968
rect 200 -71156 212 -70980
rect 246 -71156 258 -70980
rect 200 -71168 258 -71156
rect -258 -71416 -200 -71404
rect -258 -71592 -246 -71416
rect -212 -71592 -200 -71416
rect -258 -71604 -200 -71592
rect 200 -71416 258 -71404
rect 200 -71592 212 -71416
rect 246 -71592 258 -71416
rect 200 -71604 258 -71592
rect -258 -71852 -200 -71840
rect -258 -72028 -246 -71852
rect -212 -72028 -200 -71852
rect -258 -72040 -200 -72028
rect 200 -71852 258 -71840
rect 200 -72028 212 -71852
rect 246 -72028 258 -71852
rect 200 -72040 258 -72028
rect -258 -72288 -200 -72276
rect -258 -72464 -246 -72288
rect -212 -72464 -200 -72288
rect -258 -72476 -200 -72464
rect 200 -72288 258 -72276
rect 200 -72464 212 -72288
rect 246 -72464 258 -72288
rect 200 -72476 258 -72464
rect -258 -72724 -200 -72712
rect -258 -72900 -246 -72724
rect -212 -72900 -200 -72724
rect -258 -72912 -200 -72900
rect 200 -72724 258 -72712
rect 200 -72900 212 -72724
rect 246 -72900 258 -72724
rect 200 -72912 258 -72900
rect -258 -73160 -200 -73148
rect -258 -73336 -246 -73160
rect -212 -73336 -200 -73160
rect -258 -73348 -200 -73336
rect 200 -73160 258 -73148
rect 200 -73336 212 -73160
rect 246 -73336 258 -73160
rect 200 -73348 258 -73336
rect -258 -73596 -200 -73584
rect -258 -73772 -246 -73596
rect -212 -73772 -200 -73596
rect -258 -73784 -200 -73772
rect 200 -73596 258 -73584
rect 200 -73772 212 -73596
rect 246 -73772 258 -73596
rect 200 -73784 258 -73772
rect -258 -74032 -200 -74020
rect -258 -74208 -246 -74032
rect -212 -74208 -200 -74032
rect -258 -74220 -200 -74208
rect 200 -74032 258 -74020
rect 200 -74208 212 -74032
rect 246 -74208 258 -74032
rect 200 -74220 258 -74208
rect -258 -74468 -200 -74456
rect -258 -74644 -246 -74468
rect -212 -74644 -200 -74468
rect -258 -74656 -200 -74644
rect 200 -74468 258 -74456
rect 200 -74644 212 -74468
rect 246 -74644 258 -74468
rect 200 -74656 258 -74644
rect -258 -74904 -200 -74892
rect -258 -75080 -246 -74904
rect -212 -75080 -200 -74904
rect -258 -75092 -200 -75080
rect 200 -74904 258 -74892
rect 200 -75080 212 -74904
rect 246 -75080 258 -74904
rect 200 -75092 258 -75080
rect -258 -75340 -200 -75328
rect -258 -75516 -246 -75340
rect -212 -75516 -200 -75340
rect -258 -75528 -200 -75516
rect 200 -75340 258 -75328
rect 200 -75516 212 -75340
rect 246 -75516 258 -75340
rect 200 -75528 258 -75516
rect -258 -75776 -200 -75764
rect -258 -75952 -246 -75776
rect -212 -75952 -200 -75776
rect -258 -75964 -200 -75952
rect 200 -75776 258 -75764
rect 200 -75952 212 -75776
rect 246 -75952 258 -75776
rect 200 -75964 258 -75952
rect -258 -76212 -200 -76200
rect -258 -76388 -246 -76212
rect -212 -76388 -200 -76212
rect -258 -76400 -200 -76388
rect 200 -76212 258 -76200
rect 200 -76388 212 -76212
rect 246 -76388 258 -76212
rect 200 -76400 258 -76388
rect -258 -76648 -200 -76636
rect -258 -76824 -246 -76648
rect -212 -76824 -200 -76648
rect -258 -76836 -200 -76824
rect 200 -76648 258 -76636
rect 200 -76824 212 -76648
rect 246 -76824 258 -76648
rect 200 -76836 258 -76824
rect -258 -77084 -200 -77072
rect -258 -77260 -246 -77084
rect -212 -77260 -200 -77084
rect -258 -77272 -200 -77260
rect 200 -77084 258 -77072
rect 200 -77260 212 -77084
rect 246 -77260 258 -77084
rect 200 -77272 258 -77260
rect -258 -77520 -200 -77508
rect -258 -77696 -246 -77520
rect -212 -77696 -200 -77520
rect -258 -77708 -200 -77696
rect 200 -77520 258 -77508
rect 200 -77696 212 -77520
rect 246 -77696 258 -77520
rect 200 -77708 258 -77696
rect -258 -77956 -200 -77944
rect -258 -78132 -246 -77956
rect -212 -78132 -200 -77956
rect -258 -78144 -200 -78132
rect 200 -77956 258 -77944
rect 200 -78132 212 -77956
rect 246 -78132 258 -77956
rect 200 -78144 258 -78132
rect -258 -78392 -200 -78380
rect -258 -78568 -246 -78392
rect -212 -78568 -200 -78392
rect -258 -78580 -200 -78568
rect 200 -78392 258 -78380
rect 200 -78568 212 -78392
rect 246 -78568 258 -78392
rect 200 -78580 258 -78568
rect -258 -78828 -200 -78816
rect -258 -79004 -246 -78828
rect -212 -79004 -200 -78828
rect -258 -79016 -200 -79004
rect 200 -78828 258 -78816
rect 200 -79004 212 -78828
rect 246 -79004 258 -78828
rect 200 -79016 258 -79004
rect -258 -79264 -200 -79252
rect -258 -79440 -246 -79264
rect -212 -79440 -200 -79264
rect -258 -79452 -200 -79440
rect 200 -79264 258 -79252
rect 200 -79440 212 -79264
rect 246 -79440 258 -79264
rect 200 -79452 258 -79440
rect -258 -79700 -200 -79688
rect -258 -79876 -246 -79700
rect -212 -79876 -200 -79700
rect -258 -79888 -200 -79876
rect 200 -79700 258 -79688
rect 200 -79876 212 -79700
rect 246 -79876 258 -79700
rect 200 -79888 258 -79876
rect -258 -80136 -200 -80124
rect -258 -80312 -246 -80136
rect -212 -80312 -200 -80136
rect -258 -80324 -200 -80312
rect 200 -80136 258 -80124
rect 200 -80312 212 -80136
rect 246 -80312 258 -80136
rect 200 -80324 258 -80312
rect -258 -80572 -200 -80560
rect -258 -80748 -246 -80572
rect -212 -80748 -200 -80572
rect -258 -80760 -200 -80748
rect 200 -80572 258 -80560
rect 200 -80748 212 -80572
rect 246 -80748 258 -80572
rect 200 -80760 258 -80748
rect -258 -81008 -200 -80996
rect -258 -81184 -246 -81008
rect -212 -81184 -200 -81008
rect -258 -81196 -200 -81184
rect 200 -81008 258 -80996
rect 200 -81184 212 -81008
rect 246 -81184 258 -81008
rect 200 -81196 258 -81184
rect -258 -81444 -200 -81432
rect -258 -81620 -246 -81444
rect -212 -81620 -200 -81444
rect -258 -81632 -200 -81620
rect 200 -81444 258 -81432
rect 200 -81620 212 -81444
rect 246 -81620 258 -81444
rect 200 -81632 258 -81620
rect -258 -81880 -200 -81868
rect -258 -82056 -246 -81880
rect -212 -82056 -200 -81880
rect -258 -82068 -200 -82056
rect 200 -81880 258 -81868
rect 200 -82056 212 -81880
rect 246 -82056 258 -81880
rect 200 -82068 258 -82056
rect -258 -82316 -200 -82304
rect -258 -82492 -246 -82316
rect -212 -82492 -200 -82316
rect -258 -82504 -200 -82492
rect 200 -82316 258 -82304
rect 200 -82492 212 -82316
rect 246 -82492 258 -82316
rect 200 -82504 258 -82492
rect -258 -82752 -200 -82740
rect -258 -82928 -246 -82752
rect -212 -82928 -200 -82752
rect -258 -82940 -200 -82928
rect 200 -82752 258 -82740
rect 200 -82928 212 -82752
rect 246 -82928 258 -82752
rect 200 -82940 258 -82928
rect -258 -83188 -200 -83176
rect -258 -83364 -246 -83188
rect -212 -83364 -200 -83188
rect -258 -83376 -200 -83364
rect 200 -83188 258 -83176
rect 200 -83364 212 -83188
rect 246 -83364 258 -83188
rect 200 -83376 258 -83364
rect -258 -83624 -200 -83612
rect -258 -83800 -246 -83624
rect -212 -83800 -200 -83624
rect -258 -83812 -200 -83800
rect 200 -83624 258 -83612
rect 200 -83800 212 -83624
rect 246 -83800 258 -83624
rect 200 -83812 258 -83800
rect -258 -84060 -200 -84048
rect -258 -84236 -246 -84060
rect -212 -84236 -200 -84060
rect -258 -84248 -200 -84236
rect 200 -84060 258 -84048
rect 200 -84236 212 -84060
rect 246 -84236 258 -84060
rect 200 -84248 258 -84236
<< pdiffc >>
rect -246 84060 -212 84236
rect 212 84060 246 84236
rect -246 83624 -212 83800
rect 212 83624 246 83800
rect -246 83188 -212 83364
rect 212 83188 246 83364
rect -246 82752 -212 82928
rect 212 82752 246 82928
rect -246 82316 -212 82492
rect 212 82316 246 82492
rect -246 81880 -212 82056
rect 212 81880 246 82056
rect -246 81444 -212 81620
rect 212 81444 246 81620
rect -246 81008 -212 81184
rect 212 81008 246 81184
rect -246 80572 -212 80748
rect 212 80572 246 80748
rect -246 80136 -212 80312
rect 212 80136 246 80312
rect -246 79700 -212 79876
rect 212 79700 246 79876
rect -246 79264 -212 79440
rect 212 79264 246 79440
rect -246 78828 -212 79004
rect 212 78828 246 79004
rect -246 78392 -212 78568
rect 212 78392 246 78568
rect -246 77956 -212 78132
rect 212 77956 246 78132
rect -246 77520 -212 77696
rect 212 77520 246 77696
rect -246 77084 -212 77260
rect 212 77084 246 77260
rect -246 76648 -212 76824
rect 212 76648 246 76824
rect -246 76212 -212 76388
rect 212 76212 246 76388
rect -246 75776 -212 75952
rect 212 75776 246 75952
rect -246 75340 -212 75516
rect 212 75340 246 75516
rect -246 74904 -212 75080
rect 212 74904 246 75080
rect -246 74468 -212 74644
rect 212 74468 246 74644
rect -246 74032 -212 74208
rect 212 74032 246 74208
rect -246 73596 -212 73772
rect 212 73596 246 73772
rect -246 73160 -212 73336
rect 212 73160 246 73336
rect -246 72724 -212 72900
rect 212 72724 246 72900
rect -246 72288 -212 72464
rect 212 72288 246 72464
rect -246 71852 -212 72028
rect 212 71852 246 72028
rect -246 71416 -212 71592
rect 212 71416 246 71592
rect -246 70980 -212 71156
rect 212 70980 246 71156
rect -246 70544 -212 70720
rect 212 70544 246 70720
rect -246 70108 -212 70284
rect 212 70108 246 70284
rect -246 69672 -212 69848
rect 212 69672 246 69848
rect -246 69236 -212 69412
rect 212 69236 246 69412
rect -246 68800 -212 68976
rect 212 68800 246 68976
rect -246 68364 -212 68540
rect 212 68364 246 68540
rect -246 67928 -212 68104
rect 212 67928 246 68104
rect -246 67492 -212 67668
rect 212 67492 246 67668
rect -246 67056 -212 67232
rect 212 67056 246 67232
rect -246 66620 -212 66796
rect 212 66620 246 66796
rect -246 66184 -212 66360
rect 212 66184 246 66360
rect -246 65748 -212 65924
rect 212 65748 246 65924
rect -246 65312 -212 65488
rect 212 65312 246 65488
rect -246 64876 -212 65052
rect 212 64876 246 65052
rect -246 64440 -212 64616
rect 212 64440 246 64616
rect -246 64004 -212 64180
rect 212 64004 246 64180
rect -246 63568 -212 63744
rect 212 63568 246 63744
rect -246 63132 -212 63308
rect 212 63132 246 63308
rect -246 62696 -212 62872
rect 212 62696 246 62872
rect -246 62260 -212 62436
rect 212 62260 246 62436
rect -246 61824 -212 62000
rect 212 61824 246 62000
rect -246 61388 -212 61564
rect 212 61388 246 61564
rect -246 60952 -212 61128
rect 212 60952 246 61128
rect -246 60516 -212 60692
rect 212 60516 246 60692
rect -246 60080 -212 60256
rect 212 60080 246 60256
rect -246 59644 -212 59820
rect 212 59644 246 59820
rect -246 59208 -212 59384
rect 212 59208 246 59384
rect -246 58772 -212 58948
rect 212 58772 246 58948
rect -246 58336 -212 58512
rect 212 58336 246 58512
rect -246 57900 -212 58076
rect 212 57900 246 58076
rect -246 57464 -212 57640
rect 212 57464 246 57640
rect -246 57028 -212 57204
rect 212 57028 246 57204
rect -246 56592 -212 56768
rect 212 56592 246 56768
rect -246 56156 -212 56332
rect 212 56156 246 56332
rect -246 55720 -212 55896
rect 212 55720 246 55896
rect -246 55284 -212 55460
rect 212 55284 246 55460
rect -246 54848 -212 55024
rect 212 54848 246 55024
rect -246 54412 -212 54588
rect 212 54412 246 54588
rect -246 53976 -212 54152
rect 212 53976 246 54152
rect -246 53540 -212 53716
rect 212 53540 246 53716
rect -246 53104 -212 53280
rect 212 53104 246 53280
rect -246 52668 -212 52844
rect 212 52668 246 52844
rect -246 52232 -212 52408
rect 212 52232 246 52408
rect -246 51796 -212 51972
rect 212 51796 246 51972
rect -246 51360 -212 51536
rect 212 51360 246 51536
rect -246 50924 -212 51100
rect 212 50924 246 51100
rect -246 50488 -212 50664
rect 212 50488 246 50664
rect -246 50052 -212 50228
rect 212 50052 246 50228
rect -246 49616 -212 49792
rect 212 49616 246 49792
rect -246 49180 -212 49356
rect 212 49180 246 49356
rect -246 48744 -212 48920
rect 212 48744 246 48920
rect -246 48308 -212 48484
rect 212 48308 246 48484
rect -246 47872 -212 48048
rect 212 47872 246 48048
rect -246 47436 -212 47612
rect 212 47436 246 47612
rect -246 47000 -212 47176
rect 212 47000 246 47176
rect -246 46564 -212 46740
rect 212 46564 246 46740
rect -246 46128 -212 46304
rect 212 46128 246 46304
rect -246 45692 -212 45868
rect 212 45692 246 45868
rect -246 45256 -212 45432
rect 212 45256 246 45432
rect -246 44820 -212 44996
rect 212 44820 246 44996
rect -246 44384 -212 44560
rect 212 44384 246 44560
rect -246 43948 -212 44124
rect 212 43948 246 44124
rect -246 43512 -212 43688
rect 212 43512 246 43688
rect -246 43076 -212 43252
rect 212 43076 246 43252
rect -246 42640 -212 42816
rect 212 42640 246 42816
rect -246 42204 -212 42380
rect 212 42204 246 42380
rect -246 41768 -212 41944
rect 212 41768 246 41944
rect -246 41332 -212 41508
rect 212 41332 246 41508
rect -246 40896 -212 41072
rect 212 40896 246 41072
rect -246 40460 -212 40636
rect 212 40460 246 40636
rect -246 40024 -212 40200
rect 212 40024 246 40200
rect -246 39588 -212 39764
rect 212 39588 246 39764
rect -246 39152 -212 39328
rect 212 39152 246 39328
rect -246 38716 -212 38892
rect 212 38716 246 38892
rect -246 38280 -212 38456
rect 212 38280 246 38456
rect -246 37844 -212 38020
rect 212 37844 246 38020
rect -246 37408 -212 37584
rect 212 37408 246 37584
rect -246 36972 -212 37148
rect 212 36972 246 37148
rect -246 36536 -212 36712
rect 212 36536 246 36712
rect -246 36100 -212 36276
rect 212 36100 246 36276
rect -246 35664 -212 35840
rect 212 35664 246 35840
rect -246 35228 -212 35404
rect 212 35228 246 35404
rect -246 34792 -212 34968
rect 212 34792 246 34968
rect -246 34356 -212 34532
rect 212 34356 246 34532
rect -246 33920 -212 34096
rect 212 33920 246 34096
rect -246 33484 -212 33660
rect 212 33484 246 33660
rect -246 33048 -212 33224
rect 212 33048 246 33224
rect -246 32612 -212 32788
rect 212 32612 246 32788
rect -246 32176 -212 32352
rect 212 32176 246 32352
rect -246 31740 -212 31916
rect 212 31740 246 31916
rect -246 31304 -212 31480
rect 212 31304 246 31480
rect -246 30868 -212 31044
rect 212 30868 246 31044
rect -246 30432 -212 30608
rect 212 30432 246 30608
rect -246 29996 -212 30172
rect 212 29996 246 30172
rect -246 29560 -212 29736
rect 212 29560 246 29736
rect -246 29124 -212 29300
rect 212 29124 246 29300
rect -246 28688 -212 28864
rect 212 28688 246 28864
rect -246 28252 -212 28428
rect 212 28252 246 28428
rect -246 27816 -212 27992
rect 212 27816 246 27992
rect -246 27380 -212 27556
rect 212 27380 246 27556
rect -246 26944 -212 27120
rect 212 26944 246 27120
rect -246 26508 -212 26684
rect 212 26508 246 26684
rect -246 26072 -212 26248
rect 212 26072 246 26248
rect -246 25636 -212 25812
rect 212 25636 246 25812
rect -246 25200 -212 25376
rect 212 25200 246 25376
rect -246 24764 -212 24940
rect 212 24764 246 24940
rect -246 24328 -212 24504
rect 212 24328 246 24504
rect -246 23892 -212 24068
rect 212 23892 246 24068
rect -246 23456 -212 23632
rect 212 23456 246 23632
rect -246 23020 -212 23196
rect 212 23020 246 23196
rect -246 22584 -212 22760
rect 212 22584 246 22760
rect -246 22148 -212 22324
rect 212 22148 246 22324
rect -246 21712 -212 21888
rect 212 21712 246 21888
rect -246 21276 -212 21452
rect 212 21276 246 21452
rect -246 20840 -212 21016
rect 212 20840 246 21016
rect -246 20404 -212 20580
rect 212 20404 246 20580
rect -246 19968 -212 20144
rect 212 19968 246 20144
rect -246 19532 -212 19708
rect 212 19532 246 19708
rect -246 19096 -212 19272
rect 212 19096 246 19272
rect -246 18660 -212 18836
rect 212 18660 246 18836
rect -246 18224 -212 18400
rect 212 18224 246 18400
rect -246 17788 -212 17964
rect 212 17788 246 17964
rect -246 17352 -212 17528
rect 212 17352 246 17528
rect -246 16916 -212 17092
rect 212 16916 246 17092
rect -246 16480 -212 16656
rect 212 16480 246 16656
rect -246 16044 -212 16220
rect 212 16044 246 16220
rect -246 15608 -212 15784
rect 212 15608 246 15784
rect -246 15172 -212 15348
rect 212 15172 246 15348
rect -246 14736 -212 14912
rect 212 14736 246 14912
rect -246 14300 -212 14476
rect 212 14300 246 14476
rect -246 13864 -212 14040
rect 212 13864 246 14040
rect -246 13428 -212 13604
rect 212 13428 246 13604
rect -246 12992 -212 13168
rect 212 12992 246 13168
rect -246 12556 -212 12732
rect 212 12556 246 12732
rect -246 12120 -212 12296
rect 212 12120 246 12296
rect -246 11684 -212 11860
rect 212 11684 246 11860
rect -246 11248 -212 11424
rect 212 11248 246 11424
rect -246 10812 -212 10988
rect 212 10812 246 10988
rect -246 10376 -212 10552
rect 212 10376 246 10552
rect -246 9940 -212 10116
rect 212 9940 246 10116
rect -246 9504 -212 9680
rect 212 9504 246 9680
rect -246 9068 -212 9244
rect 212 9068 246 9244
rect -246 8632 -212 8808
rect 212 8632 246 8808
rect -246 8196 -212 8372
rect 212 8196 246 8372
rect -246 7760 -212 7936
rect 212 7760 246 7936
rect -246 7324 -212 7500
rect 212 7324 246 7500
rect -246 6888 -212 7064
rect 212 6888 246 7064
rect -246 6452 -212 6628
rect 212 6452 246 6628
rect -246 6016 -212 6192
rect 212 6016 246 6192
rect -246 5580 -212 5756
rect 212 5580 246 5756
rect -246 5144 -212 5320
rect 212 5144 246 5320
rect -246 4708 -212 4884
rect 212 4708 246 4884
rect -246 4272 -212 4448
rect 212 4272 246 4448
rect -246 3836 -212 4012
rect 212 3836 246 4012
rect -246 3400 -212 3576
rect 212 3400 246 3576
rect -246 2964 -212 3140
rect 212 2964 246 3140
rect -246 2528 -212 2704
rect 212 2528 246 2704
rect -246 2092 -212 2268
rect 212 2092 246 2268
rect -246 1656 -212 1832
rect 212 1656 246 1832
rect -246 1220 -212 1396
rect 212 1220 246 1396
rect -246 784 -212 960
rect 212 784 246 960
rect -246 348 -212 524
rect 212 348 246 524
rect -246 -88 -212 88
rect 212 -88 246 88
rect -246 -524 -212 -348
rect 212 -524 246 -348
rect -246 -960 -212 -784
rect 212 -960 246 -784
rect -246 -1396 -212 -1220
rect 212 -1396 246 -1220
rect -246 -1832 -212 -1656
rect 212 -1832 246 -1656
rect -246 -2268 -212 -2092
rect 212 -2268 246 -2092
rect -246 -2704 -212 -2528
rect 212 -2704 246 -2528
rect -246 -3140 -212 -2964
rect 212 -3140 246 -2964
rect -246 -3576 -212 -3400
rect 212 -3576 246 -3400
rect -246 -4012 -212 -3836
rect 212 -4012 246 -3836
rect -246 -4448 -212 -4272
rect 212 -4448 246 -4272
rect -246 -4884 -212 -4708
rect 212 -4884 246 -4708
rect -246 -5320 -212 -5144
rect 212 -5320 246 -5144
rect -246 -5756 -212 -5580
rect 212 -5756 246 -5580
rect -246 -6192 -212 -6016
rect 212 -6192 246 -6016
rect -246 -6628 -212 -6452
rect 212 -6628 246 -6452
rect -246 -7064 -212 -6888
rect 212 -7064 246 -6888
rect -246 -7500 -212 -7324
rect 212 -7500 246 -7324
rect -246 -7936 -212 -7760
rect 212 -7936 246 -7760
rect -246 -8372 -212 -8196
rect 212 -8372 246 -8196
rect -246 -8808 -212 -8632
rect 212 -8808 246 -8632
rect -246 -9244 -212 -9068
rect 212 -9244 246 -9068
rect -246 -9680 -212 -9504
rect 212 -9680 246 -9504
rect -246 -10116 -212 -9940
rect 212 -10116 246 -9940
rect -246 -10552 -212 -10376
rect 212 -10552 246 -10376
rect -246 -10988 -212 -10812
rect 212 -10988 246 -10812
rect -246 -11424 -212 -11248
rect 212 -11424 246 -11248
rect -246 -11860 -212 -11684
rect 212 -11860 246 -11684
rect -246 -12296 -212 -12120
rect 212 -12296 246 -12120
rect -246 -12732 -212 -12556
rect 212 -12732 246 -12556
rect -246 -13168 -212 -12992
rect 212 -13168 246 -12992
rect -246 -13604 -212 -13428
rect 212 -13604 246 -13428
rect -246 -14040 -212 -13864
rect 212 -14040 246 -13864
rect -246 -14476 -212 -14300
rect 212 -14476 246 -14300
rect -246 -14912 -212 -14736
rect 212 -14912 246 -14736
rect -246 -15348 -212 -15172
rect 212 -15348 246 -15172
rect -246 -15784 -212 -15608
rect 212 -15784 246 -15608
rect -246 -16220 -212 -16044
rect 212 -16220 246 -16044
rect -246 -16656 -212 -16480
rect 212 -16656 246 -16480
rect -246 -17092 -212 -16916
rect 212 -17092 246 -16916
rect -246 -17528 -212 -17352
rect 212 -17528 246 -17352
rect -246 -17964 -212 -17788
rect 212 -17964 246 -17788
rect -246 -18400 -212 -18224
rect 212 -18400 246 -18224
rect -246 -18836 -212 -18660
rect 212 -18836 246 -18660
rect -246 -19272 -212 -19096
rect 212 -19272 246 -19096
rect -246 -19708 -212 -19532
rect 212 -19708 246 -19532
rect -246 -20144 -212 -19968
rect 212 -20144 246 -19968
rect -246 -20580 -212 -20404
rect 212 -20580 246 -20404
rect -246 -21016 -212 -20840
rect 212 -21016 246 -20840
rect -246 -21452 -212 -21276
rect 212 -21452 246 -21276
rect -246 -21888 -212 -21712
rect 212 -21888 246 -21712
rect -246 -22324 -212 -22148
rect 212 -22324 246 -22148
rect -246 -22760 -212 -22584
rect 212 -22760 246 -22584
rect -246 -23196 -212 -23020
rect 212 -23196 246 -23020
rect -246 -23632 -212 -23456
rect 212 -23632 246 -23456
rect -246 -24068 -212 -23892
rect 212 -24068 246 -23892
rect -246 -24504 -212 -24328
rect 212 -24504 246 -24328
rect -246 -24940 -212 -24764
rect 212 -24940 246 -24764
rect -246 -25376 -212 -25200
rect 212 -25376 246 -25200
rect -246 -25812 -212 -25636
rect 212 -25812 246 -25636
rect -246 -26248 -212 -26072
rect 212 -26248 246 -26072
rect -246 -26684 -212 -26508
rect 212 -26684 246 -26508
rect -246 -27120 -212 -26944
rect 212 -27120 246 -26944
rect -246 -27556 -212 -27380
rect 212 -27556 246 -27380
rect -246 -27992 -212 -27816
rect 212 -27992 246 -27816
rect -246 -28428 -212 -28252
rect 212 -28428 246 -28252
rect -246 -28864 -212 -28688
rect 212 -28864 246 -28688
rect -246 -29300 -212 -29124
rect 212 -29300 246 -29124
rect -246 -29736 -212 -29560
rect 212 -29736 246 -29560
rect -246 -30172 -212 -29996
rect 212 -30172 246 -29996
rect -246 -30608 -212 -30432
rect 212 -30608 246 -30432
rect -246 -31044 -212 -30868
rect 212 -31044 246 -30868
rect -246 -31480 -212 -31304
rect 212 -31480 246 -31304
rect -246 -31916 -212 -31740
rect 212 -31916 246 -31740
rect -246 -32352 -212 -32176
rect 212 -32352 246 -32176
rect -246 -32788 -212 -32612
rect 212 -32788 246 -32612
rect -246 -33224 -212 -33048
rect 212 -33224 246 -33048
rect -246 -33660 -212 -33484
rect 212 -33660 246 -33484
rect -246 -34096 -212 -33920
rect 212 -34096 246 -33920
rect -246 -34532 -212 -34356
rect 212 -34532 246 -34356
rect -246 -34968 -212 -34792
rect 212 -34968 246 -34792
rect -246 -35404 -212 -35228
rect 212 -35404 246 -35228
rect -246 -35840 -212 -35664
rect 212 -35840 246 -35664
rect -246 -36276 -212 -36100
rect 212 -36276 246 -36100
rect -246 -36712 -212 -36536
rect 212 -36712 246 -36536
rect -246 -37148 -212 -36972
rect 212 -37148 246 -36972
rect -246 -37584 -212 -37408
rect 212 -37584 246 -37408
rect -246 -38020 -212 -37844
rect 212 -38020 246 -37844
rect -246 -38456 -212 -38280
rect 212 -38456 246 -38280
rect -246 -38892 -212 -38716
rect 212 -38892 246 -38716
rect -246 -39328 -212 -39152
rect 212 -39328 246 -39152
rect -246 -39764 -212 -39588
rect 212 -39764 246 -39588
rect -246 -40200 -212 -40024
rect 212 -40200 246 -40024
rect -246 -40636 -212 -40460
rect 212 -40636 246 -40460
rect -246 -41072 -212 -40896
rect 212 -41072 246 -40896
rect -246 -41508 -212 -41332
rect 212 -41508 246 -41332
rect -246 -41944 -212 -41768
rect 212 -41944 246 -41768
rect -246 -42380 -212 -42204
rect 212 -42380 246 -42204
rect -246 -42816 -212 -42640
rect 212 -42816 246 -42640
rect -246 -43252 -212 -43076
rect 212 -43252 246 -43076
rect -246 -43688 -212 -43512
rect 212 -43688 246 -43512
rect -246 -44124 -212 -43948
rect 212 -44124 246 -43948
rect -246 -44560 -212 -44384
rect 212 -44560 246 -44384
rect -246 -44996 -212 -44820
rect 212 -44996 246 -44820
rect -246 -45432 -212 -45256
rect 212 -45432 246 -45256
rect -246 -45868 -212 -45692
rect 212 -45868 246 -45692
rect -246 -46304 -212 -46128
rect 212 -46304 246 -46128
rect -246 -46740 -212 -46564
rect 212 -46740 246 -46564
rect -246 -47176 -212 -47000
rect 212 -47176 246 -47000
rect -246 -47612 -212 -47436
rect 212 -47612 246 -47436
rect -246 -48048 -212 -47872
rect 212 -48048 246 -47872
rect -246 -48484 -212 -48308
rect 212 -48484 246 -48308
rect -246 -48920 -212 -48744
rect 212 -48920 246 -48744
rect -246 -49356 -212 -49180
rect 212 -49356 246 -49180
rect -246 -49792 -212 -49616
rect 212 -49792 246 -49616
rect -246 -50228 -212 -50052
rect 212 -50228 246 -50052
rect -246 -50664 -212 -50488
rect 212 -50664 246 -50488
rect -246 -51100 -212 -50924
rect 212 -51100 246 -50924
rect -246 -51536 -212 -51360
rect 212 -51536 246 -51360
rect -246 -51972 -212 -51796
rect 212 -51972 246 -51796
rect -246 -52408 -212 -52232
rect 212 -52408 246 -52232
rect -246 -52844 -212 -52668
rect 212 -52844 246 -52668
rect -246 -53280 -212 -53104
rect 212 -53280 246 -53104
rect -246 -53716 -212 -53540
rect 212 -53716 246 -53540
rect -246 -54152 -212 -53976
rect 212 -54152 246 -53976
rect -246 -54588 -212 -54412
rect 212 -54588 246 -54412
rect -246 -55024 -212 -54848
rect 212 -55024 246 -54848
rect -246 -55460 -212 -55284
rect 212 -55460 246 -55284
rect -246 -55896 -212 -55720
rect 212 -55896 246 -55720
rect -246 -56332 -212 -56156
rect 212 -56332 246 -56156
rect -246 -56768 -212 -56592
rect 212 -56768 246 -56592
rect -246 -57204 -212 -57028
rect 212 -57204 246 -57028
rect -246 -57640 -212 -57464
rect 212 -57640 246 -57464
rect -246 -58076 -212 -57900
rect 212 -58076 246 -57900
rect -246 -58512 -212 -58336
rect 212 -58512 246 -58336
rect -246 -58948 -212 -58772
rect 212 -58948 246 -58772
rect -246 -59384 -212 -59208
rect 212 -59384 246 -59208
rect -246 -59820 -212 -59644
rect 212 -59820 246 -59644
rect -246 -60256 -212 -60080
rect 212 -60256 246 -60080
rect -246 -60692 -212 -60516
rect 212 -60692 246 -60516
rect -246 -61128 -212 -60952
rect 212 -61128 246 -60952
rect -246 -61564 -212 -61388
rect 212 -61564 246 -61388
rect -246 -62000 -212 -61824
rect 212 -62000 246 -61824
rect -246 -62436 -212 -62260
rect 212 -62436 246 -62260
rect -246 -62872 -212 -62696
rect 212 -62872 246 -62696
rect -246 -63308 -212 -63132
rect 212 -63308 246 -63132
rect -246 -63744 -212 -63568
rect 212 -63744 246 -63568
rect -246 -64180 -212 -64004
rect 212 -64180 246 -64004
rect -246 -64616 -212 -64440
rect 212 -64616 246 -64440
rect -246 -65052 -212 -64876
rect 212 -65052 246 -64876
rect -246 -65488 -212 -65312
rect 212 -65488 246 -65312
rect -246 -65924 -212 -65748
rect 212 -65924 246 -65748
rect -246 -66360 -212 -66184
rect 212 -66360 246 -66184
rect -246 -66796 -212 -66620
rect 212 -66796 246 -66620
rect -246 -67232 -212 -67056
rect 212 -67232 246 -67056
rect -246 -67668 -212 -67492
rect 212 -67668 246 -67492
rect -246 -68104 -212 -67928
rect 212 -68104 246 -67928
rect -246 -68540 -212 -68364
rect 212 -68540 246 -68364
rect -246 -68976 -212 -68800
rect 212 -68976 246 -68800
rect -246 -69412 -212 -69236
rect 212 -69412 246 -69236
rect -246 -69848 -212 -69672
rect 212 -69848 246 -69672
rect -246 -70284 -212 -70108
rect 212 -70284 246 -70108
rect -246 -70720 -212 -70544
rect 212 -70720 246 -70544
rect -246 -71156 -212 -70980
rect 212 -71156 246 -70980
rect -246 -71592 -212 -71416
rect 212 -71592 246 -71416
rect -246 -72028 -212 -71852
rect 212 -72028 246 -71852
rect -246 -72464 -212 -72288
rect 212 -72464 246 -72288
rect -246 -72900 -212 -72724
rect 212 -72900 246 -72724
rect -246 -73336 -212 -73160
rect 212 -73336 246 -73160
rect -246 -73772 -212 -73596
rect 212 -73772 246 -73596
rect -246 -74208 -212 -74032
rect 212 -74208 246 -74032
rect -246 -74644 -212 -74468
rect 212 -74644 246 -74468
rect -246 -75080 -212 -74904
rect 212 -75080 246 -74904
rect -246 -75516 -212 -75340
rect 212 -75516 246 -75340
rect -246 -75952 -212 -75776
rect 212 -75952 246 -75776
rect -246 -76388 -212 -76212
rect 212 -76388 246 -76212
rect -246 -76824 -212 -76648
rect 212 -76824 246 -76648
rect -246 -77260 -212 -77084
rect 212 -77260 246 -77084
rect -246 -77696 -212 -77520
rect 212 -77696 246 -77520
rect -246 -78132 -212 -77956
rect 212 -78132 246 -77956
rect -246 -78568 -212 -78392
rect 212 -78568 246 -78392
rect -246 -79004 -212 -78828
rect 212 -79004 246 -78828
rect -246 -79440 -212 -79264
rect 212 -79440 246 -79264
rect -246 -79876 -212 -79700
rect 212 -79876 246 -79700
rect -246 -80312 -212 -80136
rect 212 -80312 246 -80136
rect -246 -80748 -212 -80572
rect 212 -80748 246 -80572
rect -246 -81184 -212 -81008
rect 212 -81184 246 -81008
rect -246 -81620 -212 -81444
rect 212 -81620 246 -81444
rect -246 -82056 -212 -81880
rect 212 -82056 246 -81880
rect -246 -82492 -212 -82316
rect 212 -82492 246 -82316
rect -246 -82928 -212 -82752
rect 212 -82928 246 -82752
rect -246 -83364 -212 -83188
rect 212 -83364 246 -83188
rect -246 -83800 -212 -83624
rect 212 -83800 246 -83624
rect -246 -84236 -212 -84060
rect 212 -84236 246 -84060
<< nsubdiff >>
rect -360 84397 -264 84431
rect 264 84397 360 84431
rect -360 84335 -326 84397
rect 326 84335 360 84397
rect -360 -84397 -326 -84335
rect 326 -84397 360 -84335
rect -360 -84431 -264 -84397
rect 264 -84431 360 -84397
<< nsubdiffcont >>
rect -264 84397 264 84431
rect -360 -84335 -326 84335
rect 326 -84335 360 84335
rect -264 -84431 264 -84397
<< poly >>
rect -200 84329 200 84345
rect -200 84295 -184 84329
rect 184 84295 200 84329
rect -200 84248 200 84295
rect -200 84001 200 84048
rect -200 83967 -184 84001
rect 184 83967 200 84001
rect -200 83951 200 83967
rect -200 83893 200 83909
rect -200 83859 -184 83893
rect 184 83859 200 83893
rect -200 83812 200 83859
rect -200 83565 200 83612
rect -200 83531 -184 83565
rect 184 83531 200 83565
rect -200 83515 200 83531
rect -200 83457 200 83473
rect -200 83423 -184 83457
rect 184 83423 200 83457
rect -200 83376 200 83423
rect -200 83129 200 83176
rect -200 83095 -184 83129
rect 184 83095 200 83129
rect -200 83079 200 83095
rect -200 83021 200 83037
rect -200 82987 -184 83021
rect 184 82987 200 83021
rect -200 82940 200 82987
rect -200 82693 200 82740
rect -200 82659 -184 82693
rect 184 82659 200 82693
rect -200 82643 200 82659
rect -200 82585 200 82601
rect -200 82551 -184 82585
rect 184 82551 200 82585
rect -200 82504 200 82551
rect -200 82257 200 82304
rect -200 82223 -184 82257
rect 184 82223 200 82257
rect -200 82207 200 82223
rect -200 82149 200 82165
rect -200 82115 -184 82149
rect 184 82115 200 82149
rect -200 82068 200 82115
rect -200 81821 200 81868
rect -200 81787 -184 81821
rect 184 81787 200 81821
rect -200 81771 200 81787
rect -200 81713 200 81729
rect -200 81679 -184 81713
rect 184 81679 200 81713
rect -200 81632 200 81679
rect -200 81385 200 81432
rect -200 81351 -184 81385
rect 184 81351 200 81385
rect -200 81335 200 81351
rect -200 81277 200 81293
rect -200 81243 -184 81277
rect 184 81243 200 81277
rect -200 81196 200 81243
rect -200 80949 200 80996
rect -200 80915 -184 80949
rect 184 80915 200 80949
rect -200 80899 200 80915
rect -200 80841 200 80857
rect -200 80807 -184 80841
rect 184 80807 200 80841
rect -200 80760 200 80807
rect -200 80513 200 80560
rect -200 80479 -184 80513
rect 184 80479 200 80513
rect -200 80463 200 80479
rect -200 80405 200 80421
rect -200 80371 -184 80405
rect 184 80371 200 80405
rect -200 80324 200 80371
rect -200 80077 200 80124
rect -200 80043 -184 80077
rect 184 80043 200 80077
rect -200 80027 200 80043
rect -200 79969 200 79985
rect -200 79935 -184 79969
rect 184 79935 200 79969
rect -200 79888 200 79935
rect -200 79641 200 79688
rect -200 79607 -184 79641
rect 184 79607 200 79641
rect -200 79591 200 79607
rect -200 79533 200 79549
rect -200 79499 -184 79533
rect 184 79499 200 79533
rect -200 79452 200 79499
rect -200 79205 200 79252
rect -200 79171 -184 79205
rect 184 79171 200 79205
rect -200 79155 200 79171
rect -200 79097 200 79113
rect -200 79063 -184 79097
rect 184 79063 200 79097
rect -200 79016 200 79063
rect -200 78769 200 78816
rect -200 78735 -184 78769
rect 184 78735 200 78769
rect -200 78719 200 78735
rect -200 78661 200 78677
rect -200 78627 -184 78661
rect 184 78627 200 78661
rect -200 78580 200 78627
rect -200 78333 200 78380
rect -200 78299 -184 78333
rect 184 78299 200 78333
rect -200 78283 200 78299
rect -200 78225 200 78241
rect -200 78191 -184 78225
rect 184 78191 200 78225
rect -200 78144 200 78191
rect -200 77897 200 77944
rect -200 77863 -184 77897
rect 184 77863 200 77897
rect -200 77847 200 77863
rect -200 77789 200 77805
rect -200 77755 -184 77789
rect 184 77755 200 77789
rect -200 77708 200 77755
rect -200 77461 200 77508
rect -200 77427 -184 77461
rect 184 77427 200 77461
rect -200 77411 200 77427
rect -200 77353 200 77369
rect -200 77319 -184 77353
rect 184 77319 200 77353
rect -200 77272 200 77319
rect -200 77025 200 77072
rect -200 76991 -184 77025
rect 184 76991 200 77025
rect -200 76975 200 76991
rect -200 76917 200 76933
rect -200 76883 -184 76917
rect 184 76883 200 76917
rect -200 76836 200 76883
rect -200 76589 200 76636
rect -200 76555 -184 76589
rect 184 76555 200 76589
rect -200 76539 200 76555
rect -200 76481 200 76497
rect -200 76447 -184 76481
rect 184 76447 200 76481
rect -200 76400 200 76447
rect -200 76153 200 76200
rect -200 76119 -184 76153
rect 184 76119 200 76153
rect -200 76103 200 76119
rect -200 76045 200 76061
rect -200 76011 -184 76045
rect 184 76011 200 76045
rect -200 75964 200 76011
rect -200 75717 200 75764
rect -200 75683 -184 75717
rect 184 75683 200 75717
rect -200 75667 200 75683
rect -200 75609 200 75625
rect -200 75575 -184 75609
rect 184 75575 200 75609
rect -200 75528 200 75575
rect -200 75281 200 75328
rect -200 75247 -184 75281
rect 184 75247 200 75281
rect -200 75231 200 75247
rect -200 75173 200 75189
rect -200 75139 -184 75173
rect 184 75139 200 75173
rect -200 75092 200 75139
rect -200 74845 200 74892
rect -200 74811 -184 74845
rect 184 74811 200 74845
rect -200 74795 200 74811
rect -200 74737 200 74753
rect -200 74703 -184 74737
rect 184 74703 200 74737
rect -200 74656 200 74703
rect -200 74409 200 74456
rect -200 74375 -184 74409
rect 184 74375 200 74409
rect -200 74359 200 74375
rect -200 74301 200 74317
rect -200 74267 -184 74301
rect 184 74267 200 74301
rect -200 74220 200 74267
rect -200 73973 200 74020
rect -200 73939 -184 73973
rect 184 73939 200 73973
rect -200 73923 200 73939
rect -200 73865 200 73881
rect -200 73831 -184 73865
rect 184 73831 200 73865
rect -200 73784 200 73831
rect -200 73537 200 73584
rect -200 73503 -184 73537
rect 184 73503 200 73537
rect -200 73487 200 73503
rect -200 73429 200 73445
rect -200 73395 -184 73429
rect 184 73395 200 73429
rect -200 73348 200 73395
rect -200 73101 200 73148
rect -200 73067 -184 73101
rect 184 73067 200 73101
rect -200 73051 200 73067
rect -200 72993 200 73009
rect -200 72959 -184 72993
rect 184 72959 200 72993
rect -200 72912 200 72959
rect -200 72665 200 72712
rect -200 72631 -184 72665
rect 184 72631 200 72665
rect -200 72615 200 72631
rect -200 72557 200 72573
rect -200 72523 -184 72557
rect 184 72523 200 72557
rect -200 72476 200 72523
rect -200 72229 200 72276
rect -200 72195 -184 72229
rect 184 72195 200 72229
rect -200 72179 200 72195
rect -200 72121 200 72137
rect -200 72087 -184 72121
rect 184 72087 200 72121
rect -200 72040 200 72087
rect -200 71793 200 71840
rect -200 71759 -184 71793
rect 184 71759 200 71793
rect -200 71743 200 71759
rect -200 71685 200 71701
rect -200 71651 -184 71685
rect 184 71651 200 71685
rect -200 71604 200 71651
rect -200 71357 200 71404
rect -200 71323 -184 71357
rect 184 71323 200 71357
rect -200 71307 200 71323
rect -200 71249 200 71265
rect -200 71215 -184 71249
rect 184 71215 200 71249
rect -200 71168 200 71215
rect -200 70921 200 70968
rect -200 70887 -184 70921
rect 184 70887 200 70921
rect -200 70871 200 70887
rect -200 70813 200 70829
rect -200 70779 -184 70813
rect 184 70779 200 70813
rect -200 70732 200 70779
rect -200 70485 200 70532
rect -200 70451 -184 70485
rect 184 70451 200 70485
rect -200 70435 200 70451
rect -200 70377 200 70393
rect -200 70343 -184 70377
rect 184 70343 200 70377
rect -200 70296 200 70343
rect -200 70049 200 70096
rect -200 70015 -184 70049
rect 184 70015 200 70049
rect -200 69999 200 70015
rect -200 69941 200 69957
rect -200 69907 -184 69941
rect 184 69907 200 69941
rect -200 69860 200 69907
rect -200 69613 200 69660
rect -200 69579 -184 69613
rect 184 69579 200 69613
rect -200 69563 200 69579
rect -200 69505 200 69521
rect -200 69471 -184 69505
rect 184 69471 200 69505
rect -200 69424 200 69471
rect -200 69177 200 69224
rect -200 69143 -184 69177
rect 184 69143 200 69177
rect -200 69127 200 69143
rect -200 69069 200 69085
rect -200 69035 -184 69069
rect 184 69035 200 69069
rect -200 68988 200 69035
rect -200 68741 200 68788
rect -200 68707 -184 68741
rect 184 68707 200 68741
rect -200 68691 200 68707
rect -200 68633 200 68649
rect -200 68599 -184 68633
rect 184 68599 200 68633
rect -200 68552 200 68599
rect -200 68305 200 68352
rect -200 68271 -184 68305
rect 184 68271 200 68305
rect -200 68255 200 68271
rect -200 68197 200 68213
rect -200 68163 -184 68197
rect 184 68163 200 68197
rect -200 68116 200 68163
rect -200 67869 200 67916
rect -200 67835 -184 67869
rect 184 67835 200 67869
rect -200 67819 200 67835
rect -200 67761 200 67777
rect -200 67727 -184 67761
rect 184 67727 200 67761
rect -200 67680 200 67727
rect -200 67433 200 67480
rect -200 67399 -184 67433
rect 184 67399 200 67433
rect -200 67383 200 67399
rect -200 67325 200 67341
rect -200 67291 -184 67325
rect 184 67291 200 67325
rect -200 67244 200 67291
rect -200 66997 200 67044
rect -200 66963 -184 66997
rect 184 66963 200 66997
rect -200 66947 200 66963
rect -200 66889 200 66905
rect -200 66855 -184 66889
rect 184 66855 200 66889
rect -200 66808 200 66855
rect -200 66561 200 66608
rect -200 66527 -184 66561
rect 184 66527 200 66561
rect -200 66511 200 66527
rect -200 66453 200 66469
rect -200 66419 -184 66453
rect 184 66419 200 66453
rect -200 66372 200 66419
rect -200 66125 200 66172
rect -200 66091 -184 66125
rect 184 66091 200 66125
rect -200 66075 200 66091
rect -200 66017 200 66033
rect -200 65983 -184 66017
rect 184 65983 200 66017
rect -200 65936 200 65983
rect -200 65689 200 65736
rect -200 65655 -184 65689
rect 184 65655 200 65689
rect -200 65639 200 65655
rect -200 65581 200 65597
rect -200 65547 -184 65581
rect 184 65547 200 65581
rect -200 65500 200 65547
rect -200 65253 200 65300
rect -200 65219 -184 65253
rect 184 65219 200 65253
rect -200 65203 200 65219
rect -200 65145 200 65161
rect -200 65111 -184 65145
rect 184 65111 200 65145
rect -200 65064 200 65111
rect -200 64817 200 64864
rect -200 64783 -184 64817
rect 184 64783 200 64817
rect -200 64767 200 64783
rect -200 64709 200 64725
rect -200 64675 -184 64709
rect 184 64675 200 64709
rect -200 64628 200 64675
rect -200 64381 200 64428
rect -200 64347 -184 64381
rect 184 64347 200 64381
rect -200 64331 200 64347
rect -200 64273 200 64289
rect -200 64239 -184 64273
rect 184 64239 200 64273
rect -200 64192 200 64239
rect -200 63945 200 63992
rect -200 63911 -184 63945
rect 184 63911 200 63945
rect -200 63895 200 63911
rect -200 63837 200 63853
rect -200 63803 -184 63837
rect 184 63803 200 63837
rect -200 63756 200 63803
rect -200 63509 200 63556
rect -200 63475 -184 63509
rect 184 63475 200 63509
rect -200 63459 200 63475
rect -200 63401 200 63417
rect -200 63367 -184 63401
rect 184 63367 200 63401
rect -200 63320 200 63367
rect -200 63073 200 63120
rect -200 63039 -184 63073
rect 184 63039 200 63073
rect -200 63023 200 63039
rect -200 62965 200 62981
rect -200 62931 -184 62965
rect 184 62931 200 62965
rect -200 62884 200 62931
rect -200 62637 200 62684
rect -200 62603 -184 62637
rect 184 62603 200 62637
rect -200 62587 200 62603
rect -200 62529 200 62545
rect -200 62495 -184 62529
rect 184 62495 200 62529
rect -200 62448 200 62495
rect -200 62201 200 62248
rect -200 62167 -184 62201
rect 184 62167 200 62201
rect -200 62151 200 62167
rect -200 62093 200 62109
rect -200 62059 -184 62093
rect 184 62059 200 62093
rect -200 62012 200 62059
rect -200 61765 200 61812
rect -200 61731 -184 61765
rect 184 61731 200 61765
rect -200 61715 200 61731
rect -200 61657 200 61673
rect -200 61623 -184 61657
rect 184 61623 200 61657
rect -200 61576 200 61623
rect -200 61329 200 61376
rect -200 61295 -184 61329
rect 184 61295 200 61329
rect -200 61279 200 61295
rect -200 61221 200 61237
rect -200 61187 -184 61221
rect 184 61187 200 61221
rect -200 61140 200 61187
rect -200 60893 200 60940
rect -200 60859 -184 60893
rect 184 60859 200 60893
rect -200 60843 200 60859
rect -200 60785 200 60801
rect -200 60751 -184 60785
rect 184 60751 200 60785
rect -200 60704 200 60751
rect -200 60457 200 60504
rect -200 60423 -184 60457
rect 184 60423 200 60457
rect -200 60407 200 60423
rect -200 60349 200 60365
rect -200 60315 -184 60349
rect 184 60315 200 60349
rect -200 60268 200 60315
rect -200 60021 200 60068
rect -200 59987 -184 60021
rect 184 59987 200 60021
rect -200 59971 200 59987
rect -200 59913 200 59929
rect -200 59879 -184 59913
rect 184 59879 200 59913
rect -200 59832 200 59879
rect -200 59585 200 59632
rect -200 59551 -184 59585
rect 184 59551 200 59585
rect -200 59535 200 59551
rect -200 59477 200 59493
rect -200 59443 -184 59477
rect 184 59443 200 59477
rect -200 59396 200 59443
rect -200 59149 200 59196
rect -200 59115 -184 59149
rect 184 59115 200 59149
rect -200 59099 200 59115
rect -200 59041 200 59057
rect -200 59007 -184 59041
rect 184 59007 200 59041
rect -200 58960 200 59007
rect -200 58713 200 58760
rect -200 58679 -184 58713
rect 184 58679 200 58713
rect -200 58663 200 58679
rect -200 58605 200 58621
rect -200 58571 -184 58605
rect 184 58571 200 58605
rect -200 58524 200 58571
rect -200 58277 200 58324
rect -200 58243 -184 58277
rect 184 58243 200 58277
rect -200 58227 200 58243
rect -200 58169 200 58185
rect -200 58135 -184 58169
rect 184 58135 200 58169
rect -200 58088 200 58135
rect -200 57841 200 57888
rect -200 57807 -184 57841
rect 184 57807 200 57841
rect -200 57791 200 57807
rect -200 57733 200 57749
rect -200 57699 -184 57733
rect 184 57699 200 57733
rect -200 57652 200 57699
rect -200 57405 200 57452
rect -200 57371 -184 57405
rect 184 57371 200 57405
rect -200 57355 200 57371
rect -200 57297 200 57313
rect -200 57263 -184 57297
rect 184 57263 200 57297
rect -200 57216 200 57263
rect -200 56969 200 57016
rect -200 56935 -184 56969
rect 184 56935 200 56969
rect -200 56919 200 56935
rect -200 56861 200 56877
rect -200 56827 -184 56861
rect 184 56827 200 56861
rect -200 56780 200 56827
rect -200 56533 200 56580
rect -200 56499 -184 56533
rect 184 56499 200 56533
rect -200 56483 200 56499
rect -200 56425 200 56441
rect -200 56391 -184 56425
rect 184 56391 200 56425
rect -200 56344 200 56391
rect -200 56097 200 56144
rect -200 56063 -184 56097
rect 184 56063 200 56097
rect -200 56047 200 56063
rect -200 55989 200 56005
rect -200 55955 -184 55989
rect 184 55955 200 55989
rect -200 55908 200 55955
rect -200 55661 200 55708
rect -200 55627 -184 55661
rect 184 55627 200 55661
rect -200 55611 200 55627
rect -200 55553 200 55569
rect -200 55519 -184 55553
rect 184 55519 200 55553
rect -200 55472 200 55519
rect -200 55225 200 55272
rect -200 55191 -184 55225
rect 184 55191 200 55225
rect -200 55175 200 55191
rect -200 55117 200 55133
rect -200 55083 -184 55117
rect 184 55083 200 55117
rect -200 55036 200 55083
rect -200 54789 200 54836
rect -200 54755 -184 54789
rect 184 54755 200 54789
rect -200 54739 200 54755
rect -200 54681 200 54697
rect -200 54647 -184 54681
rect 184 54647 200 54681
rect -200 54600 200 54647
rect -200 54353 200 54400
rect -200 54319 -184 54353
rect 184 54319 200 54353
rect -200 54303 200 54319
rect -200 54245 200 54261
rect -200 54211 -184 54245
rect 184 54211 200 54245
rect -200 54164 200 54211
rect -200 53917 200 53964
rect -200 53883 -184 53917
rect 184 53883 200 53917
rect -200 53867 200 53883
rect -200 53809 200 53825
rect -200 53775 -184 53809
rect 184 53775 200 53809
rect -200 53728 200 53775
rect -200 53481 200 53528
rect -200 53447 -184 53481
rect 184 53447 200 53481
rect -200 53431 200 53447
rect -200 53373 200 53389
rect -200 53339 -184 53373
rect 184 53339 200 53373
rect -200 53292 200 53339
rect -200 53045 200 53092
rect -200 53011 -184 53045
rect 184 53011 200 53045
rect -200 52995 200 53011
rect -200 52937 200 52953
rect -200 52903 -184 52937
rect 184 52903 200 52937
rect -200 52856 200 52903
rect -200 52609 200 52656
rect -200 52575 -184 52609
rect 184 52575 200 52609
rect -200 52559 200 52575
rect -200 52501 200 52517
rect -200 52467 -184 52501
rect 184 52467 200 52501
rect -200 52420 200 52467
rect -200 52173 200 52220
rect -200 52139 -184 52173
rect 184 52139 200 52173
rect -200 52123 200 52139
rect -200 52065 200 52081
rect -200 52031 -184 52065
rect 184 52031 200 52065
rect -200 51984 200 52031
rect -200 51737 200 51784
rect -200 51703 -184 51737
rect 184 51703 200 51737
rect -200 51687 200 51703
rect -200 51629 200 51645
rect -200 51595 -184 51629
rect 184 51595 200 51629
rect -200 51548 200 51595
rect -200 51301 200 51348
rect -200 51267 -184 51301
rect 184 51267 200 51301
rect -200 51251 200 51267
rect -200 51193 200 51209
rect -200 51159 -184 51193
rect 184 51159 200 51193
rect -200 51112 200 51159
rect -200 50865 200 50912
rect -200 50831 -184 50865
rect 184 50831 200 50865
rect -200 50815 200 50831
rect -200 50757 200 50773
rect -200 50723 -184 50757
rect 184 50723 200 50757
rect -200 50676 200 50723
rect -200 50429 200 50476
rect -200 50395 -184 50429
rect 184 50395 200 50429
rect -200 50379 200 50395
rect -200 50321 200 50337
rect -200 50287 -184 50321
rect 184 50287 200 50321
rect -200 50240 200 50287
rect -200 49993 200 50040
rect -200 49959 -184 49993
rect 184 49959 200 49993
rect -200 49943 200 49959
rect -200 49885 200 49901
rect -200 49851 -184 49885
rect 184 49851 200 49885
rect -200 49804 200 49851
rect -200 49557 200 49604
rect -200 49523 -184 49557
rect 184 49523 200 49557
rect -200 49507 200 49523
rect -200 49449 200 49465
rect -200 49415 -184 49449
rect 184 49415 200 49449
rect -200 49368 200 49415
rect -200 49121 200 49168
rect -200 49087 -184 49121
rect 184 49087 200 49121
rect -200 49071 200 49087
rect -200 49013 200 49029
rect -200 48979 -184 49013
rect 184 48979 200 49013
rect -200 48932 200 48979
rect -200 48685 200 48732
rect -200 48651 -184 48685
rect 184 48651 200 48685
rect -200 48635 200 48651
rect -200 48577 200 48593
rect -200 48543 -184 48577
rect 184 48543 200 48577
rect -200 48496 200 48543
rect -200 48249 200 48296
rect -200 48215 -184 48249
rect 184 48215 200 48249
rect -200 48199 200 48215
rect -200 48141 200 48157
rect -200 48107 -184 48141
rect 184 48107 200 48141
rect -200 48060 200 48107
rect -200 47813 200 47860
rect -200 47779 -184 47813
rect 184 47779 200 47813
rect -200 47763 200 47779
rect -200 47705 200 47721
rect -200 47671 -184 47705
rect 184 47671 200 47705
rect -200 47624 200 47671
rect -200 47377 200 47424
rect -200 47343 -184 47377
rect 184 47343 200 47377
rect -200 47327 200 47343
rect -200 47269 200 47285
rect -200 47235 -184 47269
rect 184 47235 200 47269
rect -200 47188 200 47235
rect -200 46941 200 46988
rect -200 46907 -184 46941
rect 184 46907 200 46941
rect -200 46891 200 46907
rect -200 46833 200 46849
rect -200 46799 -184 46833
rect 184 46799 200 46833
rect -200 46752 200 46799
rect -200 46505 200 46552
rect -200 46471 -184 46505
rect 184 46471 200 46505
rect -200 46455 200 46471
rect -200 46397 200 46413
rect -200 46363 -184 46397
rect 184 46363 200 46397
rect -200 46316 200 46363
rect -200 46069 200 46116
rect -200 46035 -184 46069
rect 184 46035 200 46069
rect -200 46019 200 46035
rect -200 45961 200 45977
rect -200 45927 -184 45961
rect 184 45927 200 45961
rect -200 45880 200 45927
rect -200 45633 200 45680
rect -200 45599 -184 45633
rect 184 45599 200 45633
rect -200 45583 200 45599
rect -200 45525 200 45541
rect -200 45491 -184 45525
rect 184 45491 200 45525
rect -200 45444 200 45491
rect -200 45197 200 45244
rect -200 45163 -184 45197
rect 184 45163 200 45197
rect -200 45147 200 45163
rect -200 45089 200 45105
rect -200 45055 -184 45089
rect 184 45055 200 45089
rect -200 45008 200 45055
rect -200 44761 200 44808
rect -200 44727 -184 44761
rect 184 44727 200 44761
rect -200 44711 200 44727
rect -200 44653 200 44669
rect -200 44619 -184 44653
rect 184 44619 200 44653
rect -200 44572 200 44619
rect -200 44325 200 44372
rect -200 44291 -184 44325
rect 184 44291 200 44325
rect -200 44275 200 44291
rect -200 44217 200 44233
rect -200 44183 -184 44217
rect 184 44183 200 44217
rect -200 44136 200 44183
rect -200 43889 200 43936
rect -200 43855 -184 43889
rect 184 43855 200 43889
rect -200 43839 200 43855
rect -200 43781 200 43797
rect -200 43747 -184 43781
rect 184 43747 200 43781
rect -200 43700 200 43747
rect -200 43453 200 43500
rect -200 43419 -184 43453
rect 184 43419 200 43453
rect -200 43403 200 43419
rect -200 43345 200 43361
rect -200 43311 -184 43345
rect 184 43311 200 43345
rect -200 43264 200 43311
rect -200 43017 200 43064
rect -200 42983 -184 43017
rect 184 42983 200 43017
rect -200 42967 200 42983
rect -200 42909 200 42925
rect -200 42875 -184 42909
rect 184 42875 200 42909
rect -200 42828 200 42875
rect -200 42581 200 42628
rect -200 42547 -184 42581
rect 184 42547 200 42581
rect -200 42531 200 42547
rect -200 42473 200 42489
rect -200 42439 -184 42473
rect 184 42439 200 42473
rect -200 42392 200 42439
rect -200 42145 200 42192
rect -200 42111 -184 42145
rect 184 42111 200 42145
rect -200 42095 200 42111
rect -200 42037 200 42053
rect -200 42003 -184 42037
rect 184 42003 200 42037
rect -200 41956 200 42003
rect -200 41709 200 41756
rect -200 41675 -184 41709
rect 184 41675 200 41709
rect -200 41659 200 41675
rect -200 41601 200 41617
rect -200 41567 -184 41601
rect 184 41567 200 41601
rect -200 41520 200 41567
rect -200 41273 200 41320
rect -200 41239 -184 41273
rect 184 41239 200 41273
rect -200 41223 200 41239
rect -200 41165 200 41181
rect -200 41131 -184 41165
rect 184 41131 200 41165
rect -200 41084 200 41131
rect -200 40837 200 40884
rect -200 40803 -184 40837
rect 184 40803 200 40837
rect -200 40787 200 40803
rect -200 40729 200 40745
rect -200 40695 -184 40729
rect 184 40695 200 40729
rect -200 40648 200 40695
rect -200 40401 200 40448
rect -200 40367 -184 40401
rect 184 40367 200 40401
rect -200 40351 200 40367
rect -200 40293 200 40309
rect -200 40259 -184 40293
rect 184 40259 200 40293
rect -200 40212 200 40259
rect -200 39965 200 40012
rect -200 39931 -184 39965
rect 184 39931 200 39965
rect -200 39915 200 39931
rect -200 39857 200 39873
rect -200 39823 -184 39857
rect 184 39823 200 39857
rect -200 39776 200 39823
rect -200 39529 200 39576
rect -200 39495 -184 39529
rect 184 39495 200 39529
rect -200 39479 200 39495
rect -200 39421 200 39437
rect -200 39387 -184 39421
rect 184 39387 200 39421
rect -200 39340 200 39387
rect -200 39093 200 39140
rect -200 39059 -184 39093
rect 184 39059 200 39093
rect -200 39043 200 39059
rect -200 38985 200 39001
rect -200 38951 -184 38985
rect 184 38951 200 38985
rect -200 38904 200 38951
rect -200 38657 200 38704
rect -200 38623 -184 38657
rect 184 38623 200 38657
rect -200 38607 200 38623
rect -200 38549 200 38565
rect -200 38515 -184 38549
rect 184 38515 200 38549
rect -200 38468 200 38515
rect -200 38221 200 38268
rect -200 38187 -184 38221
rect 184 38187 200 38221
rect -200 38171 200 38187
rect -200 38113 200 38129
rect -200 38079 -184 38113
rect 184 38079 200 38113
rect -200 38032 200 38079
rect -200 37785 200 37832
rect -200 37751 -184 37785
rect 184 37751 200 37785
rect -200 37735 200 37751
rect -200 37677 200 37693
rect -200 37643 -184 37677
rect 184 37643 200 37677
rect -200 37596 200 37643
rect -200 37349 200 37396
rect -200 37315 -184 37349
rect 184 37315 200 37349
rect -200 37299 200 37315
rect -200 37241 200 37257
rect -200 37207 -184 37241
rect 184 37207 200 37241
rect -200 37160 200 37207
rect -200 36913 200 36960
rect -200 36879 -184 36913
rect 184 36879 200 36913
rect -200 36863 200 36879
rect -200 36805 200 36821
rect -200 36771 -184 36805
rect 184 36771 200 36805
rect -200 36724 200 36771
rect -200 36477 200 36524
rect -200 36443 -184 36477
rect 184 36443 200 36477
rect -200 36427 200 36443
rect -200 36369 200 36385
rect -200 36335 -184 36369
rect 184 36335 200 36369
rect -200 36288 200 36335
rect -200 36041 200 36088
rect -200 36007 -184 36041
rect 184 36007 200 36041
rect -200 35991 200 36007
rect -200 35933 200 35949
rect -200 35899 -184 35933
rect 184 35899 200 35933
rect -200 35852 200 35899
rect -200 35605 200 35652
rect -200 35571 -184 35605
rect 184 35571 200 35605
rect -200 35555 200 35571
rect -200 35497 200 35513
rect -200 35463 -184 35497
rect 184 35463 200 35497
rect -200 35416 200 35463
rect -200 35169 200 35216
rect -200 35135 -184 35169
rect 184 35135 200 35169
rect -200 35119 200 35135
rect -200 35061 200 35077
rect -200 35027 -184 35061
rect 184 35027 200 35061
rect -200 34980 200 35027
rect -200 34733 200 34780
rect -200 34699 -184 34733
rect 184 34699 200 34733
rect -200 34683 200 34699
rect -200 34625 200 34641
rect -200 34591 -184 34625
rect 184 34591 200 34625
rect -200 34544 200 34591
rect -200 34297 200 34344
rect -200 34263 -184 34297
rect 184 34263 200 34297
rect -200 34247 200 34263
rect -200 34189 200 34205
rect -200 34155 -184 34189
rect 184 34155 200 34189
rect -200 34108 200 34155
rect -200 33861 200 33908
rect -200 33827 -184 33861
rect 184 33827 200 33861
rect -200 33811 200 33827
rect -200 33753 200 33769
rect -200 33719 -184 33753
rect 184 33719 200 33753
rect -200 33672 200 33719
rect -200 33425 200 33472
rect -200 33391 -184 33425
rect 184 33391 200 33425
rect -200 33375 200 33391
rect -200 33317 200 33333
rect -200 33283 -184 33317
rect 184 33283 200 33317
rect -200 33236 200 33283
rect -200 32989 200 33036
rect -200 32955 -184 32989
rect 184 32955 200 32989
rect -200 32939 200 32955
rect -200 32881 200 32897
rect -200 32847 -184 32881
rect 184 32847 200 32881
rect -200 32800 200 32847
rect -200 32553 200 32600
rect -200 32519 -184 32553
rect 184 32519 200 32553
rect -200 32503 200 32519
rect -200 32445 200 32461
rect -200 32411 -184 32445
rect 184 32411 200 32445
rect -200 32364 200 32411
rect -200 32117 200 32164
rect -200 32083 -184 32117
rect 184 32083 200 32117
rect -200 32067 200 32083
rect -200 32009 200 32025
rect -200 31975 -184 32009
rect 184 31975 200 32009
rect -200 31928 200 31975
rect -200 31681 200 31728
rect -200 31647 -184 31681
rect 184 31647 200 31681
rect -200 31631 200 31647
rect -200 31573 200 31589
rect -200 31539 -184 31573
rect 184 31539 200 31573
rect -200 31492 200 31539
rect -200 31245 200 31292
rect -200 31211 -184 31245
rect 184 31211 200 31245
rect -200 31195 200 31211
rect -200 31137 200 31153
rect -200 31103 -184 31137
rect 184 31103 200 31137
rect -200 31056 200 31103
rect -200 30809 200 30856
rect -200 30775 -184 30809
rect 184 30775 200 30809
rect -200 30759 200 30775
rect -200 30701 200 30717
rect -200 30667 -184 30701
rect 184 30667 200 30701
rect -200 30620 200 30667
rect -200 30373 200 30420
rect -200 30339 -184 30373
rect 184 30339 200 30373
rect -200 30323 200 30339
rect -200 30265 200 30281
rect -200 30231 -184 30265
rect 184 30231 200 30265
rect -200 30184 200 30231
rect -200 29937 200 29984
rect -200 29903 -184 29937
rect 184 29903 200 29937
rect -200 29887 200 29903
rect -200 29829 200 29845
rect -200 29795 -184 29829
rect 184 29795 200 29829
rect -200 29748 200 29795
rect -200 29501 200 29548
rect -200 29467 -184 29501
rect 184 29467 200 29501
rect -200 29451 200 29467
rect -200 29393 200 29409
rect -200 29359 -184 29393
rect 184 29359 200 29393
rect -200 29312 200 29359
rect -200 29065 200 29112
rect -200 29031 -184 29065
rect 184 29031 200 29065
rect -200 29015 200 29031
rect -200 28957 200 28973
rect -200 28923 -184 28957
rect 184 28923 200 28957
rect -200 28876 200 28923
rect -200 28629 200 28676
rect -200 28595 -184 28629
rect 184 28595 200 28629
rect -200 28579 200 28595
rect -200 28521 200 28537
rect -200 28487 -184 28521
rect 184 28487 200 28521
rect -200 28440 200 28487
rect -200 28193 200 28240
rect -200 28159 -184 28193
rect 184 28159 200 28193
rect -200 28143 200 28159
rect -200 28085 200 28101
rect -200 28051 -184 28085
rect 184 28051 200 28085
rect -200 28004 200 28051
rect -200 27757 200 27804
rect -200 27723 -184 27757
rect 184 27723 200 27757
rect -200 27707 200 27723
rect -200 27649 200 27665
rect -200 27615 -184 27649
rect 184 27615 200 27649
rect -200 27568 200 27615
rect -200 27321 200 27368
rect -200 27287 -184 27321
rect 184 27287 200 27321
rect -200 27271 200 27287
rect -200 27213 200 27229
rect -200 27179 -184 27213
rect 184 27179 200 27213
rect -200 27132 200 27179
rect -200 26885 200 26932
rect -200 26851 -184 26885
rect 184 26851 200 26885
rect -200 26835 200 26851
rect -200 26777 200 26793
rect -200 26743 -184 26777
rect 184 26743 200 26777
rect -200 26696 200 26743
rect -200 26449 200 26496
rect -200 26415 -184 26449
rect 184 26415 200 26449
rect -200 26399 200 26415
rect -200 26341 200 26357
rect -200 26307 -184 26341
rect 184 26307 200 26341
rect -200 26260 200 26307
rect -200 26013 200 26060
rect -200 25979 -184 26013
rect 184 25979 200 26013
rect -200 25963 200 25979
rect -200 25905 200 25921
rect -200 25871 -184 25905
rect 184 25871 200 25905
rect -200 25824 200 25871
rect -200 25577 200 25624
rect -200 25543 -184 25577
rect 184 25543 200 25577
rect -200 25527 200 25543
rect -200 25469 200 25485
rect -200 25435 -184 25469
rect 184 25435 200 25469
rect -200 25388 200 25435
rect -200 25141 200 25188
rect -200 25107 -184 25141
rect 184 25107 200 25141
rect -200 25091 200 25107
rect -200 25033 200 25049
rect -200 24999 -184 25033
rect 184 24999 200 25033
rect -200 24952 200 24999
rect -200 24705 200 24752
rect -200 24671 -184 24705
rect 184 24671 200 24705
rect -200 24655 200 24671
rect -200 24597 200 24613
rect -200 24563 -184 24597
rect 184 24563 200 24597
rect -200 24516 200 24563
rect -200 24269 200 24316
rect -200 24235 -184 24269
rect 184 24235 200 24269
rect -200 24219 200 24235
rect -200 24161 200 24177
rect -200 24127 -184 24161
rect 184 24127 200 24161
rect -200 24080 200 24127
rect -200 23833 200 23880
rect -200 23799 -184 23833
rect 184 23799 200 23833
rect -200 23783 200 23799
rect -200 23725 200 23741
rect -200 23691 -184 23725
rect 184 23691 200 23725
rect -200 23644 200 23691
rect -200 23397 200 23444
rect -200 23363 -184 23397
rect 184 23363 200 23397
rect -200 23347 200 23363
rect -200 23289 200 23305
rect -200 23255 -184 23289
rect 184 23255 200 23289
rect -200 23208 200 23255
rect -200 22961 200 23008
rect -200 22927 -184 22961
rect 184 22927 200 22961
rect -200 22911 200 22927
rect -200 22853 200 22869
rect -200 22819 -184 22853
rect 184 22819 200 22853
rect -200 22772 200 22819
rect -200 22525 200 22572
rect -200 22491 -184 22525
rect 184 22491 200 22525
rect -200 22475 200 22491
rect -200 22417 200 22433
rect -200 22383 -184 22417
rect 184 22383 200 22417
rect -200 22336 200 22383
rect -200 22089 200 22136
rect -200 22055 -184 22089
rect 184 22055 200 22089
rect -200 22039 200 22055
rect -200 21981 200 21997
rect -200 21947 -184 21981
rect 184 21947 200 21981
rect -200 21900 200 21947
rect -200 21653 200 21700
rect -200 21619 -184 21653
rect 184 21619 200 21653
rect -200 21603 200 21619
rect -200 21545 200 21561
rect -200 21511 -184 21545
rect 184 21511 200 21545
rect -200 21464 200 21511
rect -200 21217 200 21264
rect -200 21183 -184 21217
rect 184 21183 200 21217
rect -200 21167 200 21183
rect -200 21109 200 21125
rect -200 21075 -184 21109
rect 184 21075 200 21109
rect -200 21028 200 21075
rect -200 20781 200 20828
rect -200 20747 -184 20781
rect 184 20747 200 20781
rect -200 20731 200 20747
rect -200 20673 200 20689
rect -200 20639 -184 20673
rect 184 20639 200 20673
rect -200 20592 200 20639
rect -200 20345 200 20392
rect -200 20311 -184 20345
rect 184 20311 200 20345
rect -200 20295 200 20311
rect -200 20237 200 20253
rect -200 20203 -184 20237
rect 184 20203 200 20237
rect -200 20156 200 20203
rect -200 19909 200 19956
rect -200 19875 -184 19909
rect 184 19875 200 19909
rect -200 19859 200 19875
rect -200 19801 200 19817
rect -200 19767 -184 19801
rect 184 19767 200 19801
rect -200 19720 200 19767
rect -200 19473 200 19520
rect -200 19439 -184 19473
rect 184 19439 200 19473
rect -200 19423 200 19439
rect -200 19365 200 19381
rect -200 19331 -184 19365
rect 184 19331 200 19365
rect -200 19284 200 19331
rect -200 19037 200 19084
rect -200 19003 -184 19037
rect 184 19003 200 19037
rect -200 18987 200 19003
rect -200 18929 200 18945
rect -200 18895 -184 18929
rect 184 18895 200 18929
rect -200 18848 200 18895
rect -200 18601 200 18648
rect -200 18567 -184 18601
rect 184 18567 200 18601
rect -200 18551 200 18567
rect -200 18493 200 18509
rect -200 18459 -184 18493
rect 184 18459 200 18493
rect -200 18412 200 18459
rect -200 18165 200 18212
rect -200 18131 -184 18165
rect 184 18131 200 18165
rect -200 18115 200 18131
rect -200 18057 200 18073
rect -200 18023 -184 18057
rect 184 18023 200 18057
rect -200 17976 200 18023
rect -200 17729 200 17776
rect -200 17695 -184 17729
rect 184 17695 200 17729
rect -200 17679 200 17695
rect -200 17621 200 17637
rect -200 17587 -184 17621
rect 184 17587 200 17621
rect -200 17540 200 17587
rect -200 17293 200 17340
rect -200 17259 -184 17293
rect 184 17259 200 17293
rect -200 17243 200 17259
rect -200 17185 200 17201
rect -200 17151 -184 17185
rect 184 17151 200 17185
rect -200 17104 200 17151
rect -200 16857 200 16904
rect -200 16823 -184 16857
rect 184 16823 200 16857
rect -200 16807 200 16823
rect -200 16749 200 16765
rect -200 16715 -184 16749
rect 184 16715 200 16749
rect -200 16668 200 16715
rect -200 16421 200 16468
rect -200 16387 -184 16421
rect 184 16387 200 16421
rect -200 16371 200 16387
rect -200 16313 200 16329
rect -200 16279 -184 16313
rect 184 16279 200 16313
rect -200 16232 200 16279
rect -200 15985 200 16032
rect -200 15951 -184 15985
rect 184 15951 200 15985
rect -200 15935 200 15951
rect -200 15877 200 15893
rect -200 15843 -184 15877
rect 184 15843 200 15877
rect -200 15796 200 15843
rect -200 15549 200 15596
rect -200 15515 -184 15549
rect 184 15515 200 15549
rect -200 15499 200 15515
rect -200 15441 200 15457
rect -200 15407 -184 15441
rect 184 15407 200 15441
rect -200 15360 200 15407
rect -200 15113 200 15160
rect -200 15079 -184 15113
rect 184 15079 200 15113
rect -200 15063 200 15079
rect -200 15005 200 15021
rect -200 14971 -184 15005
rect 184 14971 200 15005
rect -200 14924 200 14971
rect -200 14677 200 14724
rect -200 14643 -184 14677
rect 184 14643 200 14677
rect -200 14627 200 14643
rect -200 14569 200 14585
rect -200 14535 -184 14569
rect 184 14535 200 14569
rect -200 14488 200 14535
rect -200 14241 200 14288
rect -200 14207 -184 14241
rect 184 14207 200 14241
rect -200 14191 200 14207
rect -200 14133 200 14149
rect -200 14099 -184 14133
rect 184 14099 200 14133
rect -200 14052 200 14099
rect -200 13805 200 13852
rect -200 13771 -184 13805
rect 184 13771 200 13805
rect -200 13755 200 13771
rect -200 13697 200 13713
rect -200 13663 -184 13697
rect 184 13663 200 13697
rect -200 13616 200 13663
rect -200 13369 200 13416
rect -200 13335 -184 13369
rect 184 13335 200 13369
rect -200 13319 200 13335
rect -200 13261 200 13277
rect -200 13227 -184 13261
rect 184 13227 200 13261
rect -200 13180 200 13227
rect -200 12933 200 12980
rect -200 12899 -184 12933
rect 184 12899 200 12933
rect -200 12883 200 12899
rect -200 12825 200 12841
rect -200 12791 -184 12825
rect 184 12791 200 12825
rect -200 12744 200 12791
rect -200 12497 200 12544
rect -200 12463 -184 12497
rect 184 12463 200 12497
rect -200 12447 200 12463
rect -200 12389 200 12405
rect -200 12355 -184 12389
rect 184 12355 200 12389
rect -200 12308 200 12355
rect -200 12061 200 12108
rect -200 12027 -184 12061
rect 184 12027 200 12061
rect -200 12011 200 12027
rect -200 11953 200 11969
rect -200 11919 -184 11953
rect 184 11919 200 11953
rect -200 11872 200 11919
rect -200 11625 200 11672
rect -200 11591 -184 11625
rect 184 11591 200 11625
rect -200 11575 200 11591
rect -200 11517 200 11533
rect -200 11483 -184 11517
rect 184 11483 200 11517
rect -200 11436 200 11483
rect -200 11189 200 11236
rect -200 11155 -184 11189
rect 184 11155 200 11189
rect -200 11139 200 11155
rect -200 11081 200 11097
rect -200 11047 -184 11081
rect 184 11047 200 11081
rect -200 11000 200 11047
rect -200 10753 200 10800
rect -200 10719 -184 10753
rect 184 10719 200 10753
rect -200 10703 200 10719
rect -200 10645 200 10661
rect -200 10611 -184 10645
rect 184 10611 200 10645
rect -200 10564 200 10611
rect -200 10317 200 10364
rect -200 10283 -184 10317
rect 184 10283 200 10317
rect -200 10267 200 10283
rect -200 10209 200 10225
rect -200 10175 -184 10209
rect 184 10175 200 10209
rect -200 10128 200 10175
rect -200 9881 200 9928
rect -200 9847 -184 9881
rect 184 9847 200 9881
rect -200 9831 200 9847
rect -200 9773 200 9789
rect -200 9739 -184 9773
rect 184 9739 200 9773
rect -200 9692 200 9739
rect -200 9445 200 9492
rect -200 9411 -184 9445
rect 184 9411 200 9445
rect -200 9395 200 9411
rect -200 9337 200 9353
rect -200 9303 -184 9337
rect 184 9303 200 9337
rect -200 9256 200 9303
rect -200 9009 200 9056
rect -200 8975 -184 9009
rect 184 8975 200 9009
rect -200 8959 200 8975
rect -200 8901 200 8917
rect -200 8867 -184 8901
rect 184 8867 200 8901
rect -200 8820 200 8867
rect -200 8573 200 8620
rect -200 8539 -184 8573
rect 184 8539 200 8573
rect -200 8523 200 8539
rect -200 8465 200 8481
rect -200 8431 -184 8465
rect 184 8431 200 8465
rect -200 8384 200 8431
rect -200 8137 200 8184
rect -200 8103 -184 8137
rect 184 8103 200 8137
rect -200 8087 200 8103
rect -200 8029 200 8045
rect -200 7995 -184 8029
rect 184 7995 200 8029
rect -200 7948 200 7995
rect -200 7701 200 7748
rect -200 7667 -184 7701
rect 184 7667 200 7701
rect -200 7651 200 7667
rect -200 7593 200 7609
rect -200 7559 -184 7593
rect 184 7559 200 7593
rect -200 7512 200 7559
rect -200 7265 200 7312
rect -200 7231 -184 7265
rect 184 7231 200 7265
rect -200 7215 200 7231
rect -200 7157 200 7173
rect -200 7123 -184 7157
rect 184 7123 200 7157
rect -200 7076 200 7123
rect -200 6829 200 6876
rect -200 6795 -184 6829
rect 184 6795 200 6829
rect -200 6779 200 6795
rect -200 6721 200 6737
rect -200 6687 -184 6721
rect 184 6687 200 6721
rect -200 6640 200 6687
rect -200 6393 200 6440
rect -200 6359 -184 6393
rect 184 6359 200 6393
rect -200 6343 200 6359
rect -200 6285 200 6301
rect -200 6251 -184 6285
rect 184 6251 200 6285
rect -200 6204 200 6251
rect -200 5957 200 6004
rect -200 5923 -184 5957
rect 184 5923 200 5957
rect -200 5907 200 5923
rect -200 5849 200 5865
rect -200 5815 -184 5849
rect 184 5815 200 5849
rect -200 5768 200 5815
rect -200 5521 200 5568
rect -200 5487 -184 5521
rect 184 5487 200 5521
rect -200 5471 200 5487
rect -200 5413 200 5429
rect -200 5379 -184 5413
rect 184 5379 200 5413
rect -200 5332 200 5379
rect -200 5085 200 5132
rect -200 5051 -184 5085
rect 184 5051 200 5085
rect -200 5035 200 5051
rect -200 4977 200 4993
rect -200 4943 -184 4977
rect 184 4943 200 4977
rect -200 4896 200 4943
rect -200 4649 200 4696
rect -200 4615 -184 4649
rect 184 4615 200 4649
rect -200 4599 200 4615
rect -200 4541 200 4557
rect -200 4507 -184 4541
rect 184 4507 200 4541
rect -200 4460 200 4507
rect -200 4213 200 4260
rect -200 4179 -184 4213
rect 184 4179 200 4213
rect -200 4163 200 4179
rect -200 4105 200 4121
rect -200 4071 -184 4105
rect 184 4071 200 4105
rect -200 4024 200 4071
rect -200 3777 200 3824
rect -200 3743 -184 3777
rect 184 3743 200 3777
rect -200 3727 200 3743
rect -200 3669 200 3685
rect -200 3635 -184 3669
rect 184 3635 200 3669
rect -200 3588 200 3635
rect -200 3341 200 3388
rect -200 3307 -184 3341
rect 184 3307 200 3341
rect -200 3291 200 3307
rect -200 3233 200 3249
rect -200 3199 -184 3233
rect 184 3199 200 3233
rect -200 3152 200 3199
rect -200 2905 200 2952
rect -200 2871 -184 2905
rect 184 2871 200 2905
rect -200 2855 200 2871
rect -200 2797 200 2813
rect -200 2763 -184 2797
rect 184 2763 200 2797
rect -200 2716 200 2763
rect -200 2469 200 2516
rect -200 2435 -184 2469
rect 184 2435 200 2469
rect -200 2419 200 2435
rect -200 2361 200 2377
rect -200 2327 -184 2361
rect 184 2327 200 2361
rect -200 2280 200 2327
rect -200 2033 200 2080
rect -200 1999 -184 2033
rect 184 1999 200 2033
rect -200 1983 200 1999
rect -200 1925 200 1941
rect -200 1891 -184 1925
rect 184 1891 200 1925
rect -200 1844 200 1891
rect -200 1597 200 1644
rect -200 1563 -184 1597
rect 184 1563 200 1597
rect -200 1547 200 1563
rect -200 1489 200 1505
rect -200 1455 -184 1489
rect 184 1455 200 1489
rect -200 1408 200 1455
rect -200 1161 200 1208
rect -200 1127 -184 1161
rect 184 1127 200 1161
rect -200 1111 200 1127
rect -200 1053 200 1069
rect -200 1019 -184 1053
rect 184 1019 200 1053
rect -200 972 200 1019
rect -200 725 200 772
rect -200 691 -184 725
rect 184 691 200 725
rect -200 675 200 691
rect -200 617 200 633
rect -200 583 -184 617
rect 184 583 200 617
rect -200 536 200 583
rect -200 289 200 336
rect -200 255 -184 289
rect 184 255 200 289
rect -200 239 200 255
rect -200 181 200 197
rect -200 147 -184 181
rect 184 147 200 181
rect -200 100 200 147
rect -200 -147 200 -100
rect -200 -181 -184 -147
rect 184 -181 200 -147
rect -200 -197 200 -181
rect -200 -255 200 -239
rect -200 -289 -184 -255
rect 184 -289 200 -255
rect -200 -336 200 -289
rect -200 -583 200 -536
rect -200 -617 -184 -583
rect 184 -617 200 -583
rect -200 -633 200 -617
rect -200 -691 200 -675
rect -200 -725 -184 -691
rect 184 -725 200 -691
rect -200 -772 200 -725
rect -200 -1019 200 -972
rect -200 -1053 -184 -1019
rect 184 -1053 200 -1019
rect -200 -1069 200 -1053
rect -200 -1127 200 -1111
rect -200 -1161 -184 -1127
rect 184 -1161 200 -1127
rect -200 -1208 200 -1161
rect -200 -1455 200 -1408
rect -200 -1489 -184 -1455
rect 184 -1489 200 -1455
rect -200 -1505 200 -1489
rect -200 -1563 200 -1547
rect -200 -1597 -184 -1563
rect 184 -1597 200 -1563
rect -200 -1644 200 -1597
rect -200 -1891 200 -1844
rect -200 -1925 -184 -1891
rect 184 -1925 200 -1891
rect -200 -1941 200 -1925
rect -200 -1999 200 -1983
rect -200 -2033 -184 -1999
rect 184 -2033 200 -1999
rect -200 -2080 200 -2033
rect -200 -2327 200 -2280
rect -200 -2361 -184 -2327
rect 184 -2361 200 -2327
rect -200 -2377 200 -2361
rect -200 -2435 200 -2419
rect -200 -2469 -184 -2435
rect 184 -2469 200 -2435
rect -200 -2516 200 -2469
rect -200 -2763 200 -2716
rect -200 -2797 -184 -2763
rect 184 -2797 200 -2763
rect -200 -2813 200 -2797
rect -200 -2871 200 -2855
rect -200 -2905 -184 -2871
rect 184 -2905 200 -2871
rect -200 -2952 200 -2905
rect -200 -3199 200 -3152
rect -200 -3233 -184 -3199
rect 184 -3233 200 -3199
rect -200 -3249 200 -3233
rect -200 -3307 200 -3291
rect -200 -3341 -184 -3307
rect 184 -3341 200 -3307
rect -200 -3388 200 -3341
rect -200 -3635 200 -3588
rect -200 -3669 -184 -3635
rect 184 -3669 200 -3635
rect -200 -3685 200 -3669
rect -200 -3743 200 -3727
rect -200 -3777 -184 -3743
rect 184 -3777 200 -3743
rect -200 -3824 200 -3777
rect -200 -4071 200 -4024
rect -200 -4105 -184 -4071
rect 184 -4105 200 -4071
rect -200 -4121 200 -4105
rect -200 -4179 200 -4163
rect -200 -4213 -184 -4179
rect 184 -4213 200 -4179
rect -200 -4260 200 -4213
rect -200 -4507 200 -4460
rect -200 -4541 -184 -4507
rect 184 -4541 200 -4507
rect -200 -4557 200 -4541
rect -200 -4615 200 -4599
rect -200 -4649 -184 -4615
rect 184 -4649 200 -4615
rect -200 -4696 200 -4649
rect -200 -4943 200 -4896
rect -200 -4977 -184 -4943
rect 184 -4977 200 -4943
rect -200 -4993 200 -4977
rect -200 -5051 200 -5035
rect -200 -5085 -184 -5051
rect 184 -5085 200 -5051
rect -200 -5132 200 -5085
rect -200 -5379 200 -5332
rect -200 -5413 -184 -5379
rect 184 -5413 200 -5379
rect -200 -5429 200 -5413
rect -200 -5487 200 -5471
rect -200 -5521 -184 -5487
rect 184 -5521 200 -5487
rect -200 -5568 200 -5521
rect -200 -5815 200 -5768
rect -200 -5849 -184 -5815
rect 184 -5849 200 -5815
rect -200 -5865 200 -5849
rect -200 -5923 200 -5907
rect -200 -5957 -184 -5923
rect 184 -5957 200 -5923
rect -200 -6004 200 -5957
rect -200 -6251 200 -6204
rect -200 -6285 -184 -6251
rect 184 -6285 200 -6251
rect -200 -6301 200 -6285
rect -200 -6359 200 -6343
rect -200 -6393 -184 -6359
rect 184 -6393 200 -6359
rect -200 -6440 200 -6393
rect -200 -6687 200 -6640
rect -200 -6721 -184 -6687
rect 184 -6721 200 -6687
rect -200 -6737 200 -6721
rect -200 -6795 200 -6779
rect -200 -6829 -184 -6795
rect 184 -6829 200 -6795
rect -200 -6876 200 -6829
rect -200 -7123 200 -7076
rect -200 -7157 -184 -7123
rect 184 -7157 200 -7123
rect -200 -7173 200 -7157
rect -200 -7231 200 -7215
rect -200 -7265 -184 -7231
rect 184 -7265 200 -7231
rect -200 -7312 200 -7265
rect -200 -7559 200 -7512
rect -200 -7593 -184 -7559
rect 184 -7593 200 -7559
rect -200 -7609 200 -7593
rect -200 -7667 200 -7651
rect -200 -7701 -184 -7667
rect 184 -7701 200 -7667
rect -200 -7748 200 -7701
rect -200 -7995 200 -7948
rect -200 -8029 -184 -7995
rect 184 -8029 200 -7995
rect -200 -8045 200 -8029
rect -200 -8103 200 -8087
rect -200 -8137 -184 -8103
rect 184 -8137 200 -8103
rect -200 -8184 200 -8137
rect -200 -8431 200 -8384
rect -200 -8465 -184 -8431
rect 184 -8465 200 -8431
rect -200 -8481 200 -8465
rect -200 -8539 200 -8523
rect -200 -8573 -184 -8539
rect 184 -8573 200 -8539
rect -200 -8620 200 -8573
rect -200 -8867 200 -8820
rect -200 -8901 -184 -8867
rect 184 -8901 200 -8867
rect -200 -8917 200 -8901
rect -200 -8975 200 -8959
rect -200 -9009 -184 -8975
rect 184 -9009 200 -8975
rect -200 -9056 200 -9009
rect -200 -9303 200 -9256
rect -200 -9337 -184 -9303
rect 184 -9337 200 -9303
rect -200 -9353 200 -9337
rect -200 -9411 200 -9395
rect -200 -9445 -184 -9411
rect 184 -9445 200 -9411
rect -200 -9492 200 -9445
rect -200 -9739 200 -9692
rect -200 -9773 -184 -9739
rect 184 -9773 200 -9739
rect -200 -9789 200 -9773
rect -200 -9847 200 -9831
rect -200 -9881 -184 -9847
rect 184 -9881 200 -9847
rect -200 -9928 200 -9881
rect -200 -10175 200 -10128
rect -200 -10209 -184 -10175
rect 184 -10209 200 -10175
rect -200 -10225 200 -10209
rect -200 -10283 200 -10267
rect -200 -10317 -184 -10283
rect 184 -10317 200 -10283
rect -200 -10364 200 -10317
rect -200 -10611 200 -10564
rect -200 -10645 -184 -10611
rect 184 -10645 200 -10611
rect -200 -10661 200 -10645
rect -200 -10719 200 -10703
rect -200 -10753 -184 -10719
rect 184 -10753 200 -10719
rect -200 -10800 200 -10753
rect -200 -11047 200 -11000
rect -200 -11081 -184 -11047
rect 184 -11081 200 -11047
rect -200 -11097 200 -11081
rect -200 -11155 200 -11139
rect -200 -11189 -184 -11155
rect 184 -11189 200 -11155
rect -200 -11236 200 -11189
rect -200 -11483 200 -11436
rect -200 -11517 -184 -11483
rect 184 -11517 200 -11483
rect -200 -11533 200 -11517
rect -200 -11591 200 -11575
rect -200 -11625 -184 -11591
rect 184 -11625 200 -11591
rect -200 -11672 200 -11625
rect -200 -11919 200 -11872
rect -200 -11953 -184 -11919
rect 184 -11953 200 -11919
rect -200 -11969 200 -11953
rect -200 -12027 200 -12011
rect -200 -12061 -184 -12027
rect 184 -12061 200 -12027
rect -200 -12108 200 -12061
rect -200 -12355 200 -12308
rect -200 -12389 -184 -12355
rect 184 -12389 200 -12355
rect -200 -12405 200 -12389
rect -200 -12463 200 -12447
rect -200 -12497 -184 -12463
rect 184 -12497 200 -12463
rect -200 -12544 200 -12497
rect -200 -12791 200 -12744
rect -200 -12825 -184 -12791
rect 184 -12825 200 -12791
rect -200 -12841 200 -12825
rect -200 -12899 200 -12883
rect -200 -12933 -184 -12899
rect 184 -12933 200 -12899
rect -200 -12980 200 -12933
rect -200 -13227 200 -13180
rect -200 -13261 -184 -13227
rect 184 -13261 200 -13227
rect -200 -13277 200 -13261
rect -200 -13335 200 -13319
rect -200 -13369 -184 -13335
rect 184 -13369 200 -13335
rect -200 -13416 200 -13369
rect -200 -13663 200 -13616
rect -200 -13697 -184 -13663
rect 184 -13697 200 -13663
rect -200 -13713 200 -13697
rect -200 -13771 200 -13755
rect -200 -13805 -184 -13771
rect 184 -13805 200 -13771
rect -200 -13852 200 -13805
rect -200 -14099 200 -14052
rect -200 -14133 -184 -14099
rect 184 -14133 200 -14099
rect -200 -14149 200 -14133
rect -200 -14207 200 -14191
rect -200 -14241 -184 -14207
rect 184 -14241 200 -14207
rect -200 -14288 200 -14241
rect -200 -14535 200 -14488
rect -200 -14569 -184 -14535
rect 184 -14569 200 -14535
rect -200 -14585 200 -14569
rect -200 -14643 200 -14627
rect -200 -14677 -184 -14643
rect 184 -14677 200 -14643
rect -200 -14724 200 -14677
rect -200 -14971 200 -14924
rect -200 -15005 -184 -14971
rect 184 -15005 200 -14971
rect -200 -15021 200 -15005
rect -200 -15079 200 -15063
rect -200 -15113 -184 -15079
rect 184 -15113 200 -15079
rect -200 -15160 200 -15113
rect -200 -15407 200 -15360
rect -200 -15441 -184 -15407
rect 184 -15441 200 -15407
rect -200 -15457 200 -15441
rect -200 -15515 200 -15499
rect -200 -15549 -184 -15515
rect 184 -15549 200 -15515
rect -200 -15596 200 -15549
rect -200 -15843 200 -15796
rect -200 -15877 -184 -15843
rect 184 -15877 200 -15843
rect -200 -15893 200 -15877
rect -200 -15951 200 -15935
rect -200 -15985 -184 -15951
rect 184 -15985 200 -15951
rect -200 -16032 200 -15985
rect -200 -16279 200 -16232
rect -200 -16313 -184 -16279
rect 184 -16313 200 -16279
rect -200 -16329 200 -16313
rect -200 -16387 200 -16371
rect -200 -16421 -184 -16387
rect 184 -16421 200 -16387
rect -200 -16468 200 -16421
rect -200 -16715 200 -16668
rect -200 -16749 -184 -16715
rect 184 -16749 200 -16715
rect -200 -16765 200 -16749
rect -200 -16823 200 -16807
rect -200 -16857 -184 -16823
rect 184 -16857 200 -16823
rect -200 -16904 200 -16857
rect -200 -17151 200 -17104
rect -200 -17185 -184 -17151
rect 184 -17185 200 -17151
rect -200 -17201 200 -17185
rect -200 -17259 200 -17243
rect -200 -17293 -184 -17259
rect 184 -17293 200 -17259
rect -200 -17340 200 -17293
rect -200 -17587 200 -17540
rect -200 -17621 -184 -17587
rect 184 -17621 200 -17587
rect -200 -17637 200 -17621
rect -200 -17695 200 -17679
rect -200 -17729 -184 -17695
rect 184 -17729 200 -17695
rect -200 -17776 200 -17729
rect -200 -18023 200 -17976
rect -200 -18057 -184 -18023
rect 184 -18057 200 -18023
rect -200 -18073 200 -18057
rect -200 -18131 200 -18115
rect -200 -18165 -184 -18131
rect 184 -18165 200 -18131
rect -200 -18212 200 -18165
rect -200 -18459 200 -18412
rect -200 -18493 -184 -18459
rect 184 -18493 200 -18459
rect -200 -18509 200 -18493
rect -200 -18567 200 -18551
rect -200 -18601 -184 -18567
rect 184 -18601 200 -18567
rect -200 -18648 200 -18601
rect -200 -18895 200 -18848
rect -200 -18929 -184 -18895
rect 184 -18929 200 -18895
rect -200 -18945 200 -18929
rect -200 -19003 200 -18987
rect -200 -19037 -184 -19003
rect 184 -19037 200 -19003
rect -200 -19084 200 -19037
rect -200 -19331 200 -19284
rect -200 -19365 -184 -19331
rect 184 -19365 200 -19331
rect -200 -19381 200 -19365
rect -200 -19439 200 -19423
rect -200 -19473 -184 -19439
rect 184 -19473 200 -19439
rect -200 -19520 200 -19473
rect -200 -19767 200 -19720
rect -200 -19801 -184 -19767
rect 184 -19801 200 -19767
rect -200 -19817 200 -19801
rect -200 -19875 200 -19859
rect -200 -19909 -184 -19875
rect 184 -19909 200 -19875
rect -200 -19956 200 -19909
rect -200 -20203 200 -20156
rect -200 -20237 -184 -20203
rect 184 -20237 200 -20203
rect -200 -20253 200 -20237
rect -200 -20311 200 -20295
rect -200 -20345 -184 -20311
rect 184 -20345 200 -20311
rect -200 -20392 200 -20345
rect -200 -20639 200 -20592
rect -200 -20673 -184 -20639
rect 184 -20673 200 -20639
rect -200 -20689 200 -20673
rect -200 -20747 200 -20731
rect -200 -20781 -184 -20747
rect 184 -20781 200 -20747
rect -200 -20828 200 -20781
rect -200 -21075 200 -21028
rect -200 -21109 -184 -21075
rect 184 -21109 200 -21075
rect -200 -21125 200 -21109
rect -200 -21183 200 -21167
rect -200 -21217 -184 -21183
rect 184 -21217 200 -21183
rect -200 -21264 200 -21217
rect -200 -21511 200 -21464
rect -200 -21545 -184 -21511
rect 184 -21545 200 -21511
rect -200 -21561 200 -21545
rect -200 -21619 200 -21603
rect -200 -21653 -184 -21619
rect 184 -21653 200 -21619
rect -200 -21700 200 -21653
rect -200 -21947 200 -21900
rect -200 -21981 -184 -21947
rect 184 -21981 200 -21947
rect -200 -21997 200 -21981
rect -200 -22055 200 -22039
rect -200 -22089 -184 -22055
rect 184 -22089 200 -22055
rect -200 -22136 200 -22089
rect -200 -22383 200 -22336
rect -200 -22417 -184 -22383
rect 184 -22417 200 -22383
rect -200 -22433 200 -22417
rect -200 -22491 200 -22475
rect -200 -22525 -184 -22491
rect 184 -22525 200 -22491
rect -200 -22572 200 -22525
rect -200 -22819 200 -22772
rect -200 -22853 -184 -22819
rect 184 -22853 200 -22819
rect -200 -22869 200 -22853
rect -200 -22927 200 -22911
rect -200 -22961 -184 -22927
rect 184 -22961 200 -22927
rect -200 -23008 200 -22961
rect -200 -23255 200 -23208
rect -200 -23289 -184 -23255
rect 184 -23289 200 -23255
rect -200 -23305 200 -23289
rect -200 -23363 200 -23347
rect -200 -23397 -184 -23363
rect 184 -23397 200 -23363
rect -200 -23444 200 -23397
rect -200 -23691 200 -23644
rect -200 -23725 -184 -23691
rect 184 -23725 200 -23691
rect -200 -23741 200 -23725
rect -200 -23799 200 -23783
rect -200 -23833 -184 -23799
rect 184 -23833 200 -23799
rect -200 -23880 200 -23833
rect -200 -24127 200 -24080
rect -200 -24161 -184 -24127
rect 184 -24161 200 -24127
rect -200 -24177 200 -24161
rect -200 -24235 200 -24219
rect -200 -24269 -184 -24235
rect 184 -24269 200 -24235
rect -200 -24316 200 -24269
rect -200 -24563 200 -24516
rect -200 -24597 -184 -24563
rect 184 -24597 200 -24563
rect -200 -24613 200 -24597
rect -200 -24671 200 -24655
rect -200 -24705 -184 -24671
rect 184 -24705 200 -24671
rect -200 -24752 200 -24705
rect -200 -24999 200 -24952
rect -200 -25033 -184 -24999
rect 184 -25033 200 -24999
rect -200 -25049 200 -25033
rect -200 -25107 200 -25091
rect -200 -25141 -184 -25107
rect 184 -25141 200 -25107
rect -200 -25188 200 -25141
rect -200 -25435 200 -25388
rect -200 -25469 -184 -25435
rect 184 -25469 200 -25435
rect -200 -25485 200 -25469
rect -200 -25543 200 -25527
rect -200 -25577 -184 -25543
rect 184 -25577 200 -25543
rect -200 -25624 200 -25577
rect -200 -25871 200 -25824
rect -200 -25905 -184 -25871
rect 184 -25905 200 -25871
rect -200 -25921 200 -25905
rect -200 -25979 200 -25963
rect -200 -26013 -184 -25979
rect 184 -26013 200 -25979
rect -200 -26060 200 -26013
rect -200 -26307 200 -26260
rect -200 -26341 -184 -26307
rect 184 -26341 200 -26307
rect -200 -26357 200 -26341
rect -200 -26415 200 -26399
rect -200 -26449 -184 -26415
rect 184 -26449 200 -26415
rect -200 -26496 200 -26449
rect -200 -26743 200 -26696
rect -200 -26777 -184 -26743
rect 184 -26777 200 -26743
rect -200 -26793 200 -26777
rect -200 -26851 200 -26835
rect -200 -26885 -184 -26851
rect 184 -26885 200 -26851
rect -200 -26932 200 -26885
rect -200 -27179 200 -27132
rect -200 -27213 -184 -27179
rect 184 -27213 200 -27179
rect -200 -27229 200 -27213
rect -200 -27287 200 -27271
rect -200 -27321 -184 -27287
rect 184 -27321 200 -27287
rect -200 -27368 200 -27321
rect -200 -27615 200 -27568
rect -200 -27649 -184 -27615
rect 184 -27649 200 -27615
rect -200 -27665 200 -27649
rect -200 -27723 200 -27707
rect -200 -27757 -184 -27723
rect 184 -27757 200 -27723
rect -200 -27804 200 -27757
rect -200 -28051 200 -28004
rect -200 -28085 -184 -28051
rect 184 -28085 200 -28051
rect -200 -28101 200 -28085
rect -200 -28159 200 -28143
rect -200 -28193 -184 -28159
rect 184 -28193 200 -28159
rect -200 -28240 200 -28193
rect -200 -28487 200 -28440
rect -200 -28521 -184 -28487
rect 184 -28521 200 -28487
rect -200 -28537 200 -28521
rect -200 -28595 200 -28579
rect -200 -28629 -184 -28595
rect 184 -28629 200 -28595
rect -200 -28676 200 -28629
rect -200 -28923 200 -28876
rect -200 -28957 -184 -28923
rect 184 -28957 200 -28923
rect -200 -28973 200 -28957
rect -200 -29031 200 -29015
rect -200 -29065 -184 -29031
rect 184 -29065 200 -29031
rect -200 -29112 200 -29065
rect -200 -29359 200 -29312
rect -200 -29393 -184 -29359
rect 184 -29393 200 -29359
rect -200 -29409 200 -29393
rect -200 -29467 200 -29451
rect -200 -29501 -184 -29467
rect 184 -29501 200 -29467
rect -200 -29548 200 -29501
rect -200 -29795 200 -29748
rect -200 -29829 -184 -29795
rect 184 -29829 200 -29795
rect -200 -29845 200 -29829
rect -200 -29903 200 -29887
rect -200 -29937 -184 -29903
rect 184 -29937 200 -29903
rect -200 -29984 200 -29937
rect -200 -30231 200 -30184
rect -200 -30265 -184 -30231
rect 184 -30265 200 -30231
rect -200 -30281 200 -30265
rect -200 -30339 200 -30323
rect -200 -30373 -184 -30339
rect 184 -30373 200 -30339
rect -200 -30420 200 -30373
rect -200 -30667 200 -30620
rect -200 -30701 -184 -30667
rect 184 -30701 200 -30667
rect -200 -30717 200 -30701
rect -200 -30775 200 -30759
rect -200 -30809 -184 -30775
rect 184 -30809 200 -30775
rect -200 -30856 200 -30809
rect -200 -31103 200 -31056
rect -200 -31137 -184 -31103
rect 184 -31137 200 -31103
rect -200 -31153 200 -31137
rect -200 -31211 200 -31195
rect -200 -31245 -184 -31211
rect 184 -31245 200 -31211
rect -200 -31292 200 -31245
rect -200 -31539 200 -31492
rect -200 -31573 -184 -31539
rect 184 -31573 200 -31539
rect -200 -31589 200 -31573
rect -200 -31647 200 -31631
rect -200 -31681 -184 -31647
rect 184 -31681 200 -31647
rect -200 -31728 200 -31681
rect -200 -31975 200 -31928
rect -200 -32009 -184 -31975
rect 184 -32009 200 -31975
rect -200 -32025 200 -32009
rect -200 -32083 200 -32067
rect -200 -32117 -184 -32083
rect 184 -32117 200 -32083
rect -200 -32164 200 -32117
rect -200 -32411 200 -32364
rect -200 -32445 -184 -32411
rect 184 -32445 200 -32411
rect -200 -32461 200 -32445
rect -200 -32519 200 -32503
rect -200 -32553 -184 -32519
rect 184 -32553 200 -32519
rect -200 -32600 200 -32553
rect -200 -32847 200 -32800
rect -200 -32881 -184 -32847
rect 184 -32881 200 -32847
rect -200 -32897 200 -32881
rect -200 -32955 200 -32939
rect -200 -32989 -184 -32955
rect 184 -32989 200 -32955
rect -200 -33036 200 -32989
rect -200 -33283 200 -33236
rect -200 -33317 -184 -33283
rect 184 -33317 200 -33283
rect -200 -33333 200 -33317
rect -200 -33391 200 -33375
rect -200 -33425 -184 -33391
rect 184 -33425 200 -33391
rect -200 -33472 200 -33425
rect -200 -33719 200 -33672
rect -200 -33753 -184 -33719
rect 184 -33753 200 -33719
rect -200 -33769 200 -33753
rect -200 -33827 200 -33811
rect -200 -33861 -184 -33827
rect 184 -33861 200 -33827
rect -200 -33908 200 -33861
rect -200 -34155 200 -34108
rect -200 -34189 -184 -34155
rect 184 -34189 200 -34155
rect -200 -34205 200 -34189
rect -200 -34263 200 -34247
rect -200 -34297 -184 -34263
rect 184 -34297 200 -34263
rect -200 -34344 200 -34297
rect -200 -34591 200 -34544
rect -200 -34625 -184 -34591
rect 184 -34625 200 -34591
rect -200 -34641 200 -34625
rect -200 -34699 200 -34683
rect -200 -34733 -184 -34699
rect 184 -34733 200 -34699
rect -200 -34780 200 -34733
rect -200 -35027 200 -34980
rect -200 -35061 -184 -35027
rect 184 -35061 200 -35027
rect -200 -35077 200 -35061
rect -200 -35135 200 -35119
rect -200 -35169 -184 -35135
rect 184 -35169 200 -35135
rect -200 -35216 200 -35169
rect -200 -35463 200 -35416
rect -200 -35497 -184 -35463
rect 184 -35497 200 -35463
rect -200 -35513 200 -35497
rect -200 -35571 200 -35555
rect -200 -35605 -184 -35571
rect 184 -35605 200 -35571
rect -200 -35652 200 -35605
rect -200 -35899 200 -35852
rect -200 -35933 -184 -35899
rect 184 -35933 200 -35899
rect -200 -35949 200 -35933
rect -200 -36007 200 -35991
rect -200 -36041 -184 -36007
rect 184 -36041 200 -36007
rect -200 -36088 200 -36041
rect -200 -36335 200 -36288
rect -200 -36369 -184 -36335
rect 184 -36369 200 -36335
rect -200 -36385 200 -36369
rect -200 -36443 200 -36427
rect -200 -36477 -184 -36443
rect 184 -36477 200 -36443
rect -200 -36524 200 -36477
rect -200 -36771 200 -36724
rect -200 -36805 -184 -36771
rect 184 -36805 200 -36771
rect -200 -36821 200 -36805
rect -200 -36879 200 -36863
rect -200 -36913 -184 -36879
rect 184 -36913 200 -36879
rect -200 -36960 200 -36913
rect -200 -37207 200 -37160
rect -200 -37241 -184 -37207
rect 184 -37241 200 -37207
rect -200 -37257 200 -37241
rect -200 -37315 200 -37299
rect -200 -37349 -184 -37315
rect 184 -37349 200 -37315
rect -200 -37396 200 -37349
rect -200 -37643 200 -37596
rect -200 -37677 -184 -37643
rect 184 -37677 200 -37643
rect -200 -37693 200 -37677
rect -200 -37751 200 -37735
rect -200 -37785 -184 -37751
rect 184 -37785 200 -37751
rect -200 -37832 200 -37785
rect -200 -38079 200 -38032
rect -200 -38113 -184 -38079
rect 184 -38113 200 -38079
rect -200 -38129 200 -38113
rect -200 -38187 200 -38171
rect -200 -38221 -184 -38187
rect 184 -38221 200 -38187
rect -200 -38268 200 -38221
rect -200 -38515 200 -38468
rect -200 -38549 -184 -38515
rect 184 -38549 200 -38515
rect -200 -38565 200 -38549
rect -200 -38623 200 -38607
rect -200 -38657 -184 -38623
rect 184 -38657 200 -38623
rect -200 -38704 200 -38657
rect -200 -38951 200 -38904
rect -200 -38985 -184 -38951
rect 184 -38985 200 -38951
rect -200 -39001 200 -38985
rect -200 -39059 200 -39043
rect -200 -39093 -184 -39059
rect 184 -39093 200 -39059
rect -200 -39140 200 -39093
rect -200 -39387 200 -39340
rect -200 -39421 -184 -39387
rect 184 -39421 200 -39387
rect -200 -39437 200 -39421
rect -200 -39495 200 -39479
rect -200 -39529 -184 -39495
rect 184 -39529 200 -39495
rect -200 -39576 200 -39529
rect -200 -39823 200 -39776
rect -200 -39857 -184 -39823
rect 184 -39857 200 -39823
rect -200 -39873 200 -39857
rect -200 -39931 200 -39915
rect -200 -39965 -184 -39931
rect 184 -39965 200 -39931
rect -200 -40012 200 -39965
rect -200 -40259 200 -40212
rect -200 -40293 -184 -40259
rect 184 -40293 200 -40259
rect -200 -40309 200 -40293
rect -200 -40367 200 -40351
rect -200 -40401 -184 -40367
rect 184 -40401 200 -40367
rect -200 -40448 200 -40401
rect -200 -40695 200 -40648
rect -200 -40729 -184 -40695
rect 184 -40729 200 -40695
rect -200 -40745 200 -40729
rect -200 -40803 200 -40787
rect -200 -40837 -184 -40803
rect 184 -40837 200 -40803
rect -200 -40884 200 -40837
rect -200 -41131 200 -41084
rect -200 -41165 -184 -41131
rect 184 -41165 200 -41131
rect -200 -41181 200 -41165
rect -200 -41239 200 -41223
rect -200 -41273 -184 -41239
rect 184 -41273 200 -41239
rect -200 -41320 200 -41273
rect -200 -41567 200 -41520
rect -200 -41601 -184 -41567
rect 184 -41601 200 -41567
rect -200 -41617 200 -41601
rect -200 -41675 200 -41659
rect -200 -41709 -184 -41675
rect 184 -41709 200 -41675
rect -200 -41756 200 -41709
rect -200 -42003 200 -41956
rect -200 -42037 -184 -42003
rect 184 -42037 200 -42003
rect -200 -42053 200 -42037
rect -200 -42111 200 -42095
rect -200 -42145 -184 -42111
rect 184 -42145 200 -42111
rect -200 -42192 200 -42145
rect -200 -42439 200 -42392
rect -200 -42473 -184 -42439
rect 184 -42473 200 -42439
rect -200 -42489 200 -42473
rect -200 -42547 200 -42531
rect -200 -42581 -184 -42547
rect 184 -42581 200 -42547
rect -200 -42628 200 -42581
rect -200 -42875 200 -42828
rect -200 -42909 -184 -42875
rect 184 -42909 200 -42875
rect -200 -42925 200 -42909
rect -200 -42983 200 -42967
rect -200 -43017 -184 -42983
rect 184 -43017 200 -42983
rect -200 -43064 200 -43017
rect -200 -43311 200 -43264
rect -200 -43345 -184 -43311
rect 184 -43345 200 -43311
rect -200 -43361 200 -43345
rect -200 -43419 200 -43403
rect -200 -43453 -184 -43419
rect 184 -43453 200 -43419
rect -200 -43500 200 -43453
rect -200 -43747 200 -43700
rect -200 -43781 -184 -43747
rect 184 -43781 200 -43747
rect -200 -43797 200 -43781
rect -200 -43855 200 -43839
rect -200 -43889 -184 -43855
rect 184 -43889 200 -43855
rect -200 -43936 200 -43889
rect -200 -44183 200 -44136
rect -200 -44217 -184 -44183
rect 184 -44217 200 -44183
rect -200 -44233 200 -44217
rect -200 -44291 200 -44275
rect -200 -44325 -184 -44291
rect 184 -44325 200 -44291
rect -200 -44372 200 -44325
rect -200 -44619 200 -44572
rect -200 -44653 -184 -44619
rect 184 -44653 200 -44619
rect -200 -44669 200 -44653
rect -200 -44727 200 -44711
rect -200 -44761 -184 -44727
rect 184 -44761 200 -44727
rect -200 -44808 200 -44761
rect -200 -45055 200 -45008
rect -200 -45089 -184 -45055
rect 184 -45089 200 -45055
rect -200 -45105 200 -45089
rect -200 -45163 200 -45147
rect -200 -45197 -184 -45163
rect 184 -45197 200 -45163
rect -200 -45244 200 -45197
rect -200 -45491 200 -45444
rect -200 -45525 -184 -45491
rect 184 -45525 200 -45491
rect -200 -45541 200 -45525
rect -200 -45599 200 -45583
rect -200 -45633 -184 -45599
rect 184 -45633 200 -45599
rect -200 -45680 200 -45633
rect -200 -45927 200 -45880
rect -200 -45961 -184 -45927
rect 184 -45961 200 -45927
rect -200 -45977 200 -45961
rect -200 -46035 200 -46019
rect -200 -46069 -184 -46035
rect 184 -46069 200 -46035
rect -200 -46116 200 -46069
rect -200 -46363 200 -46316
rect -200 -46397 -184 -46363
rect 184 -46397 200 -46363
rect -200 -46413 200 -46397
rect -200 -46471 200 -46455
rect -200 -46505 -184 -46471
rect 184 -46505 200 -46471
rect -200 -46552 200 -46505
rect -200 -46799 200 -46752
rect -200 -46833 -184 -46799
rect 184 -46833 200 -46799
rect -200 -46849 200 -46833
rect -200 -46907 200 -46891
rect -200 -46941 -184 -46907
rect 184 -46941 200 -46907
rect -200 -46988 200 -46941
rect -200 -47235 200 -47188
rect -200 -47269 -184 -47235
rect 184 -47269 200 -47235
rect -200 -47285 200 -47269
rect -200 -47343 200 -47327
rect -200 -47377 -184 -47343
rect 184 -47377 200 -47343
rect -200 -47424 200 -47377
rect -200 -47671 200 -47624
rect -200 -47705 -184 -47671
rect 184 -47705 200 -47671
rect -200 -47721 200 -47705
rect -200 -47779 200 -47763
rect -200 -47813 -184 -47779
rect 184 -47813 200 -47779
rect -200 -47860 200 -47813
rect -200 -48107 200 -48060
rect -200 -48141 -184 -48107
rect 184 -48141 200 -48107
rect -200 -48157 200 -48141
rect -200 -48215 200 -48199
rect -200 -48249 -184 -48215
rect 184 -48249 200 -48215
rect -200 -48296 200 -48249
rect -200 -48543 200 -48496
rect -200 -48577 -184 -48543
rect 184 -48577 200 -48543
rect -200 -48593 200 -48577
rect -200 -48651 200 -48635
rect -200 -48685 -184 -48651
rect 184 -48685 200 -48651
rect -200 -48732 200 -48685
rect -200 -48979 200 -48932
rect -200 -49013 -184 -48979
rect 184 -49013 200 -48979
rect -200 -49029 200 -49013
rect -200 -49087 200 -49071
rect -200 -49121 -184 -49087
rect 184 -49121 200 -49087
rect -200 -49168 200 -49121
rect -200 -49415 200 -49368
rect -200 -49449 -184 -49415
rect 184 -49449 200 -49415
rect -200 -49465 200 -49449
rect -200 -49523 200 -49507
rect -200 -49557 -184 -49523
rect 184 -49557 200 -49523
rect -200 -49604 200 -49557
rect -200 -49851 200 -49804
rect -200 -49885 -184 -49851
rect 184 -49885 200 -49851
rect -200 -49901 200 -49885
rect -200 -49959 200 -49943
rect -200 -49993 -184 -49959
rect 184 -49993 200 -49959
rect -200 -50040 200 -49993
rect -200 -50287 200 -50240
rect -200 -50321 -184 -50287
rect 184 -50321 200 -50287
rect -200 -50337 200 -50321
rect -200 -50395 200 -50379
rect -200 -50429 -184 -50395
rect 184 -50429 200 -50395
rect -200 -50476 200 -50429
rect -200 -50723 200 -50676
rect -200 -50757 -184 -50723
rect 184 -50757 200 -50723
rect -200 -50773 200 -50757
rect -200 -50831 200 -50815
rect -200 -50865 -184 -50831
rect 184 -50865 200 -50831
rect -200 -50912 200 -50865
rect -200 -51159 200 -51112
rect -200 -51193 -184 -51159
rect 184 -51193 200 -51159
rect -200 -51209 200 -51193
rect -200 -51267 200 -51251
rect -200 -51301 -184 -51267
rect 184 -51301 200 -51267
rect -200 -51348 200 -51301
rect -200 -51595 200 -51548
rect -200 -51629 -184 -51595
rect 184 -51629 200 -51595
rect -200 -51645 200 -51629
rect -200 -51703 200 -51687
rect -200 -51737 -184 -51703
rect 184 -51737 200 -51703
rect -200 -51784 200 -51737
rect -200 -52031 200 -51984
rect -200 -52065 -184 -52031
rect 184 -52065 200 -52031
rect -200 -52081 200 -52065
rect -200 -52139 200 -52123
rect -200 -52173 -184 -52139
rect 184 -52173 200 -52139
rect -200 -52220 200 -52173
rect -200 -52467 200 -52420
rect -200 -52501 -184 -52467
rect 184 -52501 200 -52467
rect -200 -52517 200 -52501
rect -200 -52575 200 -52559
rect -200 -52609 -184 -52575
rect 184 -52609 200 -52575
rect -200 -52656 200 -52609
rect -200 -52903 200 -52856
rect -200 -52937 -184 -52903
rect 184 -52937 200 -52903
rect -200 -52953 200 -52937
rect -200 -53011 200 -52995
rect -200 -53045 -184 -53011
rect 184 -53045 200 -53011
rect -200 -53092 200 -53045
rect -200 -53339 200 -53292
rect -200 -53373 -184 -53339
rect 184 -53373 200 -53339
rect -200 -53389 200 -53373
rect -200 -53447 200 -53431
rect -200 -53481 -184 -53447
rect 184 -53481 200 -53447
rect -200 -53528 200 -53481
rect -200 -53775 200 -53728
rect -200 -53809 -184 -53775
rect 184 -53809 200 -53775
rect -200 -53825 200 -53809
rect -200 -53883 200 -53867
rect -200 -53917 -184 -53883
rect 184 -53917 200 -53883
rect -200 -53964 200 -53917
rect -200 -54211 200 -54164
rect -200 -54245 -184 -54211
rect 184 -54245 200 -54211
rect -200 -54261 200 -54245
rect -200 -54319 200 -54303
rect -200 -54353 -184 -54319
rect 184 -54353 200 -54319
rect -200 -54400 200 -54353
rect -200 -54647 200 -54600
rect -200 -54681 -184 -54647
rect 184 -54681 200 -54647
rect -200 -54697 200 -54681
rect -200 -54755 200 -54739
rect -200 -54789 -184 -54755
rect 184 -54789 200 -54755
rect -200 -54836 200 -54789
rect -200 -55083 200 -55036
rect -200 -55117 -184 -55083
rect 184 -55117 200 -55083
rect -200 -55133 200 -55117
rect -200 -55191 200 -55175
rect -200 -55225 -184 -55191
rect 184 -55225 200 -55191
rect -200 -55272 200 -55225
rect -200 -55519 200 -55472
rect -200 -55553 -184 -55519
rect 184 -55553 200 -55519
rect -200 -55569 200 -55553
rect -200 -55627 200 -55611
rect -200 -55661 -184 -55627
rect 184 -55661 200 -55627
rect -200 -55708 200 -55661
rect -200 -55955 200 -55908
rect -200 -55989 -184 -55955
rect 184 -55989 200 -55955
rect -200 -56005 200 -55989
rect -200 -56063 200 -56047
rect -200 -56097 -184 -56063
rect 184 -56097 200 -56063
rect -200 -56144 200 -56097
rect -200 -56391 200 -56344
rect -200 -56425 -184 -56391
rect 184 -56425 200 -56391
rect -200 -56441 200 -56425
rect -200 -56499 200 -56483
rect -200 -56533 -184 -56499
rect 184 -56533 200 -56499
rect -200 -56580 200 -56533
rect -200 -56827 200 -56780
rect -200 -56861 -184 -56827
rect 184 -56861 200 -56827
rect -200 -56877 200 -56861
rect -200 -56935 200 -56919
rect -200 -56969 -184 -56935
rect 184 -56969 200 -56935
rect -200 -57016 200 -56969
rect -200 -57263 200 -57216
rect -200 -57297 -184 -57263
rect 184 -57297 200 -57263
rect -200 -57313 200 -57297
rect -200 -57371 200 -57355
rect -200 -57405 -184 -57371
rect 184 -57405 200 -57371
rect -200 -57452 200 -57405
rect -200 -57699 200 -57652
rect -200 -57733 -184 -57699
rect 184 -57733 200 -57699
rect -200 -57749 200 -57733
rect -200 -57807 200 -57791
rect -200 -57841 -184 -57807
rect 184 -57841 200 -57807
rect -200 -57888 200 -57841
rect -200 -58135 200 -58088
rect -200 -58169 -184 -58135
rect 184 -58169 200 -58135
rect -200 -58185 200 -58169
rect -200 -58243 200 -58227
rect -200 -58277 -184 -58243
rect 184 -58277 200 -58243
rect -200 -58324 200 -58277
rect -200 -58571 200 -58524
rect -200 -58605 -184 -58571
rect 184 -58605 200 -58571
rect -200 -58621 200 -58605
rect -200 -58679 200 -58663
rect -200 -58713 -184 -58679
rect 184 -58713 200 -58679
rect -200 -58760 200 -58713
rect -200 -59007 200 -58960
rect -200 -59041 -184 -59007
rect 184 -59041 200 -59007
rect -200 -59057 200 -59041
rect -200 -59115 200 -59099
rect -200 -59149 -184 -59115
rect 184 -59149 200 -59115
rect -200 -59196 200 -59149
rect -200 -59443 200 -59396
rect -200 -59477 -184 -59443
rect 184 -59477 200 -59443
rect -200 -59493 200 -59477
rect -200 -59551 200 -59535
rect -200 -59585 -184 -59551
rect 184 -59585 200 -59551
rect -200 -59632 200 -59585
rect -200 -59879 200 -59832
rect -200 -59913 -184 -59879
rect 184 -59913 200 -59879
rect -200 -59929 200 -59913
rect -200 -59987 200 -59971
rect -200 -60021 -184 -59987
rect 184 -60021 200 -59987
rect -200 -60068 200 -60021
rect -200 -60315 200 -60268
rect -200 -60349 -184 -60315
rect 184 -60349 200 -60315
rect -200 -60365 200 -60349
rect -200 -60423 200 -60407
rect -200 -60457 -184 -60423
rect 184 -60457 200 -60423
rect -200 -60504 200 -60457
rect -200 -60751 200 -60704
rect -200 -60785 -184 -60751
rect 184 -60785 200 -60751
rect -200 -60801 200 -60785
rect -200 -60859 200 -60843
rect -200 -60893 -184 -60859
rect 184 -60893 200 -60859
rect -200 -60940 200 -60893
rect -200 -61187 200 -61140
rect -200 -61221 -184 -61187
rect 184 -61221 200 -61187
rect -200 -61237 200 -61221
rect -200 -61295 200 -61279
rect -200 -61329 -184 -61295
rect 184 -61329 200 -61295
rect -200 -61376 200 -61329
rect -200 -61623 200 -61576
rect -200 -61657 -184 -61623
rect 184 -61657 200 -61623
rect -200 -61673 200 -61657
rect -200 -61731 200 -61715
rect -200 -61765 -184 -61731
rect 184 -61765 200 -61731
rect -200 -61812 200 -61765
rect -200 -62059 200 -62012
rect -200 -62093 -184 -62059
rect 184 -62093 200 -62059
rect -200 -62109 200 -62093
rect -200 -62167 200 -62151
rect -200 -62201 -184 -62167
rect 184 -62201 200 -62167
rect -200 -62248 200 -62201
rect -200 -62495 200 -62448
rect -200 -62529 -184 -62495
rect 184 -62529 200 -62495
rect -200 -62545 200 -62529
rect -200 -62603 200 -62587
rect -200 -62637 -184 -62603
rect 184 -62637 200 -62603
rect -200 -62684 200 -62637
rect -200 -62931 200 -62884
rect -200 -62965 -184 -62931
rect 184 -62965 200 -62931
rect -200 -62981 200 -62965
rect -200 -63039 200 -63023
rect -200 -63073 -184 -63039
rect 184 -63073 200 -63039
rect -200 -63120 200 -63073
rect -200 -63367 200 -63320
rect -200 -63401 -184 -63367
rect 184 -63401 200 -63367
rect -200 -63417 200 -63401
rect -200 -63475 200 -63459
rect -200 -63509 -184 -63475
rect 184 -63509 200 -63475
rect -200 -63556 200 -63509
rect -200 -63803 200 -63756
rect -200 -63837 -184 -63803
rect 184 -63837 200 -63803
rect -200 -63853 200 -63837
rect -200 -63911 200 -63895
rect -200 -63945 -184 -63911
rect 184 -63945 200 -63911
rect -200 -63992 200 -63945
rect -200 -64239 200 -64192
rect -200 -64273 -184 -64239
rect 184 -64273 200 -64239
rect -200 -64289 200 -64273
rect -200 -64347 200 -64331
rect -200 -64381 -184 -64347
rect 184 -64381 200 -64347
rect -200 -64428 200 -64381
rect -200 -64675 200 -64628
rect -200 -64709 -184 -64675
rect 184 -64709 200 -64675
rect -200 -64725 200 -64709
rect -200 -64783 200 -64767
rect -200 -64817 -184 -64783
rect 184 -64817 200 -64783
rect -200 -64864 200 -64817
rect -200 -65111 200 -65064
rect -200 -65145 -184 -65111
rect 184 -65145 200 -65111
rect -200 -65161 200 -65145
rect -200 -65219 200 -65203
rect -200 -65253 -184 -65219
rect 184 -65253 200 -65219
rect -200 -65300 200 -65253
rect -200 -65547 200 -65500
rect -200 -65581 -184 -65547
rect 184 -65581 200 -65547
rect -200 -65597 200 -65581
rect -200 -65655 200 -65639
rect -200 -65689 -184 -65655
rect 184 -65689 200 -65655
rect -200 -65736 200 -65689
rect -200 -65983 200 -65936
rect -200 -66017 -184 -65983
rect 184 -66017 200 -65983
rect -200 -66033 200 -66017
rect -200 -66091 200 -66075
rect -200 -66125 -184 -66091
rect 184 -66125 200 -66091
rect -200 -66172 200 -66125
rect -200 -66419 200 -66372
rect -200 -66453 -184 -66419
rect 184 -66453 200 -66419
rect -200 -66469 200 -66453
rect -200 -66527 200 -66511
rect -200 -66561 -184 -66527
rect 184 -66561 200 -66527
rect -200 -66608 200 -66561
rect -200 -66855 200 -66808
rect -200 -66889 -184 -66855
rect 184 -66889 200 -66855
rect -200 -66905 200 -66889
rect -200 -66963 200 -66947
rect -200 -66997 -184 -66963
rect 184 -66997 200 -66963
rect -200 -67044 200 -66997
rect -200 -67291 200 -67244
rect -200 -67325 -184 -67291
rect 184 -67325 200 -67291
rect -200 -67341 200 -67325
rect -200 -67399 200 -67383
rect -200 -67433 -184 -67399
rect 184 -67433 200 -67399
rect -200 -67480 200 -67433
rect -200 -67727 200 -67680
rect -200 -67761 -184 -67727
rect 184 -67761 200 -67727
rect -200 -67777 200 -67761
rect -200 -67835 200 -67819
rect -200 -67869 -184 -67835
rect 184 -67869 200 -67835
rect -200 -67916 200 -67869
rect -200 -68163 200 -68116
rect -200 -68197 -184 -68163
rect 184 -68197 200 -68163
rect -200 -68213 200 -68197
rect -200 -68271 200 -68255
rect -200 -68305 -184 -68271
rect 184 -68305 200 -68271
rect -200 -68352 200 -68305
rect -200 -68599 200 -68552
rect -200 -68633 -184 -68599
rect 184 -68633 200 -68599
rect -200 -68649 200 -68633
rect -200 -68707 200 -68691
rect -200 -68741 -184 -68707
rect 184 -68741 200 -68707
rect -200 -68788 200 -68741
rect -200 -69035 200 -68988
rect -200 -69069 -184 -69035
rect 184 -69069 200 -69035
rect -200 -69085 200 -69069
rect -200 -69143 200 -69127
rect -200 -69177 -184 -69143
rect 184 -69177 200 -69143
rect -200 -69224 200 -69177
rect -200 -69471 200 -69424
rect -200 -69505 -184 -69471
rect 184 -69505 200 -69471
rect -200 -69521 200 -69505
rect -200 -69579 200 -69563
rect -200 -69613 -184 -69579
rect 184 -69613 200 -69579
rect -200 -69660 200 -69613
rect -200 -69907 200 -69860
rect -200 -69941 -184 -69907
rect 184 -69941 200 -69907
rect -200 -69957 200 -69941
rect -200 -70015 200 -69999
rect -200 -70049 -184 -70015
rect 184 -70049 200 -70015
rect -200 -70096 200 -70049
rect -200 -70343 200 -70296
rect -200 -70377 -184 -70343
rect 184 -70377 200 -70343
rect -200 -70393 200 -70377
rect -200 -70451 200 -70435
rect -200 -70485 -184 -70451
rect 184 -70485 200 -70451
rect -200 -70532 200 -70485
rect -200 -70779 200 -70732
rect -200 -70813 -184 -70779
rect 184 -70813 200 -70779
rect -200 -70829 200 -70813
rect -200 -70887 200 -70871
rect -200 -70921 -184 -70887
rect 184 -70921 200 -70887
rect -200 -70968 200 -70921
rect -200 -71215 200 -71168
rect -200 -71249 -184 -71215
rect 184 -71249 200 -71215
rect -200 -71265 200 -71249
rect -200 -71323 200 -71307
rect -200 -71357 -184 -71323
rect 184 -71357 200 -71323
rect -200 -71404 200 -71357
rect -200 -71651 200 -71604
rect -200 -71685 -184 -71651
rect 184 -71685 200 -71651
rect -200 -71701 200 -71685
rect -200 -71759 200 -71743
rect -200 -71793 -184 -71759
rect 184 -71793 200 -71759
rect -200 -71840 200 -71793
rect -200 -72087 200 -72040
rect -200 -72121 -184 -72087
rect 184 -72121 200 -72087
rect -200 -72137 200 -72121
rect -200 -72195 200 -72179
rect -200 -72229 -184 -72195
rect 184 -72229 200 -72195
rect -200 -72276 200 -72229
rect -200 -72523 200 -72476
rect -200 -72557 -184 -72523
rect 184 -72557 200 -72523
rect -200 -72573 200 -72557
rect -200 -72631 200 -72615
rect -200 -72665 -184 -72631
rect 184 -72665 200 -72631
rect -200 -72712 200 -72665
rect -200 -72959 200 -72912
rect -200 -72993 -184 -72959
rect 184 -72993 200 -72959
rect -200 -73009 200 -72993
rect -200 -73067 200 -73051
rect -200 -73101 -184 -73067
rect 184 -73101 200 -73067
rect -200 -73148 200 -73101
rect -200 -73395 200 -73348
rect -200 -73429 -184 -73395
rect 184 -73429 200 -73395
rect -200 -73445 200 -73429
rect -200 -73503 200 -73487
rect -200 -73537 -184 -73503
rect 184 -73537 200 -73503
rect -200 -73584 200 -73537
rect -200 -73831 200 -73784
rect -200 -73865 -184 -73831
rect 184 -73865 200 -73831
rect -200 -73881 200 -73865
rect -200 -73939 200 -73923
rect -200 -73973 -184 -73939
rect 184 -73973 200 -73939
rect -200 -74020 200 -73973
rect -200 -74267 200 -74220
rect -200 -74301 -184 -74267
rect 184 -74301 200 -74267
rect -200 -74317 200 -74301
rect -200 -74375 200 -74359
rect -200 -74409 -184 -74375
rect 184 -74409 200 -74375
rect -200 -74456 200 -74409
rect -200 -74703 200 -74656
rect -200 -74737 -184 -74703
rect 184 -74737 200 -74703
rect -200 -74753 200 -74737
rect -200 -74811 200 -74795
rect -200 -74845 -184 -74811
rect 184 -74845 200 -74811
rect -200 -74892 200 -74845
rect -200 -75139 200 -75092
rect -200 -75173 -184 -75139
rect 184 -75173 200 -75139
rect -200 -75189 200 -75173
rect -200 -75247 200 -75231
rect -200 -75281 -184 -75247
rect 184 -75281 200 -75247
rect -200 -75328 200 -75281
rect -200 -75575 200 -75528
rect -200 -75609 -184 -75575
rect 184 -75609 200 -75575
rect -200 -75625 200 -75609
rect -200 -75683 200 -75667
rect -200 -75717 -184 -75683
rect 184 -75717 200 -75683
rect -200 -75764 200 -75717
rect -200 -76011 200 -75964
rect -200 -76045 -184 -76011
rect 184 -76045 200 -76011
rect -200 -76061 200 -76045
rect -200 -76119 200 -76103
rect -200 -76153 -184 -76119
rect 184 -76153 200 -76119
rect -200 -76200 200 -76153
rect -200 -76447 200 -76400
rect -200 -76481 -184 -76447
rect 184 -76481 200 -76447
rect -200 -76497 200 -76481
rect -200 -76555 200 -76539
rect -200 -76589 -184 -76555
rect 184 -76589 200 -76555
rect -200 -76636 200 -76589
rect -200 -76883 200 -76836
rect -200 -76917 -184 -76883
rect 184 -76917 200 -76883
rect -200 -76933 200 -76917
rect -200 -76991 200 -76975
rect -200 -77025 -184 -76991
rect 184 -77025 200 -76991
rect -200 -77072 200 -77025
rect -200 -77319 200 -77272
rect -200 -77353 -184 -77319
rect 184 -77353 200 -77319
rect -200 -77369 200 -77353
rect -200 -77427 200 -77411
rect -200 -77461 -184 -77427
rect 184 -77461 200 -77427
rect -200 -77508 200 -77461
rect -200 -77755 200 -77708
rect -200 -77789 -184 -77755
rect 184 -77789 200 -77755
rect -200 -77805 200 -77789
rect -200 -77863 200 -77847
rect -200 -77897 -184 -77863
rect 184 -77897 200 -77863
rect -200 -77944 200 -77897
rect -200 -78191 200 -78144
rect -200 -78225 -184 -78191
rect 184 -78225 200 -78191
rect -200 -78241 200 -78225
rect -200 -78299 200 -78283
rect -200 -78333 -184 -78299
rect 184 -78333 200 -78299
rect -200 -78380 200 -78333
rect -200 -78627 200 -78580
rect -200 -78661 -184 -78627
rect 184 -78661 200 -78627
rect -200 -78677 200 -78661
rect -200 -78735 200 -78719
rect -200 -78769 -184 -78735
rect 184 -78769 200 -78735
rect -200 -78816 200 -78769
rect -200 -79063 200 -79016
rect -200 -79097 -184 -79063
rect 184 -79097 200 -79063
rect -200 -79113 200 -79097
rect -200 -79171 200 -79155
rect -200 -79205 -184 -79171
rect 184 -79205 200 -79171
rect -200 -79252 200 -79205
rect -200 -79499 200 -79452
rect -200 -79533 -184 -79499
rect 184 -79533 200 -79499
rect -200 -79549 200 -79533
rect -200 -79607 200 -79591
rect -200 -79641 -184 -79607
rect 184 -79641 200 -79607
rect -200 -79688 200 -79641
rect -200 -79935 200 -79888
rect -200 -79969 -184 -79935
rect 184 -79969 200 -79935
rect -200 -79985 200 -79969
rect -200 -80043 200 -80027
rect -200 -80077 -184 -80043
rect 184 -80077 200 -80043
rect -200 -80124 200 -80077
rect -200 -80371 200 -80324
rect -200 -80405 -184 -80371
rect 184 -80405 200 -80371
rect -200 -80421 200 -80405
rect -200 -80479 200 -80463
rect -200 -80513 -184 -80479
rect 184 -80513 200 -80479
rect -200 -80560 200 -80513
rect -200 -80807 200 -80760
rect -200 -80841 -184 -80807
rect 184 -80841 200 -80807
rect -200 -80857 200 -80841
rect -200 -80915 200 -80899
rect -200 -80949 -184 -80915
rect 184 -80949 200 -80915
rect -200 -80996 200 -80949
rect -200 -81243 200 -81196
rect -200 -81277 -184 -81243
rect 184 -81277 200 -81243
rect -200 -81293 200 -81277
rect -200 -81351 200 -81335
rect -200 -81385 -184 -81351
rect 184 -81385 200 -81351
rect -200 -81432 200 -81385
rect -200 -81679 200 -81632
rect -200 -81713 -184 -81679
rect 184 -81713 200 -81679
rect -200 -81729 200 -81713
rect -200 -81787 200 -81771
rect -200 -81821 -184 -81787
rect 184 -81821 200 -81787
rect -200 -81868 200 -81821
rect -200 -82115 200 -82068
rect -200 -82149 -184 -82115
rect 184 -82149 200 -82115
rect -200 -82165 200 -82149
rect -200 -82223 200 -82207
rect -200 -82257 -184 -82223
rect 184 -82257 200 -82223
rect -200 -82304 200 -82257
rect -200 -82551 200 -82504
rect -200 -82585 -184 -82551
rect 184 -82585 200 -82551
rect -200 -82601 200 -82585
rect -200 -82659 200 -82643
rect -200 -82693 -184 -82659
rect 184 -82693 200 -82659
rect -200 -82740 200 -82693
rect -200 -82987 200 -82940
rect -200 -83021 -184 -82987
rect 184 -83021 200 -82987
rect -200 -83037 200 -83021
rect -200 -83095 200 -83079
rect -200 -83129 -184 -83095
rect 184 -83129 200 -83095
rect -200 -83176 200 -83129
rect -200 -83423 200 -83376
rect -200 -83457 -184 -83423
rect 184 -83457 200 -83423
rect -200 -83473 200 -83457
rect -200 -83531 200 -83515
rect -200 -83565 -184 -83531
rect 184 -83565 200 -83531
rect -200 -83612 200 -83565
rect -200 -83859 200 -83812
rect -200 -83893 -184 -83859
rect 184 -83893 200 -83859
rect -200 -83909 200 -83893
rect -200 -83967 200 -83951
rect -200 -84001 -184 -83967
rect 184 -84001 200 -83967
rect -200 -84048 200 -84001
rect -200 -84295 200 -84248
rect -200 -84329 -184 -84295
rect 184 -84329 200 -84295
rect -200 -84345 200 -84329
<< polycont >>
rect -184 84295 184 84329
rect -184 83967 184 84001
rect -184 83859 184 83893
rect -184 83531 184 83565
rect -184 83423 184 83457
rect -184 83095 184 83129
rect -184 82987 184 83021
rect -184 82659 184 82693
rect -184 82551 184 82585
rect -184 82223 184 82257
rect -184 82115 184 82149
rect -184 81787 184 81821
rect -184 81679 184 81713
rect -184 81351 184 81385
rect -184 81243 184 81277
rect -184 80915 184 80949
rect -184 80807 184 80841
rect -184 80479 184 80513
rect -184 80371 184 80405
rect -184 80043 184 80077
rect -184 79935 184 79969
rect -184 79607 184 79641
rect -184 79499 184 79533
rect -184 79171 184 79205
rect -184 79063 184 79097
rect -184 78735 184 78769
rect -184 78627 184 78661
rect -184 78299 184 78333
rect -184 78191 184 78225
rect -184 77863 184 77897
rect -184 77755 184 77789
rect -184 77427 184 77461
rect -184 77319 184 77353
rect -184 76991 184 77025
rect -184 76883 184 76917
rect -184 76555 184 76589
rect -184 76447 184 76481
rect -184 76119 184 76153
rect -184 76011 184 76045
rect -184 75683 184 75717
rect -184 75575 184 75609
rect -184 75247 184 75281
rect -184 75139 184 75173
rect -184 74811 184 74845
rect -184 74703 184 74737
rect -184 74375 184 74409
rect -184 74267 184 74301
rect -184 73939 184 73973
rect -184 73831 184 73865
rect -184 73503 184 73537
rect -184 73395 184 73429
rect -184 73067 184 73101
rect -184 72959 184 72993
rect -184 72631 184 72665
rect -184 72523 184 72557
rect -184 72195 184 72229
rect -184 72087 184 72121
rect -184 71759 184 71793
rect -184 71651 184 71685
rect -184 71323 184 71357
rect -184 71215 184 71249
rect -184 70887 184 70921
rect -184 70779 184 70813
rect -184 70451 184 70485
rect -184 70343 184 70377
rect -184 70015 184 70049
rect -184 69907 184 69941
rect -184 69579 184 69613
rect -184 69471 184 69505
rect -184 69143 184 69177
rect -184 69035 184 69069
rect -184 68707 184 68741
rect -184 68599 184 68633
rect -184 68271 184 68305
rect -184 68163 184 68197
rect -184 67835 184 67869
rect -184 67727 184 67761
rect -184 67399 184 67433
rect -184 67291 184 67325
rect -184 66963 184 66997
rect -184 66855 184 66889
rect -184 66527 184 66561
rect -184 66419 184 66453
rect -184 66091 184 66125
rect -184 65983 184 66017
rect -184 65655 184 65689
rect -184 65547 184 65581
rect -184 65219 184 65253
rect -184 65111 184 65145
rect -184 64783 184 64817
rect -184 64675 184 64709
rect -184 64347 184 64381
rect -184 64239 184 64273
rect -184 63911 184 63945
rect -184 63803 184 63837
rect -184 63475 184 63509
rect -184 63367 184 63401
rect -184 63039 184 63073
rect -184 62931 184 62965
rect -184 62603 184 62637
rect -184 62495 184 62529
rect -184 62167 184 62201
rect -184 62059 184 62093
rect -184 61731 184 61765
rect -184 61623 184 61657
rect -184 61295 184 61329
rect -184 61187 184 61221
rect -184 60859 184 60893
rect -184 60751 184 60785
rect -184 60423 184 60457
rect -184 60315 184 60349
rect -184 59987 184 60021
rect -184 59879 184 59913
rect -184 59551 184 59585
rect -184 59443 184 59477
rect -184 59115 184 59149
rect -184 59007 184 59041
rect -184 58679 184 58713
rect -184 58571 184 58605
rect -184 58243 184 58277
rect -184 58135 184 58169
rect -184 57807 184 57841
rect -184 57699 184 57733
rect -184 57371 184 57405
rect -184 57263 184 57297
rect -184 56935 184 56969
rect -184 56827 184 56861
rect -184 56499 184 56533
rect -184 56391 184 56425
rect -184 56063 184 56097
rect -184 55955 184 55989
rect -184 55627 184 55661
rect -184 55519 184 55553
rect -184 55191 184 55225
rect -184 55083 184 55117
rect -184 54755 184 54789
rect -184 54647 184 54681
rect -184 54319 184 54353
rect -184 54211 184 54245
rect -184 53883 184 53917
rect -184 53775 184 53809
rect -184 53447 184 53481
rect -184 53339 184 53373
rect -184 53011 184 53045
rect -184 52903 184 52937
rect -184 52575 184 52609
rect -184 52467 184 52501
rect -184 52139 184 52173
rect -184 52031 184 52065
rect -184 51703 184 51737
rect -184 51595 184 51629
rect -184 51267 184 51301
rect -184 51159 184 51193
rect -184 50831 184 50865
rect -184 50723 184 50757
rect -184 50395 184 50429
rect -184 50287 184 50321
rect -184 49959 184 49993
rect -184 49851 184 49885
rect -184 49523 184 49557
rect -184 49415 184 49449
rect -184 49087 184 49121
rect -184 48979 184 49013
rect -184 48651 184 48685
rect -184 48543 184 48577
rect -184 48215 184 48249
rect -184 48107 184 48141
rect -184 47779 184 47813
rect -184 47671 184 47705
rect -184 47343 184 47377
rect -184 47235 184 47269
rect -184 46907 184 46941
rect -184 46799 184 46833
rect -184 46471 184 46505
rect -184 46363 184 46397
rect -184 46035 184 46069
rect -184 45927 184 45961
rect -184 45599 184 45633
rect -184 45491 184 45525
rect -184 45163 184 45197
rect -184 45055 184 45089
rect -184 44727 184 44761
rect -184 44619 184 44653
rect -184 44291 184 44325
rect -184 44183 184 44217
rect -184 43855 184 43889
rect -184 43747 184 43781
rect -184 43419 184 43453
rect -184 43311 184 43345
rect -184 42983 184 43017
rect -184 42875 184 42909
rect -184 42547 184 42581
rect -184 42439 184 42473
rect -184 42111 184 42145
rect -184 42003 184 42037
rect -184 41675 184 41709
rect -184 41567 184 41601
rect -184 41239 184 41273
rect -184 41131 184 41165
rect -184 40803 184 40837
rect -184 40695 184 40729
rect -184 40367 184 40401
rect -184 40259 184 40293
rect -184 39931 184 39965
rect -184 39823 184 39857
rect -184 39495 184 39529
rect -184 39387 184 39421
rect -184 39059 184 39093
rect -184 38951 184 38985
rect -184 38623 184 38657
rect -184 38515 184 38549
rect -184 38187 184 38221
rect -184 38079 184 38113
rect -184 37751 184 37785
rect -184 37643 184 37677
rect -184 37315 184 37349
rect -184 37207 184 37241
rect -184 36879 184 36913
rect -184 36771 184 36805
rect -184 36443 184 36477
rect -184 36335 184 36369
rect -184 36007 184 36041
rect -184 35899 184 35933
rect -184 35571 184 35605
rect -184 35463 184 35497
rect -184 35135 184 35169
rect -184 35027 184 35061
rect -184 34699 184 34733
rect -184 34591 184 34625
rect -184 34263 184 34297
rect -184 34155 184 34189
rect -184 33827 184 33861
rect -184 33719 184 33753
rect -184 33391 184 33425
rect -184 33283 184 33317
rect -184 32955 184 32989
rect -184 32847 184 32881
rect -184 32519 184 32553
rect -184 32411 184 32445
rect -184 32083 184 32117
rect -184 31975 184 32009
rect -184 31647 184 31681
rect -184 31539 184 31573
rect -184 31211 184 31245
rect -184 31103 184 31137
rect -184 30775 184 30809
rect -184 30667 184 30701
rect -184 30339 184 30373
rect -184 30231 184 30265
rect -184 29903 184 29937
rect -184 29795 184 29829
rect -184 29467 184 29501
rect -184 29359 184 29393
rect -184 29031 184 29065
rect -184 28923 184 28957
rect -184 28595 184 28629
rect -184 28487 184 28521
rect -184 28159 184 28193
rect -184 28051 184 28085
rect -184 27723 184 27757
rect -184 27615 184 27649
rect -184 27287 184 27321
rect -184 27179 184 27213
rect -184 26851 184 26885
rect -184 26743 184 26777
rect -184 26415 184 26449
rect -184 26307 184 26341
rect -184 25979 184 26013
rect -184 25871 184 25905
rect -184 25543 184 25577
rect -184 25435 184 25469
rect -184 25107 184 25141
rect -184 24999 184 25033
rect -184 24671 184 24705
rect -184 24563 184 24597
rect -184 24235 184 24269
rect -184 24127 184 24161
rect -184 23799 184 23833
rect -184 23691 184 23725
rect -184 23363 184 23397
rect -184 23255 184 23289
rect -184 22927 184 22961
rect -184 22819 184 22853
rect -184 22491 184 22525
rect -184 22383 184 22417
rect -184 22055 184 22089
rect -184 21947 184 21981
rect -184 21619 184 21653
rect -184 21511 184 21545
rect -184 21183 184 21217
rect -184 21075 184 21109
rect -184 20747 184 20781
rect -184 20639 184 20673
rect -184 20311 184 20345
rect -184 20203 184 20237
rect -184 19875 184 19909
rect -184 19767 184 19801
rect -184 19439 184 19473
rect -184 19331 184 19365
rect -184 19003 184 19037
rect -184 18895 184 18929
rect -184 18567 184 18601
rect -184 18459 184 18493
rect -184 18131 184 18165
rect -184 18023 184 18057
rect -184 17695 184 17729
rect -184 17587 184 17621
rect -184 17259 184 17293
rect -184 17151 184 17185
rect -184 16823 184 16857
rect -184 16715 184 16749
rect -184 16387 184 16421
rect -184 16279 184 16313
rect -184 15951 184 15985
rect -184 15843 184 15877
rect -184 15515 184 15549
rect -184 15407 184 15441
rect -184 15079 184 15113
rect -184 14971 184 15005
rect -184 14643 184 14677
rect -184 14535 184 14569
rect -184 14207 184 14241
rect -184 14099 184 14133
rect -184 13771 184 13805
rect -184 13663 184 13697
rect -184 13335 184 13369
rect -184 13227 184 13261
rect -184 12899 184 12933
rect -184 12791 184 12825
rect -184 12463 184 12497
rect -184 12355 184 12389
rect -184 12027 184 12061
rect -184 11919 184 11953
rect -184 11591 184 11625
rect -184 11483 184 11517
rect -184 11155 184 11189
rect -184 11047 184 11081
rect -184 10719 184 10753
rect -184 10611 184 10645
rect -184 10283 184 10317
rect -184 10175 184 10209
rect -184 9847 184 9881
rect -184 9739 184 9773
rect -184 9411 184 9445
rect -184 9303 184 9337
rect -184 8975 184 9009
rect -184 8867 184 8901
rect -184 8539 184 8573
rect -184 8431 184 8465
rect -184 8103 184 8137
rect -184 7995 184 8029
rect -184 7667 184 7701
rect -184 7559 184 7593
rect -184 7231 184 7265
rect -184 7123 184 7157
rect -184 6795 184 6829
rect -184 6687 184 6721
rect -184 6359 184 6393
rect -184 6251 184 6285
rect -184 5923 184 5957
rect -184 5815 184 5849
rect -184 5487 184 5521
rect -184 5379 184 5413
rect -184 5051 184 5085
rect -184 4943 184 4977
rect -184 4615 184 4649
rect -184 4507 184 4541
rect -184 4179 184 4213
rect -184 4071 184 4105
rect -184 3743 184 3777
rect -184 3635 184 3669
rect -184 3307 184 3341
rect -184 3199 184 3233
rect -184 2871 184 2905
rect -184 2763 184 2797
rect -184 2435 184 2469
rect -184 2327 184 2361
rect -184 1999 184 2033
rect -184 1891 184 1925
rect -184 1563 184 1597
rect -184 1455 184 1489
rect -184 1127 184 1161
rect -184 1019 184 1053
rect -184 691 184 725
rect -184 583 184 617
rect -184 255 184 289
rect -184 147 184 181
rect -184 -181 184 -147
rect -184 -289 184 -255
rect -184 -617 184 -583
rect -184 -725 184 -691
rect -184 -1053 184 -1019
rect -184 -1161 184 -1127
rect -184 -1489 184 -1455
rect -184 -1597 184 -1563
rect -184 -1925 184 -1891
rect -184 -2033 184 -1999
rect -184 -2361 184 -2327
rect -184 -2469 184 -2435
rect -184 -2797 184 -2763
rect -184 -2905 184 -2871
rect -184 -3233 184 -3199
rect -184 -3341 184 -3307
rect -184 -3669 184 -3635
rect -184 -3777 184 -3743
rect -184 -4105 184 -4071
rect -184 -4213 184 -4179
rect -184 -4541 184 -4507
rect -184 -4649 184 -4615
rect -184 -4977 184 -4943
rect -184 -5085 184 -5051
rect -184 -5413 184 -5379
rect -184 -5521 184 -5487
rect -184 -5849 184 -5815
rect -184 -5957 184 -5923
rect -184 -6285 184 -6251
rect -184 -6393 184 -6359
rect -184 -6721 184 -6687
rect -184 -6829 184 -6795
rect -184 -7157 184 -7123
rect -184 -7265 184 -7231
rect -184 -7593 184 -7559
rect -184 -7701 184 -7667
rect -184 -8029 184 -7995
rect -184 -8137 184 -8103
rect -184 -8465 184 -8431
rect -184 -8573 184 -8539
rect -184 -8901 184 -8867
rect -184 -9009 184 -8975
rect -184 -9337 184 -9303
rect -184 -9445 184 -9411
rect -184 -9773 184 -9739
rect -184 -9881 184 -9847
rect -184 -10209 184 -10175
rect -184 -10317 184 -10283
rect -184 -10645 184 -10611
rect -184 -10753 184 -10719
rect -184 -11081 184 -11047
rect -184 -11189 184 -11155
rect -184 -11517 184 -11483
rect -184 -11625 184 -11591
rect -184 -11953 184 -11919
rect -184 -12061 184 -12027
rect -184 -12389 184 -12355
rect -184 -12497 184 -12463
rect -184 -12825 184 -12791
rect -184 -12933 184 -12899
rect -184 -13261 184 -13227
rect -184 -13369 184 -13335
rect -184 -13697 184 -13663
rect -184 -13805 184 -13771
rect -184 -14133 184 -14099
rect -184 -14241 184 -14207
rect -184 -14569 184 -14535
rect -184 -14677 184 -14643
rect -184 -15005 184 -14971
rect -184 -15113 184 -15079
rect -184 -15441 184 -15407
rect -184 -15549 184 -15515
rect -184 -15877 184 -15843
rect -184 -15985 184 -15951
rect -184 -16313 184 -16279
rect -184 -16421 184 -16387
rect -184 -16749 184 -16715
rect -184 -16857 184 -16823
rect -184 -17185 184 -17151
rect -184 -17293 184 -17259
rect -184 -17621 184 -17587
rect -184 -17729 184 -17695
rect -184 -18057 184 -18023
rect -184 -18165 184 -18131
rect -184 -18493 184 -18459
rect -184 -18601 184 -18567
rect -184 -18929 184 -18895
rect -184 -19037 184 -19003
rect -184 -19365 184 -19331
rect -184 -19473 184 -19439
rect -184 -19801 184 -19767
rect -184 -19909 184 -19875
rect -184 -20237 184 -20203
rect -184 -20345 184 -20311
rect -184 -20673 184 -20639
rect -184 -20781 184 -20747
rect -184 -21109 184 -21075
rect -184 -21217 184 -21183
rect -184 -21545 184 -21511
rect -184 -21653 184 -21619
rect -184 -21981 184 -21947
rect -184 -22089 184 -22055
rect -184 -22417 184 -22383
rect -184 -22525 184 -22491
rect -184 -22853 184 -22819
rect -184 -22961 184 -22927
rect -184 -23289 184 -23255
rect -184 -23397 184 -23363
rect -184 -23725 184 -23691
rect -184 -23833 184 -23799
rect -184 -24161 184 -24127
rect -184 -24269 184 -24235
rect -184 -24597 184 -24563
rect -184 -24705 184 -24671
rect -184 -25033 184 -24999
rect -184 -25141 184 -25107
rect -184 -25469 184 -25435
rect -184 -25577 184 -25543
rect -184 -25905 184 -25871
rect -184 -26013 184 -25979
rect -184 -26341 184 -26307
rect -184 -26449 184 -26415
rect -184 -26777 184 -26743
rect -184 -26885 184 -26851
rect -184 -27213 184 -27179
rect -184 -27321 184 -27287
rect -184 -27649 184 -27615
rect -184 -27757 184 -27723
rect -184 -28085 184 -28051
rect -184 -28193 184 -28159
rect -184 -28521 184 -28487
rect -184 -28629 184 -28595
rect -184 -28957 184 -28923
rect -184 -29065 184 -29031
rect -184 -29393 184 -29359
rect -184 -29501 184 -29467
rect -184 -29829 184 -29795
rect -184 -29937 184 -29903
rect -184 -30265 184 -30231
rect -184 -30373 184 -30339
rect -184 -30701 184 -30667
rect -184 -30809 184 -30775
rect -184 -31137 184 -31103
rect -184 -31245 184 -31211
rect -184 -31573 184 -31539
rect -184 -31681 184 -31647
rect -184 -32009 184 -31975
rect -184 -32117 184 -32083
rect -184 -32445 184 -32411
rect -184 -32553 184 -32519
rect -184 -32881 184 -32847
rect -184 -32989 184 -32955
rect -184 -33317 184 -33283
rect -184 -33425 184 -33391
rect -184 -33753 184 -33719
rect -184 -33861 184 -33827
rect -184 -34189 184 -34155
rect -184 -34297 184 -34263
rect -184 -34625 184 -34591
rect -184 -34733 184 -34699
rect -184 -35061 184 -35027
rect -184 -35169 184 -35135
rect -184 -35497 184 -35463
rect -184 -35605 184 -35571
rect -184 -35933 184 -35899
rect -184 -36041 184 -36007
rect -184 -36369 184 -36335
rect -184 -36477 184 -36443
rect -184 -36805 184 -36771
rect -184 -36913 184 -36879
rect -184 -37241 184 -37207
rect -184 -37349 184 -37315
rect -184 -37677 184 -37643
rect -184 -37785 184 -37751
rect -184 -38113 184 -38079
rect -184 -38221 184 -38187
rect -184 -38549 184 -38515
rect -184 -38657 184 -38623
rect -184 -38985 184 -38951
rect -184 -39093 184 -39059
rect -184 -39421 184 -39387
rect -184 -39529 184 -39495
rect -184 -39857 184 -39823
rect -184 -39965 184 -39931
rect -184 -40293 184 -40259
rect -184 -40401 184 -40367
rect -184 -40729 184 -40695
rect -184 -40837 184 -40803
rect -184 -41165 184 -41131
rect -184 -41273 184 -41239
rect -184 -41601 184 -41567
rect -184 -41709 184 -41675
rect -184 -42037 184 -42003
rect -184 -42145 184 -42111
rect -184 -42473 184 -42439
rect -184 -42581 184 -42547
rect -184 -42909 184 -42875
rect -184 -43017 184 -42983
rect -184 -43345 184 -43311
rect -184 -43453 184 -43419
rect -184 -43781 184 -43747
rect -184 -43889 184 -43855
rect -184 -44217 184 -44183
rect -184 -44325 184 -44291
rect -184 -44653 184 -44619
rect -184 -44761 184 -44727
rect -184 -45089 184 -45055
rect -184 -45197 184 -45163
rect -184 -45525 184 -45491
rect -184 -45633 184 -45599
rect -184 -45961 184 -45927
rect -184 -46069 184 -46035
rect -184 -46397 184 -46363
rect -184 -46505 184 -46471
rect -184 -46833 184 -46799
rect -184 -46941 184 -46907
rect -184 -47269 184 -47235
rect -184 -47377 184 -47343
rect -184 -47705 184 -47671
rect -184 -47813 184 -47779
rect -184 -48141 184 -48107
rect -184 -48249 184 -48215
rect -184 -48577 184 -48543
rect -184 -48685 184 -48651
rect -184 -49013 184 -48979
rect -184 -49121 184 -49087
rect -184 -49449 184 -49415
rect -184 -49557 184 -49523
rect -184 -49885 184 -49851
rect -184 -49993 184 -49959
rect -184 -50321 184 -50287
rect -184 -50429 184 -50395
rect -184 -50757 184 -50723
rect -184 -50865 184 -50831
rect -184 -51193 184 -51159
rect -184 -51301 184 -51267
rect -184 -51629 184 -51595
rect -184 -51737 184 -51703
rect -184 -52065 184 -52031
rect -184 -52173 184 -52139
rect -184 -52501 184 -52467
rect -184 -52609 184 -52575
rect -184 -52937 184 -52903
rect -184 -53045 184 -53011
rect -184 -53373 184 -53339
rect -184 -53481 184 -53447
rect -184 -53809 184 -53775
rect -184 -53917 184 -53883
rect -184 -54245 184 -54211
rect -184 -54353 184 -54319
rect -184 -54681 184 -54647
rect -184 -54789 184 -54755
rect -184 -55117 184 -55083
rect -184 -55225 184 -55191
rect -184 -55553 184 -55519
rect -184 -55661 184 -55627
rect -184 -55989 184 -55955
rect -184 -56097 184 -56063
rect -184 -56425 184 -56391
rect -184 -56533 184 -56499
rect -184 -56861 184 -56827
rect -184 -56969 184 -56935
rect -184 -57297 184 -57263
rect -184 -57405 184 -57371
rect -184 -57733 184 -57699
rect -184 -57841 184 -57807
rect -184 -58169 184 -58135
rect -184 -58277 184 -58243
rect -184 -58605 184 -58571
rect -184 -58713 184 -58679
rect -184 -59041 184 -59007
rect -184 -59149 184 -59115
rect -184 -59477 184 -59443
rect -184 -59585 184 -59551
rect -184 -59913 184 -59879
rect -184 -60021 184 -59987
rect -184 -60349 184 -60315
rect -184 -60457 184 -60423
rect -184 -60785 184 -60751
rect -184 -60893 184 -60859
rect -184 -61221 184 -61187
rect -184 -61329 184 -61295
rect -184 -61657 184 -61623
rect -184 -61765 184 -61731
rect -184 -62093 184 -62059
rect -184 -62201 184 -62167
rect -184 -62529 184 -62495
rect -184 -62637 184 -62603
rect -184 -62965 184 -62931
rect -184 -63073 184 -63039
rect -184 -63401 184 -63367
rect -184 -63509 184 -63475
rect -184 -63837 184 -63803
rect -184 -63945 184 -63911
rect -184 -64273 184 -64239
rect -184 -64381 184 -64347
rect -184 -64709 184 -64675
rect -184 -64817 184 -64783
rect -184 -65145 184 -65111
rect -184 -65253 184 -65219
rect -184 -65581 184 -65547
rect -184 -65689 184 -65655
rect -184 -66017 184 -65983
rect -184 -66125 184 -66091
rect -184 -66453 184 -66419
rect -184 -66561 184 -66527
rect -184 -66889 184 -66855
rect -184 -66997 184 -66963
rect -184 -67325 184 -67291
rect -184 -67433 184 -67399
rect -184 -67761 184 -67727
rect -184 -67869 184 -67835
rect -184 -68197 184 -68163
rect -184 -68305 184 -68271
rect -184 -68633 184 -68599
rect -184 -68741 184 -68707
rect -184 -69069 184 -69035
rect -184 -69177 184 -69143
rect -184 -69505 184 -69471
rect -184 -69613 184 -69579
rect -184 -69941 184 -69907
rect -184 -70049 184 -70015
rect -184 -70377 184 -70343
rect -184 -70485 184 -70451
rect -184 -70813 184 -70779
rect -184 -70921 184 -70887
rect -184 -71249 184 -71215
rect -184 -71357 184 -71323
rect -184 -71685 184 -71651
rect -184 -71793 184 -71759
rect -184 -72121 184 -72087
rect -184 -72229 184 -72195
rect -184 -72557 184 -72523
rect -184 -72665 184 -72631
rect -184 -72993 184 -72959
rect -184 -73101 184 -73067
rect -184 -73429 184 -73395
rect -184 -73537 184 -73503
rect -184 -73865 184 -73831
rect -184 -73973 184 -73939
rect -184 -74301 184 -74267
rect -184 -74409 184 -74375
rect -184 -74737 184 -74703
rect -184 -74845 184 -74811
rect -184 -75173 184 -75139
rect -184 -75281 184 -75247
rect -184 -75609 184 -75575
rect -184 -75717 184 -75683
rect -184 -76045 184 -76011
rect -184 -76153 184 -76119
rect -184 -76481 184 -76447
rect -184 -76589 184 -76555
rect -184 -76917 184 -76883
rect -184 -77025 184 -76991
rect -184 -77353 184 -77319
rect -184 -77461 184 -77427
rect -184 -77789 184 -77755
rect -184 -77897 184 -77863
rect -184 -78225 184 -78191
rect -184 -78333 184 -78299
rect -184 -78661 184 -78627
rect -184 -78769 184 -78735
rect -184 -79097 184 -79063
rect -184 -79205 184 -79171
rect -184 -79533 184 -79499
rect -184 -79641 184 -79607
rect -184 -79969 184 -79935
rect -184 -80077 184 -80043
rect -184 -80405 184 -80371
rect -184 -80513 184 -80479
rect -184 -80841 184 -80807
rect -184 -80949 184 -80915
rect -184 -81277 184 -81243
rect -184 -81385 184 -81351
rect -184 -81713 184 -81679
rect -184 -81821 184 -81787
rect -184 -82149 184 -82115
rect -184 -82257 184 -82223
rect -184 -82585 184 -82551
rect -184 -82693 184 -82659
rect -184 -83021 184 -82987
rect -184 -83129 184 -83095
rect -184 -83457 184 -83423
rect -184 -83565 184 -83531
rect -184 -83893 184 -83859
rect -184 -84001 184 -83967
rect -184 -84329 184 -84295
<< locali >>
rect -360 84397 -264 84431
rect 264 84397 360 84431
rect -360 84335 -326 84397
rect 326 84335 360 84397
rect -200 84295 -184 84329
rect 184 84295 200 84329
rect -246 84236 -212 84252
rect -246 84044 -212 84060
rect 212 84236 246 84252
rect 212 84044 246 84060
rect -200 83967 -184 84001
rect 184 83967 200 84001
rect -200 83859 -184 83893
rect 184 83859 200 83893
rect -246 83800 -212 83816
rect -246 83608 -212 83624
rect 212 83800 246 83816
rect 212 83608 246 83624
rect -200 83531 -184 83565
rect 184 83531 200 83565
rect -200 83423 -184 83457
rect 184 83423 200 83457
rect -246 83364 -212 83380
rect -246 83172 -212 83188
rect 212 83364 246 83380
rect 212 83172 246 83188
rect -200 83095 -184 83129
rect 184 83095 200 83129
rect -200 82987 -184 83021
rect 184 82987 200 83021
rect -246 82928 -212 82944
rect -246 82736 -212 82752
rect 212 82928 246 82944
rect 212 82736 246 82752
rect -200 82659 -184 82693
rect 184 82659 200 82693
rect -200 82551 -184 82585
rect 184 82551 200 82585
rect -246 82492 -212 82508
rect -246 82300 -212 82316
rect 212 82492 246 82508
rect 212 82300 246 82316
rect -200 82223 -184 82257
rect 184 82223 200 82257
rect -200 82115 -184 82149
rect 184 82115 200 82149
rect -246 82056 -212 82072
rect -246 81864 -212 81880
rect 212 82056 246 82072
rect 212 81864 246 81880
rect -200 81787 -184 81821
rect 184 81787 200 81821
rect -200 81679 -184 81713
rect 184 81679 200 81713
rect -246 81620 -212 81636
rect -246 81428 -212 81444
rect 212 81620 246 81636
rect 212 81428 246 81444
rect -200 81351 -184 81385
rect 184 81351 200 81385
rect -200 81243 -184 81277
rect 184 81243 200 81277
rect -246 81184 -212 81200
rect -246 80992 -212 81008
rect 212 81184 246 81200
rect 212 80992 246 81008
rect -200 80915 -184 80949
rect 184 80915 200 80949
rect -200 80807 -184 80841
rect 184 80807 200 80841
rect -246 80748 -212 80764
rect -246 80556 -212 80572
rect 212 80748 246 80764
rect 212 80556 246 80572
rect -200 80479 -184 80513
rect 184 80479 200 80513
rect -200 80371 -184 80405
rect 184 80371 200 80405
rect -246 80312 -212 80328
rect -246 80120 -212 80136
rect 212 80312 246 80328
rect 212 80120 246 80136
rect -200 80043 -184 80077
rect 184 80043 200 80077
rect -200 79935 -184 79969
rect 184 79935 200 79969
rect -246 79876 -212 79892
rect -246 79684 -212 79700
rect 212 79876 246 79892
rect 212 79684 246 79700
rect -200 79607 -184 79641
rect 184 79607 200 79641
rect -200 79499 -184 79533
rect 184 79499 200 79533
rect -246 79440 -212 79456
rect -246 79248 -212 79264
rect 212 79440 246 79456
rect 212 79248 246 79264
rect -200 79171 -184 79205
rect 184 79171 200 79205
rect -200 79063 -184 79097
rect 184 79063 200 79097
rect -246 79004 -212 79020
rect -246 78812 -212 78828
rect 212 79004 246 79020
rect 212 78812 246 78828
rect -200 78735 -184 78769
rect 184 78735 200 78769
rect -200 78627 -184 78661
rect 184 78627 200 78661
rect -246 78568 -212 78584
rect -246 78376 -212 78392
rect 212 78568 246 78584
rect 212 78376 246 78392
rect -200 78299 -184 78333
rect 184 78299 200 78333
rect -200 78191 -184 78225
rect 184 78191 200 78225
rect -246 78132 -212 78148
rect -246 77940 -212 77956
rect 212 78132 246 78148
rect 212 77940 246 77956
rect -200 77863 -184 77897
rect 184 77863 200 77897
rect -200 77755 -184 77789
rect 184 77755 200 77789
rect -246 77696 -212 77712
rect -246 77504 -212 77520
rect 212 77696 246 77712
rect 212 77504 246 77520
rect -200 77427 -184 77461
rect 184 77427 200 77461
rect -200 77319 -184 77353
rect 184 77319 200 77353
rect -246 77260 -212 77276
rect -246 77068 -212 77084
rect 212 77260 246 77276
rect 212 77068 246 77084
rect -200 76991 -184 77025
rect 184 76991 200 77025
rect -200 76883 -184 76917
rect 184 76883 200 76917
rect -246 76824 -212 76840
rect -246 76632 -212 76648
rect 212 76824 246 76840
rect 212 76632 246 76648
rect -200 76555 -184 76589
rect 184 76555 200 76589
rect -200 76447 -184 76481
rect 184 76447 200 76481
rect -246 76388 -212 76404
rect -246 76196 -212 76212
rect 212 76388 246 76404
rect 212 76196 246 76212
rect -200 76119 -184 76153
rect 184 76119 200 76153
rect -200 76011 -184 76045
rect 184 76011 200 76045
rect -246 75952 -212 75968
rect -246 75760 -212 75776
rect 212 75952 246 75968
rect 212 75760 246 75776
rect -200 75683 -184 75717
rect 184 75683 200 75717
rect -200 75575 -184 75609
rect 184 75575 200 75609
rect -246 75516 -212 75532
rect -246 75324 -212 75340
rect 212 75516 246 75532
rect 212 75324 246 75340
rect -200 75247 -184 75281
rect 184 75247 200 75281
rect -200 75139 -184 75173
rect 184 75139 200 75173
rect -246 75080 -212 75096
rect -246 74888 -212 74904
rect 212 75080 246 75096
rect 212 74888 246 74904
rect -200 74811 -184 74845
rect 184 74811 200 74845
rect -200 74703 -184 74737
rect 184 74703 200 74737
rect -246 74644 -212 74660
rect -246 74452 -212 74468
rect 212 74644 246 74660
rect 212 74452 246 74468
rect -200 74375 -184 74409
rect 184 74375 200 74409
rect -200 74267 -184 74301
rect 184 74267 200 74301
rect -246 74208 -212 74224
rect -246 74016 -212 74032
rect 212 74208 246 74224
rect 212 74016 246 74032
rect -200 73939 -184 73973
rect 184 73939 200 73973
rect -200 73831 -184 73865
rect 184 73831 200 73865
rect -246 73772 -212 73788
rect -246 73580 -212 73596
rect 212 73772 246 73788
rect 212 73580 246 73596
rect -200 73503 -184 73537
rect 184 73503 200 73537
rect -200 73395 -184 73429
rect 184 73395 200 73429
rect -246 73336 -212 73352
rect -246 73144 -212 73160
rect 212 73336 246 73352
rect 212 73144 246 73160
rect -200 73067 -184 73101
rect 184 73067 200 73101
rect -200 72959 -184 72993
rect 184 72959 200 72993
rect -246 72900 -212 72916
rect -246 72708 -212 72724
rect 212 72900 246 72916
rect 212 72708 246 72724
rect -200 72631 -184 72665
rect 184 72631 200 72665
rect -200 72523 -184 72557
rect 184 72523 200 72557
rect -246 72464 -212 72480
rect -246 72272 -212 72288
rect 212 72464 246 72480
rect 212 72272 246 72288
rect -200 72195 -184 72229
rect 184 72195 200 72229
rect -200 72087 -184 72121
rect 184 72087 200 72121
rect -246 72028 -212 72044
rect -246 71836 -212 71852
rect 212 72028 246 72044
rect 212 71836 246 71852
rect -200 71759 -184 71793
rect 184 71759 200 71793
rect -200 71651 -184 71685
rect 184 71651 200 71685
rect -246 71592 -212 71608
rect -246 71400 -212 71416
rect 212 71592 246 71608
rect 212 71400 246 71416
rect -200 71323 -184 71357
rect 184 71323 200 71357
rect -200 71215 -184 71249
rect 184 71215 200 71249
rect -246 71156 -212 71172
rect -246 70964 -212 70980
rect 212 71156 246 71172
rect 212 70964 246 70980
rect -200 70887 -184 70921
rect 184 70887 200 70921
rect -200 70779 -184 70813
rect 184 70779 200 70813
rect -246 70720 -212 70736
rect -246 70528 -212 70544
rect 212 70720 246 70736
rect 212 70528 246 70544
rect -200 70451 -184 70485
rect 184 70451 200 70485
rect -200 70343 -184 70377
rect 184 70343 200 70377
rect -246 70284 -212 70300
rect -246 70092 -212 70108
rect 212 70284 246 70300
rect 212 70092 246 70108
rect -200 70015 -184 70049
rect 184 70015 200 70049
rect -200 69907 -184 69941
rect 184 69907 200 69941
rect -246 69848 -212 69864
rect -246 69656 -212 69672
rect 212 69848 246 69864
rect 212 69656 246 69672
rect -200 69579 -184 69613
rect 184 69579 200 69613
rect -200 69471 -184 69505
rect 184 69471 200 69505
rect -246 69412 -212 69428
rect -246 69220 -212 69236
rect 212 69412 246 69428
rect 212 69220 246 69236
rect -200 69143 -184 69177
rect 184 69143 200 69177
rect -200 69035 -184 69069
rect 184 69035 200 69069
rect -246 68976 -212 68992
rect -246 68784 -212 68800
rect 212 68976 246 68992
rect 212 68784 246 68800
rect -200 68707 -184 68741
rect 184 68707 200 68741
rect -200 68599 -184 68633
rect 184 68599 200 68633
rect -246 68540 -212 68556
rect -246 68348 -212 68364
rect 212 68540 246 68556
rect 212 68348 246 68364
rect -200 68271 -184 68305
rect 184 68271 200 68305
rect -200 68163 -184 68197
rect 184 68163 200 68197
rect -246 68104 -212 68120
rect -246 67912 -212 67928
rect 212 68104 246 68120
rect 212 67912 246 67928
rect -200 67835 -184 67869
rect 184 67835 200 67869
rect -200 67727 -184 67761
rect 184 67727 200 67761
rect -246 67668 -212 67684
rect -246 67476 -212 67492
rect 212 67668 246 67684
rect 212 67476 246 67492
rect -200 67399 -184 67433
rect 184 67399 200 67433
rect -200 67291 -184 67325
rect 184 67291 200 67325
rect -246 67232 -212 67248
rect -246 67040 -212 67056
rect 212 67232 246 67248
rect 212 67040 246 67056
rect -200 66963 -184 66997
rect 184 66963 200 66997
rect -200 66855 -184 66889
rect 184 66855 200 66889
rect -246 66796 -212 66812
rect -246 66604 -212 66620
rect 212 66796 246 66812
rect 212 66604 246 66620
rect -200 66527 -184 66561
rect 184 66527 200 66561
rect -200 66419 -184 66453
rect 184 66419 200 66453
rect -246 66360 -212 66376
rect -246 66168 -212 66184
rect 212 66360 246 66376
rect 212 66168 246 66184
rect -200 66091 -184 66125
rect 184 66091 200 66125
rect -200 65983 -184 66017
rect 184 65983 200 66017
rect -246 65924 -212 65940
rect -246 65732 -212 65748
rect 212 65924 246 65940
rect 212 65732 246 65748
rect -200 65655 -184 65689
rect 184 65655 200 65689
rect -200 65547 -184 65581
rect 184 65547 200 65581
rect -246 65488 -212 65504
rect -246 65296 -212 65312
rect 212 65488 246 65504
rect 212 65296 246 65312
rect -200 65219 -184 65253
rect 184 65219 200 65253
rect -200 65111 -184 65145
rect 184 65111 200 65145
rect -246 65052 -212 65068
rect -246 64860 -212 64876
rect 212 65052 246 65068
rect 212 64860 246 64876
rect -200 64783 -184 64817
rect 184 64783 200 64817
rect -200 64675 -184 64709
rect 184 64675 200 64709
rect -246 64616 -212 64632
rect -246 64424 -212 64440
rect 212 64616 246 64632
rect 212 64424 246 64440
rect -200 64347 -184 64381
rect 184 64347 200 64381
rect -200 64239 -184 64273
rect 184 64239 200 64273
rect -246 64180 -212 64196
rect -246 63988 -212 64004
rect 212 64180 246 64196
rect 212 63988 246 64004
rect -200 63911 -184 63945
rect 184 63911 200 63945
rect -200 63803 -184 63837
rect 184 63803 200 63837
rect -246 63744 -212 63760
rect -246 63552 -212 63568
rect 212 63744 246 63760
rect 212 63552 246 63568
rect -200 63475 -184 63509
rect 184 63475 200 63509
rect -200 63367 -184 63401
rect 184 63367 200 63401
rect -246 63308 -212 63324
rect -246 63116 -212 63132
rect 212 63308 246 63324
rect 212 63116 246 63132
rect -200 63039 -184 63073
rect 184 63039 200 63073
rect -200 62931 -184 62965
rect 184 62931 200 62965
rect -246 62872 -212 62888
rect -246 62680 -212 62696
rect 212 62872 246 62888
rect 212 62680 246 62696
rect -200 62603 -184 62637
rect 184 62603 200 62637
rect -200 62495 -184 62529
rect 184 62495 200 62529
rect -246 62436 -212 62452
rect -246 62244 -212 62260
rect 212 62436 246 62452
rect 212 62244 246 62260
rect -200 62167 -184 62201
rect 184 62167 200 62201
rect -200 62059 -184 62093
rect 184 62059 200 62093
rect -246 62000 -212 62016
rect -246 61808 -212 61824
rect 212 62000 246 62016
rect 212 61808 246 61824
rect -200 61731 -184 61765
rect 184 61731 200 61765
rect -200 61623 -184 61657
rect 184 61623 200 61657
rect -246 61564 -212 61580
rect -246 61372 -212 61388
rect 212 61564 246 61580
rect 212 61372 246 61388
rect -200 61295 -184 61329
rect 184 61295 200 61329
rect -200 61187 -184 61221
rect 184 61187 200 61221
rect -246 61128 -212 61144
rect -246 60936 -212 60952
rect 212 61128 246 61144
rect 212 60936 246 60952
rect -200 60859 -184 60893
rect 184 60859 200 60893
rect -200 60751 -184 60785
rect 184 60751 200 60785
rect -246 60692 -212 60708
rect -246 60500 -212 60516
rect 212 60692 246 60708
rect 212 60500 246 60516
rect -200 60423 -184 60457
rect 184 60423 200 60457
rect -200 60315 -184 60349
rect 184 60315 200 60349
rect -246 60256 -212 60272
rect -246 60064 -212 60080
rect 212 60256 246 60272
rect 212 60064 246 60080
rect -200 59987 -184 60021
rect 184 59987 200 60021
rect -200 59879 -184 59913
rect 184 59879 200 59913
rect -246 59820 -212 59836
rect -246 59628 -212 59644
rect 212 59820 246 59836
rect 212 59628 246 59644
rect -200 59551 -184 59585
rect 184 59551 200 59585
rect -200 59443 -184 59477
rect 184 59443 200 59477
rect -246 59384 -212 59400
rect -246 59192 -212 59208
rect 212 59384 246 59400
rect 212 59192 246 59208
rect -200 59115 -184 59149
rect 184 59115 200 59149
rect -200 59007 -184 59041
rect 184 59007 200 59041
rect -246 58948 -212 58964
rect -246 58756 -212 58772
rect 212 58948 246 58964
rect 212 58756 246 58772
rect -200 58679 -184 58713
rect 184 58679 200 58713
rect -200 58571 -184 58605
rect 184 58571 200 58605
rect -246 58512 -212 58528
rect -246 58320 -212 58336
rect 212 58512 246 58528
rect 212 58320 246 58336
rect -200 58243 -184 58277
rect 184 58243 200 58277
rect -200 58135 -184 58169
rect 184 58135 200 58169
rect -246 58076 -212 58092
rect -246 57884 -212 57900
rect 212 58076 246 58092
rect 212 57884 246 57900
rect -200 57807 -184 57841
rect 184 57807 200 57841
rect -200 57699 -184 57733
rect 184 57699 200 57733
rect -246 57640 -212 57656
rect -246 57448 -212 57464
rect 212 57640 246 57656
rect 212 57448 246 57464
rect -200 57371 -184 57405
rect 184 57371 200 57405
rect -200 57263 -184 57297
rect 184 57263 200 57297
rect -246 57204 -212 57220
rect -246 57012 -212 57028
rect 212 57204 246 57220
rect 212 57012 246 57028
rect -200 56935 -184 56969
rect 184 56935 200 56969
rect -200 56827 -184 56861
rect 184 56827 200 56861
rect -246 56768 -212 56784
rect -246 56576 -212 56592
rect 212 56768 246 56784
rect 212 56576 246 56592
rect -200 56499 -184 56533
rect 184 56499 200 56533
rect -200 56391 -184 56425
rect 184 56391 200 56425
rect -246 56332 -212 56348
rect -246 56140 -212 56156
rect 212 56332 246 56348
rect 212 56140 246 56156
rect -200 56063 -184 56097
rect 184 56063 200 56097
rect -200 55955 -184 55989
rect 184 55955 200 55989
rect -246 55896 -212 55912
rect -246 55704 -212 55720
rect 212 55896 246 55912
rect 212 55704 246 55720
rect -200 55627 -184 55661
rect 184 55627 200 55661
rect -200 55519 -184 55553
rect 184 55519 200 55553
rect -246 55460 -212 55476
rect -246 55268 -212 55284
rect 212 55460 246 55476
rect 212 55268 246 55284
rect -200 55191 -184 55225
rect 184 55191 200 55225
rect -200 55083 -184 55117
rect 184 55083 200 55117
rect -246 55024 -212 55040
rect -246 54832 -212 54848
rect 212 55024 246 55040
rect 212 54832 246 54848
rect -200 54755 -184 54789
rect 184 54755 200 54789
rect -200 54647 -184 54681
rect 184 54647 200 54681
rect -246 54588 -212 54604
rect -246 54396 -212 54412
rect 212 54588 246 54604
rect 212 54396 246 54412
rect -200 54319 -184 54353
rect 184 54319 200 54353
rect -200 54211 -184 54245
rect 184 54211 200 54245
rect -246 54152 -212 54168
rect -246 53960 -212 53976
rect 212 54152 246 54168
rect 212 53960 246 53976
rect -200 53883 -184 53917
rect 184 53883 200 53917
rect -200 53775 -184 53809
rect 184 53775 200 53809
rect -246 53716 -212 53732
rect -246 53524 -212 53540
rect 212 53716 246 53732
rect 212 53524 246 53540
rect -200 53447 -184 53481
rect 184 53447 200 53481
rect -200 53339 -184 53373
rect 184 53339 200 53373
rect -246 53280 -212 53296
rect -246 53088 -212 53104
rect 212 53280 246 53296
rect 212 53088 246 53104
rect -200 53011 -184 53045
rect 184 53011 200 53045
rect -200 52903 -184 52937
rect 184 52903 200 52937
rect -246 52844 -212 52860
rect -246 52652 -212 52668
rect 212 52844 246 52860
rect 212 52652 246 52668
rect -200 52575 -184 52609
rect 184 52575 200 52609
rect -200 52467 -184 52501
rect 184 52467 200 52501
rect -246 52408 -212 52424
rect -246 52216 -212 52232
rect 212 52408 246 52424
rect 212 52216 246 52232
rect -200 52139 -184 52173
rect 184 52139 200 52173
rect -200 52031 -184 52065
rect 184 52031 200 52065
rect -246 51972 -212 51988
rect -246 51780 -212 51796
rect 212 51972 246 51988
rect 212 51780 246 51796
rect -200 51703 -184 51737
rect 184 51703 200 51737
rect -200 51595 -184 51629
rect 184 51595 200 51629
rect -246 51536 -212 51552
rect -246 51344 -212 51360
rect 212 51536 246 51552
rect 212 51344 246 51360
rect -200 51267 -184 51301
rect 184 51267 200 51301
rect -200 51159 -184 51193
rect 184 51159 200 51193
rect -246 51100 -212 51116
rect -246 50908 -212 50924
rect 212 51100 246 51116
rect 212 50908 246 50924
rect -200 50831 -184 50865
rect 184 50831 200 50865
rect -200 50723 -184 50757
rect 184 50723 200 50757
rect -246 50664 -212 50680
rect -246 50472 -212 50488
rect 212 50664 246 50680
rect 212 50472 246 50488
rect -200 50395 -184 50429
rect 184 50395 200 50429
rect -200 50287 -184 50321
rect 184 50287 200 50321
rect -246 50228 -212 50244
rect -246 50036 -212 50052
rect 212 50228 246 50244
rect 212 50036 246 50052
rect -200 49959 -184 49993
rect 184 49959 200 49993
rect -200 49851 -184 49885
rect 184 49851 200 49885
rect -246 49792 -212 49808
rect -246 49600 -212 49616
rect 212 49792 246 49808
rect 212 49600 246 49616
rect -200 49523 -184 49557
rect 184 49523 200 49557
rect -200 49415 -184 49449
rect 184 49415 200 49449
rect -246 49356 -212 49372
rect -246 49164 -212 49180
rect 212 49356 246 49372
rect 212 49164 246 49180
rect -200 49087 -184 49121
rect 184 49087 200 49121
rect -200 48979 -184 49013
rect 184 48979 200 49013
rect -246 48920 -212 48936
rect -246 48728 -212 48744
rect 212 48920 246 48936
rect 212 48728 246 48744
rect -200 48651 -184 48685
rect 184 48651 200 48685
rect -200 48543 -184 48577
rect 184 48543 200 48577
rect -246 48484 -212 48500
rect -246 48292 -212 48308
rect 212 48484 246 48500
rect 212 48292 246 48308
rect -200 48215 -184 48249
rect 184 48215 200 48249
rect -200 48107 -184 48141
rect 184 48107 200 48141
rect -246 48048 -212 48064
rect -246 47856 -212 47872
rect 212 48048 246 48064
rect 212 47856 246 47872
rect -200 47779 -184 47813
rect 184 47779 200 47813
rect -200 47671 -184 47705
rect 184 47671 200 47705
rect -246 47612 -212 47628
rect -246 47420 -212 47436
rect 212 47612 246 47628
rect 212 47420 246 47436
rect -200 47343 -184 47377
rect 184 47343 200 47377
rect -200 47235 -184 47269
rect 184 47235 200 47269
rect -246 47176 -212 47192
rect -246 46984 -212 47000
rect 212 47176 246 47192
rect 212 46984 246 47000
rect -200 46907 -184 46941
rect 184 46907 200 46941
rect -200 46799 -184 46833
rect 184 46799 200 46833
rect -246 46740 -212 46756
rect -246 46548 -212 46564
rect 212 46740 246 46756
rect 212 46548 246 46564
rect -200 46471 -184 46505
rect 184 46471 200 46505
rect -200 46363 -184 46397
rect 184 46363 200 46397
rect -246 46304 -212 46320
rect -246 46112 -212 46128
rect 212 46304 246 46320
rect 212 46112 246 46128
rect -200 46035 -184 46069
rect 184 46035 200 46069
rect -200 45927 -184 45961
rect 184 45927 200 45961
rect -246 45868 -212 45884
rect -246 45676 -212 45692
rect 212 45868 246 45884
rect 212 45676 246 45692
rect -200 45599 -184 45633
rect 184 45599 200 45633
rect -200 45491 -184 45525
rect 184 45491 200 45525
rect -246 45432 -212 45448
rect -246 45240 -212 45256
rect 212 45432 246 45448
rect 212 45240 246 45256
rect -200 45163 -184 45197
rect 184 45163 200 45197
rect -200 45055 -184 45089
rect 184 45055 200 45089
rect -246 44996 -212 45012
rect -246 44804 -212 44820
rect 212 44996 246 45012
rect 212 44804 246 44820
rect -200 44727 -184 44761
rect 184 44727 200 44761
rect -200 44619 -184 44653
rect 184 44619 200 44653
rect -246 44560 -212 44576
rect -246 44368 -212 44384
rect 212 44560 246 44576
rect 212 44368 246 44384
rect -200 44291 -184 44325
rect 184 44291 200 44325
rect -200 44183 -184 44217
rect 184 44183 200 44217
rect -246 44124 -212 44140
rect -246 43932 -212 43948
rect 212 44124 246 44140
rect 212 43932 246 43948
rect -200 43855 -184 43889
rect 184 43855 200 43889
rect -200 43747 -184 43781
rect 184 43747 200 43781
rect -246 43688 -212 43704
rect -246 43496 -212 43512
rect 212 43688 246 43704
rect 212 43496 246 43512
rect -200 43419 -184 43453
rect 184 43419 200 43453
rect -200 43311 -184 43345
rect 184 43311 200 43345
rect -246 43252 -212 43268
rect -246 43060 -212 43076
rect 212 43252 246 43268
rect 212 43060 246 43076
rect -200 42983 -184 43017
rect 184 42983 200 43017
rect -200 42875 -184 42909
rect 184 42875 200 42909
rect -246 42816 -212 42832
rect -246 42624 -212 42640
rect 212 42816 246 42832
rect 212 42624 246 42640
rect -200 42547 -184 42581
rect 184 42547 200 42581
rect -200 42439 -184 42473
rect 184 42439 200 42473
rect -246 42380 -212 42396
rect -246 42188 -212 42204
rect 212 42380 246 42396
rect 212 42188 246 42204
rect -200 42111 -184 42145
rect 184 42111 200 42145
rect -200 42003 -184 42037
rect 184 42003 200 42037
rect -246 41944 -212 41960
rect -246 41752 -212 41768
rect 212 41944 246 41960
rect 212 41752 246 41768
rect -200 41675 -184 41709
rect 184 41675 200 41709
rect -200 41567 -184 41601
rect 184 41567 200 41601
rect -246 41508 -212 41524
rect -246 41316 -212 41332
rect 212 41508 246 41524
rect 212 41316 246 41332
rect -200 41239 -184 41273
rect 184 41239 200 41273
rect -200 41131 -184 41165
rect 184 41131 200 41165
rect -246 41072 -212 41088
rect -246 40880 -212 40896
rect 212 41072 246 41088
rect 212 40880 246 40896
rect -200 40803 -184 40837
rect 184 40803 200 40837
rect -200 40695 -184 40729
rect 184 40695 200 40729
rect -246 40636 -212 40652
rect -246 40444 -212 40460
rect 212 40636 246 40652
rect 212 40444 246 40460
rect -200 40367 -184 40401
rect 184 40367 200 40401
rect -200 40259 -184 40293
rect 184 40259 200 40293
rect -246 40200 -212 40216
rect -246 40008 -212 40024
rect 212 40200 246 40216
rect 212 40008 246 40024
rect -200 39931 -184 39965
rect 184 39931 200 39965
rect -200 39823 -184 39857
rect 184 39823 200 39857
rect -246 39764 -212 39780
rect -246 39572 -212 39588
rect 212 39764 246 39780
rect 212 39572 246 39588
rect -200 39495 -184 39529
rect 184 39495 200 39529
rect -200 39387 -184 39421
rect 184 39387 200 39421
rect -246 39328 -212 39344
rect -246 39136 -212 39152
rect 212 39328 246 39344
rect 212 39136 246 39152
rect -200 39059 -184 39093
rect 184 39059 200 39093
rect -200 38951 -184 38985
rect 184 38951 200 38985
rect -246 38892 -212 38908
rect -246 38700 -212 38716
rect 212 38892 246 38908
rect 212 38700 246 38716
rect -200 38623 -184 38657
rect 184 38623 200 38657
rect -200 38515 -184 38549
rect 184 38515 200 38549
rect -246 38456 -212 38472
rect -246 38264 -212 38280
rect 212 38456 246 38472
rect 212 38264 246 38280
rect -200 38187 -184 38221
rect 184 38187 200 38221
rect -200 38079 -184 38113
rect 184 38079 200 38113
rect -246 38020 -212 38036
rect -246 37828 -212 37844
rect 212 38020 246 38036
rect 212 37828 246 37844
rect -200 37751 -184 37785
rect 184 37751 200 37785
rect -200 37643 -184 37677
rect 184 37643 200 37677
rect -246 37584 -212 37600
rect -246 37392 -212 37408
rect 212 37584 246 37600
rect 212 37392 246 37408
rect -200 37315 -184 37349
rect 184 37315 200 37349
rect -200 37207 -184 37241
rect 184 37207 200 37241
rect -246 37148 -212 37164
rect -246 36956 -212 36972
rect 212 37148 246 37164
rect 212 36956 246 36972
rect -200 36879 -184 36913
rect 184 36879 200 36913
rect -200 36771 -184 36805
rect 184 36771 200 36805
rect -246 36712 -212 36728
rect -246 36520 -212 36536
rect 212 36712 246 36728
rect 212 36520 246 36536
rect -200 36443 -184 36477
rect 184 36443 200 36477
rect -200 36335 -184 36369
rect 184 36335 200 36369
rect -246 36276 -212 36292
rect -246 36084 -212 36100
rect 212 36276 246 36292
rect 212 36084 246 36100
rect -200 36007 -184 36041
rect 184 36007 200 36041
rect -200 35899 -184 35933
rect 184 35899 200 35933
rect -246 35840 -212 35856
rect -246 35648 -212 35664
rect 212 35840 246 35856
rect 212 35648 246 35664
rect -200 35571 -184 35605
rect 184 35571 200 35605
rect -200 35463 -184 35497
rect 184 35463 200 35497
rect -246 35404 -212 35420
rect -246 35212 -212 35228
rect 212 35404 246 35420
rect 212 35212 246 35228
rect -200 35135 -184 35169
rect 184 35135 200 35169
rect -200 35027 -184 35061
rect 184 35027 200 35061
rect -246 34968 -212 34984
rect -246 34776 -212 34792
rect 212 34968 246 34984
rect 212 34776 246 34792
rect -200 34699 -184 34733
rect 184 34699 200 34733
rect -200 34591 -184 34625
rect 184 34591 200 34625
rect -246 34532 -212 34548
rect -246 34340 -212 34356
rect 212 34532 246 34548
rect 212 34340 246 34356
rect -200 34263 -184 34297
rect 184 34263 200 34297
rect -200 34155 -184 34189
rect 184 34155 200 34189
rect -246 34096 -212 34112
rect -246 33904 -212 33920
rect 212 34096 246 34112
rect 212 33904 246 33920
rect -200 33827 -184 33861
rect 184 33827 200 33861
rect -200 33719 -184 33753
rect 184 33719 200 33753
rect -246 33660 -212 33676
rect -246 33468 -212 33484
rect 212 33660 246 33676
rect 212 33468 246 33484
rect -200 33391 -184 33425
rect 184 33391 200 33425
rect -200 33283 -184 33317
rect 184 33283 200 33317
rect -246 33224 -212 33240
rect -246 33032 -212 33048
rect 212 33224 246 33240
rect 212 33032 246 33048
rect -200 32955 -184 32989
rect 184 32955 200 32989
rect -200 32847 -184 32881
rect 184 32847 200 32881
rect -246 32788 -212 32804
rect -246 32596 -212 32612
rect 212 32788 246 32804
rect 212 32596 246 32612
rect -200 32519 -184 32553
rect 184 32519 200 32553
rect -200 32411 -184 32445
rect 184 32411 200 32445
rect -246 32352 -212 32368
rect -246 32160 -212 32176
rect 212 32352 246 32368
rect 212 32160 246 32176
rect -200 32083 -184 32117
rect 184 32083 200 32117
rect -200 31975 -184 32009
rect 184 31975 200 32009
rect -246 31916 -212 31932
rect -246 31724 -212 31740
rect 212 31916 246 31932
rect 212 31724 246 31740
rect -200 31647 -184 31681
rect 184 31647 200 31681
rect -200 31539 -184 31573
rect 184 31539 200 31573
rect -246 31480 -212 31496
rect -246 31288 -212 31304
rect 212 31480 246 31496
rect 212 31288 246 31304
rect -200 31211 -184 31245
rect 184 31211 200 31245
rect -200 31103 -184 31137
rect 184 31103 200 31137
rect -246 31044 -212 31060
rect -246 30852 -212 30868
rect 212 31044 246 31060
rect 212 30852 246 30868
rect -200 30775 -184 30809
rect 184 30775 200 30809
rect -200 30667 -184 30701
rect 184 30667 200 30701
rect -246 30608 -212 30624
rect -246 30416 -212 30432
rect 212 30608 246 30624
rect 212 30416 246 30432
rect -200 30339 -184 30373
rect 184 30339 200 30373
rect -200 30231 -184 30265
rect 184 30231 200 30265
rect -246 30172 -212 30188
rect -246 29980 -212 29996
rect 212 30172 246 30188
rect 212 29980 246 29996
rect -200 29903 -184 29937
rect 184 29903 200 29937
rect -200 29795 -184 29829
rect 184 29795 200 29829
rect -246 29736 -212 29752
rect -246 29544 -212 29560
rect 212 29736 246 29752
rect 212 29544 246 29560
rect -200 29467 -184 29501
rect 184 29467 200 29501
rect -200 29359 -184 29393
rect 184 29359 200 29393
rect -246 29300 -212 29316
rect -246 29108 -212 29124
rect 212 29300 246 29316
rect 212 29108 246 29124
rect -200 29031 -184 29065
rect 184 29031 200 29065
rect -200 28923 -184 28957
rect 184 28923 200 28957
rect -246 28864 -212 28880
rect -246 28672 -212 28688
rect 212 28864 246 28880
rect 212 28672 246 28688
rect -200 28595 -184 28629
rect 184 28595 200 28629
rect -200 28487 -184 28521
rect 184 28487 200 28521
rect -246 28428 -212 28444
rect -246 28236 -212 28252
rect 212 28428 246 28444
rect 212 28236 246 28252
rect -200 28159 -184 28193
rect 184 28159 200 28193
rect -200 28051 -184 28085
rect 184 28051 200 28085
rect -246 27992 -212 28008
rect -246 27800 -212 27816
rect 212 27992 246 28008
rect 212 27800 246 27816
rect -200 27723 -184 27757
rect 184 27723 200 27757
rect -200 27615 -184 27649
rect 184 27615 200 27649
rect -246 27556 -212 27572
rect -246 27364 -212 27380
rect 212 27556 246 27572
rect 212 27364 246 27380
rect -200 27287 -184 27321
rect 184 27287 200 27321
rect -200 27179 -184 27213
rect 184 27179 200 27213
rect -246 27120 -212 27136
rect -246 26928 -212 26944
rect 212 27120 246 27136
rect 212 26928 246 26944
rect -200 26851 -184 26885
rect 184 26851 200 26885
rect -200 26743 -184 26777
rect 184 26743 200 26777
rect -246 26684 -212 26700
rect -246 26492 -212 26508
rect 212 26684 246 26700
rect 212 26492 246 26508
rect -200 26415 -184 26449
rect 184 26415 200 26449
rect -200 26307 -184 26341
rect 184 26307 200 26341
rect -246 26248 -212 26264
rect -246 26056 -212 26072
rect 212 26248 246 26264
rect 212 26056 246 26072
rect -200 25979 -184 26013
rect 184 25979 200 26013
rect -200 25871 -184 25905
rect 184 25871 200 25905
rect -246 25812 -212 25828
rect -246 25620 -212 25636
rect 212 25812 246 25828
rect 212 25620 246 25636
rect -200 25543 -184 25577
rect 184 25543 200 25577
rect -200 25435 -184 25469
rect 184 25435 200 25469
rect -246 25376 -212 25392
rect -246 25184 -212 25200
rect 212 25376 246 25392
rect 212 25184 246 25200
rect -200 25107 -184 25141
rect 184 25107 200 25141
rect -200 24999 -184 25033
rect 184 24999 200 25033
rect -246 24940 -212 24956
rect -246 24748 -212 24764
rect 212 24940 246 24956
rect 212 24748 246 24764
rect -200 24671 -184 24705
rect 184 24671 200 24705
rect -200 24563 -184 24597
rect 184 24563 200 24597
rect -246 24504 -212 24520
rect -246 24312 -212 24328
rect 212 24504 246 24520
rect 212 24312 246 24328
rect -200 24235 -184 24269
rect 184 24235 200 24269
rect -200 24127 -184 24161
rect 184 24127 200 24161
rect -246 24068 -212 24084
rect -246 23876 -212 23892
rect 212 24068 246 24084
rect 212 23876 246 23892
rect -200 23799 -184 23833
rect 184 23799 200 23833
rect -200 23691 -184 23725
rect 184 23691 200 23725
rect -246 23632 -212 23648
rect -246 23440 -212 23456
rect 212 23632 246 23648
rect 212 23440 246 23456
rect -200 23363 -184 23397
rect 184 23363 200 23397
rect -200 23255 -184 23289
rect 184 23255 200 23289
rect -246 23196 -212 23212
rect -246 23004 -212 23020
rect 212 23196 246 23212
rect 212 23004 246 23020
rect -200 22927 -184 22961
rect 184 22927 200 22961
rect -200 22819 -184 22853
rect 184 22819 200 22853
rect -246 22760 -212 22776
rect -246 22568 -212 22584
rect 212 22760 246 22776
rect 212 22568 246 22584
rect -200 22491 -184 22525
rect 184 22491 200 22525
rect -200 22383 -184 22417
rect 184 22383 200 22417
rect -246 22324 -212 22340
rect -246 22132 -212 22148
rect 212 22324 246 22340
rect 212 22132 246 22148
rect -200 22055 -184 22089
rect 184 22055 200 22089
rect -200 21947 -184 21981
rect 184 21947 200 21981
rect -246 21888 -212 21904
rect -246 21696 -212 21712
rect 212 21888 246 21904
rect 212 21696 246 21712
rect -200 21619 -184 21653
rect 184 21619 200 21653
rect -200 21511 -184 21545
rect 184 21511 200 21545
rect -246 21452 -212 21468
rect -246 21260 -212 21276
rect 212 21452 246 21468
rect 212 21260 246 21276
rect -200 21183 -184 21217
rect 184 21183 200 21217
rect -200 21075 -184 21109
rect 184 21075 200 21109
rect -246 21016 -212 21032
rect -246 20824 -212 20840
rect 212 21016 246 21032
rect 212 20824 246 20840
rect -200 20747 -184 20781
rect 184 20747 200 20781
rect -200 20639 -184 20673
rect 184 20639 200 20673
rect -246 20580 -212 20596
rect -246 20388 -212 20404
rect 212 20580 246 20596
rect 212 20388 246 20404
rect -200 20311 -184 20345
rect 184 20311 200 20345
rect -200 20203 -184 20237
rect 184 20203 200 20237
rect -246 20144 -212 20160
rect -246 19952 -212 19968
rect 212 20144 246 20160
rect 212 19952 246 19968
rect -200 19875 -184 19909
rect 184 19875 200 19909
rect -200 19767 -184 19801
rect 184 19767 200 19801
rect -246 19708 -212 19724
rect -246 19516 -212 19532
rect 212 19708 246 19724
rect 212 19516 246 19532
rect -200 19439 -184 19473
rect 184 19439 200 19473
rect -200 19331 -184 19365
rect 184 19331 200 19365
rect -246 19272 -212 19288
rect -246 19080 -212 19096
rect 212 19272 246 19288
rect 212 19080 246 19096
rect -200 19003 -184 19037
rect 184 19003 200 19037
rect -200 18895 -184 18929
rect 184 18895 200 18929
rect -246 18836 -212 18852
rect -246 18644 -212 18660
rect 212 18836 246 18852
rect 212 18644 246 18660
rect -200 18567 -184 18601
rect 184 18567 200 18601
rect -200 18459 -184 18493
rect 184 18459 200 18493
rect -246 18400 -212 18416
rect -246 18208 -212 18224
rect 212 18400 246 18416
rect 212 18208 246 18224
rect -200 18131 -184 18165
rect 184 18131 200 18165
rect -200 18023 -184 18057
rect 184 18023 200 18057
rect -246 17964 -212 17980
rect -246 17772 -212 17788
rect 212 17964 246 17980
rect 212 17772 246 17788
rect -200 17695 -184 17729
rect 184 17695 200 17729
rect -200 17587 -184 17621
rect 184 17587 200 17621
rect -246 17528 -212 17544
rect -246 17336 -212 17352
rect 212 17528 246 17544
rect 212 17336 246 17352
rect -200 17259 -184 17293
rect 184 17259 200 17293
rect -200 17151 -184 17185
rect 184 17151 200 17185
rect -246 17092 -212 17108
rect -246 16900 -212 16916
rect 212 17092 246 17108
rect 212 16900 246 16916
rect -200 16823 -184 16857
rect 184 16823 200 16857
rect -200 16715 -184 16749
rect 184 16715 200 16749
rect -246 16656 -212 16672
rect -246 16464 -212 16480
rect 212 16656 246 16672
rect 212 16464 246 16480
rect -200 16387 -184 16421
rect 184 16387 200 16421
rect -200 16279 -184 16313
rect 184 16279 200 16313
rect -246 16220 -212 16236
rect -246 16028 -212 16044
rect 212 16220 246 16236
rect 212 16028 246 16044
rect -200 15951 -184 15985
rect 184 15951 200 15985
rect -200 15843 -184 15877
rect 184 15843 200 15877
rect -246 15784 -212 15800
rect -246 15592 -212 15608
rect 212 15784 246 15800
rect 212 15592 246 15608
rect -200 15515 -184 15549
rect 184 15515 200 15549
rect -200 15407 -184 15441
rect 184 15407 200 15441
rect -246 15348 -212 15364
rect -246 15156 -212 15172
rect 212 15348 246 15364
rect 212 15156 246 15172
rect -200 15079 -184 15113
rect 184 15079 200 15113
rect -200 14971 -184 15005
rect 184 14971 200 15005
rect -246 14912 -212 14928
rect -246 14720 -212 14736
rect 212 14912 246 14928
rect 212 14720 246 14736
rect -200 14643 -184 14677
rect 184 14643 200 14677
rect -200 14535 -184 14569
rect 184 14535 200 14569
rect -246 14476 -212 14492
rect -246 14284 -212 14300
rect 212 14476 246 14492
rect 212 14284 246 14300
rect -200 14207 -184 14241
rect 184 14207 200 14241
rect -200 14099 -184 14133
rect 184 14099 200 14133
rect -246 14040 -212 14056
rect -246 13848 -212 13864
rect 212 14040 246 14056
rect 212 13848 246 13864
rect -200 13771 -184 13805
rect 184 13771 200 13805
rect -200 13663 -184 13697
rect 184 13663 200 13697
rect -246 13604 -212 13620
rect -246 13412 -212 13428
rect 212 13604 246 13620
rect 212 13412 246 13428
rect -200 13335 -184 13369
rect 184 13335 200 13369
rect -200 13227 -184 13261
rect 184 13227 200 13261
rect -246 13168 -212 13184
rect -246 12976 -212 12992
rect 212 13168 246 13184
rect 212 12976 246 12992
rect -200 12899 -184 12933
rect 184 12899 200 12933
rect -200 12791 -184 12825
rect 184 12791 200 12825
rect -246 12732 -212 12748
rect -246 12540 -212 12556
rect 212 12732 246 12748
rect 212 12540 246 12556
rect -200 12463 -184 12497
rect 184 12463 200 12497
rect -200 12355 -184 12389
rect 184 12355 200 12389
rect -246 12296 -212 12312
rect -246 12104 -212 12120
rect 212 12296 246 12312
rect 212 12104 246 12120
rect -200 12027 -184 12061
rect 184 12027 200 12061
rect -200 11919 -184 11953
rect 184 11919 200 11953
rect -246 11860 -212 11876
rect -246 11668 -212 11684
rect 212 11860 246 11876
rect 212 11668 246 11684
rect -200 11591 -184 11625
rect 184 11591 200 11625
rect -200 11483 -184 11517
rect 184 11483 200 11517
rect -246 11424 -212 11440
rect -246 11232 -212 11248
rect 212 11424 246 11440
rect 212 11232 246 11248
rect -200 11155 -184 11189
rect 184 11155 200 11189
rect -200 11047 -184 11081
rect 184 11047 200 11081
rect -246 10988 -212 11004
rect -246 10796 -212 10812
rect 212 10988 246 11004
rect 212 10796 246 10812
rect -200 10719 -184 10753
rect 184 10719 200 10753
rect -200 10611 -184 10645
rect 184 10611 200 10645
rect -246 10552 -212 10568
rect -246 10360 -212 10376
rect 212 10552 246 10568
rect 212 10360 246 10376
rect -200 10283 -184 10317
rect 184 10283 200 10317
rect -200 10175 -184 10209
rect 184 10175 200 10209
rect -246 10116 -212 10132
rect -246 9924 -212 9940
rect 212 10116 246 10132
rect 212 9924 246 9940
rect -200 9847 -184 9881
rect 184 9847 200 9881
rect -200 9739 -184 9773
rect 184 9739 200 9773
rect -246 9680 -212 9696
rect -246 9488 -212 9504
rect 212 9680 246 9696
rect 212 9488 246 9504
rect -200 9411 -184 9445
rect 184 9411 200 9445
rect -200 9303 -184 9337
rect 184 9303 200 9337
rect -246 9244 -212 9260
rect -246 9052 -212 9068
rect 212 9244 246 9260
rect 212 9052 246 9068
rect -200 8975 -184 9009
rect 184 8975 200 9009
rect -200 8867 -184 8901
rect 184 8867 200 8901
rect -246 8808 -212 8824
rect -246 8616 -212 8632
rect 212 8808 246 8824
rect 212 8616 246 8632
rect -200 8539 -184 8573
rect 184 8539 200 8573
rect -200 8431 -184 8465
rect 184 8431 200 8465
rect -246 8372 -212 8388
rect -246 8180 -212 8196
rect 212 8372 246 8388
rect 212 8180 246 8196
rect -200 8103 -184 8137
rect 184 8103 200 8137
rect -200 7995 -184 8029
rect 184 7995 200 8029
rect -246 7936 -212 7952
rect -246 7744 -212 7760
rect 212 7936 246 7952
rect 212 7744 246 7760
rect -200 7667 -184 7701
rect 184 7667 200 7701
rect -200 7559 -184 7593
rect 184 7559 200 7593
rect -246 7500 -212 7516
rect -246 7308 -212 7324
rect 212 7500 246 7516
rect 212 7308 246 7324
rect -200 7231 -184 7265
rect 184 7231 200 7265
rect -200 7123 -184 7157
rect 184 7123 200 7157
rect -246 7064 -212 7080
rect -246 6872 -212 6888
rect 212 7064 246 7080
rect 212 6872 246 6888
rect -200 6795 -184 6829
rect 184 6795 200 6829
rect -200 6687 -184 6721
rect 184 6687 200 6721
rect -246 6628 -212 6644
rect -246 6436 -212 6452
rect 212 6628 246 6644
rect 212 6436 246 6452
rect -200 6359 -184 6393
rect 184 6359 200 6393
rect -200 6251 -184 6285
rect 184 6251 200 6285
rect -246 6192 -212 6208
rect -246 6000 -212 6016
rect 212 6192 246 6208
rect 212 6000 246 6016
rect -200 5923 -184 5957
rect 184 5923 200 5957
rect -200 5815 -184 5849
rect 184 5815 200 5849
rect -246 5756 -212 5772
rect -246 5564 -212 5580
rect 212 5756 246 5772
rect 212 5564 246 5580
rect -200 5487 -184 5521
rect 184 5487 200 5521
rect -200 5379 -184 5413
rect 184 5379 200 5413
rect -246 5320 -212 5336
rect -246 5128 -212 5144
rect 212 5320 246 5336
rect 212 5128 246 5144
rect -200 5051 -184 5085
rect 184 5051 200 5085
rect -200 4943 -184 4977
rect 184 4943 200 4977
rect -246 4884 -212 4900
rect -246 4692 -212 4708
rect 212 4884 246 4900
rect 212 4692 246 4708
rect -200 4615 -184 4649
rect 184 4615 200 4649
rect -200 4507 -184 4541
rect 184 4507 200 4541
rect -246 4448 -212 4464
rect -246 4256 -212 4272
rect 212 4448 246 4464
rect 212 4256 246 4272
rect -200 4179 -184 4213
rect 184 4179 200 4213
rect -200 4071 -184 4105
rect 184 4071 200 4105
rect -246 4012 -212 4028
rect -246 3820 -212 3836
rect 212 4012 246 4028
rect 212 3820 246 3836
rect -200 3743 -184 3777
rect 184 3743 200 3777
rect -200 3635 -184 3669
rect 184 3635 200 3669
rect -246 3576 -212 3592
rect -246 3384 -212 3400
rect 212 3576 246 3592
rect 212 3384 246 3400
rect -200 3307 -184 3341
rect 184 3307 200 3341
rect -200 3199 -184 3233
rect 184 3199 200 3233
rect -246 3140 -212 3156
rect -246 2948 -212 2964
rect 212 3140 246 3156
rect 212 2948 246 2964
rect -200 2871 -184 2905
rect 184 2871 200 2905
rect -200 2763 -184 2797
rect 184 2763 200 2797
rect -246 2704 -212 2720
rect -246 2512 -212 2528
rect 212 2704 246 2720
rect 212 2512 246 2528
rect -200 2435 -184 2469
rect 184 2435 200 2469
rect -200 2327 -184 2361
rect 184 2327 200 2361
rect -246 2268 -212 2284
rect -246 2076 -212 2092
rect 212 2268 246 2284
rect 212 2076 246 2092
rect -200 1999 -184 2033
rect 184 1999 200 2033
rect -200 1891 -184 1925
rect 184 1891 200 1925
rect -246 1832 -212 1848
rect -246 1640 -212 1656
rect 212 1832 246 1848
rect 212 1640 246 1656
rect -200 1563 -184 1597
rect 184 1563 200 1597
rect -200 1455 -184 1489
rect 184 1455 200 1489
rect -246 1396 -212 1412
rect -246 1204 -212 1220
rect 212 1396 246 1412
rect 212 1204 246 1220
rect -200 1127 -184 1161
rect 184 1127 200 1161
rect -200 1019 -184 1053
rect 184 1019 200 1053
rect -246 960 -212 976
rect -246 768 -212 784
rect 212 960 246 976
rect 212 768 246 784
rect -200 691 -184 725
rect 184 691 200 725
rect -200 583 -184 617
rect 184 583 200 617
rect -246 524 -212 540
rect -246 332 -212 348
rect 212 524 246 540
rect 212 332 246 348
rect -200 255 -184 289
rect 184 255 200 289
rect -200 147 -184 181
rect 184 147 200 181
rect -246 88 -212 104
rect -246 -104 -212 -88
rect 212 88 246 104
rect 212 -104 246 -88
rect -200 -181 -184 -147
rect 184 -181 200 -147
rect -200 -289 -184 -255
rect 184 -289 200 -255
rect -246 -348 -212 -332
rect -246 -540 -212 -524
rect 212 -348 246 -332
rect 212 -540 246 -524
rect -200 -617 -184 -583
rect 184 -617 200 -583
rect -200 -725 -184 -691
rect 184 -725 200 -691
rect -246 -784 -212 -768
rect -246 -976 -212 -960
rect 212 -784 246 -768
rect 212 -976 246 -960
rect -200 -1053 -184 -1019
rect 184 -1053 200 -1019
rect -200 -1161 -184 -1127
rect 184 -1161 200 -1127
rect -246 -1220 -212 -1204
rect -246 -1412 -212 -1396
rect 212 -1220 246 -1204
rect 212 -1412 246 -1396
rect -200 -1489 -184 -1455
rect 184 -1489 200 -1455
rect -200 -1597 -184 -1563
rect 184 -1597 200 -1563
rect -246 -1656 -212 -1640
rect -246 -1848 -212 -1832
rect 212 -1656 246 -1640
rect 212 -1848 246 -1832
rect -200 -1925 -184 -1891
rect 184 -1925 200 -1891
rect -200 -2033 -184 -1999
rect 184 -2033 200 -1999
rect -246 -2092 -212 -2076
rect -246 -2284 -212 -2268
rect 212 -2092 246 -2076
rect 212 -2284 246 -2268
rect -200 -2361 -184 -2327
rect 184 -2361 200 -2327
rect -200 -2469 -184 -2435
rect 184 -2469 200 -2435
rect -246 -2528 -212 -2512
rect -246 -2720 -212 -2704
rect 212 -2528 246 -2512
rect 212 -2720 246 -2704
rect -200 -2797 -184 -2763
rect 184 -2797 200 -2763
rect -200 -2905 -184 -2871
rect 184 -2905 200 -2871
rect -246 -2964 -212 -2948
rect -246 -3156 -212 -3140
rect 212 -2964 246 -2948
rect 212 -3156 246 -3140
rect -200 -3233 -184 -3199
rect 184 -3233 200 -3199
rect -200 -3341 -184 -3307
rect 184 -3341 200 -3307
rect -246 -3400 -212 -3384
rect -246 -3592 -212 -3576
rect 212 -3400 246 -3384
rect 212 -3592 246 -3576
rect -200 -3669 -184 -3635
rect 184 -3669 200 -3635
rect -200 -3777 -184 -3743
rect 184 -3777 200 -3743
rect -246 -3836 -212 -3820
rect -246 -4028 -212 -4012
rect 212 -3836 246 -3820
rect 212 -4028 246 -4012
rect -200 -4105 -184 -4071
rect 184 -4105 200 -4071
rect -200 -4213 -184 -4179
rect 184 -4213 200 -4179
rect -246 -4272 -212 -4256
rect -246 -4464 -212 -4448
rect 212 -4272 246 -4256
rect 212 -4464 246 -4448
rect -200 -4541 -184 -4507
rect 184 -4541 200 -4507
rect -200 -4649 -184 -4615
rect 184 -4649 200 -4615
rect -246 -4708 -212 -4692
rect -246 -4900 -212 -4884
rect 212 -4708 246 -4692
rect 212 -4900 246 -4884
rect -200 -4977 -184 -4943
rect 184 -4977 200 -4943
rect -200 -5085 -184 -5051
rect 184 -5085 200 -5051
rect -246 -5144 -212 -5128
rect -246 -5336 -212 -5320
rect 212 -5144 246 -5128
rect 212 -5336 246 -5320
rect -200 -5413 -184 -5379
rect 184 -5413 200 -5379
rect -200 -5521 -184 -5487
rect 184 -5521 200 -5487
rect -246 -5580 -212 -5564
rect -246 -5772 -212 -5756
rect 212 -5580 246 -5564
rect 212 -5772 246 -5756
rect -200 -5849 -184 -5815
rect 184 -5849 200 -5815
rect -200 -5957 -184 -5923
rect 184 -5957 200 -5923
rect -246 -6016 -212 -6000
rect -246 -6208 -212 -6192
rect 212 -6016 246 -6000
rect 212 -6208 246 -6192
rect -200 -6285 -184 -6251
rect 184 -6285 200 -6251
rect -200 -6393 -184 -6359
rect 184 -6393 200 -6359
rect -246 -6452 -212 -6436
rect -246 -6644 -212 -6628
rect 212 -6452 246 -6436
rect 212 -6644 246 -6628
rect -200 -6721 -184 -6687
rect 184 -6721 200 -6687
rect -200 -6829 -184 -6795
rect 184 -6829 200 -6795
rect -246 -6888 -212 -6872
rect -246 -7080 -212 -7064
rect 212 -6888 246 -6872
rect 212 -7080 246 -7064
rect -200 -7157 -184 -7123
rect 184 -7157 200 -7123
rect -200 -7265 -184 -7231
rect 184 -7265 200 -7231
rect -246 -7324 -212 -7308
rect -246 -7516 -212 -7500
rect 212 -7324 246 -7308
rect 212 -7516 246 -7500
rect -200 -7593 -184 -7559
rect 184 -7593 200 -7559
rect -200 -7701 -184 -7667
rect 184 -7701 200 -7667
rect -246 -7760 -212 -7744
rect -246 -7952 -212 -7936
rect 212 -7760 246 -7744
rect 212 -7952 246 -7936
rect -200 -8029 -184 -7995
rect 184 -8029 200 -7995
rect -200 -8137 -184 -8103
rect 184 -8137 200 -8103
rect -246 -8196 -212 -8180
rect -246 -8388 -212 -8372
rect 212 -8196 246 -8180
rect 212 -8388 246 -8372
rect -200 -8465 -184 -8431
rect 184 -8465 200 -8431
rect -200 -8573 -184 -8539
rect 184 -8573 200 -8539
rect -246 -8632 -212 -8616
rect -246 -8824 -212 -8808
rect 212 -8632 246 -8616
rect 212 -8824 246 -8808
rect -200 -8901 -184 -8867
rect 184 -8901 200 -8867
rect -200 -9009 -184 -8975
rect 184 -9009 200 -8975
rect -246 -9068 -212 -9052
rect -246 -9260 -212 -9244
rect 212 -9068 246 -9052
rect 212 -9260 246 -9244
rect -200 -9337 -184 -9303
rect 184 -9337 200 -9303
rect -200 -9445 -184 -9411
rect 184 -9445 200 -9411
rect -246 -9504 -212 -9488
rect -246 -9696 -212 -9680
rect 212 -9504 246 -9488
rect 212 -9696 246 -9680
rect -200 -9773 -184 -9739
rect 184 -9773 200 -9739
rect -200 -9881 -184 -9847
rect 184 -9881 200 -9847
rect -246 -9940 -212 -9924
rect -246 -10132 -212 -10116
rect 212 -9940 246 -9924
rect 212 -10132 246 -10116
rect -200 -10209 -184 -10175
rect 184 -10209 200 -10175
rect -200 -10317 -184 -10283
rect 184 -10317 200 -10283
rect -246 -10376 -212 -10360
rect -246 -10568 -212 -10552
rect 212 -10376 246 -10360
rect 212 -10568 246 -10552
rect -200 -10645 -184 -10611
rect 184 -10645 200 -10611
rect -200 -10753 -184 -10719
rect 184 -10753 200 -10719
rect -246 -10812 -212 -10796
rect -246 -11004 -212 -10988
rect 212 -10812 246 -10796
rect 212 -11004 246 -10988
rect -200 -11081 -184 -11047
rect 184 -11081 200 -11047
rect -200 -11189 -184 -11155
rect 184 -11189 200 -11155
rect -246 -11248 -212 -11232
rect -246 -11440 -212 -11424
rect 212 -11248 246 -11232
rect 212 -11440 246 -11424
rect -200 -11517 -184 -11483
rect 184 -11517 200 -11483
rect -200 -11625 -184 -11591
rect 184 -11625 200 -11591
rect -246 -11684 -212 -11668
rect -246 -11876 -212 -11860
rect 212 -11684 246 -11668
rect 212 -11876 246 -11860
rect -200 -11953 -184 -11919
rect 184 -11953 200 -11919
rect -200 -12061 -184 -12027
rect 184 -12061 200 -12027
rect -246 -12120 -212 -12104
rect -246 -12312 -212 -12296
rect 212 -12120 246 -12104
rect 212 -12312 246 -12296
rect -200 -12389 -184 -12355
rect 184 -12389 200 -12355
rect -200 -12497 -184 -12463
rect 184 -12497 200 -12463
rect -246 -12556 -212 -12540
rect -246 -12748 -212 -12732
rect 212 -12556 246 -12540
rect 212 -12748 246 -12732
rect -200 -12825 -184 -12791
rect 184 -12825 200 -12791
rect -200 -12933 -184 -12899
rect 184 -12933 200 -12899
rect -246 -12992 -212 -12976
rect -246 -13184 -212 -13168
rect 212 -12992 246 -12976
rect 212 -13184 246 -13168
rect -200 -13261 -184 -13227
rect 184 -13261 200 -13227
rect -200 -13369 -184 -13335
rect 184 -13369 200 -13335
rect -246 -13428 -212 -13412
rect -246 -13620 -212 -13604
rect 212 -13428 246 -13412
rect 212 -13620 246 -13604
rect -200 -13697 -184 -13663
rect 184 -13697 200 -13663
rect -200 -13805 -184 -13771
rect 184 -13805 200 -13771
rect -246 -13864 -212 -13848
rect -246 -14056 -212 -14040
rect 212 -13864 246 -13848
rect 212 -14056 246 -14040
rect -200 -14133 -184 -14099
rect 184 -14133 200 -14099
rect -200 -14241 -184 -14207
rect 184 -14241 200 -14207
rect -246 -14300 -212 -14284
rect -246 -14492 -212 -14476
rect 212 -14300 246 -14284
rect 212 -14492 246 -14476
rect -200 -14569 -184 -14535
rect 184 -14569 200 -14535
rect -200 -14677 -184 -14643
rect 184 -14677 200 -14643
rect -246 -14736 -212 -14720
rect -246 -14928 -212 -14912
rect 212 -14736 246 -14720
rect 212 -14928 246 -14912
rect -200 -15005 -184 -14971
rect 184 -15005 200 -14971
rect -200 -15113 -184 -15079
rect 184 -15113 200 -15079
rect -246 -15172 -212 -15156
rect -246 -15364 -212 -15348
rect 212 -15172 246 -15156
rect 212 -15364 246 -15348
rect -200 -15441 -184 -15407
rect 184 -15441 200 -15407
rect -200 -15549 -184 -15515
rect 184 -15549 200 -15515
rect -246 -15608 -212 -15592
rect -246 -15800 -212 -15784
rect 212 -15608 246 -15592
rect 212 -15800 246 -15784
rect -200 -15877 -184 -15843
rect 184 -15877 200 -15843
rect -200 -15985 -184 -15951
rect 184 -15985 200 -15951
rect -246 -16044 -212 -16028
rect -246 -16236 -212 -16220
rect 212 -16044 246 -16028
rect 212 -16236 246 -16220
rect -200 -16313 -184 -16279
rect 184 -16313 200 -16279
rect -200 -16421 -184 -16387
rect 184 -16421 200 -16387
rect -246 -16480 -212 -16464
rect -246 -16672 -212 -16656
rect 212 -16480 246 -16464
rect 212 -16672 246 -16656
rect -200 -16749 -184 -16715
rect 184 -16749 200 -16715
rect -200 -16857 -184 -16823
rect 184 -16857 200 -16823
rect -246 -16916 -212 -16900
rect -246 -17108 -212 -17092
rect 212 -16916 246 -16900
rect 212 -17108 246 -17092
rect -200 -17185 -184 -17151
rect 184 -17185 200 -17151
rect -200 -17293 -184 -17259
rect 184 -17293 200 -17259
rect -246 -17352 -212 -17336
rect -246 -17544 -212 -17528
rect 212 -17352 246 -17336
rect 212 -17544 246 -17528
rect -200 -17621 -184 -17587
rect 184 -17621 200 -17587
rect -200 -17729 -184 -17695
rect 184 -17729 200 -17695
rect -246 -17788 -212 -17772
rect -246 -17980 -212 -17964
rect 212 -17788 246 -17772
rect 212 -17980 246 -17964
rect -200 -18057 -184 -18023
rect 184 -18057 200 -18023
rect -200 -18165 -184 -18131
rect 184 -18165 200 -18131
rect -246 -18224 -212 -18208
rect -246 -18416 -212 -18400
rect 212 -18224 246 -18208
rect 212 -18416 246 -18400
rect -200 -18493 -184 -18459
rect 184 -18493 200 -18459
rect -200 -18601 -184 -18567
rect 184 -18601 200 -18567
rect -246 -18660 -212 -18644
rect -246 -18852 -212 -18836
rect 212 -18660 246 -18644
rect 212 -18852 246 -18836
rect -200 -18929 -184 -18895
rect 184 -18929 200 -18895
rect -200 -19037 -184 -19003
rect 184 -19037 200 -19003
rect -246 -19096 -212 -19080
rect -246 -19288 -212 -19272
rect 212 -19096 246 -19080
rect 212 -19288 246 -19272
rect -200 -19365 -184 -19331
rect 184 -19365 200 -19331
rect -200 -19473 -184 -19439
rect 184 -19473 200 -19439
rect -246 -19532 -212 -19516
rect -246 -19724 -212 -19708
rect 212 -19532 246 -19516
rect 212 -19724 246 -19708
rect -200 -19801 -184 -19767
rect 184 -19801 200 -19767
rect -200 -19909 -184 -19875
rect 184 -19909 200 -19875
rect -246 -19968 -212 -19952
rect -246 -20160 -212 -20144
rect 212 -19968 246 -19952
rect 212 -20160 246 -20144
rect -200 -20237 -184 -20203
rect 184 -20237 200 -20203
rect -200 -20345 -184 -20311
rect 184 -20345 200 -20311
rect -246 -20404 -212 -20388
rect -246 -20596 -212 -20580
rect 212 -20404 246 -20388
rect 212 -20596 246 -20580
rect -200 -20673 -184 -20639
rect 184 -20673 200 -20639
rect -200 -20781 -184 -20747
rect 184 -20781 200 -20747
rect -246 -20840 -212 -20824
rect -246 -21032 -212 -21016
rect 212 -20840 246 -20824
rect 212 -21032 246 -21016
rect -200 -21109 -184 -21075
rect 184 -21109 200 -21075
rect -200 -21217 -184 -21183
rect 184 -21217 200 -21183
rect -246 -21276 -212 -21260
rect -246 -21468 -212 -21452
rect 212 -21276 246 -21260
rect 212 -21468 246 -21452
rect -200 -21545 -184 -21511
rect 184 -21545 200 -21511
rect -200 -21653 -184 -21619
rect 184 -21653 200 -21619
rect -246 -21712 -212 -21696
rect -246 -21904 -212 -21888
rect 212 -21712 246 -21696
rect 212 -21904 246 -21888
rect -200 -21981 -184 -21947
rect 184 -21981 200 -21947
rect -200 -22089 -184 -22055
rect 184 -22089 200 -22055
rect -246 -22148 -212 -22132
rect -246 -22340 -212 -22324
rect 212 -22148 246 -22132
rect 212 -22340 246 -22324
rect -200 -22417 -184 -22383
rect 184 -22417 200 -22383
rect -200 -22525 -184 -22491
rect 184 -22525 200 -22491
rect -246 -22584 -212 -22568
rect -246 -22776 -212 -22760
rect 212 -22584 246 -22568
rect 212 -22776 246 -22760
rect -200 -22853 -184 -22819
rect 184 -22853 200 -22819
rect -200 -22961 -184 -22927
rect 184 -22961 200 -22927
rect -246 -23020 -212 -23004
rect -246 -23212 -212 -23196
rect 212 -23020 246 -23004
rect 212 -23212 246 -23196
rect -200 -23289 -184 -23255
rect 184 -23289 200 -23255
rect -200 -23397 -184 -23363
rect 184 -23397 200 -23363
rect -246 -23456 -212 -23440
rect -246 -23648 -212 -23632
rect 212 -23456 246 -23440
rect 212 -23648 246 -23632
rect -200 -23725 -184 -23691
rect 184 -23725 200 -23691
rect -200 -23833 -184 -23799
rect 184 -23833 200 -23799
rect -246 -23892 -212 -23876
rect -246 -24084 -212 -24068
rect 212 -23892 246 -23876
rect 212 -24084 246 -24068
rect -200 -24161 -184 -24127
rect 184 -24161 200 -24127
rect -200 -24269 -184 -24235
rect 184 -24269 200 -24235
rect -246 -24328 -212 -24312
rect -246 -24520 -212 -24504
rect 212 -24328 246 -24312
rect 212 -24520 246 -24504
rect -200 -24597 -184 -24563
rect 184 -24597 200 -24563
rect -200 -24705 -184 -24671
rect 184 -24705 200 -24671
rect -246 -24764 -212 -24748
rect -246 -24956 -212 -24940
rect 212 -24764 246 -24748
rect 212 -24956 246 -24940
rect -200 -25033 -184 -24999
rect 184 -25033 200 -24999
rect -200 -25141 -184 -25107
rect 184 -25141 200 -25107
rect -246 -25200 -212 -25184
rect -246 -25392 -212 -25376
rect 212 -25200 246 -25184
rect 212 -25392 246 -25376
rect -200 -25469 -184 -25435
rect 184 -25469 200 -25435
rect -200 -25577 -184 -25543
rect 184 -25577 200 -25543
rect -246 -25636 -212 -25620
rect -246 -25828 -212 -25812
rect 212 -25636 246 -25620
rect 212 -25828 246 -25812
rect -200 -25905 -184 -25871
rect 184 -25905 200 -25871
rect -200 -26013 -184 -25979
rect 184 -26013 200 -25979
rect -246 -26072 -212 -26056
rect -246 -26264 -212 -26248
rect 212 -26072 246 -26056
rect 212 -26264 246 -26248
rect -200 -26341 -184 -26307
rect 184 -26341 200 -26307
rect -200 -26449 -184 -26415
rect 184 -26449 200 -26415
rect -246 -26508 -212 -26492
rect -246 -26700 -212 -26684
rect 212 -26508 246 -26492
rect 212 -26700 246 -26684
rect -200 -26777 -184 -26743
rect 184 -26777 200 -26743
rect -200 -26885 -184 -26851
rect 184 -26885 200 -26851
rect -246 -26944 -212 -26928
rect -246 -27136 -212 -27120
rect 212 -26944 246 -26928
rect 212 -27136 246 -27120
rect -200 -27213 -184 -27179
rect 184 -27213 200 -27179
rect -200 -27321 -184 -27287
rect 184 -27321 200 -27287
rect -246 -27380 -212 -27364
rect -246 -27572 -212 -27556
rect 212 -27380 246 -27364
rect 212 -27572 246 -27556
rect -200 -27649 -184 -27615
rect 184 -27649 200 -27615
rect -200 -27757 -184 -27723
rect 184 -27757 200 -27723
rect -246 -27816 -212 -27800
rect -246 -28008 -212 -27992
rect 212 -27816 246 -27800
rect 212 -28008 246 -27992
rect -200 -28085 -184 -28051
rect 184 -28085 200 -28051
rect -200 -28193 -184 -28159
rect 184 -28193 200 -28159
rect -246 -28252 -212 -28236
rect -246 -28444 -212 -28428
rect 212 -28252 246 -28236
rect 212 -28444 246 -28428
rect -200 -28521 -184 -28487
rect 184 -28521 200 -28487
rect -200 -28629 -184 -28595
rect 184 -28629 200 -28595
rect -246 -28688 -212 -28672
rect -246 -28880 -212 -28864
rect 212 -28688 246 -28672
rect 212 -28880 246 -28864
rect -200 -28957 -184 -28923
rect 184 -28957 200 -28923
rect -200 -29065 -184 -29031
rect 184 -29065 200 -29031
rect -246 -29124 -212 -29108
rect -246 -29316 -212 -29300
rect 212 -29124 246 -29108
rect 212 -29316 246 -29300
rect -200 -29393 -184 -29359
rect 184 -29393 200 -29359
rect -200 -29501 -184 -29467
rect 184 -29501 200 -29467
rect -246 -29560 -212 -29544
rect -246 -29752 -212 -29736
rect 212 -29560 246 -29544
rect 212 -29752 246 -29736
rect -200 -29829 -184 -29795
rect 184 -29829 200 -29795
rect -200 -29937 -184 -29903
rect 184 -29937 200 -29903
rect -246 -29996 -212 -29980
rect -246 -30188 -212 -30172
rect 212 -29996 246 -29980
rect 212 -30188 246 -30172
rect -200 -30265 -184 -30231
rect 184 -30265 200 -30231
rect -200 -30373 -184 -30339
rect 184 -30373 200 -30339
rect -246 -30432 -212 -30416
rect -246 -30624 -212 -30608
rect 212 -30432 246 -30416
rect 212 -30624 246 -30608
rect -200 -30701 -184 -30667
rect 184 -30701 200 -30667
rect -200 -30809 -184 -30775
rect 184 -30809 200 -30775
rect -246 -30868 -212 -30852
rect -246 -31060 -212 -31044
rect 212 -30868 246 -30852
rect 212 -31060 246 -31044
rect -200 -31137 -184 -31103
rect 184 -31137 200 -31103
rect -200 -31245 -184 -31211
rect 184 -31245 200 -31211
rect -246 -31304 -212 -31288
rect -246 -31496 -212 -31480
rect 212 -31304 246 -31288
rect 212 -31496 246 -31480
rect -200 -31573 -184 -31539
rect 184 -31573 200 -31539
rect -200 -31681 -184 -31647
rect 184 -31681 200 -31647
rect -246 -31740 -212 -31724
rect -246 -31932 -212 -31916
rect 212 -31740 246 -31724
rect 212 -31932 246 -31916
rect -200 -32009 -184 -31975
rect 184 -32009 200 -31975
rect -200 -32117 -184 -32083
rect 184 -32117 200 -32083
rect -246 -32176 -212 -32160
rect -246 -32368 -212 -32352
rect 212 -32176 246 -32160
rect 212 -32368 246 -32352
rect -200 -32445 -184 -32411
rect 184 -32445 200 -32411
rect -200 -32553 -184 -32519
rect 184 -32553 200 -32519
rect -246 -32612 -212 -32596
rect -246 -32804 -212 -32788
rect 212 -32612 246 -32596
rect 212 -32804 246 -32788
rect -200 -32881 -184 -32847
rect 184 -32881 200 -32847
rect -200 -32989 -184 -32955
rect 184 -32989 200 -32955
rect -246 -33048 -212 -33032
rect -246 -33240 -212 -33224
rect 212 -33048 246 -33032
rect 212 -33240 246 -33224
rect -200 -33317 -184 -33283
rect 184 -33317 200 -33283
rect -200 -33425 -184 -33391
rect 184 -33425 200 -33391
rect -246 -33484 -212 -33468
rect -246 -33676 -212 -33660
rect 212 -33484 246 -33468
rect 212 -33676 246 -33660
rect -200 -33753 -184 -33719
rect 184 -33753 200 -33719
rect -200 -33861 -184 -33827
rect 184 -33861 200 -33827
rect -246 -33920 -212 -33904
rect -246 -34112 -212 -34096
rect 212 -33920 246 -33904
rect 212 -34112 246 -34096
rect -200 -34189 -184 -34155
rect 184 -34189 200 -34155
rect -200 -34297 -184 -34263
rect 184 -34297 200 -34263
rect -246 -34356 -212 -34340
rect -246 -34548 -212 -34532
rect 212 -34356 246 -34340
rect 212 -34548 246 -34532
rect -200 -34625 -184 -34591
rect 184 -34625 200 -34591
rect -200 -34733 -184 -34699
rect 184 -34733 200 -34699
rect -246 -34792 -212 -34776
rect -246 -34984 -212 -34968
rect 212 -34792 246 -34776
rect 212 -34984 246 -34968
rect -200 -35061 -184 -35027
rect 184 -35061 200 -35027
rect -200 -35169 -184 -35135
rect 184 -35169 200 -35135
rect -246 -35228 -212 -35212
rect -246 -35420 -212 -35404
rect 212 -35228 246 -35212
rect 212 -35420 246 -35404
rect -200 -35497 -184 -35463
rect 184 -35497 200 -35463
rect -200 -35605 -184 -35571
rect 184 -35605 200 -35571
rect -246 -35664 -212 -35648
rect -246 -35856 -212 -35840
rect 212 -35664 246 -35648
rect 212 -35856 246 -35840
rect -200 -35933 -184 -35899
rect 184 -35933 200 -35899
rect -200 -36041 -184 -36007
rect 184 -36041 200 -36007
rect -246 -36100 -212 -36084
rect -246 -36292 -212 -36276
rect 212 -36100 246 -36084
rect 212 -36292 246 -36276
rect -200 -36369 -184 -36335
rect 184 -36369 200 -36335
rect -200 -36477 -184 -36443
rect 184 -36477 200 -36443
rect -246 -36536 -212 -36520
rect -246 -36728 -212 -36712
rect 212 -36536 246 -36520
rect 212 -36728 246 -36712
rect -200 -36805 -184 -36771
rect 184 -36805 200 -36771
rect -200 -36913 -184 -36879
rect 184 -36913 200 -36879
rect -246 -36972 -212 -36956
rect -246 -37164 -212 -37148
rect 212 -36972 246 -36956
rect 212 -37164 246 -37148
rect -200 -37241 -184 -37207
rect 184 -37241 200 -37207
rect -200 -37349 -184 -37315
rect 184 -37349 200 -37315
rect -246 -37408 -212 -37392
rect -246 -37600 -212 -37584
rect 212 -37408 246 -37392
rect 212 -37600 246 -37584
rect -200 -37677 -184 -37643
rect 184 -37677 200 -37643
rect -200 -37785 -184 -37751
rect 184 -37785 200 -37751
rect -246 -37844 -212 -37828
rect -246 -38036 -212 -38020
rect 212 -37844 246 -37828
rect 212 -38036 246 -38020
rect -200 -38113 -184 -38079
rect 184 -38113 200 -38079
rect -200 -38221 -184 -38187
rect 184 -38221 200 -38187
rect -246 -38280 -212 -38264
rect -246 -38472 -212 -38456
rect 212 -38280 246 -38264
rect 212 -38472 246 -38456
rect -200 -38549 -184 -38515
rect 184 -38549 200 -38515
rect -200 -38657 -184 -38623
rect 184 -38657 200 -38623
rect -246 -38716 -212 -38700
rect -246 -38908 -212 -38892
rect 212 -38716 246 -38700
rect 212 -38908 246 -38892
rect -200 -38985 -184 -38951
rect 184 -38985 200 -38951
rect -200 -39093 -184 -39059
rect 184 -39093 200 -39059
rect -246 -39152 -212 -39136
rect -246 -39344 -212 -39328
rect 212 -39152 246 -39136
rect 212 -39344 246 -39328
rect -200 -39421 -184 -39387
rect 184 -39421 200 -39387
rect -200 -39529 -184 -39495
rect 184 -39529 200 -39495
rect -246 -39588 -212 -39572
rect -246 -39780 -212 -39764
rect 212 -39588 246 -39572
rect 212 -39780 246 -39764
rect -200 -39857 -184 -39823
rect 184 -39857 200 -39823
rect -200 -39965 -184 -39931
rect 184 -39965 200 -39931
rect -246 -40024 -212 -40008
rect -246 -40216 -212 -40200
rect 212 -40024 246 -40008
rect 212 -40216 246 -40200
rect -200 -40293 -184 -40259
rect 184 -40293 200 -40259
rect -200 -40401 -184 -40367
rect 184 -40401 200 -40367
rect -246 -40460 -212 -40444
rect -246 -40652 -212 -40636
rect 212 -40460 246 -40444
rect 212 -40652 246 -40636
rect -200 -40729 -184 -40695
rect 184 -40729 200 -40695
rect -200 -40837 -184 -40803
rect 184 -40837 200 -40803
rect -246 -40896 -212 -40880
rect -246 -41088 -212 -41072
rect 212 -40896 246 -40880
rect 212 -41088 246 -41072
rect -200 -41165 -184 -41131
rect 184 -41165 200 -41131
rect -200 -41273 -184 -41239
rect 184 -41273 200 -41239
rect -246 -41332 -212 -41316
rect -246 -41524 -212 -41508
rect 212 -41332 246 -41316
rect 212 -41524 246 -41508
rect -200 -41601 -184 -41567
rect 184 -41601 200 -41567
rect -200 -41709 -184 -41675
rect 184 -41709 200 -41675
rect -246 -41768 -212 -41752
rect -246 -41960 -212 -41944
rect 212 -41768 246 -41752
rect 212 -41960 246 -41944
rect -200 -42037 -184 -42003
rect 184 -42037 200 -42003
rect -200 -42145 -184 -42111
rect 184 -42145 200 -42111
rect -246 -42204 -212 -42188
rect -246 -42396 -212 -42380
rect 212 -42204 246 -42188
rect 212 -42396 246 -42380
rect -200 -42473 -184 -42439
rect 184 -42473 200 -42439
rect -200 -42581 -184 -42547
rect 184 -42581 200 -42547
rect -246 -42640 -212 -42624
rect -246 -42832 -212 -42816
rect 212 -42640 246 -42624
rect 212 -42832 246 -42816
rect -200 -42909 -184 -42875
rect 184 -42909 200 -42875
rect -200 -43017 -184 -42983
rect 184 -43017 200 -42983
rect -246 -43076 -212 -43060
rect -246 -43268 -212 -43252
rect 212 -43076 246 -43060
rect 212 -43268 246 -43252
rect -200 -43345 -184 -43311
rect 184 -43345 200 -43311
rect -200 -43453 -184 -43419
rect 184 -43453 200 -43419
rect -246 -43512 -212 -43496
rect -246 -43704 -212 -43688
rect 212 -43512 246 -43496
rect 212 -43704 246 -43688
rect -200 -43781 -184 -43747
rect 184 -43781 200 -43747
rect -200 -43889 -184 -43855
rect 184 -43889 200 -43855
rect -246 -43948 -212 -43932
rect -246 -44140 -212 -44124
rect 212 -43948 246 -43932
rect 212 -44140 246 -44124
rect -200 -44217 -184 -44183
rect 184 -44217 200 -44183
rect -200 -44325 -184 -44291
rect 184 -44325 200 -44291
rect -246 -44384 -212 -44368
rect -246 -44576 -212 -44560
rect 212 -44384 246 -44368
rect 212 -44576 246 -44560
rect -200 -44653 -184 -44619
rect 184 -44653 200 -44619
rect -200 -44761 -184 -44727
rect 184 -44761 200 -44727
rect -246 -44820 -212 -44804
rect -246 -45012 -212 -44996
rect 212 -44820 246 -44804
rect 212 -45012 246 -44996
rect -200 -45089 -184 -45055
rect 184 -45089 200 -45055
rect -200 -45197 -184 -45163
rect 184 -45197 200 -45163
rect -246 -45256 -212 -45240
rect -246 -45448 -212 -45432
rect 212 -45256 246 -45240
rect 212 -45448 246 -45432
rect -200 -45525 -184 -45491
rect 184 -45525 200 -45491
rect -200 -45633 -184 -45599
rect 184 -45633 200 -45599
rect -246 -45692 -212 -45676
rect -246 -45884 -212 -45868
rect 212 -45692 246 -45676
rect 212 -45884 246 -45868
rect -200 -45961 -184 -45927
rect 184 -45961 200 -45927
rect -200 -46069 -184 -46035
rect 184 -46069 200 -46035
rect -246 -46128 -212 -46112
rect -246 -46320 -212 -46304
rect 212 -46128 246 -46112
rect 212 -46320 246 -46304
rect -200 -46397 -184 -46363
rect 184 -46397 200 -46363
rect -200 -46505 -184 -46471
rect 184 -46505 200 -46471
rect -246 -46564 -212 -46548
rect -246 -46756 -212 -46740
rect 212 -46564 246 -46548
rect 212 -46756 246 -46740
rect -200 -46833 -184 -46799
rect 184 -46833 200 -46799
rect -200 -46941 -184 -46907
rect 184 -46941 200 -46907
rect -246 -47000 -212 -46984
rect -246 -47192 -212 -47176
rect 212 -47000 246 -46984
rect 212 -47192 246 -47176
rect -200 -47269 -184 -47235
rect 184 -47269 200 -47235
rect -200 -47377 -184 -47343
rect 184 -47377 200 -47343
rect -246 -47436 -212 -47420
rect -246 -47628 -212 -47612
rect 212 -47436 246 -47420
rect 212 -47628 246 -47612
rect -200 -47705 -184 -47671
rect 184 -47705 200 -47671
rect -200 -47813 -184 -47779
rect 184 -47813 200 -47779
rect -246 -47872 -212 -47856
rect -246 -48064 -212 -48048
rect 212 -47872 246 -47856
rect 212 -48064 246 -48048
rect -200 -48141 -184 -48107
rect 184 -48141 200 -48107
rect -200 -48249 -184 -48215
rect 184 -48249 200 -48215
rect -246 -48308 -212 -48292
rect -246 -48500 -212 -48484
rect 212 -48308 246 -48292
rect 212 -48500 246 -48484
rect -200 -48577 -184 -48543
rect 184 -48577 200 -48543
rect -200 -48685 -184 -48651
rect 184 -48685 200 -48651
rect -246 -48744 -212 -48728
rect -246 -48936 -212 -48920
rect 212 -48744 246 -48728
rect 212 -48936 246 -48920
rect -200 -49013 -184 -48979
rect 184 -49013 200 -48979
rect -200 -49121 -184 -49087
rect 184 -49121 200 -49087
rect -246 -49180 -212 -49164
rect -246 -49372 -212 -49356
rect 212 -49180 246 -49164
rect 212 -49372 246 -49356
rect -200 -49449 -184 -49415
rect 184 -49449 200 -49415
rect -200 -49557 -184 -49523
rect 184 -49557 200 -49523
rect -246 -49616 -212 -49600
rect -246 -49808 -212 -49792
rect 212 -49616 246 -49600
rect 212 -49808 246 -49792
rect -200 -49885 -184 -49851
rect 184 -49885 200 -49851
rect -200 -49993 -184 -49959
rect 184 -49993 200 -49959
rect -246 -50052 -212 -50036
rect -246 -50244 -212 -50228
rect 212 -50052 246 -50036
rect 212 -50244 246 -50228
rect -200 -50321 -184 -50287
rect 184 -50321 200 -50287
rect -200 -50429 -184 -50395
rect 184 -50429 200 -50395
rect -246 -50488 -212 -50472
rect -246 -50680 -212 -50664
rect 212 -50488 246 -50472
rect 212 -50680 246 -50664
rect -200 -50757 -184 -50723
rect 184 -50757 200 -50723
rect -200 -50865 -184 -50831
rect 184 -50865 200 -50831
rect -246 -50924 -212 -50908
rect -246 -51116 -212 -51100
rect 212 -50924 246 -50908
rect 212 -51116 246 -51100
rect -200 -51193 -184 -51159
rect 184 -51193 200 -51159
rect -200 -51301 -184 -51267
rect 184 -51301 200 -51267
rect -246 -51360 -212 -51344
rect -246 -51552 -212 -51536
rect 212 -51360 246 -51344
rect 212 -51552 246 -51536
rect -200 -51629 -184 -51595
rect 184 -51629 200 -51595
rect -200 -51737 -184 -51703
rect 184 -51737 200 -51703
rect -246 -51796 -212 -51780
rect -246 -51988 -212 -51972
rect 212 -51796 246 -51780
rect 212 -51988 246 -51972
rect -200 -52065 -184 -52031
rect 184 -52065 200 -52031
rect -200 -52173 -184 -52139
rect 184 -52173 200 -52139
rect -246 -52232 -212 -52216
rect -246 -52424 -212 -52408
rect 212 -52232 246 -52216
rect 212 -52424 246 -52408
rect -200 -52501 -184 -52467
rect 184 -52501 200 -52467
rect -200 -52609 -184 -52575
rect 184 -52609 200 -52575
rect -246 -52668 -212 -52652
rect -246 -52860 -212 -52844
rect 212 -52668 246 -52652
rect 212 -52860 246 -52844
rect -200 -52937 -184 -52903
rect 184 -52937 200 -52903
rect -200 -53045 -184 -53011
rect 184 -53045 200 -53011
rect -246 -53104 -212 -53088
rect -246 -53296 -212 -53280
rect 212 -53104 246 -53088
rect 212 -53296 246 -53280
rect -200 -53373 -184 -53339
rect 184 -53373 200 -53339
rect -200 -53481 -184 -53447
rect 184 -53481 200 -53447
rect -246 -53540 -212 -53524
rect -246 -53732 -212 -53716
rect 212 -53540 246 -53524
rect 212 -53732 246 -53716
rect -200 -53809 -184 -53775
rect 184 -53809 200 -53775
rect -200 -53917 -184 -53883
rect 184 -53917 200 -53883
rect -246 -53976 -212 -53960
rect -246 -54168 -212 -54152
rect 212 -53976 246 -53960
rect 212 -54168 246 -54152
rect -200 -54245 -184 -54211
rect 184 -54245 200 -54211
rect -200 -54353 -184 -54319
rect 184 -54353 200 -54319
rect -246 -54412 -212 -54396
rect -246 -54604 -212 -54588
rect 212 -54412 246 -54396
rect 212 -54604 246 -54588
rect -200 -54681 -184 -54647
rect 184 -54681 200 -54647
rect -200 -54789 -184 -54755
rect 184 -54789 200 -54755
rect -246 -54848 -212 -54832
rect -246 -55040 -212 -55024
rect 212 -54848 246 -54832
rect 212 -55040 246 -55024
rect -200 -55117 -184 -55083
rect 184 -55117 200 -55083
rect -200 -55225 -184 -55191
rect 184 -55225 200 -55191
rect -246 -55284 -212 -55268
rect -246 -55476 -212 -55460
rect 212 -55284 246 -55268
rect 212 -55476 246 -55460
rect -200 -55553 -184 -55519
rect 184 -55553 200 -55519
rect -200 -55661 -184 -55627
rect 184 -55661 200 -55627
rect -246 -55720 -212 -55704
rect -246 -55912 -212 -55896
rect 212 -55720 246 -55704
rect 212 -55912 246 -55896
rect -200 -55989 -184 -55955
rect 184 -55989 200 -55955
rect -200 -56097 -184 -56063
rect 184 -56097 200 -56063
rect -246 -56156 -212 -56140
rect -246 -56348 -212 -56332
rect 212 -56156 246 -56140
rect 212 -56348 246 -56332
rect -200 -56425 -184 -56391
rect 184 -56425 200 -56391
rect -200 -56533 -184 -56499
rect 184 -56533 200 -56499
rect -246 -56592 -212 -56576
rect -246 -56784 -212 -56768
rect 212 -56592 246 -56576
rect 212 -56784 246 -56768
rect -200 -56861 -184 -56827
rect 184 -56861 200 -56827
rect -200 -56969 -184 -56935
rect 184 -56969 200 -56935
rect -246 -57028 -212 -57012
rect -246 -57220 -212 -57204
rect 212 -57028 246 -57012
rect 212 -57220 246 -57204
rect -200 -57297 -184 -57263
rect 184 -57297 200 -57263
rect -200 -57405 -184 -57371
rect 184 -57405 200 -57371
rect -246 -57464 -212 -57448
rect -246 -57656 -212 -57640
rect 212 -57464 246 -57448
rect 212 -57656 246 -57640
rect -200 -57733 -184 -57699
rect 184 -57733 200 -57699
rect -200 -57841 -184 -57807
rect 184 -57841 200 -57807
rect -246 -57900 -212 -57884
rect -246 -58092 -212 -58076
rect 212 -57900 246 -57884
rect 212 -58092 246 -58076
rect -200 -58169 -184 -58135
rect 184 -58169 200 -58135
rect -200 -58277 -184 -58243
rect 184 -58277 200 -58243
rect -246 -58336 -212 -58320
rect -246 -58528 -212 -58512
rect 212 -58336 246 -58320
rect 212 -58528 246 -58512
rect -200 -58605 -184 -58571
rect 184 -58605 200 -58571
rect -200 -58713 -184 -58679
rect 184 -58713 200 -58679
rect -246 -58772 -212 -58756
rect -246 -58964 -212 -58948
rect 212 -58772 246 -58756
rect 212 -58964 246 -58948
rect -200 -59041 -184 -59007
rect 184 -59041 200 -59007
rect -200 -59149 -184 -59115
rect 184 -59149 200 -59115
rect -246 -59208 -212 -59192
rect -246 -59400 -212 -59384
rect 212 -59208 246 -59192
rect 212 -59400 246 -59384
rect -200 -59477 -184 -59443
rect 184 -59477 200 -59443
rect -200 -59585 -184 -59551
rect 184 -59585 200 -59551
rect -246 -59644 -212 -59628
rect -246 -59836 -212 -59820
rect 212 -59644 246 -59628
rect 212 -59836 246 -59820
rect -200 -59913 -184 -59879
rect 184 -59913 200 -59879
rect -200 -60021 -184 -59987
rect 184 -60021 200 -59987
rect -246 -60080 -212 -60064
rect -246 -60272 -212 -60256
rect 212 -60080 246 -60064
rect 212 -60272 246 -60256
rect -200 -60349 -184 -60315
rect 184 -60349 200 -60315
rect -200 -60457 -184 -60423
rect 184 -60457 200 -60423
rect -246 -60516 -212 -60500
rect -246 -60708 -212 -60692
rect 212 -60516 246 -60500
rect 212 -60708 246 -60692
rect -200 -60785 -184 -60751
rect 184 -60785 200 -60751
rect -200 -60893 -184 -60859
rect 184 -60893 200 -60859
rect -246 -60952 -212 -60936
rect -246 -61144 -212 -61128
rect 212 -60952 246 -60936
rect 212 -61144 246 -61128
rect -200 -61221 -184 -61187
rect 184 -61221 200 -61187
rect -200 -61329 -184 -61295
rect 184 -61329 200 -61295
rect -246 -61388 -212 -61372
rect -246 -61580 -212 -61564
rect 212 -61388 246 -61372
rect 212 -61580 246 -61564
rect -200 -61657 -184 -61623
rect 184 -61657 200 -61623
rect -200 -61765 -184 -61731
rect 184 -61765 200 -61731
rect -246 -61824 -212 -61808
rect -246 -62016 -212 -62000
rect 212 -61824 246 -61808
rect 212 -62016 246 -62000
rect -200 -62093 -184 -62059
rect 184 -62093 200 -62059
rect -200 -62201 -184 -62167
rect 184 -62201 200 -62167
rect -246 -62260 -212 -62244
rect -246 -62452 -212 -62436
rect 212 -62260 246 -62244
rect 212 -62452 246 -62436
rect -200 -62529 -184 -62495
rect 184 -62529 200 -62495
rect -200 -62637 -184 -62603
rect 184 -62637 200 -62603
rect -246 -62696 -212 -62680
rect -246 -62888 -212 -62872
rect 212 -62696 246 -62680
rect 212 -62888 246 -62872
rect -200 -62965 -184 -62931
rect 184 -62965 200 -62931
rect -200 -63073 -184 -63039
rect 184 -63073 200 -63039
rect -246 -63132 -212 -63116
rect -246 -63324 -212 -63308
rect 212 -63132 246 -63116
rect 212 -63324 246 -63308
rect -200 -63401 -184 -63367
rect 184 -63401 200 -63367
rect -200 -63509 -184 -63475
rect 184 -63509 200 -63475
rect -246 -63568 -212 -63552
rect -246 -63760 -212 -63744
rect 212 -63568 246 -63552
rect 212 -63760 246 -63744
rect -200 -63837 -184 -63803
rect 184 -63837 200 -63803
rect -200 -63945 -184 -63911
rect 184 -63945 200 -63911
rect -246 -64004 -212 -63988
rect -246 -64196 -212 -64180
rect 212 -64004 246 -63988
rect 212 -64196 246 -64180
rect -200 -64273 -184 -64239
rect 184 -64273 200 -64239
rect -200 -64381 -184 -64347
rect 184 -64381 200 -64347
rect -246 -64440 -212 -64424
rect -246 -64632 -212 -64616
rect 212 -64440 246 -64424
rect 212 -64632 246 -64616
rect -200 -64709 -184 -64675
rect 184 -64709 200 -64675
rect -200 -64817 -184 -64783
rect 184 -64817 200 -64783
rect -246 -64876 -212 -64860
rect -246 -65068 -212 -65052
rect 212 -64876 246 -64860
rect 212 -65068 246 -65052
rect -200 -65145 -184 -65111
rect 184 -65145 200 -65111
rect -200 -65253 -184 -65219
rect 184 -65253 200 -65219
rect -246 -65312 -212 -65296
rect -246 -65504 -212 -65488
rect 212 -65312 246 -65296
rect 212 -65504 246 -65488
rect -200 -65581 -184 -65547
rect 184 -65581 200 -65547
rect -200 -65689 -184 -65655
rect 184 -65689 200 -65655
rect -246 -65748 -212 -65732
rect -246 -65940 -212 -65924
rect 212 -65748 246 -65732
rect 212 -65940 246 -65924
rect -200 -66017 -184 -65983
rect 184 -66017 200 -65983
rect -200 -66125 -184 -66091
rect 184 -66125 200 -66091
rect -246 -66184 -212 -66168
rect -246 -66376 -212 -66360
rect 212 -66184 246 -66168
rect 212 -66376 246 -66360
rect -200 -66453 -184 -66419
rect 184 -66453 200 -66419
rect -200 -66561 -184 -66527
rect 184 -66561 200 -66527
rect -246 -66620 -212 -66604
rect -246 -66812 -212 -66796
rect 212 -66620 246 -66604
rect 212 -66812 246 -66796
rect -200 -66889 -184 -66855
rect 184 -66889 200 -66855
rect -200 -66997 -184 -66963
rect 184 -66997 200 -66963
rect -246 -67056 -212 -67040
rect -246 -67248 -212 -67232
rect 212 -67056 246 -67040
rect 212 -67248 246 -67232
rect -200 -67325 -184 -67291
rect 184 -67325 200 -67291
rect -200 -67433 -184 -67399
rect 184 -67433 200 -67399
rect -246 -67492 -212 -67476
rect -246 -67684 -212 -67668
rect 212 -67492 246 -67476
rect 212 -67684 246 -67668
rect -200 -67761 -184 -67727
rect 184 -67761 200 -67727
rect -200 -67869 -184 -67835
rect 184 -67869 200 -67835
rect -246 -67928 -212 -67912
rect -246 -68120 -212 -68104
rect 212 -67928 246 -67912
rect 212 -68120 246 -68104
rect -200 -68197 -184 -68163
rect 184 -68197 200 -68163
rect -200 -68305 -184 -68271
rect 184 -68305 200 -68271
rect -246 -68364 -212 -68348
rect -246 -68556 -212 -68540
rect 212 -68364 246 -68348
rect 212 -68556 246 -68540
rect -200 -68633 -184 -68599
rect 184 -68633 200 -68599
rect -200 -68741 -184 -68707
rect 184 -68741 200 -68707
rect -246 -68800 -212 -68784
rect -246 -68992 -212 -68976
rect 212 -68800 246 -68784
rect 212 -68992 246 -68976
rect -200 -69069 -184 -69035
rect 184 -69069 200 -69035
rect -200 -69177 -184 -69143
rect 184 -69177 200 -69143
rect -246 -69236 -212 -69220
rect -246 -69428 -212 -69412
rect 212 -69236 246 -69220
rect 212 -69428 246 -69412
rect -200 -69505 -184 -69471
rect 184 -69505 200 -69471
rect -200 -69613 -184 -69579
rect 184 -69613 200 -69579
rect -246 -69672 -212 -69656
rect -246 -69864 -212 -69848
rect 212 -69672 246 -69656
rect 212 -69864 246 -69848
rect -200 -69941 -184 -69907
rect 184 -69941 200 -69907
rect -200 -70049 -184 -70015
rect 184 -70049 200 -70015
rect -246 -70108 -212 -70092
rect -246 -70300 -212 -70284
rect 212 -70108 246 -70092
rect 212 -70300 246 -70284
rect -200 -70377 -184 -70343
rect 184 -70377 200 -70343
rect -200 -70485 -184 -70451
rect 184 -70485 200 -70451
rect -246 -70544 -212 -70528
rect -246 -70736 -212 -70720
rect 212 -70544 246 -70528
rect 212 -70736 246 -70720
rect -200 -70813 -184 -70779
rect 184 -70813 200 -70779
rect -200 -70921 -184 -70887
rect 184 -70921 200 -70887
rect -246 -70980 -212 -70964
rect -246 -71172 -212 -71156
rect 212 -70980 246 -70964
rect 212 -71172 246 -71156
rect -200 -71249 -184 -71215
rect 184 -71249 200 -71215
rect -200 -71357 -184 -71323
rect 184 -71357 200 -71323
rect -246 -71416 -212 -71400
rect -246 -71608 -212 -71592
rect 212 -71416 246 -71400
rect 212 -71608 246 -71592
rect -200 -71685 -184 -71651
rect 184 -71685 200 -71651
rect -200 -71793 -184 -71759
rect 184 -71793 200 -71759
rect -246 -71852 -212 -71836
rect -246 -72044 -212 -72028
rect 212 -71852 246 -71836
rect 212 -72044 246 -72028
rect -200 -72121 -184 -72087
rect 184 -72121 200 -72087
rect -200 -72229 -184 -72195
rect 184 -72229 200 -72195
rect -246 -72288 -212 -72272
rect -246 -72480 -212 -72464
rect 212 -72288 246 -72272
rect 212 -72480 246 -72464
rect -200 -72557 -184 -72523
rect 184 -72557 200 -72523
rect -200 -72665 -184 -72631
rect 184 -72665 200 -72631
rect -246 -72724 -212 -72708
rect -246 -72916 -212 -72900
rect 212 -72724 246 -72708
rect 212 -72916 246 -72900
rect -200 -72993 -184 -72959
rect 184 -72993 200 -72959
rect -200 -73101 -184 -73067
rect 184 -73101 200 -73067
rect -246 -73160 -212 -73144
rect -246 -73352 -212 -73336
rect 212 -73160 246 -73144
rect 212 -73352 246 -73336
rect -200 -73429 -184 -73395
rect 184 -73429 200 -73395
rect -200 -73537 -184 -73503
rect 184 -73537 200 -73503
rect -246 -73596 -212 -73580
rect -246 -73788 -212 -73772
rect 212 -73596 246 -73580
rect 212 -73788 246 -73772
rect -200 -73865 -184 -73831
rect 184 -73865 200 -73831
rect -200 -73973 -184 -73939
rect 184 -73973 200 -73939
rect -246 -74032 -212 -74016
rect -246 -74224 -212 -74208
rect 212 -74032 246 -74016
rect 212 -74224 246 -74208
rect -200 -74301 -184 -74267
rect 184 -74301 200 -74267
rect -200 -74409 -184 -74375
rect 184 -74409 200 -74375
rect -246 -74468 -212 -74452
rect -246 -74660 -212 -74644
rect 212 -74468 246 -74452
rect 212 -74660 246 -74644
rect -200 -74737 -184 -74703
rect 184 -74737 200 -74703
rect -200 -74845 -184 -74811
rect 184 -74845 200 -74811
rect -246 -74904 -212 -74888
rect -246 -75096 -212 -75080
rect 212 -74904 246 -74888
rect 212 -75096 246 -75080
rect -200 -75173 -184 -75139
rect 184 -75173 200 -75139
rect -200 -75281 -184 -75247
rect 184 -75281 200 -75247
rect -246 -75340 -212 -75324
rect -246 -75532 -212 -75516
rect 212 -75340 246 -75324
rect 212 -75532 246 -75516
rect -200 -75609 -184 -75575
rect 184 -75609 200 -75575
rect -200 -75717 -184 -75683
rect 184 -75717 200 -75683
rect -246 -75776 -212 -75760
rect -246 -75968 -212 -75952
rect 212 -75776 246 -75760
rect 212 -75968 246 -75952
rect -200 -76045 -184 -76011
rect 184 -76045 200 -76011
rect -200 -76153 -184 -76119
rect 184 -76153 200 -76119
rect -246 -76212 -212 -76196
rect -246 -76404 -212 -76388
rect 212 -76212 246 -76196
rect 212 -76404 246 -76388
rect -200 -76481 -184 -76447
rect 184 -76481 200 -76447
rect -200 -76589 -184 -76555
rect 184 -76589 200 -76555
rect -246 -76648 -212 -76632
rect -246 -76840 -212 -76824
rect 212 -76648 246 -76632
rect 212 -76840 246 -76824
rect -200 -76917 -184 -76883
rect 184 -76917 200 -76883
rect -200 -77025 -184 -76991
rect 184 -77025 200 -76991
rect -246 -77084 -212 -77068
rect -246 -77276 -212 -77260
rect 212 -77084 246 -77068
rect 212 -77276 246 -77260
rect -200 -77353 -184 -77319
rect 184 -77353 200 -77319
rect -200 -77461 -184 -77427
rect 184 -77461 200 -77427
rect -246 -77520 -212 -77504
rect -246 -77712 -212 -77696
rect 212 -77520 246 -77504
rect 212 -77712 246 -77696
rect -200 -77789 -184 -77755
rect 184 -77789 200 -77755
rect -200 -77897 -184 -77863
rect 184 -77897 200 -77863
rect -246 -77956 -212 -77940
rect -246 -78148 -212 -78132
rect 212 -77956 246 -77940
rect 212 -78148 246 -78132
rect -200 -78225 -184 -78191
rect 184 -78225 200 -78191
rect -200 -78333 -184 -78299
rect 184 -78333 200 -78299
rect -246 -78392 -212 -78376
rect -246 -78584 -212 -78568
rect 212 -78392 246 -78376
rect 212 -78584 246 -78568
rect -200 -78661 -184 -78627
rect 184 -78661 200 -78627
rect -200 -78769 -184 -78735
rect 184 -78769 200 -78735
rect -246 -78828 -212 -78812
rect -246 -79020 -212 -79004
rect 212 -78828 246 -78812
rect 212 -79020 246 -79004
rect -200 -79097 -184 -79063
rect 184 -79097 200 -79063
rect -200 -79205 -184 -79171
rect 184 -79205 200 -79171
rect -246 -79264 -212 -79248
rect -246 -79456 -212 -79440
rect 212 -79264 246 -79248
rect 212 -79456 246 -79440
rect -200 -79533 -184 -79499
rect 184 -79533 200 -79499
rect -200 -79641 -184 -79607
rect 184 -79641 200 -79607
rect -246 -79700 -212 -79684
rect -246 -79892 -212 -79876
rect 212 -79700 246 -79684
rect 212 -79892 246 -79876
rect -200 -79969 -184 -79935
rect 184 -79969 200 -79935
rect -200 -80077 -184 -80043
rect 184 -80077 200 -80043
rect -246 -80136 -212 -80120
rect -246 -80328 -212 -80312
rect 212 -80136 246 -80120
rect 212 -80328 246 -80312
rect -200 -80405 -184 -80371
rect 184 -80405 200 -80371
rect -200 -80513 -184 -80479
rect 184 -80513 200 -80479
rect -246 -80572 -212 -80556
rect -246 -80764 -212 -80748
rect 212 -80572 246 -80556
rect 212 -80764 246 -80748
rect -200 -80841 -184 -80807
rect 184 -80841 200 -80807
rect -200 -80949 -184 -80915
rect 184 -80949 200 -80915
rect -246 -81008 -212 -80992
rect -246 -81200 -212 -81184
rect 212 -81008 246 -80992
rect 212 -81200 246 -81184
rect -200 -81277 -184 -81243
rect 184 -81277 200 -81243
rect -200 -81385 -184 -81351
rect 184 -81385 200 -81351
rect -246 -81444 -212 -81428
rect -246 -81636 -212 -81620
rect 212 -81444 246 -81428
rect 212 -81636 246 -81620
rect -200 -81713 -184 -81679
rect 184 -81713 200 -81679
rect -200 -81821 -184 -81787
rect 184 -81821 200 -81787
rect -246 -81880 -212 -81864
rect -246 -82072 -212 -82056
rect 212 -81880 246 -81864
rect 212 -82072 246 -82056
rect -200 -82149 -184 -82115
rect 184 -82149 200 -82115
rect -200 -82257 -184 -82223
rect 184 -82257 200 -82223
rect -246 -82316 -212 -82300
rect -246 -82508 -212 -82492
rect 212 -82316 246 -82300
rect 212 -82508 246 -82492
rect -200 -82585 -184 -82551
rect 184 -82585 200 -82551
rect -200 -82693 -184 -82659
rect 184 -82693 200 -82659
rect -246 -82752 -212 -82736
rect -246 -82944 -212 -82928
rect 212 -82752 246 -82736
rect 212 -82944 246 -82928
rect -200 -83021 -184 -82987
rect 184 -83021 200 -82987
rect -200 -83129 -184 -83095
rect 184 -83129 200 -83095
rect -246 -83188 -212 -83172
rect -246 -83380 -212 -83364
rect 212 -83188 246 -83172
rect 212 -83380 246 -83364
rect -200 -83457 -184 -83423
rect 184 -83457 200 -83423
rect -200 -83565 -184 -83531
rect 184 -83565 200 -83531
rect -246 -83624 -212 -83608
rect -246 -83816 -212 -83800
rect 212 -83624 246 -83608
rect 212 -83816 246 -83800
rect -200 -83893 -184 -83859
rect 184 -83893 200 -83859
rect -200 -84001 -184 -83967
rect 184 -84001 200 -83967
rect -246 -84060 -212 -84044
rect -246 -84252 -212 -84236
rect 212 -84060 246 -84044
rect 212 -84252 246 -84236
rect -200 -84329 -184 -84295
rect 184 -84329 200 -84295
rect -360 -84397 -326 -84335
rect 326 -84397 360 -84335
rect -360 -84431 -264 -84397
rect 264 -84431 360 -84397
<< viali >>
rect -184 84295 184 84329
rect -246 84060 -212 84236
rect 212 84060 246 84236
rect -184 83967 184 84001
rect -184 83859 184 83893
rect -246 83624 -212 83800
rect 212 83624 246 83800
rect -184 83531 184 83565
rect -184 83423 184 83457
rect -246 83188 -212 83364
rect 212 83188 246 83364
rect -184 83095 184 83129
rect -184 82987 184 83021
rect -246 82752 -212 82928
rect 212 82752 246 82928
rect -184 82659 184 82693
rect -184 82551 184 82585
rect -246 82316 -212 82492
rect 212 82316 246 82492
rect -184 82223 184 82257
rect -184 82115 184 82149
rect -246 81880 -212 82056
rect 212 81880 246 82056
rect -184 81787 184 81821
rect -184 81679 184 81713
rect -246 81444 -212 81620
rect 212 81444 246 81620
rect -184 81351 184 81385
rect -184 81243 184 81277
rect -246 81008 -212 81184
rect 212 81008 246 81184
rect -184 80915 184 80949
rect -184 80807 184 80841
rect -246 80572 -212 80748
rect 212 80572 246 80748
rect -184 80479 184 80513
rect -184 80371 184 80405
rect -246 80136 -212 80312
rect 212 80136 246 80312
rect -184 80043 184 80077
rect -184 79935 184 79969
rect -246 79700 -212 79876
rect 212 79700 246 79876
rect -184 79607 184 79641
rect -184 79499 184 79533
rect -246 79264 -212 79440
rect 212 79264 246 79440
rect -184 79171 184 79205
rect -184 79063 184 79097
rect -246 78828 -212 79004
rect 212 78828 246 79004
rect -184 78735 184 78769
rect -184 78627 184 78661
rect -246 78392 -212 78568
rect 212 78392 246 78568
rect -184 78299 184 78333
rect -184 78191 184 78225
rect -246 77956 -212 78132
rect 212 77956 246 78132
rect -184 77863 184 77897
rect -184 77755 184 77789
rect -246 77520 -212 77696
rect 212 77520 246 77696
rect -184 77427 184 77461
rect -184 77319 184 77353
rect -246 77084 -212 77260
rect 212 77084 246 77260
rect -184 76991 184 77025
rect -184 76883 184 76917
rect -246 76648 -212 76824
rect 212 76648 246 76824
rect -184 76555 184 76589
rect -184 76447 184 76481
rect -246 76212 -212 76388
rect 212 76212 246 76388
rect -184 76119 184 76153
rect -184 76011 184 76045
rect -246 75776 -212 75952
rect 212 75776 246 75952
rect -184 75683 184 75717
rect -184 75575 184 75609
rect -246 75340 -212 75516
rect 212 75340 246 75516
rect -184 75247 184 75281
rect -184 75139 184 75173
rect -246 74904 -212 75080
rect 212 74904 246 75080
rect -184 74811 184 74845
rect -184 74703 184 74737
rect -246 74468 -212 74644
rect 212 74468 246 74644
rect -184 74375 184 74409
rect -184 74267 184 74301
rect -246 74032 -212 74208
rect 212 74032 246 74208
rect -184 73939 184 73973
rect -184 73831 184 73865
rect -246 73596 -212 73772
rect 212 73596 246 73772
rect -184 73503 184 73537
rect -184 73395 184 73429
rect -246 73160 -212 73336
rect 212 73160 246 73336
rect -184 73067 184 73101
rect -184 72959 184 72993
rect -246 72724 -212 72900
rect 212 72724 246 72900
rect -184 72631 184 72665
rect -184 72523 184 72557
rect -246 72288 -212 72464
rect 212 72288 246 72464
rect -184 72195 184 72229
rect -184 72087 184 72121
rect -246 71852 -212 72028
rect 212 71852 246 72028
rect -184 71759 184 71793
rect -184 71651 184 71685
rect -246 71416 -212 71592
rect 212 71416 246 71592
rect -184 71323 184 71357
rect -184 71215 184 71249
rect -246 70980 -212 71156
rect 212 70980 246 71156
rect -184 70887 184 70921
rect -184 70779 184 70813
rect -246 70544 -212 70720
rect 212 70544 246 70720
rect -184 70451 184 70485
rect -184 70343 184 70377
rect -246 70108 -212 70284
rect 212 70108 246 70284
rect -184 70015 184 70049
rect -184 69907 184 69941
rect -246 69672 -212 69848
rect 212 69672 246 69848
rect -184 69579 184 69613
rect -184 69471 184 69505
rect -246 69236 -212 69412
rect 212 69236 246 69412
rect -184 69143 184 69177
rect -184 69035 184 69069
rect -246 68800 -212 68976
rect 212 68800 246 68976
rect -184 68707 184 68741
rect -184 68599 184 68633
rect -246 68364 -212 68540
rect 212 68364 246 68540
rect -184 68271 184 68305
rect -184 68163 184 68197
rect -246 67928 -212 68104
rect 212 67928 246 68104
rect -184 67835 184 67869
rect -184 67727 184 67761
rect -246 67492 -212 67668
rect 212 67492 246 67668
rect -184 67399 184 67433
rect -184 67291 184 67325
rect -246 67056 -212 67232
rect 212 67056 246 67232
rect -184 66963 184 66997
rect -184 66855 184 66889
rect -246 66620 -212 66796
rect 212 66620 246 66796
rect -184 66527 184 66561
rect -184 66419 184 66453
rect -246 66184 -212 66360
rect 212 66184 246 66360
rect -184 66091 184 66125
rect -184 65983 184 66017
rect -246 65748 -212 65924
rect 212 65748 246 65924
rect -184 65655 184 65689
rect -184 65547 184 65581
rect -246 65312 -212 65488
rect 212 65312 246 65488
rect -184 65219 184 65253
rect -184 65111 184 65145
rect -246 64876 -212 65052
rect 212 64876 246 65052
rect -184 64783 184 64817
rect -184 64675 184 64709
rect -246 64440 -212 64616
rect 212 64440 246 64616
rect -184 64347 184 64381
rect -184 64239 184 64273
rect -246 64004 -212 64180
rect 212 64004 246 64180
rect -184 63911 184 63945
rect -184 63803 184 63837
rect -246 63568 -212 63744
rect 212 63568 246 63744
rect -184 63475 184 63509
rect -184 63367 184 63401
rect -246 63132 -212 63308
rect 212 63132 246 63308
rect -184 63039 184 63073
rect -184 62931 184 62965
rect -246 62696 -212 62872
rect 212 62696 246 62872
rect -184 62603 184 62637
rect -184 62495 184 62529
rect -246 62260 -212 62436
rect 212 62260 246 62436
rect -184 62167 184 62201
rect -184 62059 184 62093
rect -246 61824 -212 62000
rect 212 61824 246 62000
rect -184 61731 184 61765
rect -184 61623 184 61657
rect -246 61388 -212 61564
rect 212 61388 246 61564
rect -184 61295 184 61329
rect -184 61187 184 61221
rect -246 60952 -212 61128
rect 212 60952 246 61128
rect -184 60859 184 60893
rect -184 60751 184 60785
rect -246 60516 -212 60692
rect 212 60516 246 60692
rect -184 60423 184 60457
rect -184 60315 184 60349
rect -246 60080 -212 60256
rect 212 60080 246 60256
rect -184 59987 184 60021
rect -184 59879 184 59913
rect -246 59644 -212 59820
rect 212 59644 246 59820
rect -184 59551 184 59585
rect -184 59443 184 59477
rect -246 59208 -212 59384
rect 212 59208 246 59384
rect -184 59115 184 59149
rect -184 59007 184 59041
rect -246 58772 -212 58948
rect 212 58772 246 58948
rect -184 58679 184 58713
rect -184 58571 184 58605
rect -246 58336 -212 58512
rect 212 58336 246 58512
rect -184 58243 184 58277
rect -184 58135 184 58169
rect -246 57900 -212 58076
rect 212 57900 246 58076
rect -184 57807 184 57841
rect -184 57699 184 57733
rect -246 57464 -212 57640
rect 212 57464 246 57640
rect -184 57371 184 57405
rect -184 57263 184 57297
rect -246 57028 -212 57204
rect 212 57028 246 57204
rect -184 56935 184 56969
rect -184 56827 184 56861
rect -246 56592 -212 56768
rect 212 56592 246 56768
rect -184 56499 184 56533
rect -184 56391 184 56425
rect -246 56156 -212 56332
rect 212 56156 246 56332
rect -184 56063 184 56097
rect -184 55955 184 55989
rect -246 55720 -212 55896
rect 212 55720 246 55896
rect -184 55627 184 55661
rect -184 55519 184 55553
rect -246 55284 -212 55460
rect 212 55284 246 55460
rect -184 55191 184 55225
rect -184 55083 184 55117
rect -246 54848 -212 55024
rect 212 54848 246 55024
rect -184 54755 184 54789
rect -184 54647 184 54681
rect -246 54412 -212 54588
rect 212 54412 246 54588
rect -184 54319 184 54353
rect -184 54211 184 54245
rect -246 53976 -212 54152
rect 212 53976 246 54152
rect -184 53883 184 53917
rect -184 53775 184 53809
rect -246 53540 -212 53716
rect 212 53540 246 53716
rect -184 53447 184 53481
rect -184 53339 184 53373
rect -246 53104 -212 53280
rect 212 53104 246 53280
rect -184 53011 184 53045
rect -184 52903 184 52937
rect -246 52668 -212 52844
rect 212 52668 246 52844
rect -184 52575 184 52609
rect -184 52467 184 52501
rect -246 52232 -212 52408
rect 212 52232 246 52408
rect -184 52139 184 52173
rect -184 52031 184 52065
rect -246 51796 -212 51972
rect 212 51796 246 51972
rect -184 51703 184 51737
rect -184 51595 184 51629
rect -246 51360 -212 51536
rect 212 51360 246 51536
rect -184 51267 184 51301
rect -184 51159 184 51193
rect -246 50924 -212 51100
rect 212 50924 246 51100
rect -184 50831 184 50865
rect -184 50723 184 50757
rect -246 50488 -212 50664
rect 212 50488 246 50664
rect -184 50395 184 50429
rect -184 50287 184 50321
rect -246 50052 -212 50228
rect 212 50052 246 50228
rect -184 49959 184 49993
rect -184 49851 184 49885
rect -246 49616 -212 49792
rect 212 49616 246 49792
rect -184 49523 184 49557
rect -184 49415 184 49449
rect -246 49180 -212 49356
rect 212 49180 246 49356
rect -184 49087 184 49121
rect -184 48979 184 49013
rect -246 48744 -212 48920
rect 212 48744 246 48920
rect -184 48651 184 48685
rect -184 48543 184 48577
rect -246 48308 -212 48484
rect 212 48308 246 48484
rect -184 48215 184 48249
rect -184 48107 184 48141
rect -246 47872 -212 48048
rect 212 47872 246 48048
rect -184 47779 184 47813
rect -184 47671 184 47705
rect -246 47436 -212 47612
rect 212 47436 246 47612
rect -184 47343 184 47377
rect -184 47235 184 47269
rect -246 47000 -212 47176
rect 212 47000 246 47176
rect -184 46907 184 46941
rect -184 46799 184 46833
rect -246 46564 -212 46740
rect 212 46564 246 46740
rect -184 46471 184 46505
rect -184 46363 184 46397
rect -246 46128 -212 46304
rect 212 46128 246 46304
rect -184 46035 184 46069
rect -184 45927 184 45961
rect -246 45692 -212 45868
rect 212 45692 246 45868
rect -184 45599 184 45633
rect -184 45491 184 45525
rect -246 45256 -212 45432
rect 212 45256 246 45432
rect -184 45163 184 45197
rect -184 45055 184 45089
rect -246 44820 -212 44996
rect 212 44820 246 44996
rect -184 44727 184 44761
rect -184 44619 184 44653
rect -246 44384 -212 44560
rect 212 44384 246 44560
rect -184 44291 184 44325
rect -184 44183 184 44217
rect -246 43948 -212 44124
rect 212 43948 246 44124
rect -184 43855 184 43889
rect -184 43747 184 43781
rect -246 43512 -212 43688
rect 212 43512 246 43688
rect -184 43419 184 43453
rect -184 43311 184 43345
rect -246 43076 -212 43252
rect 212 43076 246 43252
rect -184 42983 184 43017
rect -184 42875 184 42909
rect -246 42640 -212 42816
rect 212 42640 246 42816
rect -184 42547 184 42581
rect -184 42439 184 42473
rect -246 42204 -212 42380
rect 212 42204 246 42380
rect -184 42111 184 42145
rect -184 42003 184 42037
rect -246 41768 -212 41944
rect 212 41768 246 41944
rect -184 41675 184 41709
rect -184 41567 184 41601
rect -246 41332 -212 41508
rect 212 41332 246 41508
rect -184 41239 184 41273
rect -184 41131 184 41165
rect -246 40896 -212 41072
rect 212 40896 246 41072
rect -184 40803 184 40837
rect -184 40695 184 40729
rect -246 40460 -212 40636
rect 212 40460 246 40636
rect -184 40367 184 40401
rect -184 40259 184 40293
rect -246 40024 -212 40200
rect 212 40024 246 40200
rect -184 39931 184 39965
rect -184 39823 184 39857
rect -246 39588 -212 39764
rect 212 39588 246 39764
rect -184 39495 184 39529
rect -184 39387 184 39421
rect -246 39152 -212 39328
rect 212 39152 246 39328
rect -184 39059 184 39093
rect -184 38951 184 38985
rect -246 38716 -212 38892
rect 212 38716 246 38892
rect -184 38623 184 38657
rect -184 38515 184 38549
rect -246 38280 -212 38456
rect 212 38280 246 38456
rect -184 38187 184 38221
rect -184 38079 184 38113
rect -246 37844 -212 38020
rect 212 37844 246 38020
rect -184 37751 184 37785
rect -184 37643 184 37677
rect -246 37408 -212 37584
rect 212 37408 246 37584
rect -184 37315 184 37349
rect -184 37207 184 37241
rect -246 36972 -212 37148
rect 212 36972 246 37148
rect -184 36879 184 36913
rect -184 36771 184 36805
rect -246 36536 -212 36712
rect 212 36536 246 36712
rect -184 36443 184 36477
rect -184 36335 184 36369
rect -246 36100 -212 36276
rect 212 36100 246 36276
rect -184 36007 184 36041
rect -184 35899 184 35933
rect -246 35664 -212 35840
rect 212 35664 246 35840
rect -184 35571 184 35605
rect -184 35463 184 35497
rect -246 35228 -212 35404
rect 212 35228 246 35404
rect -184 35135 184 35169
rect -184 35027 184 35061
rect -246 34792 -212 34968
rect 212 34792 246 34968
rect -184 34699 184 34733
rect -184 34591 184 34625
rect -246 34356 -212 34532
rect 212 34356 246 34532
rect -184 34263 184 34297
rect -184 34155 184 34189
rect -246 33920 -212 34096
rect 212 33920 246 34096
rect -184 33827 184 33861
rect -184 33719 184 33753
rect -246 33484 -212 33660
rect 212 33484 246 33660
rect -184 33391 184 33425
rect -184 33283 184 33317
rect -246 33048 -212 33224
rect 212 33048 246 33224
rect -184 32955 184 32989
rect -184 32847 184 32881
rect -246 32612 -212 32788
rect 212 32612 246 32788
rect -184 32519 184 32553
rect -184 32411 184 32445
rect -246 32176 -212 32352
rect 212 32176 246 32352
rect -184 32083 184 32117
rect -184 31975 184 32009
rect -246 31740 -212 31916
rect 212 31740 246 31916
rect -184 31647 184 31681
rect -184 31539 184 31573
rect -246 31304 -212 31480
rect 212 31304 246 31480
rect -184 31211 184 31245
rect -184 31103 184 31137
rect -246 30868 -212 31044
rect 212 30868 246 31044
rect -184 30775 184 30809
rect -184 30667 184 30701
rect -246 30432 -212 30608
rect 212 30432 246 30608
rect -184 30339 184 30373
rect -184 30231 184 30265
rect -246 29996 -212 30172
rect 212 29996 246 30172
rect -184 29903 184 29937
rect -184 29795 184 29829
rect -246 29560 -212 29736
rect 212 29560 246 29736
rect -184 29467 184 29501
rect -184 29359 184 29393
rect -246 29124 -212 29300
rect 212 29124 246 29300
rect -184 29031 184 29065
rect -184 28923 184 28957
rect -246 28688 -212 28864
rect 212 28688 246 28864
rect -184 28595 184 28629
rect -184 28487 184 28521
rect -246 28252 -212 28428
rect 212 28252 246 28428
rect -184 28159 184 28193
rect -184 28051 184 28085
rect -246 27816 -212 27992
rect 212 27816 246 27992
rect -184 27723 184 27757
rect -184 27615 184 27649
rect -246 27380 -212 27556
rect 212 27380 246 27556
rect -184 27287 184 27321
rect -184 27179 184 27213
rect -246 26944 -212 27120
rect 212 26944 246 27120
rect -184 26851 184 26885
rect -184 26743 184 26777
rect -246 26508 -212 26684
rect 212 26508 246 26684
rect -184 26415 184 26449
rect -184 26307 184 26341
rect -246 26072 -212 26248
rect 212 26072 246 26248
rect -184 25979 184 26013
rect -184 25871 184 25905
rect -246 25636 -212 25812
rect 212 25636 246 25812
rect -184 25543 184 25577
rect -184 25435 184 25469
rect -246 25200 -212 25376
rect 212 25200 246 25376
rect -184 25107 184 25141
rect -184 24999 184 25033
rect -246 24764 -212 24940
rect 212 24764 246 24940
rect -184 24671 184 24705
rect -184 24563 184 24597
rect -246 24328 -212 24504
rect 212 24328 246 24504
rect -184 24235 184 24269
rect -184 24127 184 24161
rect -246 23892 -212 24068
rect 212 23892 246 24068
rect -184 23799 184 23833
rect -184 23691 184 23725
rect -246 23456 -212 23632
rect 212 23456 246 23632
rect -184 23363 184 23397
rect -184 23255 184 23289
rect -246 23020 -212 23196
rect 212 23020 246 23196
rect -184 22927 184 22961
rect -184 22819 184 22853
rect -246 22584 -212 22760
rect 212 22584 246 22760
rect -184 22491 184 22525
rect -184 22383 184 22417
rect -246 22148 -212 22324
rect 212 22148 246 22324
rect -184 22055 184 22089
rect -184 21947 184 21981
rect -246 21712 -212 21888
rect 212 21712 246 21888
rect -184 21619 184 21653
rect -184 21511 184 21545
rect -246 21276 -212 21452
rect 212 21276 246 21452
rect -184 21183 184 21217
rect -184 21075 184 21109
rect -246 20840 -212 21016
rect 212 20840 246 21016
rect -184 20747 184 20781
rect -184 20639 184 20673
rect -246 20404 -212 20580
rect 212 20404 246 20580
rect -184 20311 184 20345
rect -184 20203 184 20237
rect -246 19968 -212 20144
rect 212 19968 246 20144
rect -184 19875 184 19909
rect -184 19767 184 19801
rect -246 19532 -212 19708
rect 212 19532 246 19708
rect -184 19439 184 19473
rect -184 19331 184 19365
rect -246 19096 -212 19272
rect 212 19096 246 19272
rect -184 19003 184 19037
rect -184 18895 184 18929
rect -246 18660 -212 18836
rect 212 18660 246 18836
rect -184 18567 184 18601
rect -184 18459 184 18493
rect -246 18224 -212 18400
rect 212 18224 246 18400
rect -184 18131 184 18165
rect -184 18023 184 18057
rect -246 17788 -212 17964
rect 212 17788 246 17964
rect -184 17695 184 17729
rect -184 17587 184 17621
rect -246 17352 -212 17528
rect 212 17352 246 17528
rect -184 17259 184 17293
rect -184 17151 184 17185
rect -246 16916 -212 17092
rect 212 16916 246 17092
rect -184 16823 184 16857
rect -184 16715 184 16749
rect -246 16480 -212 16656
rect 212 16480 246 16656
rect -184 16387 184 16421
rect -184 16279 184 16313
rect -246 16044 -212 16220
rect 212 16044 246 16220
rect -184 15951 184 15985
rect -184 15843 184 15877
rect -246 15608 -212 15784
rect 212 15608 246 15784
rect -184 15515 184 15549
rect -184 15407 184 15441
rect -246 15172 -212 15348
rect 212 15172 246 15348
rect -184 15079 184 15113
rect -184 14971 184 15005
rect -246 14736 -212 14912
rect 212 14736 246 14912
rect -184 14643 184 14677
rect -184 14535 184 14569
rect -246 14300 -212 14476
rect 212 14300 246 14476
rect -184 14207 184 14241
rect -184 14099 184 14133
rect -246 13864 -212 14040
rect 212 13864 246 14040
rect -184 13771 184 13805
rect -184 13663 184 13697
rect -246 13428 -212 13604
rect 212 13428 246 13604
rect -184 13335 184 13369
rect -184 13227 184 13261
rect -246 12992 -212 13168
rect 212 12992 246 13168
rect -184 12899 184 12933
rect -184 12791 184 12825
rect -246 12556 -212 12732
rect 212 12556 246 12732
rect -184 12463 184 12497
rect -184 12355 184 12389
rect -246 12120 -212 12296
rect 212 12120 246 12296
rect -184 12027 184 12061
rect -184 11919 184 11953
rect -246 11684 -212 11860
rect 212 11684 246 11860
rect -184 11591 184 11625
rect -184 11483 184 11517
rect -246 11248 -212 11424
rect 212 11248 246 11424
rect -184 11155 184 11189
rect -184 11047 184 11081
rect -246 10812 -212 10988
rect 212 10812 246 10988
rect -184 10719 184 10753
rect -184 10611 184 10645
rect -246 10376 -212 10552
rect 212 10376 246 10552
rect -184 10283 184 10317
rect -184 10175 184 10209
rect -246 9940 -212 10116
rect 212 9940 246 10116
rect -184 9847 184 9881
rect -184 9739 184 9773
rect -246 9504 -212 9680
rect 212 9504 246 9680
rect -184 9411 184 9445
rect -184 9303 184 9337
rect -246 9068 -212 9244
rect 212 9068 246 9244
rect -184 8975 184 9009
rect -184 8867 184 8901
rect -246 8632 -212 8808
rect 212 8632 246 8808
rect -184 8539 184 8573
rect -184 8431 184 8465
rect -246 8196 -212 8372
rect 212 8196 246 8372
rect -184 8103 184 8137
rect -184 7995 184 8029
rect -246 7760 -212 7936
rect 212 7760 246 7936
rect -184 7667 184 7701
rect -184 7559 184 7593
rect -246 7324 -212 7500
rect 212 7324 246 7500
rect -184 7231 184 7265
rect -184 7123 184 7157
rect -246 6888 -212 7064
rect 212 6888 246 7064
rect -184 6795 184 6829
rect -184 6687 184 6721
rect -246 6452 -212 6628
rect 212 6452 246 6628
rect -184 6359 184 6393
rect -184 6251 184 6285
rect -246 6016 -212 6192
rect 212 6016 246 6192
rect -184 5923 184 5957
rect -184 5815 184 5849
rect -246 5580 -212 5756
rect 212 5580 246 5756
rect -184 5487 184 5521
rect -184 5379 184 5413
rect -246 5144 -212 5320
rect 212 5144 246 5320
rect -184 5051 184 5085
rect -184 4943 184 4977
rect -246 4708 -212 4884
rect 212 4708 246 4884
rect -184 4615 184 4649
rect -184 4507 184 4541
rect -246 4272 -212 4448
rect 212 4272 246 4448
rect -184 4179 184 4213
rect -184 4071 184 4105
rect -246 3836 -212 4012
rect 212 3836 246 4012
rect -184 3743 184 3777
rect -184 3635 184 3669
rect -246 3400 -212 3576
rect 212 3400 246 3576
rect -184 3307 184 3341
rect -184 3199 184 3233
rect -246 2964 -212 3140
rect 212 2964 246 3140
rect -184 2871 184 2905
rect -184 2763 184 2797
rect -246 2528 -212 2704
rect 212 2528 246 2704
rect -184 2435 184 2469
rect -184 2327 184 2361
rect -246 2092 -212 2268
rect 212 2092 246 2268
rect -184 1999 184 2033
rect -184 1891 184 1925
rect -246 1656 -212 1832
rect 212 1656 246 1832
rect -184 1563 184 1597
rect -184 1455 184 1489
rect -246 1220 -212 1396
rect 212 1220 246 1396
rect -184 1127 184 1161
rect -184 1019 184 1053
rect -246 784 -212 960
rect 212 784 246 960
rect -184 691 184 725
rect -184 583 184 617
rect -246 348 -212 524
rect 212 348 246 524
rect -184 255 184 289
rect -184 147 184 181
rect -246 -88 -212 88
rect 212 -88 246 88
rect -184 -181 184 -147
rect -184 -289 184 -255
rect -246 -524 -212 -348
rect 212 -524 246 -348
rect -184 -617 184 -583
rect -184 -725 184 -691
rect -246 -960 -212 -784
rect 212 -960 246 -784
rect -184 -1053 184 -1019
rect -184 -1161 184 -1127
rect -246 -1396 -212 -1220
rect 212 -1396 246 -1220
rect -184 -1489 184 -1455
rect -184 -1597 184 -1563
rect -246 -1832 -212 -1656
rect 212 -1832 246 -1656
rect -184 -1925 184 -1891
rect -184 -2033 184 -1999
rect -246 -2268 -212 -2092
rect 212 -2268 246 -2092
rect -184 -2361 184 -2327
rect -184 -2469 184 -2435
rect -246 -2704 -212 -2528
rect 212 -2704 246 -2528
rect -184 -2797 184 -2763
rect -184 -2905 184 -2871
rect -246 -3140 -212 -2964
rect 212 -3140 246 -2964
rect -184 -3233 184 -3199
rect -184 -3341 184 -3307
rect -246 -3576 -212 -3400
rect 212 -3576 246 -3400
rect -184 -3669 184 -3635
rect -184 -3777 184 -3743
rect -246 -4012 -212 -3836
rect 212 -4012 246 -3836
rect -184 -4105 184 -4071
rect -184 -4213 184 -4179
rect -246 -4448 -212 -4272
rect 212 -4448 246 -4272
rect -184 -4541 184 -4507
rect -184 -4649 184 -4615
rect -246 -4884 -212 -4708
rect 212 -4884 246 -4708
rect -184 -4977 184 -4943
rect -184 -5085 184 -5051
rect -246 -5320 -212 -5144
rect 212 -5320 246 -5144
rect -184 -5413 184 -5379
rect -184 -5521 184 -5487
rect -246 -5756 -212 -5580
rect 212 -5756 246 -5580
rect -184 -5849 184 -5815
rect -184 -5957 184 -5923
rect -246 -6192 -212 -6016
rect 212 -6192 246 -6016
rect -184 -6285 184 -6251
rect -184 -6393 184 -6359
rect -246 -6628 -212 -6452
rect 212 -6628 246 -6452
rect -184 -6721 184 -6687
rect -184 -6829 184 -6795
rect -246 -7064 -212 -6888
rect 212 -7064 246 -6888
rect -184 -7157 184 -7123
rect -184 -7265 184 -7231
rect -246 -7500 -212 -7324
rect 212 -7500 246 -7324
rect -184 -7593 184 -7559
rect -184 -7701 184 -7667
rect -246 -7936 -212 -7760
rect 212 -7936 246 -7760
rect -184 -8029 184 -7995
rect -184 -8137 184 -8103
rect -246 -8372 -212 -8196
rect 212 -8372 246 -8196
rect -184 -8465 184 -8431
rect -184 -8573 184 -8539
rect -246 -8808 -212 -8632
rect 212 -8808 246 -8632
rect -184 -8901 184 -8867
rect -184 -9009 184 -8975
rect -246 -9244 -212 -9068
rect 212 -9244 246 -9068
rect -184 -9337 184 -9303
rect -184 -9445 184 -9411
rect -246 -9680 -212 -9504
rect 212 -9680 246 -9504
rect -184 -9773 184 -9739
rect -184 -9881 184 -9847
rect -246 -10116 -212 -9940
rect 212 -10116 246 -9940
rect -184 -10209 184 -10175
rect -184 -10317 184 -10283
rect -246 -10552 -212 -10376
rect 212 -10552 246 -10376
rect -184 -10645 184 -10611
rect -184 -10753 184 -10719
rect -246 -10988 -212 -10812
rect 212 -10988 246 -10812
rect -184 -11081 184 -11047
rect -184 -11189 184 -11155
rect -246 -11424 -212 -11248
rect 212 -11424 246 -11248
rect -184 -11517 184 -11483
rect -184 -11625 184 -11591
rect -246 -11860 -212 -11684
rect 212 -11860 246 -11684
rect -184 -11953 184 -11919
rect -184 -12061 184 -12027
rect -246 -12296 -212 -12120
rect 212 -12296 246 -12120
rect -184 -12389 184 -12355
rect -184 -12497 184 -12463
rect -246 -12732 -212 -12556
rect 212 -12732 246 -12556
rect -184 -12825 184 -12791
rect -184 -12933 184 -12899
rect -246 -13168 -212 -12992
rect 212 -13168 246 -12992
rect -184 -13261 184 -13227
rect -184 -13369 184 -13335
rect -246 -13604 -212 -13428
rect 212 -13604 246 -13428
rect -184 -13697 184 -13663
rect -184 -13805 184 -13771
rect -246 -14040 -212 -13864
rect 212 -14040 246 -13864
rect -184 -14133 184 -14099
rect -184 -14241 184 -14207
rect -246 -14476 -212 -14300
rect 212 -14476 246 -14300
rect -184 -14569 184 -14535
rect -184 -14677 184 -14643
rect -246 -14912 -212 -14736
rect 212 -14912 246 -14736
rect -184 -15005 184 -14971
rect -184 -15113 184 -15079
rect -246 -15348 -212 -15172
rect 212 -15348 246 -15172
rect -184 -15441 184 -15407
rect -184 -15549 184 -15515
rect -246 -15784 -212 -15608
rect 212 -15784 246 -15608
rect -184 -15877 184 -15843
rect -184 -15985 184 -15951
rect -246 -16220 -212 -16044
rect 212 -16220 246 -16044
rect -184 -16313 184 -16279
rect -184 -16421 184 -16387
rect -246 -16656 -212 -16480
rect 212 -16656 246 -16480
rect -184 -16749 184 -16715
rect -184 -16857 184 -16823
rect -246 -17092 -212 -16916
rect 212 -17092 246 -16916
rect -184 -17185 184 -17151
rect -184 -17293 184 -17259
rect -246 -17528 -212 -17352
rect 212 -17528 246 -17352
rect -184 -17621 184 -17587
rect -184 -17729 184 -17695
rect -246 -17964 -212 -17788
rect 212 -17964 246 -17788
rect -184 -18057 184 -18023
rect -184 -18165 184 -18131
rect -246 -18400 -212 -18224
rect 212 -18400 246 -18224
rect -184 -18493 184 -18459
rect -184 -18601 184 -18567
rect -246 -18836 -212 -18660
rect 212 -18836 246 -18660
rect -184 -18929 184 -18895
rect -184 -19037 184 -19003
rect -246 -19272 -212 -19096
rect 212 -19272 246 -19096
rect -184 -19365 184 -19331
rect -184 -19473 184 -19439
rect -246 -19708 -212 -19532
rect 212 -19708 246 -19532
rect -184 -19801 184 -19767
rect -184 -19909 184 -19875
rect -246 -20144 -212 -19968
rect 212 -20144 246 -19968
rect -184 -20237 184 -20203
rect -184 -20345 184 -20311
rect -246 -20580 -212 -20404
rect 212 -20580 246 -20404
rect -184 -20673 184 -20639
rect -184 -20781 184 -20747
rect -246 -21016 -212 -20840
rect 212 -21016 246 -20840
rect -184 -21109 184 -21075
rect -184 -21217 184 -21183
rect -246 -21452 -212 -21276
rect 212 -21452 246 -21276
rect -184 -21545 184 -21511
rect -184 -21653 184 -21619
rect -246 -21888 -212 -21712
rect 212 -21888 246 -21712
rect -184 -21981 184 -21947
rect -184 -22089 184 -22055
rect -246 -22324 -212 -22148
rect 212 -22324 246 -22148
rect -184 -22417 184 -22383
rect -184 -22525 184 -22491
rect -246 -22760 -212 -22584
rect 212 -22760 246 -22584
rect -184 -22853 184 -22819
rect -184 -22961 184 -22927
rect -246 -23196 -212 -23020
rect 212 -23196 246 -23020
rect -184 -23289 184 -23255
rect -184 -23397 184 -23363
rect -246 -23632 -212 -23456
rect 212 -23632 246 -23456
rect -184 -23725 184 -23691
rect -184 -23833 184 -23799
rect -246 -24068 -212 -23892
rect 212 -24068 246 -23892
rect -184 -24161 184 -24127
rect -184 -24269 184 -24235
rect -246 -24504 -212 -24328
rect 212 -24504 246 -24328
rect -184 -24597 184 -24563
rect -184 -24705 184 -24671
rect -246 -24940 -212 -24764
rect 212 -24940 246 -24764
rect -184 -25033 184 -24999
rect -184 -25141 184 -25107
rect -246 -25376 -212 -25200
rect 212 -25376 246 -25200
rect -184 -25469 184 -25435
rect -184 -25577 184 -25543
rect -246 -25812 -212 -25636
rect 212 -25812 246 -25636
rect -184 -25905 184 -25871
rect -184 -26013 184 -25979
rect -246 -26248 -212 -26072
rect 212 -26248 246 -26072
rect -184 -26341 184 -26307
rect -184 -26449 184 -26415
rect -246 -26684 -212 -26508
rect 212 -26684 246 -26508
rect -184 -26777 184 -26743
rect -184 -26885 184 -26851
rect -246 -27120 -212 -26944
rect 212 -27120 246 -26944
rect -184 -27213 184 -27179
rect -184 -27321 184 -27287
rect -246 -27556 -212 -27380
rect 212 -27556 246 -27380
rect -184 -27649 184 -27615
rect -184 -27757 184 -27723
rect -246 -27992 -212 -27816
rect 212 -27992 246 -27816
rect -184 -28085 184 -28051
rect -184 -28193 184 -28159
rect -246 -28428 -212 -28252
rect 212 -28428 246 -28252
rect -184 -28521 184 -28487
rect -184 -28629 184 -28595
rect -246 -28864 -212 -28688
rect 212 -28864 246 -28688
rect -184 -28957 184 -28923
rect -184 -29065 184 -29031
rect -246 -29300 -212 -29124
rect 212 -29300 246 -29124
rect -184 -29393 184 -29359
rect -184 -29501 184 -29467
rect -246 -29736 -212 -29560
rect 212 -29736 246 -29560
rect -184 -29829 184 -29795
rect -184 -29937 184 -29903
rect -246 -30172 -212 -29996
rect 212 -30172 246 -29996
rect -184 -30265 184 -30231
rect -184 -30373 184 -30339
rect -246 -30608 -212 -30432
rect 212 -30608 246 -30432
rect -184 -30701 184 -30667
rect -184 -30809 184 -30775
rect -246 -31044 -212 -30868
rect 212 -31044 246 -30868
rect -184 -31137 184 -31103
rect -184 -31245 184 -31211
rect -246 -31480 -212 -31304
rect 212 -31480 246 -31304
rect -184 -31573 184 -31539
rect -184 -31681 184 -31647
rect -246 -31916 -212 -31740
rect 212 -31916 246 -31740
rect -184 -32009 184 -31975
rect -184 -32117 184 -32083
rect -246 -32352 -212 -32176
rect 212 -32352 246 -32176
rect -184 -32445 184 -32411
rect -184 -32553 184 -32519
rect -246 -32788 -212 -32612
rect 212 -32788 246 -32612
rect -184 -32881 184 -32847
rect -184 -32989 184 -32955
rect -246 -33224 -212 -33048
rect 212 -33224 246 -33048
rect -184 -33317 184 -33283
rect -184 -33425 184 -33391
rect -246 -33660 -212 -33484
rect 212 -33660 246 -33484
rect -184 -33753 184 -33719
rect -184 -33861 184 -33827
rect -246 -34096 -212 -33920
rect 212 -34096 246 -33920
rect -184 -34189 184 -34155
rect -184 -34297 184 -34263
rect -246 -34532 -212 -34356
rect 212 -34532 246 -34356
rect -184 -34625 184 -34591
rect -184 -34733 184 -34699
rect -246 -34968 -212 -34792
rect 212 -34968 246 -34792
rect -184 -35061 184 -35027
rect -184 -35169 184 -35135
rect -246 -35404 -212 -35228
rect 212 -35404 246 -35228
rect -184 -35497 184 -35463
rect -184 -35605 184 -35571
rect -246 -35840 -212 -35664
rect 212 -35840 246 -35664
rect -184 -35933 184 -35899
rect -184 -36041 184 -36007
rect -246 -36276 -212 -36100
rect 212 -36276 246 -36100
rect -184 -36369 184 -36335
rect -184 -36477 184 -36443
rect -246 -36712 -212 -36536
rect 212 -36712 246 -36536
rect -184 -36805 184 -36771
rect -184 -36913 184 -36879
rect -246 -37148 -212 -36972
rect 212 -37148 246 -36972
rect -184 -37241 184 -37207
rect -184 -37349 184 -37315
rect -246 -37584 -212 -37408
rect 212 -37584 246 -37408
rect -184 -37677 184 -37643
rect -184 -37785 184 -37751
rect -246 -38020 -212 -37844
rect 212 -38020 246 -37844
rect -184 -38113 184 -38079
rect -184 -38221 184 -38187
rect -246 -38456 -212 -38280
rect 212 -38456 246 -38280
rect -184 -38549 184 -38515
rect -184 -38657 184 -38623
rect -246 -38892 -212 -38716
rect 212 -38892 246 -38716
rect -184 -38985 184 -38951
rect -184 -39093 184 -39059
rect -246 -39328 -212 -39152
rect 212 -39328 246 -39152
rect -184 -39421 184 -39387
rect -184 -39529 184 -39495
rect -246 -39764 -212 -39588
rect 212 -39764 246 -39588
rect -184 -39857 184 -39823
rect -184 -39965 184 -39931
rect -246 -40200 -212 -40024
rect 212 -40200 246 -40024
rect -184 -40293 184 -40259
rect -184 -40401 184 -40367
rect -246 -40636 -212 -40460
rect 212 -40636 246 -40460
rect -184 -40729 184 -40695
rect -184 -40837 184 -40803
rect -246 -41072 -212 -40896
rect 212 -41072 246 -40896
rect -184 -41165 184 -41131
rect -184 -41273 184 -41239
rect -246 -41508 -212 -41332
rect 212 -41508 246 -41332
rect -184 -41601 184 -41567
rect -184 -41709 184 -41675
rect -246 -41944 -212 -41768
rect 212 -41944 246 -41768
rect -184 -42037 184 -42003
rect -184 -42145 184 -42111
rect -246 -42380 -212 -42204
rect 212 -42380 246 -42204
rect -184 -42473 184 -42439
rect -184 -42581 184 -42547
rect -246 -42816 -212 -42640
rect 212 -42816 246 -42640
rect -184 -42909 184 -42875
rect -184 -43017 184 -42983
rect -246 -43252 -212 -43076
rect 212 -43252 246 -43076
rect -184 -43345 184 -43311
rect -184 -43453 184 -43419
rect -246 -43688 -212 -43512
rect 212 -43688 246 -43512
rect -184 -43781 184 -43747
rect -184 -43889 184 -43855
rect -246 -44124 -212 -43948
rect 212 -44124 246 -43948
rect -184 -44217 184 -44183
rect -184 -44325 184 -44291
rect -246 -44560 -212 -44384
rect 212 -44560 246 -44384
rect -184 -44653 184 -44619
rect -184 -44761 184 -44727
rect -246 -44996 -212 -44820
rect 212 -44996 246 -44820
rect -184 -45089 184 -45055
rect -184 -45197 184 -45163
rect -246 -45432 -212 -45256
rect 212 -45432 246 -45256
rect -184 -45525 184 -45491
rect -184 -45633 184 -45599
rect -246 -45868 -212 -45692
rect 212 -45868 246 -45692
rect -184 -45961 184 -45927
rect -184 -46069 184 -46035
rect -246 -46304 -212 -46128
rect 212 -46304 246 -46128
rect -184 -46397 184 -46363
rect -184 -46505 184 -46471
rect -246 -46740 -212 -46564
rect 212 -46740 246 -46564
rect -184 -46833 184 -46799
rect -184 -46941 184 -46907
rect -246 -47176 -212 -47000
rect 212 -47176 246 -47000
rect -184 -47269 184 -47235
rect -184 -47377 184 -47343
rect -246 -47612 -212 -47436
rect 212 -47612 246 -47436
rect -184 -47705 184 -47671
rect -184 -47813 184 -47779
rect -246 -48048 -212 -47872
rect 212 -48048 246 -47872
rect -184 -48141 184 -48107
rect -184 -48249 184 -48215
rect -246 -48484 -212 -48308
rect 212 -48484 246 -48308
rect -184 -48577 184 -48543
rect -184 -48685 184 -48651
rect -246 -48920 -212 -48744
rect 212 -48920 246 -48744
rect -184 -49013 184 -48979
rect -184 -49121 184 -49087
rect -246 -49356 -212 -49180
rect 212 -49356 246 -49180
rect -184 -49449 184 -49415
rect -184 -49557 184 -49523
rect -246 -49792 -212 -49616
rect 212 -49792 246 -49616
rect -184 -49885 184 -49851
rect -184 -49993 184 -49959
rect -246 -50228 -212 -50052
rect 212 -50228 246 -50052
rect -184 -50321 184 -50287
rect -184 -50429 184 -50395
rect -246 -50664 -212 -50488
rect 212 -50664 246 -50488
rect -184 -50757 184 -50723
rect -184 -50865 184 -50831
rect -246 -51100 -212 -50924
rect 212 -51100 246 -50924
rect -184 -51193 184 -51159
rect -184 -51301 184 -51267
rect -246 -51536 -212 -51360
rect 212 -51536 246 -51360
rect -184 -51629 184 -51595
rect -184 -51737 184 -51703
rect -246 -51972 -212 -51796
rect 212 -51972 246 -51796
rect -184 -52065 184 -52031
rect -184 -52173 184 -52139
rect -246 -52408 -212 -52232
rect 212 -52408 246 -52232
rect -184 -52501 184 -52467
rect -184 -52609 184 -52575
rect -246 -52844 -212 -52668
rect 212 -52844 246 -52668
rect -184 -52937 184 -52903
rect -184 -53045 184 -53011
rect -246 -53280 -212 -53104
rect 212 -53280 246 -53104
rect -184 -53373 184 -53339
rect -184 -53481 184 -53447
rect -246 -53716 -212 -53540
rect 212 -53716 246 -53540
rect -184 -53809 184 -53775
rect -184 -53917 184 -53883
rect -246 -54152 -212 -53976
rect 212 -54152 246 -53976
rect -184 -54245 184 -54211
rect -184 -54353 184 -54319
rect -246 -54588 -212 -54412
rect 212 -54588 246 -54412
rect -184 -54681 184 -54647
rect -184 -54789 184 -54755
rect -246 -55024 -212 -54848
rect 212 -55024 246 -54848
rect -184 -55117 184 -55083
rect -184 -55225 184 -55191
rect -246 -55460 -212 -55284
rect 212 -55460 246 -55284
rect -184 -55553 184 -55519
rect -184 -55661 184 -55627
rect -246 -55896 -212 -55720
rect 212 -55896 246 -55720
rect -184 -55989 184 -55955
rect -184 -56097 184 -56063
rect -246 -56332 -212 -56156
rect 212 -56332 246 -56156
rect -184 -56425 184 -56391
rect -184 -56533 184 -56499
rect -246 -56768 -212 -56592
rect 212 -56768 246 -56592
rect -184 -56861 184 -56827
rect -184 -56969 184 -56935
rect -246 -57204 -212 -57028
rect 212 -57204 246 -57028
rect -184 -57297 184 -57263
rect -184 -57405 184 -57371
rect -246 -57640 -212 -57464
rect 212 -57640 246 -57464
rect -184 -57733 184 -57699
rect -184 -57841 184 -57807
rect -246 -58076 -212 -57900
rect 212 -58076 246 -57900
rect -184 -58169 184 -58135
rect -184 -58277 184 -58243
rect -246 -58512 -212 -58336
rect 212 -58512 246 -58336
rect -184 -58605 184 -58571
rect -184 -58713 184 -58679
rect -246 -58948 -212 -58772
rect 212 -58948 246 -58772
rect -184 -59041 184 -59007
rect -184 -59149 184 -59115
rect -246 -59384 -212 -59208
rect 212 -59384 246 -59208
rect -184 -59477 184 -59443
rect -184 -59585 184 -59551
rect -246 -59820 -212 -59644
rect 212 -59820 246 -59644
rect -184 -59913 184 -59879
rect -184 -60021 184 -59987
rect -246 -60256 -212 -60080
rect 212 -60256 246 -60080
rect -184 -60349 184 -60315
rect -184 -60457 184 -60423
rect -246 -60692 -212 -60516
rect 212 -60692 246 -60516
rect -184 -60785 184 -60751
rect -184 -60893 184 -60859
rect -246 -61128 -212 -60952
rect 212 -61128 246 -60952
rect -184 -61221 184 -61187
rect -184 -61329 184 -61295
rect -246 -61564 -212 -61388
rect 212 -61564 246 -61388
rect -184 -61657 184 -61623
rect -184 -61765 184 -61731
rect -246 -62000 -212 -61824
rect 212 -62000 246 -61824
rect -184 -62093 184 -62059
rect -184 -62201 184 -62167
rect -246 -62436 -212 -62260
rect 212 -62436 246 -62260
rect -184 -62529 184 -62495
rect -184 -62637 184 -62603
rect -246 -62872 -212 -62696
rect 212 -62872 246 -62696
rect -184 -62965 184 -62931
rect -184 -63073 184 -63039
rect -246 -63308 -212 -63132
rect 212 -63308 246 -63132
rect -184 -63401 184 -63367
rect -184 -63509 184 -63475
rect -246 -63744 -212 -63568
rect 212 -63744 246 -63568
rect -184 -63837 184 -63803
rect -184 -63945 184 -63911
rect -246 -64180 -212 -64004
rect 212 -64180 246 -64004
rect -184 -64273 184 -64239
rect -184 -64381 184 -64347
rect -246 -64616 -212 -64440
rect 212 -64616 246 -64440
rect -184 -64709 184 -64675
rect -184 -64817 184 -64783
rect -246 -65052 -212 -64876
rect 212 -65052 246 -64876
rect -184 -65145 184 -65111
rect -184 -65253 184 -65219
rect -246 -65488 -212 -65312
rect 212 -65488 246 -65312
rect -184 -65581 184 -65547
rect -184 -65689 184 -65655
rect -246 -65924 -212 -65748
rect 212 -65924 246 -65748
rect -184 -66017 184 -65983
rect -184 -66125 184 -66091
rect -246 -66360 -212 -66184
rect 212 -66360 246 -66184
rect -184 -66453 184 -66419
rect -184 -66561 184 -66527
rect -246 -66796 -212 -66620
rect 212 -66796 246 -66620
rect -184 -66889 184 -66855
rect -184 -66997 184 -66963
rect -246 -67232 -212 -67056
rect 212 -67232 246 -67056
rect -184 -67325 184 -67291
rect -184 -67433 184 -67399
rect -246 -67668 -212 -67492
rect 212 -67668 246 -67492
rect -184 -67761 184 -67727
rect -184 -67869 184 -67835
rect -246 -68104 -212 -67928
rect 212 -68104 246 -67928
rect -184 -68197 184 -68163
rect -184 -68305 184 -68271
rect -246 -68540 -212 -68364
rect 212 -68540 246 -68364
rect -184 -68633 184 -68599
rect -184 -68741 184 -68707
rect -246 -68976 -212 -68800
rect 212 -68976 246 -68800
rect -184 -69069 184 -69035
rect -184 -69177 184 -69143
rect -246 -69412 -212 -69236
rect 212 -69412 246 -69236
rect -184 -69505 184 -69471
rect -184 -69613 184 -69579
rect -246 -69848 -212 -69672
rect 212 -69848 246 -69672
rect -184 -69941 184 -69907
rect -184 -70049 184 -70015
rect -246 -70284 -212 -70108
rect 212 -70284 246 -70108
rect -184 -70377 184 -70343
rect -184 -70485 184 -70451
rect -246 -70720 -212 -70544
rect 212 -70720 246 -70544
rect -184 -70813 184 -70779
rect -184 -70921 184 -70887
rect -246 -71156 -212 -70980
rect 212 -71156 246 -70980
rect -184 -71249 184 -71215
rect -184 -71357 184 -71323
rect -246 -71592 -212 -71416
rect 212 -71592 246 -71416
rect -184 -71685 184 -71651
rect -184 -71793 184 -71759
rect -246 -72028 -212 -71852
rect 212 -72028 246 -71852
rect -184 -72121 184 -72087
rect -184 -72229 184 -72195
rect -246 -72464 -212 -72288
rect 212 -72464 246 -72288
rect -184 -72557 184 -72523
rect -184 -72665 184 -72631
rect -246 -72900 -212 -72724
rect 212 -72900 246 -72724
rect -184 -72993 184 -72959
rect -184 -73101 184 -73067
rect -246 -73336 -212 -73160
rect 212 -73336 246 -73160
rect -184 -73429 184 -73395
rect -184 -73537 184 -73503
rect -246 -73772 -212 -73596
rect 212 -73772 246 -73596
rect -184 -73865 184 -73831
rect -184 -73973 184 -73939
rect -246 -74208 -212 -74032
rect 212 -74208 246 -74032
rect -184 -74301 184 -74267
rect -184 -74409 184 -74375
rect -246 -74644 -212 -74468
rect 212 -74644 246 -74468
rect -184 -74737 184 -74703
rect -184 -74845 184 -74811
rect -246 -75080 -212 -74904
rect 212 -75080 246 -74904
rect -184 -75173 184 -75139
rect -184 -75281 184 -75247
rect -246 -75516 -212 -75340
rect 212 -75516 246 -75340
rect -184 -75609 184 -75575
rect -184 -75717 184 -75683
rect -246 -75952 -212 -75776
rect 212 -75952 246 -75776
rect -184 -76045 184 -76011
rect -184 -76153 184 -76119
rect -246 -76388 -212 -76212
rect 212 -76388 246 -76212
rect -184 -76481 184 -76447
rect -184 -76589 184 -76555
rect -246 -76824 -212 -76648
rect 212 -76824 246 -76648
rect -184 -76917 184 -76883
rect -184 -77025 184 -76991
rect -246 -77260 -212 -77084
rect 212 -77260 246 -77084
rect -184 -77353 184 -77319
rect -184 -77461 184 -77427
rect -246 -77696 -212 -77520
rect 212 -77696 246 -77520
rect -184 -77789 184 -77755
rect -184 -77897 184 -77863
rect -246 -78132 -212 -77956
rect 212 -78132 246 -77956
rect -184 -78225 184 -78191
rect -184 -78333 184 -78299
rect -246 -78568 -212 -78392
rect 212 -78568 246 -78392
rect -184 -78661 184 -78627
rect -184 -78769 184 -78735
rect -246 -79004 -212 -78828
rect 212 -79004 246 -78828
rect -184 -79097 184 -79063
rect -184 -79205 184 -79171
rect -246 -79440 -212 -79264
rect 212 -79440 246 -79264
rect -184 -79533 184 -79499
rect -184 -79641 184 -79607
rect -246 -79876 -212 -79700
rect 212 -79876 246 -79700
rect -184 -79969 184 -79935
rect -184 -80077 184 -80043
rect -246 -80312 -212 -80136
rect 212 -80312 246 -80136
rect -184 -80405 184 -80371
rect -184 -80513 184 -80479
rect -246 -80748 -212 -80572
rect 212 -80748 246 -80572
rect -184 -80841 184 -80807
rect -184 -80949 184 -80915
rect -246 -81184 -212 -81008
rect 212 -81184 246 -81008
rect -184 -81277 184 -81243
rect -184 -81385 184 -81351
rect -246 -81620 -212 -81444
rect 212 -81620 246 -81444
rect -184 -81713 184 -81679
rect -184 -81821 184 -81787
rect -246 -82056 -212 -81880
rect 212 -82056 246 -81880
rect -184 -82149 184 -82115
rect -184 -82257 184 -82223
rect -246 -82492 -212 -82316
rect 212 -82492 246 -82316
rect -184 -82585 184 -82551
rect -184 -82693 184 -82659
rect -246 -82928 -212 -82752
rect 212 -82928 246 -82752
rect -184 -83021 184 -82987
rect -184 -83129 184 -83095
rect -246 -83364 -212 -83188
rect 212 -83364 246 -83188
rect -184 -83457 184 -83423
rect -184 -83565 184 -83531
rect -246 -83800 -212 -83624
rect 212 -83800 246 -83624
rect -184 -83893 184 -83859
rect -184 -84001 184 -83967
rect -246 -84236 -212 -84060
rect 212 -84236 246 -84060
rect -184 -84329 184 -84295
<< metal1 >>
rect -196 84329 196 84335
rect -196 84295 -184 84329
rect 184 84295 196 84329
rect -196 84289 196 84295
rect -252 84236 -206 84248
rect -252 84060 -246 84236
rect -212 84060 -206 84236
rect -252 84048 -206 84060
rect 206 84236 252 84248
rect 206 84060 212 84236
rect 246 84060 252 84236
rect 206 84048 252 84060
rect -196 84001 196 84007
rect -196 83967 -184 84001
rect 184 83967 196 84001
rect -196 83961 196 83967
rect -196 83893 196 83899
rect -196 83859 -184 83893
rect 184 83859 196 83893
rect -196 83853 196 83859
rect -252 83800 -206 83812
rect -252 83624 -246 83800
rect -212 83624 -206 83800
rect -252 83612 -206 83624
rect 206 83800 252 83812
rect 206 83624 212 83800
rect 246 83624 252 83800
rect 206 83612 252 83624
rect -196 83565 196 83571
rect -196 83531 -184 83565
rect 184 83531 196 83565
rect -196 83525 196 83531
rect -196 83457 196 83463
rect -196 83423 -184 83457
rect 184 83423 196 83457
rect -196 83417 196 83423
rect -252 83364 -206 83376
rect -252 83188 -246 83364
rect -212 83188 -206 83364
rect -252 83176 -206 83188
rect 206 83364 252 83376
rect 206 83188 212 83364
rect 246 83188 252 83364
rect 206 83176 252 83188
rect -196 83129 196 83135
rect -196 83095 -184 83129
rect 184 83095 196 83129
rect -196 83089 196 83095
rect -196 83021 196 83027
rect -196 82987 -184 83021
rect 184 82987 196 83021
rect -196 82981 196 82987
rect -252 82928 -206 82940
rect -252 82752 -246 82928
rect -212 82752 -206 82928
rect -252 82740 -206 82752
rect 206 82928 252 82940
rect 206 82752 212 82928
rect 246 82752 252 82928
rect 206 82740 252 82752
rect -196 82693 196 82699
rect -196 82659 -184 82693
rect 184 82659 196 82693
rect -196 82653 196 82659
rect -196 82585 196 82591
rect -196 82551 -184 82585
rect 184 82551 196 82585
rect -196 82545 196 82551
rect -252 82492 -206 82504
rect -252 82316 -246 82492
rect -212 82316 -206 82492
rect -252 82304 -206 82316
rect 206 82492 252 82504
rect 206 82316 212 82492
rect 246 82316 252 82492
rect 206 82304 252 82316
rect -196 82257 196 82263
rect -196 82223 -184 82257
rect 184 82223 196 82257
rect -196 82217 196 82223
rect -196 82149 196 82155
rect -196 82115 -184 82149
rect 184 82115 196 82149
rect -196 82109 196 82115
rect -252 82056 -206 82068
rect -252 81880 -246 82056
rect -212 81880 -206 82056
rect -252 81868 -206 81880
rect 206 82056 252 82068
rect 206 81880 212 82056
rect 246 81880 252 82056
rect 206 81868 252 81880
rect -196 81821 196 81827
rect -196 81787 -184 81821
rect 184 81787 196 81821
rect -196 81781 196 81787
rect -196 81713 196 81719
rect -196 81679 -184 81713
rect 184 81679 196 81713
rect -196 81673 196 81679
rect -252 81620 -206 81632
rect -252 81444 -246 81620
rect -212 81444 -206 81620
rect -252 81432 -206 81444
rect 206 81620 252 81632
rect 206 81444 212 81620
rect 246 81444 252 81620
rect 206 81432 252 81444
rect -196 81385 196 81391
rect -196 81351 -184 81385
rect 184 81351 196 81385
rect -196 81345 196 81351
rect -196 81277 196 81283
rect -196 81243 -184 81277
rect 184 81243 196 81277
rect -196 81237 196 81243
rect -252 81184 -206 81196
rect -252 81008 -246 81184
rect -212 81008 -206 81184
rect -252 80996 -206 81008
rect 206 81184 252 81196
rect 206 81008 212 81184
rect 246 81008 252 81184
rect 206 80996 252 81008
rect -196 80949 196 80955
rect -196 80915 -184 80949
rect 184 80915 196 80949
rect -196 80909 196 80915
rect -196 80841 196 80847
rect -196 80807 -184 80841
rect 184 80807 196 80841
rect -196 80801 196 80807
rect -252 80748 -206 80760
rect -252 80572 -246 80748
rect -212 80572 -206 80748
rect -252 80560 -206 80572
rect 206 80748 252 80760
rect 206 80572 212 80748
rect 246 80572 252 80748
rect 206 80560 252 80572
rect -196 80513 196 80519
rect -196 80479 -184 80513
rect 184 80479 196 80513
rect -196 80473 196 80479
rect -196 80405 196 80411
rect -196 80371 -184 80405
rect 184 80371 196 80405
rect -196 80365 196 80371
rect -252 80312 -206 80324
rect -252 80136 -246 80312
rect -212 80136 -206 80312
rect -252 80124 -206 80136
rect 206 80312 252 80324
rect 206 80136 212 80312
rect 246 80136 252 80312
rect 206 80124 252 80136
rect -196 80077 196 80083
rect -196 80043 -184 80077
rect 184 80043 196 80077
rect -196 80037 196 80043
rect -196 79969 196 79975
rect -196 79935 -184 79969
rect 184 79935 196 79969
rect -196 79929 196 79935
rect -252 79876 -206 79888
rect -252 79700 -246 79876
rect -212 79700 -206 79876
rect -252 79688 -206 79700
rect 206 79876 252 79888
rect 206 79700 212 79876
rect 246 79700 252 79876
rect 206 79688 252 79700
rect -196 79641 196 79647
rect -196 79607 -184 79641
rect 184 79607 196 79641
rect -196 79601 196 79607
rect -196 79533 196 79539
rect -196 79499 -184 79533
rect 184 79499 196 79533
rect -196 79493 196 79499
rect -252 79440 -206 79452
rect -252 79264 -246 79440
rect -212 79264 -206 79440
rect -252 79252 -206 79264
rect 206 79440 252 79452
rect 206 79264 212 79440
rect 246 79264 252 79440
rect 206 79252 252 79264
rect -196 79205 196 79211
rect -196 79171 -184 79205
rect 184 79171 196 79205
rect -196 79165 196 79171
rect -196 79097 196 79103
rect -196 79063 -184 79097
rect 184 79063 196 79097
rect -196 79057 196 79063
rect -252 79004 -206 79016
rect -252 78828 -246 79004
rect -212 78828 -206 79004
rect -252 78816 -206 78828
rect 206 79004 252 79016
rect 206 78828 212 79004
rect 246 78828 252 79004
rect 206 78816 252 78828
rect -196 78769 196 78775
rect -196 78735 -184 78769
rect 184 78735 196 78769
rect -196 78729 196 78735
rect -196 78661 196 78667
rect -196 78627 -184 78661
rect 184 78627 196 78661
rect -196 78621 196 78627
rect -252 78568 -206 78580
rect -252 78392 -246 78568
rect -212 78392 -206 78568
rect -252 78380 -206 78392
rect 206 78568 252 78580
rect 206 78392 212 78568
rect 246 78392 252 78568
rect 206 78380 252 78392
rect -196 78333 196 78339
rect -196 78299 -184 78333
rect 184 78299 196 78333
rect -196 78293 196 78299
rect -196 78225 196 78231
rect -196 78191 -184 78225
rect 184 78191 196 78225
rect -196 78185 196 78191
rect -252 78132 -206 78144
rect -252 77956 -246 78132
rect -212 77956 -206 78132
rect -252 77944 -206 77956
rect 206 78132 252 78144
rect 206 77956 212 78132
rect 246 77956 252 78132
rect 206 77944 252 77956
rect -196 77897 196 77903
rect -196 77863 -184 77897
rect 184 77863 196 77897
rect -196 77857 196 77863
rect -196 77789 196 77795
rect -196 77755 -184 77789
rect 184 77755 196 77789
rect -196 77749 196 77755
rect -252 77696 -206 77708
rect -252 77520 -246 77696
rect -212 77520 -206 77696
rect -252 77508 -206 77520
rect 206 77696 252 77708
rect 206 77520 212 77696
rect 246 77520 252 77696
rect 206 77508 252 77520
rect -196 77461 196 77467
rect -196 77427 -184 77461
rect 184 77427 196 77461
rect -196 77421 196 77427
rect -196 77353 196 77359
rect -196 77319 -184 77353
rect 184 77319 196 77353
rect -196 77313 196 77319
rect -252 77260 -206 77272
rect -252 77084 -246 77260
rect -212 77084 -206 77260
rect -252 77072 -206 77084
rect 206 77260 252 77272
rect 206 77084 212 77260
rect 246 77084 252 77260
rect 206 77072 252 77084
rect -196 77025 196 77031
rect -196 76991 -184 77025
rect 184 76991 196 77025
rect -196 76985 196 76991
rect -196 76917 196 76923
rect -196 76883 -184 76917
rect 184 76883 196 76917
rect -196 76877 196 76883
rect -252 76824 -206 76836
rect -252 76648 -246 76824
rect -212 76648 -206 76824
rect -252 76636 -206 76648
rect 206 76824 252 76836
rect 206 76648 212 76824
rect 246 76648 252 76824
rect 206 76636 252 76648
rect -196 76589 196 76595
rect -196 76555 -184 76589
rect 184 76555 196 76589
rect -196 76549 196 76555
rect -196 76481 196 76487
rect -196 76447 -184 76481
rect 184 76447 196 76481
rect -196 76441 196 76447
rect -252 76388 -206 76400
rect -252 76212 -246 76388
rect -212 76212 -206 76388
rect -252 76200 -206 76212
rect 206 76388 252 76400
rect 206 76212 212 76388
rect 246 76212 252 76388
rect 206 76200 252 76212
rect -196 76153 196 76159
rect -196 76119 -184 76153
rect 184 76119 196 76153
rect -196 76113 196 76119
rect -196 76045 196 76051
rect -196 76011 -184 76045
rect 184 76011 196 76045
rect -196 76005 196 76011
rect -252 75952 -206 75964
rect -252 75776 -246 75952
rect -212 75776 -206 75952
rect -252 75764 -206 75776
rect 206 75952 252 75964
rect 206 75776 212 75952
rect 246 75776 252 75952
rect 206 75764 252 75776
rect -196 75717 196 75723
rect -196 75683 -184 75717
rect 184 75683 196 75717
rect -196 75677 196 75683
rect -196 75609 196 75615
rect -196 75575 -184 75609
rect 184 75575 196 75609
rect -196 75569 196 75575
rect -252 75516 -206 75528
rect -252 75340 -246 75516
rect -212 75340 -206 75516
rect -252 75328 -206 75340
rect 206 75516 252 75528
rect 206 75340 212 75516
rect 246 75340 252 75516
rect 206 75328 252 75340
rect -196 75281 196 75287
rect -196 75247 -184 75281
rect 184 75247 196 75281
rect -196 75241 196 75247
rect -196 75173 196 75179
rect -196 75139 -184 75173
rect 184 75139 196 75173
rect -196 75133 196 75139
rect -252 75080 -206 75092
rect -252 74904 -246 75080
rect -212 74904 -206 75080
rect -252 74892 -206 74904
rect 206 75080 252 75092
rect 206 74904 212 75080
rect 246 74904 252 75080
rect 206 74892 252 74904
rect -196 74845 196 74851
rect -196 74811 -184 74845
rect 184 74811 196 74845
rect -196 74805 196 74811
rect -196 74737 196 74743
rect -196 74703 -184 74737
rect 184 74703 196 74737
rect -196 74697 196 74703
rect -252 74644 -206 74656
rect -252 74468 -246 74644
rect -212 74468 -206 74644
rect -252 74456 -206 74468
rect 206 74644 252 74656
rect 206 74468 212 74644
rect 246 74468 252 74644
rect 206 74456 252 74468
rect -196 74409 196 74415
rect -196 74375 -184 74409
rect 184 74375 196 74409
rect -196 74369 196 74375
rect -196 74301 196 74307
rect -196 74267 -184 74301
rect 184 74267 196 74301
rect -196 74261 196 74267
rect -252 74208 -206 74220
rect -252 74032 -246 74208
rect -212 74032 -206 74208
rect -252 74020 -206 74032
rect 206 74208 252 74220
rect 206 74032 212 74208
rect 246 74032 252 74208
rect 206 74020 252 74032
rect -196 73973 196 73979
rect -196 73939 -184 73973
rect 184 73939 196 73973
rect -196 73933 196 73939
rect -196 73865 196 73871
rect -196 73831 -184 73865
rect 184 73831 196 73865
rect -196 73825 196 73831
rect -252 73772 -206 73784
rect -252 73596 -246 73772
rect -212 73596 -206 73772
rect -252 73584 -206 73596
rect 206 73772 252 73784
rect 206 73596 212 73772
rect 246 73596 252 73772
rect 206 73584 252 73596
rect -196 73537 196 73543
rect -196 73503 -184 73537
rect 184 73503 196 73537
rect -196 73497 196 73503
rect -196 73429 196 73435
rect -196 73395 -184 73429
rect 184 73395 196 73429
rect -196 73389 196 73395
rect -252 73336 -206 73348
rect -252 73160 -246 73336
rect -212 73160 -206 73336
rect -252 73148 -206 73160
rect 206 73336 252 73348
rect 206 73160 212 73336
rect 246 73160 252 73336
rect 206 73148 252 73160
rect -196 73101 196 73107
rect -196 73067 -184 73101
rect 184 73067 196 73101
rect -196 73061 196 73067
rect -196 72993 196 72999
rect -196 72959 -184 72993
rect 184 72959 196 72993
rect -196 72953 196 72959
rect -252 72900 -206 72912
rect -252 72724 -246 72900
rect -212 72724 -206 72900
rect -252 72712 -206 72724
rect 206 72900 252 72912
rect 206 72724 212 72900
rect 246 72724 252 72900
rect 206 72712 252 72724
rect -196 72665 196 72671
rect -196 72631 -184 72665
rect 184 72631 196 72665
rect -196 72625 196 72631
rect -196 72557 196 72563
rect -196 72523 -184 72557
rect 184 72523 196 72557
rect -196 72517 196 72523
rect -252 72464 -206 72476
rect -252 72288 -246 72464
rect -212 72288 -206 72464
rect -252 72276 -206 72288
rect 206 72464 252 72476
rect 206 72288 212 72464
rect 246 72288 252 72464
rect 206 72276 252 72288
rect -196 72229 196 72235
rect -196 72195 -184 72229
rect 184 72195 196 72229
rect -196 72189 196 72195
rect -196 72121 196 72127
rect -196 72087 -184 72121
rect 184 72087 196 72121
rect -196 72081 196 72087
rect -252 72028 -206 72040
rect -252 71852 -246 72028
rect -212 71852 -206 72028
rect -252 71840 -206 71852
rect 206 72028 252 72040
rect 206 71852 212 72028
rect 246 71852 252 72028
rect 206 71840 252 71852
rect -196 71793 196 71799
rect -196 71759 -184 71793
rect 184 71759 196 71793
rect -196 71753 196 71759
rect -196 71685 196 71691
rect -196 71651 -184 71685
rect 184 71651 196 71685
rect -196 71645 196 71651
rect -252 71592 -206 71604
rect -252 71416 -246 71592
rect -212 71416 -206 71592
rect -252 71404 -206 71416
rect 206 71592 252 71604
rect 206 71416 212 71592
rect 246 71416 252 71592
rect 206 71404 252 71416
rect -196 71357 196 71363
rect -196 71323 -184 71357
rect 184 71323 196 71357
rect -196 71317 196 71323
rect -196 71249 196 71255
rect -196 71215 -184 71249
rect 184 71215 196 71249
rect -196 71209 196 71215
rect -252 71156 -206 71168
rect -252 70980 -246 71156
rect -212 70980 -206 71156
rect -252 70968 -206 70980
rect 206 71156 252 71168
rect 206 70980 212 71156
rect 246 70980 252 71156
rect 206 70968 252 70980
rect -196 70921 196 70927
rect -196 70887 -184 70921
rect 184 70887 196 70921
rect -196 70881 196 70887
rect -196 70813 196 70819
rect -196 70779 -184 70813
rect 184 70779 196 70813
rect -196 70773 196 70779
rect -252 70720 -206 70732
rect -252 70544 -246 70720
rect -212 70544 -206 70720
rect -252 70532 -206 70544
rect 206 70720 252 70732
rect 206 70544 212 70720
rect 246 70544 252 70720
rect 206 70532 252 70544
rect -196 70485 196 70491
rect -196 70451 -184 70485
rect 184 70451 196 70485
rect -196 70445 196 70451
rect -196 70377 196 70383
rect -196 70343 -184 70377
rect 184 70343 196 70377
rect -196 70337 196 70343
rect -252 70284 -206 70296
rect -252 70108 -246 70284
rect -212 70108 -206 70284
rect -252 70096 -206 70108
rect 206 70284 252 70296
rect 206 70108 212 70284
rect 246 70108 252 70284
rect 206 70096 252 70108
rect -196 70049 196 70055
rect -196 70015 -184 70049
rect 184 70015 196 70049
rect -196 70009 196 70015
rect -196 69941 196 69947
rect -196 69907 -184 69941
rect 184 69907 196 69941
rect -196 69901 196 69907
rect -252 69848 -206 69860
rect -252 69672 -246 69848
rect -212 69672 -206 69848
rect -252 69660 -206 69672
rect 206 69848 252 69860
rect 206 69672 212 69848
rect 246 69672 252 69848
rect 206 69660 252 69672
rect -196 69613 196 69619
rect -196 69579 -184 69613
rect 184 69579 196 69613
rect -196 69573 196 69579
rect -196 69505 196 69511
rect -196 69471 -184 69505
rect 184 69471 196 69505
rect -196 69465 196 69471
rect -252 69412 -206 69424
rect -252 69236 -246 69412
rect -212 69236 -206 69412
rect -252 69224 -206 69236
rect 206 69412 252 69424
rect 206 69236 212 69412
rect 246 69236 252 69412
rect 206 69224 252 69236
rect -196 69177 196 69183
rect -196 69143 -184 69177
rect 184 69143 196 69177
rect -196 69137 196 69143
rect -196 69069 196 69075
rect -196 69035 -184 69069
rect 184 69035 196 69069
rect -196 69029 196 69035
rect -252 68976 -206 68988
rect -252 68800 -246 68976
rect -212 68800 -206 68976
rect -252 68788 -206 68800
rect 206 68976 252 68988
rect 206 68800 212 68976
rect 246 68800 252 68976
rect 206 68788 252 68800
rect -196 68741 196 68747
rect -196 68707 -184 68741
rect 184 68707 196 68741
rect -196 68701 196 68707
rect -196 68633 196 68639
rect -196 68599 -184 68633
rect 184 68599 196 68633
rect -196 68593 196 68599
rect -252 68540 -206 68552
rect -252 68364 -246 68540
rect -212 68364 -206 68540
rect -252 68352 -206 68364
rect 206 68540 252 68552
rect 206 68364 212 68540
rect 246 68364 252 68540
rect 206 68352 252 68364
rect -196 68305 196 68311
rect -196 68271 -184 68305
rect 184 68271 196 68305
rect -196 68265 196 68271
rect -196 68197 196 68203
rect -196 68163 -184 68197
rect 184 68163 196 68197
rect -196 68157 196 68163
rect -252 68104 -206 68116
rect -252 67928 -246 68104
rect -212 67928 -206 68104
rect -252 67916 -206 67928
rect 206 68104 252 68116
rect 206 67928 212 68104
rect 246 67928 252 68104
rect 206 67916 252 67928
rect -196 67869 196 67875
rect -196 67835 -184 67869
rect 184 67835 196 67869
rect -196 67829 196 67835
rect -196 67761 196 67767
rect -196 67727 -184 67761
rect 184 67727 196 67761
rect -196 67721 196 67727
rect -252 67668 -206 67680
rect -252 67492 -246 67668
rect -212 67492 -206 67668
rect -252 67480 -206 67492
rect 206 67668 252 67680
rect 206 67492 212 67668
rect 246 67492 252 67668
rect 206 67480 252 67492
rect -196 67433 196 67439
rect -196 67399 -184 67433
rect 184 67399 196 67433
rect -196 67393 196 67399
rect -196 67325 196 67331
rect -196 67291 -184 67325
rect 184 67291 196 67325
rect -196 67285 196 67291
rect -252 67232 -206 67244
rect -252 67056 -246 67232
rect -212 67056 -206 67232
rect -252 67044 -206 67056
rect 206 67232 252 67244
rect 206 67056 212 67232
rect 246 67056 252 67232
rect 206 67044 252 67056
rect -196 66997 196 67003
rect -196 66963 -184 66997
rect 184 66963 196 66997
rect -196 66957 196 66963
rect -196 66889 196 66895
rect -196 66855 -184 66889
rect 184 66855 196 66889
rect -196 66849 196 66855
rect -252 66796 -206 66808
rect -252 66620 -246 66796
rect -212 66620 -206 66796
rect -252 66608 -206 66620
rect 206 66796 252 66808
rect 206 66620 212 66796
rect 246 66620 252 66796
rect 206 66608 252 66620
rect -196 66561 196 66567
rect -196 66527 -184 66561
rect 184 66527 196 66561
rect -196 66521 196 66527
rect -196 66453 196 66459
rect -196 66419 -184 66453
rect 184 66419 196 66453
rect -196 66413 196 66419
rect -252 66360 -206 66372
rect -252 66184 -246 66360
rect -212 66184 -206 66360
rect -252 66172 -206 66184
rect 206 66360 252 66372
rect 206 66184 212 66360
rect 246 66184 252 66360
rect 206 66172 252 66184
rect -196 66125 196 66131
rect -196 66091 -184 66125
rect 184 66091 196 66125
rect -196 66085 196 66091
rect -196 66017 196 66023
rect -196 65983 -184 66017
rect 184 65983 196 66017
rect -196 65977 196 65983
rect -252 65924 -206 65936
rect -252 65748 -246 65924
rect -212 65748 -206 65924
rect -252 65736 -206 65748
rect 206 65924 252 65936
rect 206 65748 212 65924
rect 246 65748 252 65924
rect 206 65736 252 65748
rect -196 65689 196 65695
rect -196 65655 -184 65689
rect 184 65655 196 65689
rect -196 65649 196 65655
rect -196 65581 196 65587
rect -196 65547 -184 65581
rect 184 65547 196 65581
rect -196 65541 196 65547
rect -252 65488 -206 65500
rect -252 65312 -246 65488
rect -212 65312 -206 65488
rect -252 65300 -206 65312
rect 206 65488 252 65500
rect 206 65312 212 65488
rect 246 65312 252 65488
rect 206 65300 252 65312
rect -196 65253 196 65259
rect -196 65219 -184 65253
rect 184 65219 196 65253
rect -196 65213 196 65219
rect -196 65145 196 65151
rect -196 65111 -184 65145
rect 184 65111 196 65145
rect -196 65105 196 65111
rect -252 65052 -206 65064
rect -252 64876 -246 65052
rect -212 64876 -206 65052
rect -252 64864 -206 64876
rect 206 65052 252 65064
rect 206 64876 212 65052
rect 246 64876 252 65052
rect 206 64864 252 64876
rect -196 64817 196 64823
rect -196 64783 -184 64817
rect 184 64783 196 64817
rect -196 64777 196 64783
rect -196 64709 196 64715
rect -196 64675 -184 64709
rect 184 64675 196 64709
rect -196 64669 196 64675
rect -252 64616 -206 64628
rect -252 64440 -246 64616
rect -212 64440 -206 64616
rect -252 64428 -206 64440
rect 206 64616 252 64628
rect 206 64440 212 64616
rect 246 64440 252 64616
rect 206 64428 252 64440
rect -196 64381 196 64387
rect -196 64347 -184 64381
rect 184 64347 196 64381
rect -196 64341 196 64347
rect -196 64273 196 64279
rect -196 64239 -184 64273
rect 184 64239 196 64273
rect -196 64233 196 64239
rect -252 64180 -206 64192
rect -252 64004 -246 64180
rect -212 64004 -206 64180
rect -252 63992 -206 64004
rect 206 64180 252 64192
rect 206 64004 212 64180
rect 246 64004 252 64180
rect 206 63992 252 64004
rect -196 63945 196 63951
rect -196 63911 -184 63945
rect 184 63911 196 63945
rect -196 63905 196 63911
rect -196 63837 196 63843
rect -196 63803 -184 63837
rect 184 63803 196 63837
rect -196 63797 196 63803
rect -252 63744 -206 63756
rect -252 63568 -246 63744
rect -212 63568 -206 63744
rect -252 63556 -206 63568
rect 206 63744 252 63756
rect 206 63568 212 63744
rect 246 63568 252 63744
rect 206 63556 252 63568
rect -196 63509 196 63515
rect -196 63475 -184 63509
rect 184 63475 196 63509
rect -196 63469 196 63475
rect -196 63401 196 63407
rect -196 63367 -184 63401
rect 184 63367 196 63401
rect -196 63361 196 63367
rect -252 63308 -206 63320
rect -252 63132 -246 63308
rect -212 63132 -206 63308
rect -252 63120 -206 63132
rect 206 63308 252 63320
rect 206 63132 212 63308
rect 246 63132 252 63308
rect 206 63120 252 63132
rect -196 63073 196 63079
rect -196 63039 -184 63073
rect 184 63039 196 63073
rect -196 63033 196 63039
rect -196 62965 196 62971
rect -196 62931 -184 62965
rect 184 62931 196 62965
rect -196 62925 196 62931
rect -252 62872 -206 62884
rect -252 62696 -246 62872
rect -212 62696 -206 62872
rect -252 62684 -206 62696
rect 206 62872 252 62884
rect 206 62696 212 62872
rect 246 62696 252 62872
rect 206 62684 252 62696
rect -196 62637 196 62643
rect -196 62603 -184 62637
rect 184 62603 196 62637
rect -196 62597 196 62603
rect -196 62529 196 62535
rect -196 62495 -184 62529
rect 184 62495 196 62529
rect -196 62489 196 62495
rect -252 62436 -206 62448
rect -252 62260 -246 62436
rect -212 62260 -206 62436
rect -252 62248 -206 62260
rect 206 62436 252 62448
rect 206 62260 212 62436
rect 246 62260 252 62436
rect 206 62248 252 62260
rect -196 62201 196 62207
rect -196 62167 -184 62201
rect 184 62167 196 62201
rect -196 62161 196 62167
rect -196 62093 196 62099
rect -196 62059 -184 62093
rect 184 62059 196 62093
rect -196 62053 196 62059
rect -252 62000 -206 62012
rect -252 61824 -246 62000
rect -212 61824 -206 62000
rect -252 61812 -206 61824
rect 206 62000 252 62012
rect 206 61824 212 62000
rect 246 61824 252 62000
rect 206 61812 252 61824
rect -196 61765 196 61771
rect -196 61731 -184 61765
rect 184 61731 196 61765
rect -196 61725 196 61731
rect -196 61657 196 61663
rect -196 61623 -184 61657
rect 184 61623 196 61657
rect -196 61617 196 61623
rect -252 61564 -206 61576
rect -252 61388 -246 61564
rect -212 61388 -206 61564
rect -252 61376 -206 61388
rect 206 61564 252 61576
rect 206 61388 212 61564
rect 246 61388 252 61564
rect 206 61376 252 61388
rect -196 61329 196 61335
rect -196 61295 -184 61329
rect 184 61295 196 61329
rect -196 61289 196 61295
rect -196 61221 196 61227
rect -196 61187 -184 61221
rect 184 61187 196 61221
rect -196 61181 196 61187
rect -252 61128 -206 61140
rect -252 60952 -246 61128
rect -212 60952 -206 61128
rect -252 60940 -206 60952
rect 206 61128 252 61140
rect 206 60952 212 61128
rect 246 60952 252 61128
rect 206 60940 252 60952
rect -196 60893 196 60899
rect -196 60859 -184 60893
rect 184 60859 196 60893
rect -196 60853 196 60859
rect -196 60785 196 60791
rect -196 60751 -184 60785
rect 184 60751 196 60785
rect -196 60745 196 60751
rect -252 60692 -206 60704
rect -252 60516 -246 60692
rect -212 60516 -206 60692
rect -252 60504 -206 60516
rect 206 60692 252 60704
rect 206 60516 212 60692
rect 246 60516 252 60692
rect 206 60504 252 60516
rect -196 60457 196 60463
rect -196 60423 -184 60457
rect 184 60423 196 60457
rect -196 60417 196 60423
rect -196 60349 196 60355
rect -196 60315 -184 60349
rect 184 60315 196 60349
rect -196 60309 196 60315
rect -252 60256 -206 60268
rect -252 60080 -246 60256
rect -212 60080 -206 60256
rect -252 60068 -206 60080
rect 206 60256 252 60268
rect 206 60080 212 60256
rect 246 60080 252 60256
rect 206 60068 252 60080
rect -196 60021 196 60027
rect -196 59987 -184 60021
rect 184 59987 196 60021
rect -196 59981 196 59987
rect -196 59913 196 59919
rect -196 59879 -184 59913
rect 184 59879 196 59913
rect -196 59873 196 59879
rect -252 59820 -206 59832
rect -252 59644 -246 59820
rect -212 59644 -206 59820
rect -252 59632 -206 59644
rect 206 59820 252 59832
rect 206 59644 212 59820
rect 246 59644 252 59820
rect 206 59632 252 59644
rect -196 59585 196 59591
rect -196 59551 -184 59585
rect 184 59551 196 59585
rect -196 59545 196 59551
rect -196 59477 196 59483
rect -196 59443 -184 59477
rect 184 59443 196 59477
rect -196 59437 196 59443
rect -252 59384 -206 59396
rect -252 59208 -246 59384
rect -212 59208 -206 59384
rect -252 59196 -206 59208
rect 206 59384 252 59396
rect 206 59208 212 59384
rect 246 59208 252 59384
rect 206 59196 252 59208
rect -196 59149 196 59155
rect -196 59115 -184 59149
rect 184 59115 196 59149
rect -196 59109 196 59115
rect -196 59041 196 59047
rect -196 59007 -184 59041
rect 184 59007 196 59041
rect -196 59001 196 59007
rect -252 58948 -206 58960
rect -252 58772 -246 58948
rect -212 58772 -206 58948
rect -252 58760 -206 58772
rect 206 58948 252 58960
rect 206 58772 212 58948
rect 246 58772 252 58948
rect 206 58760 252 58772
rect -196 58713 196 58719
rect -196 58679 -184 58713
rect 184 58679 196 58713
rect -196 58673 196 58679
rect -196 58605 196 58611
rect -196 58571 -184 58605
rect 184 58571 196 58605
rect -196 58565 196 58571
rect -252 58512 -206 58524
rect -252 58336 -246 58512
rect -212 58336 -206 58512
rect -252 58324 -206 58336
rect 206 58512 252 58524
rect 206 58336 212 58512
rect 246 58336 252 58512
rect 206 58324 252 58336
rect -196 58277 196 58283
rect -196 58243 -184 58277
rect 184 58243 196 58277
rect -196 58237 196 58243
rect -196 58169 196 58175
rect -196 58135 -184 58169
rect 184 58135 196 58169
rect -196 58129 196 58135
rect -252 58076 -206 58088
rect -252 57900 -246 58076
rect -212 57900 -206 58076
rect -252 57888 -206 57900
rect 206 58076 252 58088
rect 206 57900 212 58076
rect 246 57900 252 58076
rect 206 57888 252 57900
rect -196 57841 196 57847
rect -196 57807 -184 57841
rect 184 57807 196 57841
rect -196 57801 196 57807
rect -196 57733 196 57739
rect -196 57699 -184 57733
rect 184 57699 196 57733
rect -196 57693 196 57699
rect -252 57640 -206 57652
rect -252 57464 -246 57640
rect -212 57464 -206 57640
rect -252 57452 -206 57464
rect 206 57640 252 57652
rect 206 57464 212 57640
rect 246 57464 252 57640
rect 206 57452 252 57464
rect -196 57405 196 57411
rect -196 57371 -184 57405
rect 184 57371 196 57405
rect -196 57365 196 57371
rect -196 57297 196 57303
rect -196 57263 -184 57297
rect 184 57263 196 57297
rect -196 57257 196 57263
rect -252 57204 -206 57216
rect -252 57028 -246 57204
rect -212 57028 -206 57204
rect -252 57016 -206 57028
rect 206 57204 252 57216
rect 206 57028 212 57204
rect 246 57028 252 57204
rect 206 57016 252 57028
rect -196 56969 196 56975
rect -196 56935 -184 56969
rect 184 56935 196 56969
rect -196 56929 196 56935
rect -196 56861 196 56867
rect -196 56827 -184 56861
rect 184 56827 196 56861
rect -196 56821 196 56827
rect -252 56768 -206 56780
rect -252 56592 -246 56768
rect -212 56592 -206 56768
rect -252 56580 -206 56592
rect 206 56768 252 56780
rect 206 56592 212 56768
rect 246 56592 252 56768
rect 206 56580 252 56592
rect -196 56533 196 56539
rect -196 56499 -184 56533
rect 184 56499 196 56533
rect -196 56493 196 56499
rect -196 56425 196 56431
rect -196 56391 -184 56425
rect 184 56391 196 56425
rect -196 56385 196 56391
rect -252 56332 -206 56344
rect -252 56156 -246 56332
rect -212 56156 -206 56332
rect -252 56144 -206 56156
rect 206 56332 252 56344
rect 206 56156 212 56332
rect 246 56156 252 56332
rect 206 56144 252 56156
rect -196 56097 196 56103
rect -196 56063 -184 56097
rect 184 56063 196 56097
rect -196 56057 196 56063
rect -196 55989 196 55995
rect -196 55955 -184 55989
rect 184 55955 196 55989
rect -196 55949 196 55955
rect -252 55896 -206 55908
rect -252 55720 -246 55896
rect -212 55720 -206 55896
rect -252 55708 -206 55720
rect 206 55896 252 55908
rect 206 55720 212 55896
rect 246 55720 252 55896
rect 206 55708 252 55720
rect -196 55661 196 55667
rect -196 55627 -184 55661
rect 184 55627 196 55661
rect -196 55621 196 55627
rect -196 55553 196 55559
rect -196 55519 -184 55553
rect 184 55519 196 55553
rect -196 55513 196 55519
rect -252 55460 -206 55472
rect -252 55284 -246 55460
rect -212 55284 -206 55460
rect -252 55272 -206 55284
rect 206 55460 252 55472
rect 206 55284 212 55460
rect 246 55284 252 55460
rect 206 55272 252 55284
rect -196 55225 196 55231
rect -196 55191 -184 55225
rect 184 55191 196 55225
rect -196 55185 196 55191
rect -196 55117 196 55123
rect -196 55083 -184 55117
rect 184 55083 196 55117
rect -196 55077 196 55083
rect -252 55024 -206 55036
rect -252 54848 -246 55024
rect -212 54848 -206 55024
rect -252 54836 -206 54848
rect 206 55024 252 55036
rect 206 54848 212 55024
rect 246 54848 252 55024
rect 206 54836 252 54848
rect -196 54789 196 54795
rect -196 54755 -184 54789
rect 184 54755 196 54789
rect -196 54749 196 54755
rect -196 54681 196 54687
rect -196 54647 -184 54681
rect 184 54647 196 54681
rect -196 54641 196 54647
rect -252 54588 -206 54600
rect -252 54412 -246 54588
rect -212 54412 -206 54588
rect -252 54400 -206 54412
rect 206 54588 252 54600
rect 206 54412 212 54588
rect 246 54412 252 54588
rect 206 54400 252 54412
rect -196 54353 196 54359
rect -196 54319 -184 54353
rect 184 54319 196 54353
rect -196 54313 196 54319
rect -196 54245 196 54251
rect -196 54211 -184 54245
rect 184 54211 196 54245
rect -196 54205 196 54211
rect -252 54152 -206 54164
rect -252 53976 -246 54152
rect -212 53976 -206 54152
rect -252 53964 -206 53976
rect 206 54152 252 54164
rect 206 53976 212 54152
rect 246 53976 252 54152
rect 206 53964 252 53976
rect -196 53917 196 53923
rect -196 53883 -184 53917
rect 184 53883 196 53917
rect -196 53877 196 53883
rect -196 53809 196 53815
rect -196 53775 -184 53809
rect 184 53775 196 53809
rect -196 53769 196 53775
rect -252 53716 -206 53728
rect -252 53540 -246 53716
rect -212 53540 -206 53716
rect -252 53528 -206 53540
rect 206 53716 252 53728
rect 206 53540 212 53716
rect 246 53540 252 53716
rect 206 53528 252 53540
rect -196 53481 196 53487
rect -196 53447 -184 53481
rect 184 53447 196 53481
rect -196 53441 196 53447
rect -196 53373 196 53379
rect -196 53339 -184 53373
rect 184 53339 196 53373
rect -196 53333 196 53339
rect -252 53280 -206 53292
rect -252 53104 -246 53280
rect -212 53104 -206 53280
rect -252 53092 -206 53104
rect 206 53280 252 53292
rect 206 53104 212 53280
rect 246 53104 252 53280
rect 206 53092 252 53104
rect -196 53045 196 53051
rect -196 53011 -184 53045
rect 184 53011 196 53045
rect -196 53005 196 53011
rect -196 52937 196 52943
rect -196 52903 -184 52937
rect 184 52903 196 52937
rect -196 52897 196 52903
rect -252 52844 -206 52856
rect -252 52668 -246 52844
rect -212 52668 -206 52844
rect -252 52656 -206 52668
rect 206 52844 252 52856
rect 206 52668 212 52844
rect 246 52668 252 52844
rect 206 52656 252 52668
rect -196 52609 196 52615
rect -196 52575 -184 52609
rect 184 52575 196 52609
rect -196 52569 196 52575
rect -196 52501 196 52507
rect -196 52467 -184 52501
rect 184 52467 196 52501
rect -196 52461 196 52467
rect -252 52408 -206 52420
rect -252 52232 -246 52408
rect -212 52232 -206 52408
rect -252 52220 -206 52232
rect 206 52408 252 52420
rect 206 52232 212 52408
rect 246 52232 252 52408
rect 206 52220 252 52232
rect -196 52173 196 52179
rect -196 52139 -184 52173
rect 184 52139 196 52173
rect -196 52133 196 52139
rect -196 52065 196 52071
rect -196 52031 -184 52065
rect 184 52031 196 52065
rect -196 52025 196 52031
rect -252 51972 -206 51984
rect -252 51796 -246 51972
rect -212 51796 -206 51972
rect -252 51784 -206 51796
rect 206 51972 252 51984
rect 206 51796 212 51972
rect 246 51796 252 51972
rect 206 51784 252 51796
rect -196 51737 196 51743
rect -196 51703 -184 51737
rect 184 51703 196 51737
rect -196 51697 196 51703
rect -196 51629 196 51635
rect -196 51595 -184 51629
rect 184 51595 196 51629
rect -196 51589 196 51595
rect -252 51536 -206 51548
rect -252 51360 -246 51536
rect -212 51360 -206 51536
rect -252 51348 -206 51360
rect 206 51536 252 51548
rect 206 51360 212 51536
rect 246 51360 252 51536
rect 206 51348 252 51360
rect -196 51301 196 51307
rect -196 51267 -184 51301
rect 184 51267 196 51301
rect -196 51261 196 51267
rect -196 51193 196 51199
rect -196 51159 -184 51193
rect 184 51159 196 51193
rect -196 51153 196 51159
rect -252 51100 -206 51112
rect -252 50924 -246 51100
rect -212 50924 -206 51100
rect -252 50912 -206 50924
rect 206 51100 252 51112
rect 206 50924 212 51100
rect 246 50924 252 51100
rect 206 50912 252 50924
rect -196 50865 196 50871
rect -196 50831 -184 50865
rect 184 50831 196 50865
rect -196 50825 196 50831
rect -196 50757 196 50763
rect -196 50723 -184 50757
rect 184 50723 196 50757
rect -196 50717 196 50723
rect -252 50664 -206 50676
rect -252 50488 -246 50664
rect -212 50488 -206 50664
rect -252 50476 -206 50488
rect 206 50664 252 50676
rect 206 50488 212 50664
rect 246 50488 252 50664
rect 206 50476 252 50488
rect -196 50429 196 50435
rect -196 50395 -184 50429
rect 184 50395 196 50429
rect -196 50389 196 50395
rect -196 50321 196 50327
rect -196 50287 -184 50321
rect 184 50287 196 50321
rect -196 50281 196 50287
rect -252 50228 -206 50240
rect -252 50052 -246 50228
rect -212 50052 -206 50228
rect -252 50040 -206 50052
rect 206 50228 252 50240
rect 206 50052 212 50228
rect 246 50052 252 50228
rect 206 50040 252 50052
rect -196 49993 196 49999
rect -196 49959 -184 49993
rect 184 49959 196 49993
rect -196 49953 196 49959
rect -196 49885 196 49891
rect -196 49851 -184 49885
rect 184 49851 196 49885
rect -196 49845 196 49851
rect -252 49792 -206 49804
rect -252 49616 -246 49792
rect -212 49616 -206 49792
rect -252 49604 -206 49616
rect 206 49792 252 49804
rect 206 49616 212 49792
rect 246 49616 252 49792
rect 206 49604 252 49616
rect -196 49557 196 49563
rect -196 49523 -184 49557
rect 184 49523 196 49557
rect -196 49517 196 49523
rect -196 49449 196 49455
rect -196 49415 -184 49449
rect 184 49415 196 49449
rect -196 49409 196 49415
rect -252 49356 -206 49368
rect -252 49180 -246 49356
rect -212 49180 -206 49356
rect -252 49168 -206 49180
rect 206 49356 252 49368
rect 206 49180 212 49356
rect 246 49180 252 49356
rect 206 49168 252 49180
rect -196 49121 196 49127
rect -196 49087 -184 49121
rect 184 49087 196 49121
rect -196 49081 196 49087
rect -196 49013 196 49019
rect -196 48979 -184 49013
rect 184 48979 196 49013
rect -196 48973 196 48979
rect -252 48920 -206 48932
rect -252 48744 -246 48920
rect -212 48744 -206 48920
rect -252 48732 -206 48744
rect 206 48920 252 48932
rect 206 48744 212 48920
rect 246 48744 252 48920
rect 206 48732 252 48744
rect -196 48685 196 48691
rect -196 48651 -184 48685
rect 184 48651 196 48685
rect -196 48645 196 48651
rect -196 48577 196 48583
rect -196 48543 -184 48577
rect 184 48543 196 48577
rect -196 48537 196 48543
rect -252 48484 -206 48496
rect -252 48308 -246 48484
rect -212 48308 -206 48484
rect -252 48296 -206 48308
rect 206 48484 252 48496
rect 206 48308 212 48484
rect 246 48308 252 48484
rect 206 48296 252 48308
rect -196 48249 196 48255
rect -196 48215 -184 48249
rect 184 48215 196 48249
rect -196 48209 196 48215
rect -196 48141 196 48147
rect -196 48107 -184 48141
rect 184 48107 196 48141
rect -196 48101 196 48107
rect -252 48048 -206 48060
rect -252 47872 -246 48048
rect -212 47872 -206 48048
rect -252 47860 -206 47872
rect 206 48048 252 48060
rect 206 47872 212 48048
rect 246 47872 252 48048
rect 206 47860 252 47872
rect -196 47813 196 47819
rect -196 47779 -184 47813
rect 184 47779 196 47813
rect -196 47773 196 47779
rect -196 47705 196 47711
rect -196 47671 -184 47705
rect 184 47671 196 47705
rect -196 47665 196 47671
rect -252 47612 -206 47624
rect -252 47436 -246 47612
rect -212 47436 -206 47612
rect -252 47424 -206 47436
rect 206 47612 252 47624
rect 206 47436 212 47612
rect 246 47436 252 47612
rect 206 47424 252 47436
rect -196 47377 196 47383
rect -196 47343 -184 47377
rect 184 47343 196 47377
rect -196 47337 196 47343
rect -196 47269 196 47275
rect -196 47235 -184 47269
rect 184 47235 196 47269
rect -196 47229 196 47235
rect -252 47176 -206 47188
rect -252 47000 -246 47176
rect -212 47000 -206 47176
rect -252 46988 -206 47000
rect 206 47176 252 47188
rect 206 47000 212 47176
rect 246 47000 252 47176
rect 206 46988 252 47000
rect -196 46941 196 46947
rect -196 46907 -184 46941
rect 184 46907 196 46941
rect -196 46901 196 46907
rect -196 46833 196 46839
rect -196 46799 -184 46833
rect 184 46799 196 46833
rect -196 46793 196 46799
rect -252 46740 -206 46752
rect -252 46564 -246 46740
rect -212 46564 -206 46740
rect -252 46552 -206 46564
rect 206 46740 252 46752
rect 206 46564 212 46740
rect 246 46564 252 46740
rect 206 46552 252 46564
rect -196 46505 196 46511
rect -196 46471 -184 46505
rect 184 46471 196 46505
rect -196 46465 196 46471
rect -196 46397 196 46403
rect -196 46363 -184 46397
rect 184 46363 196 46397
rect -196 46357 196 46363
rect -252 46304 -206 46316
rect -252 46128 -246 46304
rect -212 46128 -206 46304
rect -252 46116 -206 46128
rect 206 46304 252 46316
rect 206 46128 212 46304
rect 246 46128 252 46304
rect 206 46116 252 46128
rect -196 46069 196 46075
rect -196 46035 -184 46069
rect 184 46035 196 46069
rect -196 46029 196 46035
rect -196 45961 196 45967
rect -196 45927 -184 45961
rect 184 45927 196 45961
rect -196 45921 196 45927
rect -252 45868 -206 45880
rect -252 45692 -246 45868
rect -212 45692 -206 45868
rect -252 45680 -206 45692
rect 206 45868 252 45880
rect 206 45692 212 45868
rect 246 45692 252 45868
rect 206 45680 252 45692
rect -196 45633 196 45639
rect -196 45599 -184 45633
rect 184 45599 196 45633
rect -196 45593 196 45599
rect -196 45525 196 45531
rect -196 45491 -184 45525
rect 184 45491 196 45525
rect -196 45485 196 45491
rect -252 45432 -206 45444
rect -252 45256 -246 45432
rect -212 45256 -206 45432
rect -252 45244 -206 45256
rect 206 45432 252 45444
rect 206 45256 212 45432
rect 246 45256 252 45432
rect 206 45244 252 45256
rect -196 45197 196 45203
rect -196 45163 -184 45197
rect 184 45163 196 45197
rect -196 45157 196 45163
rect -196 45089 196 45095
rect -196 45055 -184 45089
rect 184 45055 196 45089
rect -196 45049 196 45055
rect -252 44996 -206 45008
rect -252 44820 -246 44996
rect -212 44820 -206 44996
rect -252 44808 -206 44820
rect 206 44996 252 45008
rect 206 44820 212 44996
rect 246 44820 252 44996
rect 206 44808 252 44820
rect -196 44761 196 44767
rect -196 44727 -184 44761
rect 184 44727 196 44761
rect -196 44721 196 44727
rect -196 44653 196 44659
rect -196 44619 -184 44653
rect 184 44619 196 44653
rect -196 44613 196 44619
rect -252 44560 -206 44572
rect -252 44384 -246 44560
rect -212 44384 -206 44560
rect -252 44372 -206 44384
rect 206 44560 252 44572
rect 206 44384 212 44560
rect 246 44384 252 44560
rect 206 44372 252 44384
rect -196 44325 196 44331
rect -196 44291 -184 44325
rect 184 44291 196 44325
rect -196 44285 196 44291
rect -196 44217 196 44223
rect -196 44183 -184 44217
rect 184 44183 196 44217
rect -196 44177 196 44183
rect -252 44124 -206 44136
rect -252 43948 -246 44124
rect -212 43948 -206 44124
rect -252 43936 -206 43948
rect 206 44124 252 44136
rect 206 43948 212 44124
rect 246 43948 252 44124
rect 206 43936 252 43948
rect -196 43889 196 43895
rect -196 43855 -184 43889
rect 184 43855 196 43889
rect -196 43849 196 43855
rect -196 43781 196 43787
rect -196 43747 -184 43781
rect 184 43747 196 43781
rect -196 43741 196 43747
rect -252 43688 -206 43700
rect -252 43512 -246 43688
rect -212 43512 -206 43688
rect -252 43500 -206 43512
rect 206 43688 252 43700
rect 206 43512 212 43688
rect 246 43512 252 43688
rect 206 43500 252 43512
rect -196 43453 196 43459
rect -196 43419 -184 43453
rect 184 43419 196 43453
rect -196 43413 196 43419
rect -196 43345 196 43351
rect -196 43311 -184 43345
rect 184 43311 196 43345
rect -196 43305 196 43311
rect -252 43252 -206 43264
rect -252 43076 -246 43252
rect -212 43076 -206 43252
rect -252 43064 -206 43076
rect 206 43252 252 43264
rect 206 43076 212 43252
rect 246 43076 252 43252
rect 206 43064 252 43076
rect -196 43017 196 43023
rect -196 42983 -184 43017
rect 184 42983 196 43017
rect -196 42977 196 42983
rect -196 42909 196 42915
rect -196 42875 -184 42909
rect 184 42875 196 42909
rect -196 42869 196 42875
rect -252 42816 -206 42828
rect -252 42640 -246 42816
rect -212 42640 -206 42816
rect -252 42628 -206 42640
rect 206 42816 252 42828
rect 206 42640 212 42816
rect 246 42640 252 42816
rect 206 42628 252 42640
rect -196 42581 196 42587
rect -196 42547 -184 42581
rect 184 42547 196 42581
rect -196 42541 196 42547
rect -196 42473 196 42479
rect -196 42439 -184 42473
rect 184 42439 196 42473
rect -196 42433 196 42439
rect -252 42380 -206 42392
rect -252 42204 -246 42380
rect -212 42204 -206 42380
rect -252 42192 -206 42204
rect 206 42380 252 42392
rect 206 42204 212 42380
rect 246 42204 252 42380
rect 206 42192 252 42204
rect -196 42145 196 42151
rect -196 42111 -184 42145
rect 184 42111 196 42145
rect -196 42105 196 42111
rect -196 42037 196 42043
rect -196 42003 -184 42037
rect 184 42003 196 42037
rect -196 41997 196 42003
rect -252 41944 -206 41956
rect -252 41768 -246 41944
rect -212 41768 -206 41944
rect -252 41756 -206 41768
rect 206 41944 252 41956
rect 206 41768 212 41944
rect 246 41768 252 41944
rect 206 41756 252 41768
rect -196 41709 196 41715
rect -196 41675 -184 41709
rect 184 41675 196 41709
rect -196 41669 196 41675
rect -196 41601 196 41607
rect -196 41567 -184 41601
rect 184 41567 196 41601
rect -196 41561 196 41567
rect -252 41508 -206 41520
rect -252 41332 -246 41508
rect -212 41332 -206 41508
rect -252 41320 -206 41332
rect 206 41508 252 41520
rect 206 41332 212 41508
rect 246 41332 252 41508
rect 206 41320 252 41332
rect -196 41273 196 41279
rect -196 41239 -184 41273
rect 184 41239 196 41273
rect -196 41233 196 41239
rect -196 41165 196 41171
rect -196 41131 -184 41165
rect 184 41131 196 41165
rect -196 41125 196 41131
rect -252 41072 -206 41084
rect -252 40896 -246 41072
rect -212 40896 -206 41072
rect -252 40884 -206 40896
rect 206 41072 252 41084
rect 206 40896 212 41072
rect 246 40896 252 41072
rect 206 40884 252 40896
rect -196 40837 196 40843
rect -196 40803 -184 40837
rect 184 40803 196 40837
rect -196 40797 196 40803
rect -196 40729 196 40735
rect -196 40695 -184 40729
rect 184 40695 196 40729
rect -196 40689 196 40695
rect -252 40636 -206 40648
rect -252 40460 -246 40636
rect -212 40460 -206 40636
rect -252 40448 -206 40460
rect 206 40636 252 40648
rect 206 40460 212 40636
rect 246 40460 252 40636
rect 206 40448 252 40460
rect -196 40401 196 40407
rect -196 40367 -184 40401
rect 184 40367 196 40401
rect -196 40361 196 40367
rect -196 40293 196 40299
rect -196 40259 -184 40293
rect 184 40259 196 40293
rect -196 40253 196 40259
rect -252 40200 -206 40212
rect -252 40024 -246 40200
rect -212 40024 -206 40200
rect -252 40012 -206 40024
rect 206 40200 252 40212
rect 206 40024 212 40200
rect 246 40024 252 40200
rect 206 40012 252 40024
rect -196 39965 196 39971
rect -196 39931 -184 39965
rect 184 39931 196 39965
rect -196 39925 196 39931
rect -196 39857 196 39863
rect -196 39823 -184 39857
rect 184 39823 196 39857
rect -196 39817 196 39823
rect -252 39764 -206 39776
rect -252 39588 -246 39764
rect -212 39588 -206 39764
rect -252 39576 -206 39588
rect 206 39764 252 39776
rect 206 39588 212 39764
rect 246 39588 252 39764
rect 206 39576 252 39588
rect -196 39529 196 39535
rect -196 39495 -184 39529
rect 184 39495 196 39529
rect -196 39489 196 39495
rect -196 39421 196 39427
rect -196 39387 -184 39421
rect 184 39387 196 39421
rect -196 39381 196 39387
rect -252 39328 -206 39340
rect -252 39152 -246 39328
rect -212 39152 -206 39328
rect -252 39140 -206 39152
rect 206 39328 252 39340
rect 206 39152 212 39328
rect 246 39152 252 39328
rect 206 39140 252 39152
rect -196 39093 196 39099
rect -196 39059 -184 39093
rect 184 39059 196 39093
rect -196 39053 196 39059
rect -196 38985 196 38991
rect -196 38951 -184 38985
rect 184 38951 196 38985
rect -196 38945 196 38951
rect -252 38892 -206 38904
rect -252 38716 -246 38892
rect -212 38716 -206 38892
rect -252 38704 -206 38716
rect 206 38892 252 38904
rect 206 38716 212 38892
rect 246 38716 252 38892
rect 206 38704 252 38716
rect -196 38657 196 38663
rect -196 38623 -184 38657
rect 184 38623 196 38657
rect -196 38617 196 38623
rect -196 38549 196 38555
rect -196 38515 -184 38549
rect 184 38515 196 38549
rect -196 38509 196 38515
rect -252 38456 -206 38468
rect -252 38280 -246 38456
rect -212 38280 -206 38456
rect -252 38268 -206 38280
rect 206 38456 252 38468
rect 206 38280 212 38456
rect 246 38280 252 38456
rect 206 38268 252 38280
rect -196 38221 196 38227
rect -196 38187 -184 38221
rect 184 38187 196 38221
rect -196 38181 196 38187
rect -196 38113 196 38119
rect -196 38079 -184 38113
rect 184 38079 196 38113
rect -196 38073 196 38079
rect -252 38020 -206 38032
rect -252 37844 -246 38020
rect -212 37844 -206 38020
rect -252 37832 -206 37844
rect 206 38020 252 38032
rect 206 37844 212 38020
rect 246 37844 252 38020
rect 206 37832 252 37844
rect -196 37785 196 37791
rect -196 37751 -184 37785
rect 184 37751 196 37785
rect -196 37745 196 37751
rect -196 37677 196 37683
rect -196 37643 -184 37677
rect 184 37643 196 37677
rect -196 37637 196 37643
rect -252 37584 -206 37596
rect -252 37408 -246 37584
rect -212 37408 -206 37584
rect -252 37396 -206 37408
rect 206 37584 252 37596
rect 206 37408 212 37584
rect 246 37408 252 37584
rect 206 37396 252 37408
rect -196 37349 196 37355
rect -196 37315 -184 37349
rect 184 37315 196 37349
rect -196 37309 196 37315
rect -196 37241 196 37247
rect -196 37207 -184 37241
rect 184 37207 196 37241
rect -196 37201 196 37207
rect -252 37148 -206 37160
rect -252 36972 -246 37148
rect -212 36972 -206 37148
rect -252 36960 -206 36972
rect 206 37148 252 37160
rect 206 36972 212 37148
rect 246 36972 252 37148
rect 206 36960 252 36972
rect -196 36913 196 36919
rect -196 36879 -184 36913
rect 184 36879 196 36913
rect -196 36873 196 36879
rect -196 36805 196 36811
rect -196 36771 -184 36805
rect 184 36771 196 36805
rect -196 36765 196 36771
rect -252 36712 -206 36724
rect -252 36536 -246 36712
rect -212 36536 -206 36712
rect -252 36524 -206 36536
rect 206 36712 252 36724
rect 206 36536 212 36712
rect 246 36536 252 36712
rect 206 36524 252 36536
rect -196 36477 196 36483
rect -196 36443 -184 36477
rect 184 36443 196 36477
rect -196 36437 196 36443
rect -196 36369 196 36375
rect -196 36335 -184 36369
rect 184 36335 196 36369
rect -196 36329 196 36335
rect -252 36276 -206 36288
rect -252 36100 -246 36276
rect -212 36100 -206 36276
rect -252 36088 -206 36100
rect 206 36276 252 36288
rect 206 36100 212 36276
rect 246 36100 252 36276
rect 206 36088 252 36100
rect -196 36041 196 36047
rect -196 36007 -184 36041
rect 184 36007 196 36041
rect -196 36001 196 36007
rect -196 35933 196 35939
rect -196 35899 -184 35933
rect 184 35899 196 35933
rect -196 35893 196 35899
rect -252 35840 -206 35852
rect -252 35664 -246 35840
rect -212 35664 -206 35840
rect -252 35652 -206 35664
rect 206 35840 252 35852
rect 206 35664 212 35840
rect 246 35664 252 35840
rect 206 35652 252 35664
rect -196 35605 196 35611
rect -196 35571 -184 35605
rect 184 35571 196 35605
rect -196 35565 196 35571
rect -196 35497 196 35503
rect -196 35463 -184 35497
rect 184 35463 196 35497
rect -196 35457 196 35463
rect -252 35404 -206 35416
rect -252 35228 -246 35404
rect -212 35228 -206 35404
rect -252 35216 -206 35228
rect 206 35404 252 35416
rect 206 35228 212 35404
rect 246 35228 252 35404
rect 206 35216 252 35228
rect -196 35169 196 35175
rect -196 35135 -184 35169
rect 184 35135 196 35169
rect -196 35129 196 35135
rect -196 35061 196 35067
rect -196 35027 -184 35061
rect 184 35027 196 35061
rect -196 35021 196 35027
rect -252 34968 -206 34980
rect -252 34792 -246 34968
rect -212 34792 -206 34968
rect -252 34780 -206 34792
rect 206 34968 252 34980
rect 206 34792 212 34968
rect 246 34792 252 34968
rect 206 34780 252 34792
rect -196 34733 196 34739
rect -196 34699 -184 34733
rect 184 34699 196 34733
rect -196 34693 196 34699
rect -196 34625 196 34631
rect -196 34591 -184 34625
rect 184 34591 196 34625
rect -196 34585 196 34591
rect -252 34532 -206 34544
rect -252 34356 -246 34532
rect -212 34356 -206 34532
rect -252 34344 -206 34356
rect 206 34532 252 34544
rect 206 34356 212 34532
rect 246 34356 252 34532
rect 206 34344 252 34356
rect -196 34297 196 34303
rect -196 34263 -184 34297
rect 184 34263 196 34297
rect -196 34257 196 34263
rect -196 34189 196 34195
rect -196 34155 -184 34189
rect 184 34155 196 34189
rect -196 34149 196 34155
rect -252 34096 -206 34108
rect -252 33920 -246 34096
rect -212 33920 -206 34096
rect -252 33908 -206 33920
rect 206 34096 252 34108
rect 206 33920 212 34096
rect 246 33920 252 34096
rect 206 33908 252 33920
rect -196 33861 196 33867
rect -196 33827 -184 33861
rect 184 33827 196 33861
rect -196 33821 196 33827
rect -196 33753 196 33759
rect -196 33719 -184 33753
rect 184 33719 196 33753
rect -196 33713 196 33719
rect -252 33660 -206 33672
rect -252 33484 -246 33660
rect -212 33484 -206 33660
rect -252 33472 -206 33484
rect 206 33660 252 33672
rect 206 33484 212 33660
rect 246 33484 252 33660
rect 206 33472 252 33484
rect -196 33425 196 33431
rect -196 33391 -184 33425
rect 184 33391 196 33425
rect -196 33385 196 33391
rect -196 33317 196 33323
rect -196 33283 -184 33317
rect 184 33283 196 33317
rect -196 33277 196 33283
rect -252 33224 -206 33236
rect -252 33048 -246 33224
rect -212 33048 -206 33224
rect -252 33036 -206 33048
rect 206 33224 252 33236
rect 206 33048 212 33224
rect 246 33048 252 33224
rect 206 33036 252 33048
rect -196 32989 196 32995
rect -196 32955 -184 32989
rect 184 32955 196 32989
rect -196 32949 196 32955
rect -196 32881 196 32887
rect -196 32847 -184 32881
rect 184 32847 196 32881
rect -196 32841 196 32847
rect -252 32788 -206 32800
rect -252 32612 -246 32788
rect -212 32612 -206 32788
rect -252 32600 -206 32612
rect 206 32788 252 32800
rect 206 32612 212 32788
rect 246 32612 252 32788
rect 206 32600 252 32612
rect -196 32553 196 32559
rect -196 32519 -184 32553
rect 184 32519 196 32553
rect -196 32513 196 32519
rect -196 32445 196 32451
rect -196 32411 -184 32445
rect 184 32411 196 32445
rect -196 32405 196 32411
rect -252 32352 -206 32364
rect -252 32176 -246 32352
rect -212 32176 -206 32352
rect -252 32164 -206 32176
rect 206 32352 252 32364
rect 206 32176 212 32352
rect 246 32176 252 32352
rect 206 32164 252 32176
rect -196 32117 196 32123
rect -196 32083 -184 32117
rect 184 32083 196 32117
rect -196 32077 196 32083
rect -196 32009 196 32015
rect -196 31975 -184 32009
rect 184 31975 196 32009
rect -196 31969 196 31975
rect -252 31916 -206 31928
rect -252 31740 -246 31916
rect -212 31740 -206 31916
rect -252 31728 -206 31740
rect 206 31916 252 31928
rect 206 31740 212 31916
rect 246 31740 252 31916
rect 206 31728 252 31740
rect -196 31681 196 31687
rect -196 31647 -184 31681
rect 184 31647 196 31681
rect -196 31641 196 31647
rect -196 31573 196 31579
rect -196 31539 -184 31573
rect 184 31539 196 31573
rect -196 31533 196 31539
rect -252 31480 -206 31492
rect -252 31304 -246 31480
rect -212 31304 -206 31480
rect -252 31292 -206 31304
rect 206 31480 252 31492
rect 206 31304 212 31480
rect 246 31304 252 31480
rect 206 31292 252 31304
rect -196 31245 196 31251
rect -196 31211 -184 31245
rect 184 31211 196 31245
rect -196 31205 196 31211
rect -196 31137 196 31143
rect -196 31103 -184 31137
rect 184 31103 196 31137
rect -196 31097 196 31103
rect -252 31044 -206 31056
rect -252 30868 -246 31044
rect -212 30868 -206 31044
rect -252 30856 -206 30868
rect 206 31044 252 31056
rect 206 30868 212 31044
rect 246 30868 252 31044
rect 206 30856 252 30868
rect -196 30809 196 30815
rect -196 30775 -184 30809
rect 184 30775 196 30809
rect -196 30769 196 30775
rect -196 30701 196 30707
rect -196 30667 -184 30701
rect 184 30667 196 30701
rect -196 30661 196 30667
rect -252 30608 -206 30620
rect -252 30432 -246 30608
rect -212 30432 -206 30608
rect -252 30420 -206 30432
rect 206 30608 252 30620
rect 206 30432 212 30608
rect 246 30432 252 30608
rect 206 30420 252 30432
rect -196 30373 196 30379
rect -196 30339 -184 30373
rect 184 30339 196 30373
rect -196 30333 196 30339
rect -196 30265 196 30271
rect -196 30231 -184 30265
rect 184 30231 196 30265
rect -196 30225 196 30231
rect -252 30172 -206 30184
rect -252 29996 -246 30172
rect -212 29996 -206 30172
rect -252 29984 -206 29996
rect 206 30172 252 30184
rect 206 29996 212 30172
rect 246 29996 252 30172
rect 206 29984 252 29996
rect -196 29937 196 29943
rect -196 29903 -184 29937
rect 184 29903 196 29937
rect -196 29897 196 29903
rect -196 29829 196 29835
rect -196 29795 -184 29829
rect 184 29795 196 29829
rect -196 29789 196 29795
rect -252 29736 -206 29748
rect -252 29560 -246 29736
rect -212 29560 -206 29736
rect -252 29548 -206 29560
rect 206 29736 252 29748
rect 206 29560 212 29736
rect 246 29560 252 29736
rect 206 29548 252 29560
rect -196 29501 196 29507
rect -196 29467 -184 29501
rect 184 29467 196 29501
rect -196 29461 196 29467
rect -196 29393 196 29399
rect -196 29359 -184 29393
rect 184 29359 196 29393
rect -196 29353 196 29359
rect -252 29300 -206 29312
rect -252 29124 -246 29300
rect -212 29124 -206 29300
rect -252 29112 -206 29124
rect 206 29300 252 29312
rect 206 29124 212 29300
rect 246 29124 252 29300
rect 206 29112 252 29124
rect -196 29065 196 29071
rect -196 29031 -184 29065
rect 184 29031 196 29065
rect -196 29025 196 29031
rect -196 28957 196 28963
rect -196 28923 -184 28957
rect 184 28923 196 28957
rect -196 28917 196 28923
rect -252 28864 -206 28876
rect -252 28688 -246 28864
rect -212 28688 -206 28864
rect -252 28676 -206 28688
rect 206 28864 252 28876
rect 206 28688 212 28864
rect 246 28688 252 28864
rect 206 28676 252 28688
rect -196 28629 196 28635
rect -196 28595 -184 28629
rect 184 28595 196 28629
rect -196 28589 196 28595
rect -196 28521 196 28527
rect -196 28487 -184 28521
rect 184 28487 196 28521
rect -196 28481 196 28487
rect -252 28428 -206 28440
rect -252 28252 -246 28428
rect -212 28252 -206 28428
rect -252 28240 -206 28252
rect 206 28428 252 28440
rect 206 28252 212 28428
rect 246 28252 252 28428
rect 206 28240 252 28252
rect -196 28193 196 28199
rect -196 28159 -184 28193
rect 184 28159 196 28193
rect -196 28153 196 28159
rect -196 28085 196 28091
rect -196 28051 -184 28085
rect 184 28051 196 28085
rect -196 28045 196 28051
rect -252 27992 -206 28004
rect -252 27816 -246 27992
rect -212 27816 -206 27992
rect -252 27804 -206 27816
rect 206 27992 252 28004
rect 206 27816 212 27992
rect 246 27816 252 27992
rect 206 27804 252 27816
rect -196 27757 196 27763
rect -196 27723 -184 27757
rect 184 27723 196 27757
rect -196 27717 196 27723
rect -196 27649 196 27655
rect -196 27615 -184 27649
rect 184 27615 196 27649
rect -196 27609 196 27615
rect -252 27556 -206 27568
rect -252 27380 -246 27556
rect -212 27380 -206 27556
rect -252 27368 -206 27380
rect 206 27556 252 27568
rect 206 27380 212 27556
rect 246 27380 252 27556
rect 206 27368 252 27380
rect -196 27321 196 27327
rect -196 27287 -184 27321
rect 184 27287 196 27321
rect -196 27281 196 27287
rect -196 27213 196 27219
rect -196 27179 -184 27213
rect 184 27179 196 27213
rect -196 27173 196 27179
rect -252 27120 -206 27132
rect -252 26944 -246 27120
rect -212 26944 -206 27120
rect -252 26932 -206 26944
rect 206 27120 252 27132
rect 206 26944 212 27120
rect 246 26944 252 27120
rect 206 26932 252 26944
rect -196 26885 196 26891
rect -196 26851 -184 26885
rect 184 26851 196 26885
rect -196 26845 196 26851
rect -196 26777 196 26783
rect -196 26743 -184 26777
rect 184 26743 196 26777
rect -196 26737 196 26743
rect -252 26684 -206 26696
rect -252 26508 -246 26684
rect -212 26508 -206 26684
rect -252 26496 -206 26508
rect 206 26684 252 26696
rect 206 26508 212 26684
rect 246 26508 252 26684
rect 206 26496 252 26508
rect -196 26449 196 26455
rect -196 26415 -184 26449
rect 184 26415 196 26449
rect -196 26409 196 26415
rect -196 26341 196 26347
rect -196 26307 -184 26341
rect 184 26307 196 26341
rect -196 26301 196 26307
rect -252 26248 -206 26260
rect -252 26072 -246 26248
rect -212 26072 -206 26248
rect -252 26060 -206 26072
rect 206 26248 252 26260
rect 206 26072 212 26248
rect 246 26072 252 26248
rect 206 26060 252 26072
rect -196 26013 196 26019
rect -196 25979 -184 26013
rect 184 25979 196 26013
rect -196 25973 196 25979
rect -196 25905 196 25911
rect -196 25871 -184 25905
rect 184 25871 196 25905
rect -196 25865 196 25871
rect -252 25812 -206 25824
rect -252 25636 -246 25812
rect -212 25636 -206 25812
rect -252 25624 -206 25636
rect 206 25812 252 25824
rect 206 25636 212 25812
rect 246 25636 252 25812
rect 206 25624 252 25636
rect -196 25577 196 25583
rect -196 25543 -184 25577
rect 184 25543 196 25577
rect -196 25537 196 25543
rect -196 25469 196 25475
rect -196 25435 -184 25469
rect 184 25435 196 25469
rect -196 25429 196 25435
rect -252 25376 -206 25388
rect -252 25200 -246 25376
rect -212 25200 -206 25376
rect -252 25188 -206 25200
rect 206 25376 252 25388
rect 206 25200 212 25376
rect 246 25200 252 25376
rect 206 25188 252 25200
rect -196 25141 196 25147
rect -196 25107 -184 25141
rect 184 25107 196 25141
rect -196 25101 196 25107
rect -196 25033 196 25039
rect -196 24999 -184 25033
rect 184 24999 196 25033
rect -196 24993 196 24999
rect -252 24940 -206 24952
rect -252 24764 -246 24940
rect -212 24764 -206 24940
rect -252 24752 -206 24764
rect 206 24940 252 24952
rect 206 24764 212 24940
rect 246 24764 252 24940
rect 206 24752 252 24764
rect -196 24705 196 24711
rect -196 24671 -184 24705
rect 184 24671 196 24705
rect -196 24665 196 24671
rect -196 24597 196 24603
rect -196 24563 -184 24597
rect 184 24563 196 24597
rect -196 24557 196 24563
rect -252 24504 -206 24516
rect -252 24328 -246 24504
rect -212 24328 -206 24504
rect -252 24316 -206 24328
rect 206 24504 252 24516
rect 206 24328 212 24504
rect 246 24328 252 24504
rect 206 24316 252 24328
rect -196 24269 196 24275
rect -196 24235 -184 24269
rect 184 24235 196 24269
rect -196 24229 196 24235
rect -196 24161 196 24167
rect -196 24127 -184 24161
rect 184 24127 196 24161
rect -196 24121 196 24127
rect -252 24068 -206 24080
rect -252 23892 -246 24068
rect -212 23892 -206 24068
rect -252 23880 -206 23892
rect 206 24068 252 24080
rect 206 23892 212 24068
rect 246 23892 252 24068
rect 206 23880 252 23892
rect -196 23833 196 23839
rect -196 23799 -184 23833
rect 184 23799 196 23833
rect -196 23793 196 23799
rect -196 23725 196 23731
rect -196 23691 -184 23725
rect 184 23691 196 23725
rect -196 23685 196 23691
rect -252 23632 -206 23644
rect -252 23456 -246 23632
rect -212 23456 -206 23632
rect -252 23444 -206 23456
rect 206 23632 252 23644
rect 206 23456 212 23632
rect 246 23456 252 23632
rect 206 23444 252 23456
rect -196 23397 196 23403
rect -196 23363 -184 23397
rect 184 23363 196 23397
rect -196 23357 196 23363
rect -196 23289 196 23295
rect -196 23255 -184 23289
rect 184 23255 196 23289
rect -196 23249 196 23255
rect -252 23196 -206 23208
rect -252 23020 -246 23196
rect -212 23020 -206 23196
rect -252 23008 -206 23020
rect 206 23196 252 23208
rect 206 23020 212 23196
rect 246 23020 252 23196
rect 206 23008 252 23020
rect -196 22961 196 22967
rect -196 22927 -184 22961
rect 184 22927 196 22961
rect -196 22921 196 22927
rect -196 22853 196 22859
rect -196 22819 -184 22853
rect 184 22819 196 22853
rect -196 22813 196 22819
rect -252 22760 -206 22772
rect -252 22584 -246 22760
rect -212 22584 -206 22760
rect -252 22572 -206 22584
rect 206 22760 252 22772
rect 206 22584 212 22760
rect 246 22584 252 22760
rect 206 22572 252 22584
rect -196 22525 196 22531
rect -196 22491 -184 22525
rect 184 22491 196 22525
rect -196 22485 196 22491
rect -196 22417 196 22423
rect -196 22383 -184 22417
rect 184 22383 196 22417
rect -196 22377 196 22383
rect -252 22324 -206 22336
rect -252 22148 -246 22324
rect -212 22148 -206 22324
rect -252 22136 -206 22148
rect 206 22324 252 22336
rect 206 22148 212 22324
rect 246 22148 252 22324
rect 206 22136 252 22148
rect -196 22089 196 22095
rect -196 22055 -184 22089
rect 184 22055 196 22089
rect -196 22049 196 22055
rect -196 21981 196 21987
rect -196 21947 -184 21981
rect 184 21947 196 21981
rect -196 21941 196 21947
rect -252 21888 -206 21900
rect -252 21712 -246 21888
rect -212 21712 -206 21888
rect -252 21700 -206 21712
rect 206 21888 252 21900
rect 206 21712 212 21888
rect 246 21712 252 21888
rect 206 21700 252 21712
rect -196 21653 196 21659
rect -196 21619 -184 21653
rect 184 21619 196 21653
rect -196 21613 196 21619
rect -196 21545 196 21551
rect -196 21511 -184 21545
rect 184 21511 196 21545
rect -196 21505 196 21511
rect -252 21452 -206 21464
rect -252 21276 -246 21452
rect -212 21276 -206 21452
rect -252 21264 -206 21276
rect 206 21452 252 21464
rect 206 21276 212 21452
rect 246 21276 252 21452
rect 206 21264 252 21276
rect -196 21217 196 21223
rect -196 21183 -184 21217
rect 184 21183 196 21217
rect -196 21177 196 21183
rect -196 21109 196 21115
rect -196 21075 -184 21109
rect 184 21075 196 21109
rect -196 21069 196 21075
rect -252 21016 -206 21028
rect -252 20840 -246 21016
rect -212 20840 -206 21016
rect -252 20828 -206 20840
rect 206 21016 252 21028
rect 206 20840 212 21016
rect 246 20840 252 21016
rect 206 20828 252 20840
rect -196 20781 196 20787
rect -196 20747 -184 20781
rect 184 20747 196 20781
rect -196 20741 196 20747
rect -196 20673 196 20679
rect -196 20639 -184 20673
rect 184 20639 196 20673
rect -196 20633 196 20639
rect -252 20580 -206 20592
rect -252 20404 -246 20580
rect -212 20404 -206 20580
rect -252 20392 -206 20404
rect 206 20580 252 20592
rect 206 20404 212 20580
rect 246 20404 252 20580
rect 206 20392 252 20404
rect -196 20345 196 20351
rect -196 20311 -184 20345
rect 184 20311 196 20345
rect -196 20305 196 20311
rect -196 20237 196 20243
rect -196 20203 -184 20237
rect 184 20203 196 20237
rect -196 20197 196 20203
rect -252 20144 -206 20156
rect -252 19968 -246 20144
rect -212 19968 -206 20144
rect -252 19956 -206 19968
rect 206 20144 252 20156
rect 206 19968 212 20144
rect 246 19968 252 20144
rect 206 19956 252 19968
rect -196 19909 196 19915
rect -196 19875 -184 19909
rect 184 19875 196 19909
rect -196 19869 196 19875
rect -196 19801 196 19807
rect -196 19767 -184 19801
rect 184 19767 196 19801
rect -196 19761 196 19767
rect -252 19708 -206 19720
rect -252 19532 -246 19708
rect -212 19532 -206 19708
rect -252 19520 -206 19532
rect 206 19708 252 19720
rect 206 19532 212 19708
rect 246 19532 252 19708
rect 206 19520 252 19532
rect -196 19473 196 19479
rect -196 19439 -184 19473
rect 184 19439 196 19473
rect -196 19433 196 19439
rect -196 19365 196 19371
rect -196 19331 -184 19365
rect 184 19331 196 19365
rect -196 19325 196 19331
rect -252 19272 -206 19284
rect -252 19096 -246 19272
rect -212 19096 -206 19272
rect -252 19084 -206 19096
rect 206 19272 252 19284
rect 206 19096 212 19272
rect 246 19096 252 19272
rect 206 19084 252 19096
rect -196 19037 196 19043
rect -196 19003 -184 19037
rect 184 19003 196 19037
rect -196 18997 196 19003
rect -196 18929 196 18935
rect -196 18895 -184 18929
rect 184 18895 196 18929
rect -196 18889 196 18895
rect -252 18836 -206 18848
rect -252 18660 -246 18836
rect -212 18660 -206 18836
rect -252 18648 -206 18660
rect 206 18836 252 18848
rect 206 18660 212 18836
rect 246 18660 252 18836
rect 206 18648 252 18660
rect -196 18601 196 18607
rect -196 18567 -184 18601
rect 184 18567 196 18601
rect -196 18561 196 18567
rect -196 18493 196 18499
rect -196 18459 -184 18493
rect 184 18459 196 18493
rect -196 18453 196 18459
rect -252 18400 -206 18412
rect -252 18224 -246 18400
rect -212 18224 -206 18400
rect -252 18212 -206 18224
rect 206 18400 252 18412
rect 206 18224 212 18400
rect 246 18224 252 18400
rect 206 18212 252 18224
rect -196 18165 196 18171
rect -196 18131 -184 18165
rect 184 18131 196 18165
rect -196 18125 196 18131
rect -196 18057 196 18063
rect -196 18023 -184 18057
rect 184 18023 196 18057
rect -196 18017 196 18023
rect -252 17964 -206 17976
rect -252 17788 -246 17964
rect -212 17788 -206 17964
rect -252 17776 -206 17788
rect 206 17964 252 17976
rect 206 17788 212 17964
rect 246 17788 252 17964
rect 206 17776 252 17788
rect -196 17729 196 17735
rect -196 17695 -184 17729
rect 184 17695 196 17729
rect -196 17689 196 17695
rect -196 17621 196 17627
rect -196 17587 -184 17621
rect 184 17587 196 17621
rect -196 17581 196 17587
rect -252 17528 -206 17540
rect -252 17352 -246 17528
rect -212 17352 -206 17528
rect -252 17340 -206 17352
rect 206 17528 252 17540
rect 206 17352 212 17528
rect 246 17352 252 17528
rect 206 17340 252 17352
rect -196 17293 196 17299
rect -196 17259 -184 17293
rect 184 17259 196 17293
rect -196 17253 196 17259
rect -196 17185 196 17191
rect -196 17151 -184 17185
rect 184 17151 196 17185
rect -196 17145 196 17151
rect -252 17092 -206 17104
rect -252 16916 -246 17092
rect -212 16916 -206 17092
rect -252 16904 -206 16916
rect 206 17092 252 17104
rect 206 16916 212 17092
rect 246 16916 252 17092
rect 206 16904 252 16916
rect -196 16857 196 16863
rect -196 16823 -184 16857
rect 184 16823 196 16857
rect -196 16817 196 16823
rect -196 16749 196 16755
rect -196 16715 -184 16749
rect 184 16715 196 16749
rect -196 16709 196 16715
rect -252 16656 -206 16668
rect -252 16480 -246 16656
rect -212 16480 -206 16656
rect -252 16468 -206 16480
rect 206 16656 252 16668
rect 206 16480 212 16656
rect 246 16480 252 16656
rect 206 16468 252 16480
rect -196 16421 196 16427
rect -196 16387 -184 16421
rect 184 16387 196 16421
rect -196 16381 196 16387
rect -196 16313 196 16319
rect -196 16279 -184 16313
rect 184 16279 196 16313
rect -196 16273 196 16279
rect -252 16220 -206 16232
rect -252 16044 -246 16220
rect -212 16044 -206 16220
rect -252 16032 -206 16044
rect 206 16220 252 16232
rect 206 16044 212 16220
rect 246 16044 252 16220
rect 206 16032 252 16044
rect -196 15985 196 15991
rect -196 15951 -184 15985
rect 184 15951 196 15985
rect -196 15945 196 15951
rect -196 15877 196 15883
rect -196 15843 -184 15877
rect 184 15843 196 15877
rect -196 15837 196 15843
rect -252 15784 -206 15796
rect -252 15608 -246 15784
rect -212 15608 -206 15784
rect -252 15596 -206 15608
rect 206 15784 252 15796
rect 206 15608 212 15784
rect 246 15608 252 15784
rect 206 15596 252 15608
rect -196 15549 196 15555
rect -196 15515 -184 15549
rect 184 15515 196 15549
rect -196 15509 196 15515
rect -196 15441 196 15447
rect -196 15407 -184 15441
rect 184 15407 196 15441
rect -196 15401 196 15407
rect -252 15348 -206 15360
rect -252 15172 -246 15348
rect -212 15172 -206 15348
rect -252 15160 -206 15172
rect 206 15348 252 15360
rect 206 15172 212 15348
rect 246 15172 252 15348
rect 206 15160 252 15172
rect -196 15113 196 15119
rect -196 15079 -184 15113
rect 184 15079 196 15113
rect -196 15073 196 15079
rect -196 15005 196 15011
rect -196 14971 -184 15005
rect 184 14971 196 15005
rect -196 14965 196 14971
rect -252 14912 -206 14924
rect -252 14736 -246 14912
rect -212 14736 -206 14912
rect -252 14724 -206 14736
rect 206 14912 252 14924
rect 206 14736 212 14912
rect 246 14736 252 14912
rect 206 14724 252 14736
rect -196 14677 196 14683
rect -196 14643 -184 14677
rect 184 14643 196 14677
rect -196 14637 196 14643
rect -196 14569 196 14575
rect -196 14535 -184 14569
rect 184 14535 196 14569
rect -196 14529 196 14535
rect -252 14476 -206 14488
rect -252 14300 -246 14476
rect -212 14300 -206 14476
rect -252 14288 -206 14300
rect 206 14476 252 14488
rect 206 14300 212 14476
rect 246 14300 252 14476
rect 206 14288 252 14300
rect -196 14241 196 14247
rect -196 14207 -184 14241
rect 184 14207 196 14241
rect -196 14201 196 14207
rect -196 14133 196 14139
rect -196 14099 -184 14133
rect 184 14099 196 14133
rect -196 14093 196 14099
rect -252 14040 -206 14052
rect -252 13864 -246 14040
rect -212 13864 -206 14040
rect -252 13852 -206 13864
rect 206 14040 252 14052
rect 206 13864 212 14040
rect 246 13864 252 14040
rect 206 13852 252 13864
rect -196 13805 196 13811
rect -196 13771 -184 13805
rect 184 13771 196 13805
rect -196 13765 196 13771
rect -196 13697 196 13703
rect -196 13663 -184 13697
rect 184 13663 196 13697
rect -196 13657 196 13663
rect -252 13604 -206 13616
rect -252 13428 -246 13604
rect -212 13428 -206 13604
rect -252 13416 -206 13428
rect 206 13604 252 13616
rect 206 13428 212 13604
rect 246 13428 252 13604
rect 206 13416 252 13428
rect -196 13369 196 13375
rect -196 13335 -184 13369
rect 184 13335 196 13369
rect -196 13329 196 13335
rect -196 13261 196 13267
rect -196 13227 -184 13261
rect 184 13227 196 13261
rect -196 13221 196 13227
rect -252 13168 -206 13180
rect -252 12992 -246 13168
rect -212 12992 -206 13168
rect -252 12980 -206 12992
rect 206 13168 252 13180
rect 206 12992 212 13168
rect 246 12992 252 13168
rect 206 12980 252 12992
rect -196 12933 196 12939
rect -196 12899 -184 12933
rect 184 12899 196 12933
rect -196 12893 196 12899
rect -196 12825 196 12831
rect -196 12791 -184 12825
rect 184 12791 196 12825
rect -196 12785 196 12791
rect -252 12732 -206 12744
rect -252 12556 -246 12732
rect -212 12556 -206 12732
rect -252 12544 -206 12556
rect 206 12732 252 12744
rect 206 12556 212 12732
rect 246 12556 252 12732
rect 206 12544 252 12556
rect -196 12497 196 12503
rect -196 12463 -184 12497
rect 184 12463 196 12497
rect -196 12457 196 12463
rect -196 12389 196 12395
rect -196 12355 -184 12389
rect 184 12355 196 12389
rect -196 12349 196 12355
rect -252 12296 -206 12308
rect -252 12120 -246 12296
rect -212 12120 -206 12296
rect -252 12108 -206 12120
rect 206 12296 252 12308
rect 206 12120 212 12296
rect 246 12120 252 12296
rect 206 12108 252 12120
rect -196 12061 196 12067
rect -196 12027 -184 12061
rect 184 12027 196 12061
rect -196 12021 196 12027
rect -196 11953 196 11959
rect -196 11919 -184 11953
rect 184 11919 196 11953
rect -196 11913 196 11919
rect -252 11860 -206 11872
rect -252 11684 -246 11860
rect -212 11684 -206 11860
rect -252 11672 -206 11684
rect 206 11860 252 11872
rect 206 11684 212 11860
rect 246 11684 252 11860
rect 206 11672 252 11684
rect -196 11625 196 11631
rect -196 11591 -184 11625
rect 184 11591 196 11625
rect -196 11585 196 11591
rect -196 11517 196 11523
rect -196 11483 -184 11517
rect 184 11483 196 11517
rect -196 11477 196 11483
rect -252 11424 -206 11436
rect -252 11248 -246 11424
rect -212 11248 -206 11424
rect -252 11236 -206 11248
rect 206 11424 252 11436
rect 206 11248 212 11424
rect 246 11248 252 11424
rect 206 11236 252 11248
rect -196 11189 196 11195
rect -196 11155 -184 11189
rect 184 11155 196 11189
rect -196 11149 196 11155
rect -196 11081 196 11087
rect -196 11047 -184 11081
rect 184 11047 196 11081
rect -196 11041 196 11047
rect -252 10988 -206 11000
rect -252 10812 -246 10988
rect -212 10812 -206 10988
rect -252 10800 -206 10812
rect 206 10988 252 11000
rect 206 10812 212 10988
rect 246 10812 252 10988
rect 206 10800 252 10812
rect -196 10753 196 10759
rect -196 10719 -184 10753
rect 184 10719 196 10753
rect -196 10713 196 10719
rect -196 10645 196 10651
rect -196 10611 -184 10645
rect 184 10611 196 10645
rect -196 10605 196 10611
rect -252 10552 -206 10564
rect -252 10376 -246 10552
rect -212 10376 -206 10552
rect -252 10364 -206 10376
rect 206 10552 252 10564
rect 206 10376 212 10552
rect 246 10376 252 10552
rect 206 10364 252 10376
rect -196 10317 196 10323
rect -196 10283 -184 10317
rect 184 10283 196 10317
rect -196 10277 196 10283
rect -196 10209 196 10215
rect -196 10175 -184 10209
rect 184 10175 196 10209
rect -196 10169 196 10175
rect -252 10116 -206 10128
rect -252 9940 -246 10116
rect -212 9940 -206 10116
rect -252 9928 -206 9940
rect 206 10116 252 10128
rect 206 9940 212 10116
rect 246 9940 252 10116
rect 206 9928 252 9940
rect -196 9881 196 9887
rect -196 9847 -184 9881
rect 184 9847 196 9881
rect -196 9841 196 9847
rect -196 9773 196 9779
rect -196 9739 -184 9773
rect 184 9739 196 9773
rect -196 9733 196 9739
rect -252 9680 -206 9692
rect -252 9504 -246 9680
rect -212 9504 -206 9680
rect -252 9492 -206 9504
rect 206 9680 252 9692
rect 206 9504 212 9680
rect 246 9504 252 9680
rect 206 9492 252 9504
rect -196 9445 196 9451
rect -196 9411 -184 9445
rect 184 9411 196 9445
rect -196 9405 196 9411
rect -196 9337 196 9343
rect -196 9303 -184 9337
rect 184 9303 196 9337
rect -196 9297 196 9303
rect -252 9244 -206 9256
rect -252 9068 -246 9244
rect -212 9068 -206 9244
rect -252 9056 -206 9068
rect 206 9244 252 9256
rect 206 9068 212 9244
rect 246 9068 252 9244
rect 206 9056 252 9068
rect -196 9009 196 9015
rect -196 8975 -184 9009
rect 184 8975 196 9009
rect -196 8969 196 8975
rect -196 8901 196 8907
rect -196 8867 -184 8901
rect 184 8867 196 8901
rect -196 8861 196 8867
rect -252 8808 -206 8820
rect -252 8632 -246 8808
rect -212 8632 -206 8808
rect -252 8620 -206 8632
rect 206 8808 252 8820
rect 206 8632 212 8808
rect 246 8632 252 8808
rect 206 8620 252 8632
rect -196 8573 196 8579
rect -196 8539 -184 8573
rect 184 8539 196 8573
rect -196 8533 196 8539
rect -196 8465 196 8471
rect -196 8431 -184 8465
rect 184 8431 196 8465
rect -196 8425 196 8431
rect -252 8372 -206 8384
rect -252 8196 -246 8372
rect -212 8196 -206 8372
rect -252 8184 -206 8196
rect 206 8372 252 8384
rect 206 8196 212 8372
rect 246 8196 252 8372
rect 206 8184 252 8196
rect -196 8137 196 8143
rect -196 8103 -184 8137
rect 184 8103 196 8137
rect -196 8097 196 8103
rect -196 8029 196 8035
rect -196 7995 -184 8029
rect 184 7995 196 8029
rect -196 7989 196 7995
rect -252 7936 -206 7948
rect -252 7760 -246 7936
rect -212 7760 -206 7936
rect -252 7748 -206 7760
rect 206 7936 252 7948
rect 206 7760 212 7936
rect 246 7760 252 7936
rect 206 7748 252 7760
rect -196 7701 196 7707
rect -196 7667 -184 7701
rect 184 7667 196 7701
rect -196 7661 196 7667
rect -196 7593 196 7599
rect -196 7559 -184 7593
rect 184 7559 196 7593
rect -196 7553 196 7559
rect -252 7500 -206 7512
rect -252 7324 -246 7500
rect -212 7324 -206 7500
rect -252 7312 -206 7324
rect 206 7500 252 7512
rect 206 7324 212 7500
rect 246 7324 252 7500
rect 206 7312 252 7324
rect -196 7265 196 7271
rect -196 7231 -184 7265
rect 184 7231 196 7265
rect -196 7225 196 7231
rect -196 7157 196 7163
rect -196 7123 -184 7157
rect 184 7123 196 7157
rect -196 7117 196 7123
rect -252 7064 -206 7076
rect -252 6888 -246 7064
rect -212 6888 -206 7064
rect -252 6876 -206 6888
rect 206 7064 252 7076
rect 206 6888 212 7064
rect 246 6888 252 7064
rect 206 6876 252 6888
rect -196 6829 196 6835
rect -196 6795 -184 6829
rect 184 6795 196 6829
rect -196 6789 196 6795
rect -196 6721 196 6727
rect -196 6687 -184 6721
rect 184 6687 196 6721
rect -196 6681 196 6687
rect -252 6628 -206 6640
rect -252 6452 -246 6628
rect -212 6452 -206 6628
rect -252 6440 -206 6452
rect 206 6628 252 6640
rect 206 6452 212 6628
rect 246 6452 252 6628
rect 206 6440 252 6452
rect -196 6393 196 6399
rect -196 6359 -184 6393
rect 184 6359 196 6393
rect -196 6353 196 6359
rect -196 6285 196 6291
rect -196 6251 -184 6285
rect 184 6251 196 6285
rect -196 6245 196 6251
rect -252 6192 -206 6204
rect -252 6016 -246 6192
rect -212 6016 -206 6192
rect -252 6004 -206 6016
rect 206 6192 252 6204
rect 206 6016 212 6192
rect 246 6016 252 6192
rect 206 6004 252 6016
rect -196 5957 196 5963
rect -196 5923 -184 5957
rect 184 5923 196 5957
rect -196 5917 196 5923
rect -196 5849 196 5855
rect -196 5815 -184 5849
rect 184 5815 196 5849
rect -196 5809 196 5815
rect -252 5756 -206 5768
rect -252 5580 -246 5756
rect -212 5580 -206 5756
rect -252 5568 -206 5580
rect 206 5756 252 5768
rect 206 5580 212 5756
rect 246 5580 252 5756
rect 206 5568 252 5580
rect -196 5521 196 5527
rect -196 5487 -184 5521
rect 184 5487 196 5521
rect -196 5481 196 5487
rect -196 5413 196 5419
rect -196 5379 -184 5413
rect 184 5379 196 5413
rect -196 5373 196 5379
rect -252 5320 -206 5332
rect -252 5144 -246 5320
rect -212 5144 -206 5320
rect -252 5132 -206 5144
rect 206 5320 252 5332
rect 206 5144 212 5320
rect 246 5144 252 5320
rect 206 5132 252 5144
rect -196 5085 196 5091
rect -196 5051 -184 5085
rect 184 5051 196 5085
rect -196 5045 196 5051
rect -196 4977 196 4983
rect -196 4943 -184 4977
rect 184 4943 196 4977
rect -196 4937 196 4943
rect -252 4884 -206 4896
rect -252 4708 -246 4884
rect -212 4708 -206 4884
rect -252 4696 -206 4708
rect 206 4884 252 4896
rect 206 4708 212 4884
rect 246 4708 252 4884
rect 206 4696 252 4708
rect -196 4649 196 4655
rect -196 4615 -184 4649
rect 184 4615 196 4649
rect -196 4609 196 4615
rect -196 4541 196 4547
rect -196 4507 -184 4541
rect 184 4507 196 4541
rect -196 4501 196 4507
rect -252 4448 -206 4460
rect -252 4272 -246 4448
rect -212 4272 -206 4448
rect -252 4260 -206 4272
rect 206 4448 252 4460
rect 206 4272 212 4448
rect 246 4272 252 4448
rect 206 4260 252 4272
rect -196 4213 196 4219
rect -196 4179 -184 4213
rect 184 4179 196 4213
rect -196 4173 196 4179
rect -196 4105 196 4111
rect -196 4071 -184 4105
rect 184 4071 196 4105
rect -196 4065 196 4071
rect -252 4012 -206 4024
rect -252 3836 -246 4012
rect -212 3836 -206 4012
rect -252 3824 -206 3836
rect 206 4012 252 4024
rect 206 3836 212 4012
rect 246 3836 252 4012
rect 206 3824 252 3836
rect -196 3777 196 3783
rect -196 3743 -184 3777
rect 184 3743 196 3777
rect -196 3737 196 3743
rect -196 3669 196 3675
rect -196 3635 -184 3669
rect 184 3635 196 3669
rect -196 3629 196 3635
rect -252 3576 -206 3588
rect -252 3400 -246 3576
rect -212 3400 -206 3576
rect -252 3388 -206 3400
rect 206 3576 252 3588
rect 206 3400 212 3576
rect 246 3400 252 3576
rect 206 3388 252 3400
rect -196 3341 196 3347
rect -196 3307 -184 3341
rect 184 3307 196 3341
rect -196 3301 196 3307
rect -196 3233 196 3239
rect -196 3199 -184 3233
rect 184 3199 196 3233
rect -196 3193 196 3199
rect -252 3140 -206 3152
rect -252 2964 -246 3140
rect -212 2964 -206 3140
rect -252 2952 -206 2964
rect 206 3140 252 3152
rect 206 2964 212 3140
rect 246 2964 252 3140
rect 206 2952 252 2964
rect -196 2905 196 2911
rect -196 2871 -184 2905
rect 184 2871 196 2905
rect -196 2865 196 2871
rect -196 2797 196 2803
rect -196 2763 -184 2797
rect 184 2763 196 2797
rect -196 2757 196 2763
rect -252 2704 -206 2716
rect -252 2528 -246 2704
rect -212 2528 -206 2704
rect -252 2516 -206 2528
rect 206 2704 252 2716
rect 206 2528 212 2704
rect 246 2528 252 2704
rect 206 2516 252 2528
rect -196 2469 196 2475
rect -196 2435 -184 2469
rect 184 2435 196 2469
rect -196 2429 196 2435
rect -196 2361 196 2367
rect -196 2327 -184 2361
rect 184 2327 196 2361
rect -196 2321 196 2327
rect -252 2268 -206 2280
rect -252 2092 -246 2268
rect -212 2092 -206 2268
rect -252 2080 -206 2092
rect 206 2268 252 2280
rect 206 2092 212 2268
rect 246 2092 252 2268
rect 206 2080 252 2092
rect -196 2033 196 2039
rect -196 1999 -184 2033
rect 184 1999 196 2033
rect -196 1993 196 1999
rect -196 1925 196 1931
rect -196 1891 -184 1925
rect 184 1891 196 1925
rect -196 1885 196 1891
rect -252 1832 -206 1844
rect -252 1656 -246 1832
rect -212 1656 -206 1832
rect -252 1644 -206 1656
rect 206 1832 252 1844
rect 206 1656 212 1832
rect 246 1656 252 1832
rect 206 1644 252 1656
rect -196 1597 196 1603
rect -196 1563 -184 1597
rect 184 1563 196 1597
rect -196 1557 196 1563
rect -196 1489 196 1495
rect -196 1455 -184 1489
rect 184 1455 196 1489
rect -196 1449 196 1455
rect -252 1396 -206 1408
rect -252 1220 -246 1396
rect -212 1220 -206 1396
rect -252 1208 -206 1220
rect 206 1396 252 1408
rect 206 1220 212 1396
rect 246 1220 252 1396
rect 206 1208 252 1220
rect -196 1161 196 1167
rect -196 1127 -184 1161
rect 184 1127 196 1161
rect -196 1121 196 1127
rect -196 1053 196 1059
rect -196 1019 -184 1053
rect 184 1019 196 1053
rect -196 1013 196 1019
rect -252 960 -206 972
rect -252 784 -246 960
rect -212 784 -206 960
rect -252 772 -206 784
rect 206 960 252 972
rect 206 784 212 960
rect 246 784 252 960
rect 206 772 252 784
rect -196 725 196 731
rect -196 691 -184 725
rect 184 691 196 725
rect -196 685 196 691
rect -196 617 196 623
rect -196 583 -184 617
rect 184 583 196 617
rect -196 577 196 583
rect -252 524 -206 536
rect -252 348 -246 524
rect -212 348 -206 524
rect -252 336 -206 348
rect 206 524 252 536
rect 206 348 212 524
rect 246 348 252 524
rect 206 336 252 348
rect -196 289 196 295
rect -196 255 -184 289
rect 184 255 196 289
rect -196 249 196 255
rect -196 181 196 187
rect -196 147 -184 181
rect 184 147 196 181
rect -196 141 196 147
rect -252 88 -206 100
rect -252 -88 -246 88
rect -212 -88 -206 88
rect -252 -100 -206 -88
rect 206 88 252 100
rect 206 -88 212 88
rect 246 -88 252 88
rect 206 -100 252 -88
rect -196 -147 196 -141
rect -196 -181 -184 -147
rect 184 -181 196 -147
rect -196 -187 196 -181
rect -196 -255 196 -249
rect -196 -289 -184 -255
rect 184 -289 196 -255
rect -196 -295 196 -289
rect -252 -348 -206 -336
rect -252 -524 -246 -348
rect -212 -524 -206 -348
rect -252 -536 -206 -524
rect 206 -348 252 -336
rect 206 -524 212 -348
rect 246 -524 252 -348
rect 206 -536 252 -524
rect -196 -583 196 -577
rect -196 -617 -184 -583
rect 184 -617 196 -583
rect -196 -623 196 -617
rect -196 -691 196 -685
rect -196 -725 -184 -691
rect 184 -725 196 -691
rect -196 -731 196 -725
rect -252 -784 -206 -772
rect -252 -960 -246 -784
rect -212 -960 -206 -784
rect -252 -972 -206 -960
rect 206 -784 252 -772
rect 206 -960 212 -784
rect 246 -960 252 -784
rect 206 -972 252 -960
rect -196 -1019 196 -1013
rect -196 -1053 -184 -1019
rect 184 -1053 196 -1019
rect -196 -1059 196 -1053
rect -196 -1127 196 -1121
rect -196 -1161 -184 -1127
rect 184 -1161 196 -1127
rect -196 -1167 196 -1161
rect -252 -1220 -206 -1208
rect -252 -1396 -246 -1220
rect -212 -1396 -206 -1220
rect -252 -1408 -206 -1396
rect 206 -1220 252 -1208
rect 206 -1396 212 -1220
rect 246 -1396 252 -1220
rect 206 -1408 252 -1396
rect -196 -1455 196 -1449
rect -196 -1489 -184 -1455
rect 184 -1489 196 -1455
rect -196 -1495 196 -1489
rect -196 -1563 196 -1557
rect -196 -1597 -184 -1563
rect 184 -1597 196 -1563
rect -196 -1603 196 -1597
rect -252 -1656 -206 -1644
rect -252 -1832 -246 -1656
rect -212 -1832 -206 -1656
rect -252 -1844 -206 -1832
rect 206 -1656 252 -1644
rect 206 -1832 212 -1656
rect 246 -1832 252 -1656
rect 206 -1844 252 -1832
rect -196 -1891 196 -1885
rect -196 -1925 -184 -1891
rect 184 -1925 196 -1891
rect -196 -1931 196 -1925
rect -196 -1999 196 -1993
rect -196 -2033 -184 -1999
rect 184 -2033 196 -1999
rect -196 -2039 196 -2033
rect -252 -2092 -206 -2080
rect -252 -2268 -246 -2092
rect -212 -2268 -206 -2092
rect -252 -2280 -206 -2268
rect 206 -2092 252 -2080
rect 206 -2268 212 -2092
rect 246 -2268 252 -2092
rect 206 -2280 252 -2268
rect -196 -2327 196 -2321
rect -196 -2361 -184 -2327
rect 184 -2361 196 -2327
rect -196 -2367 196 -2361
rect -196 -2435 196 -2429
rect -196 -2469 -184 -2435
rect 184 -2469 196 -2435
rect -196 -2475 196 -2469
rect -252 -2528 -206 -2516
rect -252 -2704 -246 -2528
rect -212 -2704 -206 -2528
rect -252 -2716 -206 -2704
rect 206 -2528 252 -2516
rect 206 -2704 212 -2528
rect 246 -2704 252 -2528
rect 206 -2716 252 -2704
rect -196 -2763 196 -2757
rect -196 -2797 -184 -2763
rect 184 -2797 196 -2763
rect -196 -2803 196 -2797
rect -196 -2871 196 -2865
rect -196 -2905 -184 -2871
rect 184 -2905 196 -2871
rect -196 -2911 196 -2905
rect -252 -2964 -206 -2952
rect -252 -3140 -246 -2964
rect -212 -3140 -206 -2964
rect -252 -3152 -206 -3140
rect 206 -2964 252 -2952
rect 206 -3140 212 -2964
rect 246 -3140 252 -2964
rect 206 -3152 252 -3140
rect -196 -3199 196 -3193
rect -196 -3233 -184 -3199
rect 184 -3233 196 -3199
rect -196 -3239 196 -3233
rect -196 -3307 196 -3301
rect -196 -3341 -184 -3307
rect 184 -3341 196 -3307
rect -196 -3347 196 -3341
rect -252 -3400 -206 -3388
rect -252 -3576 -246 -3400
rect -212 -3576 -206 -3400
rect -252 -3588 -206 -3576
rect 206 -3400 252 -3388
rect 206 -3576 212 -3400
rect 246 -3576 252 -3400
rect 206 -3588 252 -3576
rect -196 -3635 196 -3629
rect -196 -3669 -184 -3635
rect 184 -3669 196 -3635
rect -196 -3675 196 -3669
rect -196 -3743 196 -3737
rect -196 -3777 -184 -3743
rect 184 -3777 196 -3743
rect -196 -3783 196 -3777
rect -252 -3836 -206 -3824
rect -252 -4012 -246 -3836
rect -212 -4012 -206 -3836
rect -252 -4024 -206 -4012
rect 206 -3836 252 -3824
rect 206 -4012 212 -3836
rect 246 -4012 252 -3836
rect 206 -4024 252 -4012
rect -196 -4071 196 -4065
rect -196 -4105 -184 -4071
rect 184 -4105 196 -4071
rect -196 -4111 196 -4105
rect -196 -4179 196 -4173
rect -196 -4213 -184 -4179
rect 184 -4213 196 -4179
rect -196 -4219 196 -4213
rect -252 -4272 -206 -4260
rect -252 -4448 -246 -4272
rect -212 -4448 -206 -4272
rect -252 -4460 -206 -4448
rect 206 -4272 252 -4260
rect 206 -4448 212 -4272
rect 246 -4448 252 -4272
rect 206 -4460 252 -4448
rect -196 -4507 196 -4501
rect -196 -4541 -184 -4507
rect 184 -4541 196 -4507
rect -196 -4547 196 -4541
rect -196 -4615 196 -4609
rect -196 -4649 -184 -4615
rect 184 -4649 196 -4615
rect -196 -4655 196 -4649
rect -252 -4708 -206 -4696
rect -252 -4884 -246 -4708
rect -212 -4884 -206 -4708
rect -252 -4896 -206 -4884
rect 206 -4708 252 -4696
rect 206 -4884 212 -4708
rect 246 -4884 252 -4708
rect 206 -4896 252 -4884
rect -196 -4943 196 -4937
rect -196 -4977 -184 -4943
rect 184 -4977 196 -4943
rect -196 -4983 196 -4977
rect -196 -5051 196 -5045
rect -196 -5085 -184 -5051
rect 184 -5085 196 -5051
rect -196 -5091 196 -5085
rect -252 -5144 -206 -5132
rect -252 -5320 -246 -5144
rect -212 -5320 -206 -5144
rect -252 -5332 -206 -5320
rect 206 -5144 252 -5132
rect 206 -5320 212 -5144
rect 246 -5320 252 -5144
rect 206 -5332 252 -5320
rect -196 -5379 196 -5373
rect -196 -5413 -184 -5379
rect 184 -5413 196 -5379
rect -196 -5419 196 -5413
rect -196 -5487 196 -5481
rect -196 -5521 -184 -5487
rect 184 -5521 196 -5487
rect -196 -5527 196 -5521
rect -252 -5580 -206 -5568
rect -252 -5756 -246 -5580
rect -212 -5756 -206 -5580
rect -252 -5768 -206 -5756
rect 206 -5580 252 -5568
rect 206 -5756 212 -5580
rect 246 -5756 252 -5580
rect 206 -5768 252 -5756
rect -196 -5815 196 -5809
rect -196 -5849 -184 -5815
rect 184 -5849 196 -5815
rect -196 -5855 196 -5849
rect -196 -5923 196 -5917
rect -196 -5957 -184 -5923
rect 184 -5957 196 -5923
rect -196 -5963 196 -5957
rect -252 -6016 -206 -6004
rect -252 -6192 -246 -6016
rect -212 -6192 -206 -6016
rect -252 -6204 -206 -6192
rect 206 -6016 252 -6004
rect 206 -6192 212 -6016
rect 246 -6192 252 -6016
rect 206 -6204 252 -6192
rect -196 -6251 196 -6245
rect -196 -6285 -184 -6251
rect 184 -6285 196 -6251
rect -196 -6291 196 -6285
rect -196 -6359 196 -6353
rect -196 -6393 -184 -6359
rect 184 -6393 196 -6359
rect -196 -6399 196 -6393
rect -252 -6452 -206 -6440
rect -252 -6628 -246 -6452
rect -212 -6628 -206 -6452
rect -252 -6640 -206 -6628
rect 206 -6452 252 -6440
rect 206 -6628 212 -6452
rect 246 -6628 252 -6452
rect 206 -6640 252 -6628
rect -196 -6687 196 -6681
rect -196 -6721 -184 -6687
rect 184 -6721 196 -6687
rect -196 -6727 196 -6721
rect -196 -6795 196 -6789
rect -196 -6829 -184 -6795
rect 184 -6829 196 -6795
rect -196 -6835 196 -6829
rect -252 -6888 -206 -6876
rect -252 -7064 -246 -6888
rect -212 -7064 -206 -6888
rect -252 -7076 -206 -7064
rect 206 -6888 252 -6876
rect 206 -7064 212 -6888
rect 246 -7064 252 -6888
rect 206 -7076 252 -7064
rect -196 -7123 196 -7117
rect -196 -7157 -184 -7123
rect 184 -7157 196 -7123
rect -196 -7163 196 -7157
rect -196 -7231 196 -7225
rect -196 -7265 -184 -7231
rect 184 -7265 196 -7231
rect -196 -7271 196 -7265
rect -252 -7324 -206 -7312
rect -252 -7500 -246 -7324
rect -212 -7500 -206 -7324
rect -252 -7512 -206 -7500
rect 206 -7324 252 -7312
rect 206 -7500 212 -7324
rect 246 -7500 252 -7324
rect 206 -7512 252 -7500
rect -196 -7559 196 -7553
rect -196 -7593 -184 -7559
rect 184 -7593 196 -7559
rect -196 -7599 196 -7593
rect -196 -7667 196 -7661
rect -196 -7701 -184 -7667
rect 184 -7701 196 -7667
rect -196 -7707 196 -7701
rect -252 -7760 -206 -7748
rect -252 -7936 -246 -7760
rect -212 -7936 -206 -7760
rect -252 -7948 -206 -7936
rect 206 -7760 252 -7748
rect 206 -7936 212 -7760
rect 246 -7936 252 -7760
rect 206 -7948 252 -7936
rect -196 -7995 196 -7989
rect -196 -8029 -184 -7995
rect 184 -8029 196 -7995
rect -196 -8035 196 -8029
rect -196 -8103 196 -8097
rect -196 -8137 -184 -8103
rect 184 -8137 196 -8103
rect -196 -8143 196 -8137
rect -252 -8196 -206 -8184
rect -252 -8372 -246 -8196
rect -212 -8372 -206 -8196
rect -252 -8384 -206 -8372
rect 206 -8196 252 -8184
rect 206 -8372 212 -8196
rect 246 -8372 252 -8196
rect 206 -8384 252 -8372
rect -196 -8431 196 -8425
rect -196 -8465 -184 -8431
rect 184 -8465 196 -8431
rect -196 -8471 196 -8465
rect -196 -8539 196 -8533
rect -196 -8573 -184 -8539
rect 184 -8573 196 -8539
rect -196 -8579 196 -8573
rect -252 -8632 -206 -8620
rect -252 -8808 -246 -8632
rect -212 -8808 -206 -8632
rect -252 -8820 -206 -8808
rect 206 -8632 252 -8620
rect 206 -8808 212 -8632
rect 246 -8808 252 -8632
rect 206 -8820 252 -8808
rect -196 -8867 196 -8861
rect -196 -8901 -184 -8867
rect 184 -8901 196 -8867
rect -196 -8907 196 -8901
rect -196 -8975 196 -8969
rect -196 -9009 -184 -8975
rect 184 -9009 196 -8975
rect -196 -9015 196 -9009
rect -252 -9068 -206 -9056
rect -252 -9244 -246 -9068
rect -212 -9244 -206 -9068
rect -252 -9256 -206 -9244
rect 206 -9068 252 -9056
rect 206 -9244 212 -9068
rect 246 -9244 252 -9068
rect 206 -9256 252 -9244
rect -196 -9303 196 -9297
rect -196 -9337 -184 -9303
rect 184 -9337 196 -9303
rect -196 -9343 196 -9337
rect -196 -9411 196 -9405
rect -196 -9445 -184 -9411
rect 184 -9445 196 -9411
rect -196 -9451 196 -9445
rect -252 -9504 -206 -9492
rect -252 -9680 -246 -9504
rect -212 -9680 -206 -9504
rect -252 -9692 -206 -9680
rect 206 -9504 252 -9492
rect 206 -9680 212 -9504
rect 246 -9680 252 -9504
rect 206 -9692 252 -9680
rect -196 -9739 196 -9733
rect -196 -9773 -184 -9739
rect 184 -9773 196 -9739
rect -196 -9779 196 -9773
rect -196 -9847 196 -9841
rect -196 -9881 -184 -9847
rect 184 -9881 196 -9847
rect -196 -9887 196 -9881
rect -252 -9940 -206 -9928
rect -252 -10116 -246 -9940
rect -212 -10116 -206 -9940
rect -252 -10128 -206 -10116
rect 206 -9940 252 -9928
rect 206 -10116 212 -9940
rect 246 -10116 252 -9940
rect 206 -10128 252 -10116
rect -196 -10175 196 -10169
rect -196 -10209 -184 -10175
rect 184 -10209 196 -10175
rect -196 -10215 196 -10209
rect -196 -10283 196 -10277
rect -196 -10317 -184 -10283
rect 184 -10317 196 -10283
rect -196 -10323 196 -10317
rect -252 -10376 -206 -10364
rect -252 -10552 -246 -10376
rect -212 -10552 -206 -10376
rect -252 -10564 -206 -10552
rect 206 -10376 252 -10364
rect 206 -10552 212 -10376
rect 246 -10552 252 -10376
rect 206 -10564 252 -10552
rect -196 -10611 196 -10605
rect -196 -10645 -184 -10611
rect 184 -10645 196 -10611
rect -196 -10651 196 -10645
rect -196 -10719 196 -10713
rect -196 -10753 -184 -10719
rect 184 -10753 196 -10719
rect -196 -10759 196 -10753
rect -252 -10812 -206 -10800
rect -252 -10988 -246 -10812
rect -212 -10988 -206 -10812
rect -252 -11000 -206 -10988
rect 206 -10812 252 -10800
rect 206 -10988 212 -10812
rect 246 -10988 252 -10812
rect 206 -11000 252 -10988
rect -196 -11047 196 -11041
rect -196 -11081 -184 -11047
rect 184 -11081 196 -11047
rect -196 -11087 196 -11081
rect -196 -11155 196 -11149
rect -196 -11189 -184 -11155
rect 184 -11189 196 -11155
rect -196 -11195 196 -11189
rect -252 -11248 -206 -11236
rect -252 -11424 -246 -11248
rect -212 -11424 -206 -11248
rect -252 -11436 -206 -11424
rect 206 -11248 252 -11236
rect 206 -11424 212 -11248
rect 246 -11424 252 -11248
rect 206 -11436 252 -11424
rect -196 -11483 196 -11477
rect -196 -11517 -184 -11483
rect 184 -11517 196 -11483
rect -196 -11523 196 -11517
rect -196 -11591 196 -11585
rect -196 -11625 -184 -11591
rect 184 -11625 196 -11591
rect -196 -11631 196 -11625
rect -252 -11684 -206 -11672
rect -252 -11860 -246 -11684
rect -212 -11860 -206 -11684
rect -252 -11872 -206 -11860
rect 206 -11684 252 -11672
rect 206 -11860 212 -11684
rect 246 -11860 252 -11684
rect 206 -11872 252 -11860
rect -196 -11919 196 -11913
rect -196 -11953 -184 -11919
rect 184 -11953 196 -11919
rect -196 -11959 196 -11953
rect -196 -12027 196 -12021
rect -196 -12061 -184 -12027
rect 184 -12061 196 -12027
rect -196 -12067 196 -12061
rect -252 -12120 -206 -12108
rect -252 -12296 -246 -12120
rect -212 -12296 -206 -12120
rect -252 -12308 -206 -12296
rect 206 -12120 252 -12108
rect 206 -12296 212 -12120
rect 246 -12296 252 -12120
rect 206 -12308 252 -12296
rect -196 -12355 196 -12349
rect -196 -12389 -184 -12355
rect 184 -12389 196 -12355
rect -196 -12395 196 -12389
rect -196 -12463 196 -12457
rect -196 -12497 -184 -12463
rect 184 -12497 196 -12463
rect -196 -12503 196 -12497
rect -252 -12556 -206 -12544
rect -252 -12732 -246 -12556
rect -212 -12732 -206 -12556
rect -252 -12744 -206 -12732
rect 206 -12556 252 -12544
rect 206 -12732 212 -12556
rect 246 -12732 252 -12556
rect 206 -12744 252 -12732
rect -196 -12791 196 -12785
rect -196 -12825 -184 -12791
rect 184 -12825 196 -12791
rect -196 -12831 196 -12825
rect -196 -12899 196 -12893
rect -196 -12933 -184 -12899
rect 184 -12933 196 -12899
rect -196 -12939 196 -12933
rect -252 -12992 -206 -12980
rect -252 -13168 -246 -12992
rect -212 -13168 -206 -12992
rect -252 -13180 -206 -13168
rect 206 -12992 252 -12980
rect 206 -13168 212 -12992
rect 246 -13168 252 -12992
rect 206 -13180 252 -13168
rect -196 -13227 196 -13221
rect -196 -13261 -184 -13227
rect 184 -13261 196 -13227
rect -196 -13267 196 -13261
rect -196 -13335 196 -13329
rect -196 -13369 -184 -13335
rect 184 -13369 196 -13335
rect -196 -13375 196 -13369
rect -252 -13428 -206 -13416
rect -252 -13604 -246 -13428
rect -212 -13604 -206 -13428
rect -252 -13616 -206 -13604
rect 206 -13428 252 -13416
rect 206 -13604 212 -13428
rect 246 -13604 252 -13428
rect 206 -13616 252 -13604
rect -196 -13663 196 -13657
rect -196 -13697 -184 -13663
rect 184 -13697 196 -13663
rect -196 -13703 196 -13697
rect -196 -13771 196 -13765
rect -196 -13805 -184 -13771
rect 184 -13805 196 -13771
rect -196 -13811 196 -13805
rect -252 -13864 -206 -13852
rect -252 -14040 -246 -13864
rect -212 -14040 -206 -13864
rect -252 -14052 -206 -14040
rect 206 -13864 252 -13852
rect 206 -14040 212 -13864
rect 246 -14040 252 -13864
rect 206 -14052 252 -14040
rect -196 -14099 196 -14093
rect -196 -14133 -184 -14099
rect 184 -14133 196 -14099
rect -196 -14139 196 -14133
rect -196 -14207 196 -14201
rect -196 -14241 -184 -14207
rect 184 -14241 196 -14207
rect -196 -14247 196 -14241
rect -252 -14300 -206 -14288
rect -252 -14476 -246 -14300
rect -212 -14476 -206 -14300
rect -252 -14488 -206 -14476
rect 206 -14300 252 -14288
rect 206 -14476 212 -14300
rect 246 -14476 252 -14300
rect 206 -14488 252 -14476
rect -196 -14535 196 -14529
rect -196 -14569 -184 -14535
rect 184 -14569 196 -14535
rect -196 -14575 196 -14569
rect -196 -14643 196 -14637
rect -196 -14677 -184 -14643
rect 184 -14677 196 -14643
rect -196 -14683 196 -14677
rect -252 -14736 -206 -14724
rect -252 -14912 -246 -14736
rect -212 -14912 -206 -14736
rect -252 -14924 -206 -14912
rect 206 -14736 252 -14724
rect 206 -14912 212 -14736
rect 246 -14912 252 -14736
rect 206 -14924 252 -14912
rect -196 -14971 196 -14965
rect -196 -15005 -184 -14971
rect 184 -15005 196 -14971
rect -196 -15011 196 -15005
rect -196 -15079 196 -15073
rect -196 -15113 -184 -15079
rect 184 -15113 196 -15079
rect -196 -15119 196 -15113
rect -252 -15172 -206 -15160
rect -252 -15348 -246 -15172
rect -212 -15348 -206 -15172
rect -252 -15360 -206 -15348
rect 206 -15172 252 -15160
rect 206 -15348 212 -15172
rect 246 -15348 252 -15172
rect 206 -15360 252 -15348
rect -196 -15407 196 -15401
rect -196 -15441 -184 -15407
rect 184 -15441 196 -15407
rect -196 -15447 196 -15441
rect -196 -15515 196 -15509
rect -196 -15549 -184 -15515
rect 184 -15549 196 -15515
rect -196 -15555 196 -15549
rect -252 -15608 -206 -15596
rect -252 -15784 -246 -15608
rect -212 -15784 -206 -15608
rect -252 -15796 -206 -15784
rect 206 -15608 252 -15596
rect 206 -15784 212 -15608
rect 246 -15784 252 -15608
rect 206 -15796 252 -15784
rect -196 -15843 196 -15837
rect -196 -15877 -184 -15843
rect 184 -15877 196 -15843
rect -196 -15883 196 -15877
rect -196 -15951 196 -15945
rect -196 -15985 -184 -15951
rect 184 -15985 196 -15951
rect -196 -15991 196 -15985
rect -252 -16044 -206 -16032
rect -252 -16220 -246 -16044
rect -212 -16220 -206 -16044
rect -252 -16232 -206 -16220
rect 206 -16044 252 -16032
rect 206 -16220 212 -16044
rect 246 -16220 252 -16044
rect 206 -16232 252 -16220
rect -196 -16279 196 -16273
rect -196 -16313 -184 -16279
rect 184 -16313 196 -16279
rect -196 -16319 196 -16313
rect -196 -16387 196 -16381
rect -196 -16421 -184 -16387
rect 184 -16421 196 -16387
rect -196 -16427 196 -16421
rect -252 -16480 -206 -16468
rect -252 -16656 -246 -16480
rect -212 -16656 -206 -16480
rect -252 -16668 -206 -16656
rect 206 -16480 252 -16468
rect 206 -16656 212 -16480
rect 246 -16656 252 -16480
rect 206 -16668 252 -16656
rect -196 -16715 196 -16709
rect -196 -16749 -184 -16715
rect 184 -16749 196 -16715
rect -196 -16755 196 -16749
rect -196 -16823 196 -16817
rect -196 -16857 -184 -16823
rect 184 -16857 196 -16823
rect -196 -16863 196 -16857
rect -252 -16916 -206 -16904
rect -252 -17092 -246 -16916
rect -212 -17092 -206 -16916
rect -252 -17104 -206 -17092
rect 206 -16916 252 -16904
rect 206 -17092 212 -16916
rect 246 -17092 252 -16916
rect 206 -17104 252 -17092
rect -196 -17151 196 -17145
rect -196 -17185 -184 -17151
rect 184 -17185 196 -17151
rect -196 -17191 196 -17185
rect -196 -17259 196 -17253
rect -196 -17293 -184 -17259
rect 184 -17293 196 -17259
rect -196 -17299 196 -17293
rect -252 -17352 -206 -17340
rect -252 -17528 -246 -17352
rect -212 -17528 -206 -17352
rect -252 -17540 -206 -17528
rect 206 -17352 252 -17340
rect 206 -17528 212 -17352
rect 246 -17528 252 -17352
rect 206 -17540 252 -17528
rect -196 -17587 196 -17581
rect -196 -17621 -184 -17587
rect 184 -17621 196 -17587
rect -196 -17627 196 -17621
rect -196 -17695 196 -17689
rect -196 -17729 -184 -17695
rect 184 -17729 196 -17695
rect -196 -17735 196 -17729
rect -252 -17788 -206 -17776
rect -252 -17964 -246 -17788
rect -212 -17964 -206 -17788
rect -252 -17976 -206 -17964
rect 206 -17788 252 -17776
rect 206 -17964 212 -17788
rect 246 -17964 252 -17788
rect 206 -17976 252 -17964
rect -196 -18023 196 -18017
rect -196 -18057 -184 -18023
rect 184 -18057 196 -18023
rect -196 -18063 196 -18057
rect -196 -18131 196 -18125
rect -196 -18165 -184 -18131
rect 184 -18165 196 -18131
rect -196 -18171 196 -18165
rect -252 -18224 -206 -18212
rect -252 -18400 -246 -18224
rect -212 -18400 -206 -18224
rect -252 -18412 -206 -18400
rect 206 -18224 252 -18212
rect 206 -18400 212 -18224
rect 246 -18400 252 -18224
rect 206 -18412 252 -18400
rect -196 -18459 196 -18453
rect -196 -18493 -184 -18459
rect 184 -18493 196 -18459
rect -196 -18499 196 -18493
rect -196 -18567 196 -18561
rect -196 -18601 -184 -18567
rect 184 -18601 196 -18567
rect -196 -18607 196 -18601
rect -252 -18660 -206 -18648
rect -252 -18836 -246 -18660
rect -212 -18836 -206 -18660
rect -252 -18848 -206 -18836
rect 206 -18660 252 -18648
rect 206 -18836 212 -18660
rect 246 -18836 252 -18660
rect 206 -18848 252 -18836
rect -196 -18895 196 -18889
rect -196 -18929 -184 -18895
rect 184 -18929 196 -18895
rect -196 -18935 196 -18929
rect -196 -19003 196 -18997
rect -196 -19037 -184 -19003
rect 184 -19037 196 -19003
rect -196 -19043 196 -19037
rect -252 -19096 -206 -19084
rect -252 -19272 -246 -19096
rect -212 -19272 -206 -19096
rect -252 -19284 -206 -19272
rect 206 -19096 252 -19084
rect 206 -19272 212 -19096
rect 246 -19272 252 -19096
rect 206 -19284 252 -19272
rect -196 -19331 196 -19325
rect -196 -19365 -184 -19331
rect 184 -19365 196 -19331
rect -196 -19371 196 -19365
rect -196 -19439 196 -19433
rect -196 -19473 -184 -19439
rect 184 -19473 196 -19439
rect -196 -19479 196 -19473
rect -252 -19532 -206 -19520
rect -252 -19708 -246 -19532
rect -212 -19708 -206 -19532
rect -252 -19720 -206 -19708
rect 206 -19532 252 -19520
rect 206 -19708 212 -19532
rect 246 -19708 252 -19532
rect 206 -19720 252 -19708
rect -196 -19767 196 -19761
rect -196 -19801 -184 -19767
rect 184 -19801 196 -19767
rect -196 -19807 196 -19801
rect -196 -19875 196 -19869
rect -196 -19909 -184 -19875
rect 184 -19909 196 -19875
rect -196 -19915 196 -19909
rect -252 -19968 -206 -19956
rect -252 -20144 -246 -19968
rect -212 -20144 -206 -19968
rect -252 -20156 -206 -20144
rect 206 -19968 252 -19956
rect 206 -20144 212 -19968
rect 246 -20144 252 -19968
rect 206 -20156 252 -20144
rect -196 -20203 196 -20197
rect -196 -20237 -184 -20203
rect 184 -20237 196 -20203
rect -196 -20243 196 -20237
rect -196 -20311 196 -20305
rect -196 -20345 -184 -20311
rect 184 -20345 196 -20311
rect -196 -20351 196 -20345
rect -252 -20404 -206 -20392
rect -252 -20580 -246 -20404
rect -212 -20580 -206 -20404
rect -252 -20592 -206 -20580
rect 206 -20404 252 -20392
rect 206 -20580 212 -20404
rect 246 -20580 252 -20404
rect 206 -20592 252 -20580
rect -196 -20639 196 -20633
rect -196 -20673 -184 -20639
rect 184 -20673 196 -20639
rect -196 -20679 196 -20673
rect -196 -20747 196 -20741
rect -196 -20781 -184 -20747
rect 184 -20781 196 -20747
rect -196 -20787 196 -20781
rect -252 -20840 -206 -20828
rect -252 -21016 -246 -20840
rect -212 -21016 -206 -20840
rect -252 -21028 -206 -21016
rect 206 -20840 252 -20828
rect 206 -21016 212 -20840
rect 246 -21016 252 -20840
rect 206 -21028 252 -21016
rect -196 -21075 196 -21069
rect -196 -21109 -184 -21075
rect 184 -21109 196 -21075
rect -196 -21115 196 -21109
rect -196 -21183 196 -21177
rect -196 -21217 -184 -21183
rect 184 -21217 196 -21183
rect -196 -21223 196 -21217
rect -252 -21276 -206 -21264
rect -252 -21452 -246 -21276
rect -212 -21452 -206 -21276
rect -252 -21464 -206 -21452
rect 206 -21276 252 -21264
rect 206 -21452 212 -21276
rect 246 -21452 252 -21276
rect 206 -21464 252 -21452
rect -196 -21511 196 -21505
rect -196 -21545 -184 -21511
rect 184 -21545 196 -21511
rect -196 -21551 196 -21545
rect -196 -21619 196 -21613
rect -196 -21653 -184 -21619
rect 184 -21653 196 -21619
rect -196 -21659 196 -21653
rect -252 -21712 -206 -21700
rect -252 -21888 -246 -21712
rect -212 -21888 -206 -21712
rect -252 -21900 -206 -21888
rect 206 -21712 252 -21700
rect 206 -21888 212 -21712
rect 246 -21888 252 -21712
rect 206 -21900 252 -21888
rect -196 -21947 196 -21941
rect -196 -21981 -184 -21947
rect 184 -21981 196 -21947
rect -196 -21987 196 -21981
rect -196 -22055 196 -22049
rect -196 -22089 -184 -22055
rect 184 -22089 196 -22055
rect -196 -22095 196 -22089
rect -252 -22148 -206 -22136
rect -252 -22324 -246 -22148
rect -212 -22324 -206 -22148
rect -252 -22336 -206 -22324
rect 206 -22148 252 -22136
rect 206 -22324 212 -22148
rect 246 -22324 252 -22148
rect 206 -22336 252 -22324
rect -196 -22383 196 -22377
rect -196 -22417 -184 -22383
rect 184 -22417 196 -22383
rect -196 -22423 196 -22417
rect -196 -22491 196 -22485
rect -196 -22525 -184 -22491
rect 184 -22525 196 -22491
rect -196 -22531 196 -22525
rect -252 -22584 -206 -22572
rect -252 -22760 -246 -22584
rect -212 -22760 -206 -22584
rect -252 -22772 -206 -22760
rect 206 -22584 252 -22572
rect 206 -22760 212 -22584
rect 246 -22760 252 -22584
rect 206 -22772 252 -22760
rect -196 -22819 196 -22813
rect -196 -22853 -184 -22819
rect 184 -22853 196 -22819
rect -196 -22859 196 -22853
rect -196 -22927 196 -22921
rect -196 -22961 -184 -22927
rect 184 -22961 196 -22927
rect -196 -22967 196 -22961
rect -252 -23020 -206 -23008
rect -252 -23196 -246 -23020
rect -212 -23196 -206 -23020
rect -252 -23208 -206 -23196
rect 206 -23020 252 -23008
rect 206 -23196 212 -23020
rect 246 -23196 252 -23020
rect 206 -23208 252 -23196
rect -196 -23255 196 -23249
rect -196 -23289 -184 -23255
rect 184 -23289 196 -23255
rect -196 -23295 196 -23289
rect -196 -23363 196 -23357
rect -196 -23397 -184 -23363
rect 184 -23397 196 -23363
rect -196 -23403 196 -23397
rect -252 -23456 -206 -23444
rect -252 -23632 -246 -23456
rect -212 -23632 -206 -23456
rect -252 -23644 -206 -23632
rect 206 -23456 252 -23444
rect 206 -23632 212 -23456
rect 246 -23632 252 -23456
rect 206 -23644 252 -23632
rect -196 -23691 196 -23685
rect -196 -23725 -184 -23691
rect 184 -23725 196 -23691
rect -196 -23731 196 -23725
rect -196 -23799 196 -23793
rect -196 -23833 -184 -23799
rect 184 -23833 196 -23799
rect -196 -23839 196 -23833
rect -252 -23892 -206 -23880
rect -252 -24068 -246 -23892
rect -212 -24068 -206 -23892
rect -252 -24080 -206 -24068
rect 206 -23892 252 -23880
rect 206 -24068 212 -23892
rect 246 -24068 252 -23892
rect 206 -24080 252 -24068
rect -196 -24127 196 -24121
rect -196 -24161 -184 -24127
rect 184 -24161 196 -24127
rect -196 -24167 196 -24161
rect -196 -24235 196 -24229
rect -196 -24269 -184 -24235
rect 184 -24269 196 -24235
rect -196 -24275 196 -24269
rect -252 -24328 -206 -24316
rect -252 -24504 -246 -24328
rect -212 -24504 -206 -24328
rect -252 -24516 -206 -24504
rect 206 -24328 252 -24316
rect 206 -24504 212 -24328
rect 246 -24504 252 -24328
rect 206 -24516 252 -24504
rect -196 -24563 196 -24557
rect -196 -24597 -184 -24563
rect 184 -24597 196 -24563
rect -196 -24603 196 -24597
rect -196 -24671 196 -24665
rect -196 -24705 -184 -24671
rect 184 -24705 196 -24671
rect -196 -24711 196 -24705
rect -252 -24764 -206 -24752
rect -252 -24940 -246 -24764
rect -212 -24940 -206 -24764
rect -252 -24952 -206 -24940
rect 206 -24764 252 -24752
rect 206 -24940 212 -24764
rect 246 -24940 252 -24764
rect 206 -24952 252 -24940
rect -196 -24999 196 -24993
rect -196 -25033 -184 -24999
rect 184 -25033 196 -24999
rect -196 -25039 196 -25033
rect -196 -25107 196 -25101
rect -196 -25141 -184 -25107
rect 184 -25141 196 -25107
rect -196 -25147 196 -25141
rect -252 -25200 -206 -25188
rect -252 -25376 -246 -25200
rect -212 -25376 -206 -25200
rect -252 -25388 -206 -25376
rect 206 -25200 252 -25188
rect 206 -25376 212 -25200
rect 246 -25376 252 -25200
rect 206 -25388 252 -25376
rect -196 -25435 196 -25429
rect -196 -25469 -184 -25435
rect 184 -25469 196 -25435
rect -196 -25475 196 -25469
rect -196 -25543 196 -25537
rect -196 -25577 -184 -25543
rect 184 -25577 196 -25543
rect -196 -25583 196 -25577
rect -252 -25636 -206 -25624
rect -252 -25812 -246 -25636
rect -212 -25812 -206 -25636
rect -252 -25824 -206 -25812
rect 206 -25636 252 -25624
rect 206 -25812 212 -25636
rect 246 -25812 252 -25636
rect 206 -25824 252 -25812
rect -196 -25871 196 -25865
rect -196 -25905 -184 -25871
rect 184 -25905 196 -25871
rect -196 -25911 196 -25905
rect -196 -25979 196 -25973
rect -196 -26013 -184 -25979
rect 184 -26013 196 -25979
rect -196 -26019 196 -26013
rect -252 -26072 -206 -26060
rect -252 -26248 -246 -26072
rect -212 -26248 -206 -26072
rect -252 -26260 -206 -26248
rect 206 -26072 252 -26060
rect 206 -26248 212 -26072
rect 246 -26248 252 -26072
rect 206 -26260 252 -26248
rect -196 -26307 196 -26301
rect -196 -26341 -184 -26307
rect 184 -26341 196 -26307
rect -196 -26347 196 -26341
rect -196 -26415 196 -26409
rect -196 -26449 -184 -26415
rect 184 -26449 196 -26415
rect -196 -26455 196 -26449
rect -252 -26508 -206 -26496
rect -252 -26684 -246 -26508
rect -212 -26684 -206 -26508
rect -252 -26696 -206 -26684
rect 206 -26508 252 -26496
rect 206 -26684 212 -26508
rect 246 -26684 252 -26508
rect 206 -26696 252 -26684
rect -196 -26743 196 -26737
rect -196 -26777 -184 -26743
rect 184 -26777 196 -26743
rect -196 -26783 196 -26777
rect -196 -26851 196 -26845
rect -196 -26885 -184 -26851
rect 184 -26885 196 -26851
rect -196 -26891 196 -26885
rect -252 -26944 -206 -26932
rect -252 -27120 -246 -26944
rect -212 -27120 -206 -26944
rect -252 -27132 -206 -27120
rect 206 -26944 252 -26932
rect 206 -27120 212 -26944
rect 246 -27120 252 -26944
rect 206 -27132 252 -27120
rect -196 -27179 196 -27173
rect -196 -27213 -184 -27179
rect 184 -27213 196 -27179
rect -196 -27219 196 -27213
rect -196 -27287 196 -27281
rect -196 -27321 -184 -27287
rect 184 -27321 196 -27287
rect -196 -27327 196 -27321
rect -252 -27380 -206 -27368
rect -252 -27556 -246 -27380
rect -212 -27556 -206 -27380
rect -252 -27568 -206 -27556
rect 206 -27380 252 -27368
rect 206 -27556 212 -27380
rect 246 -27556 252 -27380
rect 206 -27568 252 -27556
rect -196 -27615 196 -27609
rect -196 -27649 -184 -27615
rect 184 -27649 196 -27615
rect -196 -27655 196 -27649
rect -196 -27723 196 -27717
rect -196 -27757 -184 -27723
rect 184 -27757 196 -27723
rect -196 -27763 196 -27757
rect -252 -27816 -206 -27804
rect -252 -27992 -246 -27816
rect -212 -27992 -206 -27816
rect -252 -28004 -206 -27992
rect 206 -27816 252 -27804
rect 206 -27992 212 -27816
rect 246 -27992 252 -27816
rect 206 -28004 252 -27992
rect -196 -28051 196 -28045
rect -196 -28085 -184 -28051
rect 184 -28085 196 -28051
rect -196 -28091 196 -28085
rect -196 -28159 196 -28153
rect -196 -28193 -184 -28159
rect 184 -28193 196 -28159
rect -196 -28199 196 -28193
rect -252 -28252 -206 -28240
rect -252 -28428 -246 -28252
rect -212 -28428 -206 -28252
rect -252 -28440 -206 -28428
rect 206 -28252 252 -28240
rect 206 -28428 212 -28252
rect 246 -28428 252 -28252
rect 206 -28440 252 -28428
rect -196 -28487 196 -28481
rect -196 -28521 -184 -28487
rect 184 -28521 196 -28487
rect -196 -28527 196 -28521
rect -196 -28595 196 -28589
rect -196 -28629 -184 -28595
rect 184 -28629 196 -28595
rect -196 -28635 196 -28629
rect -252 -28688 -206 -28676
rect -252 -28864 -246 -28688
rect -212 -28864 -206 -28688
rect -252 -28876 -206 -28864
rect 206 -28688 252 -28676
rect 206 -28864 212 -28688
rect 246 -28864 252 -28688
rect 206 -28876 252 -28864
rect -196 -28923 196 -28917
rect -196 -28957 -184 -28923
rect 184 -28957 196 -28923
rect -196 -28963 196 -28957
rect -196 -29031 196 -29025
rect -196 -29065 -184 -29031
rect 184 -29065 196 -29031
rect -196 -29071 196 -29065
rect -252 -29124 -206 -29112
rect -252 -29300 -246 -29124
rect -212 -29300 -206 -29124
rect -252 -29312 -206 -29300
rect 206 -29124 252 -29112
rect 206 -29300 212 -29124
rect 246 -29300 252 -29124
rect 206 -29312 252 -29300
rect -196 -29359 196 -29353
rect -196 -29393 -184 -29359
rect 184 -29393 196 -29359
rect -196 -29399 196 -29393
rect -196 -29467 196 -29461
rect -196 -29501 -184 -29467
rect 184 -29501 196 -29467
rect -196 -29507 196 -29501
rect -252 -29560 -206 -29548
rect -252 -29736 -246 -29560
rect -212 -29736 -206 -29560
rect -252 -29748 -206 -29736
rect 206 -29560 252 -29548
rect 206 -29736 212 -29560
rect 246 -29736 252 -29560
rect 206 -29748 252 -29736
rect -196 -29795 196 -29789
rect -196 -29829 -184 -29795
rect 184 -29829 196 -29795
rect -196 -29835 196 -29829
rect -196 -29903 196 -29897
rect -196 -29937 -184 -29903
rect 184 -29937 196 -29903
rect -196 -29943 196 -29937
rect -252 -29996 -206 -29984
rect -252 -30172 -246 -29996
rect -212 -30172 -206 -29996
rect -252 -30184 -206 -30172
rect 206 -29996 252 -29984
rect 206 -30172 212 -29996
rect 246 -30172 252 -29996
rect 206 -30184 252 -30172
rect -196 -30231 196 -30225
rect -196 -30265 -184 -30231
rect 184 -30265 196 -30231
rect -196 -30271 196 -30265
rect -196 -30339 196 -30333
rect -196 -30373 -184 -30339
rect 184 -30373 196 -30339
rect -196 -30379 196 -30373
rect -252 -30432 -206 -30420
rect -252 -30608 -246 -30432
rect -212 -30608 -206 -30432
rect -252 -30620 -206 -30608
rect 206 -30432 252 -30420
rect 206 -30608 212 -30432
rect 246 -30608 252 -30432
rect 206 -30620 252 -30608
rect -196 -30667 196 -30661
rect -196 -30701 -184 -30667
rect 184 -30701 196 -30667
rect -196 -30707 196 -30701
rect -196 -30775 196 -30769
rect -196 -30809 -184 -30775
rect 184 -30809 196 -30775
rect -196 -30815 196 -30809
rect -252 -30868 -206 -30856
rect -252 -31044 -246 -30868
rect -212 -31044 -206 -30868
rect -252 -31056 -206 -31044
rect 206 -30868 252 -30856
rect 206 -31044 212 -30868
rect 246 -31044 252 -30868
rect 206 -31056 252 -31044
rect -196 -31103 196 -31097
rect -196 -31137 -184 -31103
rect 184 -31137 196 -31103
rect -196 -31143 196 -31137
rect -196 -31211 196 -31205
rect -196 -31245 -184 -31211
rect 184 -31245 196 -31211
rect -196 -31251 196 -31245
rect -252 -31304 -206 -31292
rect -252 -31480 -246 -31304
rect -212 -31480 -206 -31304
rect -252 -31492 -206 -31480
rect 206 -31304 252 -31292
rect 206 -31480 212 -31304
rect 246 -31480 252 -31304
rect 206 -31492 252 -31480
rect -196 -31539 196 -31533
rect -196 -31573 -184 -31539
rect 184 -31573 196 -31539
rect -196 -31579 196 -31573
rect -196 -31647 196 -31641
rect -196 -31681 -184 -31647
rect 184 -31681 196 -31647
rect -196 -31687 196 -31681
rect -252 -31740 -206 -31728
rect -252 -31916 -246 -31740
rect -212 -31916 -206 -31740
rect -252 -31928 -206 -31916
rect 206 -31740 252 -31728
rect 206 -31916 212 -31740
rect 246 -31916 252 -31740
rect 206 -31928 252 -31916
rect -196 -31975 196 -31969
rect -196 -32009 -184 -31975
rect 184 -32009 196 -31975
rect -196 -32015 196 -32009
rect -196 -32083 196 -32077
rect -196 -32117 -184 -32083
rect 184 -32117 196 -32083
rect -196 -32123 196 -32117
rect -252 -32176 -206 -32164
rect -252 -32352 -246 -32176
rect -212 -32352 -206 -32176
rect -252 -32364 -206 -32352
rect 206 -32176 252 -32164
rect 206 -32352 212 -32176
rect 246 -32352 252 -32176
rect 206 -32364 252 -32352
rect -196 -32411 196 -32405
rect -196 -32445 -184 -32411
rect 184 -32445 196 -32411
rect -196 -32451 196 -32445
rect -196 -32519 196 -32513
rect -196 -32553 -184 -32519
rect 184 -32553 196 -32519
rect -196 -32559 196 -32553
rect -252 -32612 -206 -32600
rect -252 -32788 -246 -32612
rect -212 -32788 -206 -32612
rect -252 -32800 -206 -32788
rect 206 -32612 252 -32600
rect 206 -32788 212 -32612
rect 246 -32788 252 -32612
rect 206 -32800 252 -32788
rect -196 -32847 196 -32841
rect -196 -32881 -184 -32847
rect 184 -32881 196 -32847
rect -196 -32887 196 -32881
rect -196 -32955 196 -32949
rect -196 -32989 -184 -32955
rect 184 -32989 196 -32955
rect -196 -32995 196 -32989
rect -252 -33048 -206 -33036
rect -252 -33224 -246 -33048
rect -212 -33224 -206 -33048
rect -252 -33236 -206 -33224
rect 206 -33048 252 -33036
rect 206 -33224 212 -33048
rect 246 -33224 252 -33048
rect 206 -33236 252 -33224
rect -196 -33283 196 -33277
rect -196 -33317 -184 -33283
rect 184 -33317 196 -33283
rect -196 -33323 196 -33317
rect -196 -33391 196 -33385
rect -196 -33425 -184 -33391
rect 184 -33425 196 -33391
rect -196 -33431 196 -33425
rect -252 -33484 -206 -33472
rect -252 -33660 -246 -33484
rect -212 -33660 -206 -33484
rect -252 -33672 -206 -33660
rect 206 -33484 252 -33472
rect 206 -33660 212 -33484
rect 246 -33660 252 -33484
rect 206 -33672 252 -33660
rect -196 -33719 196 -33713
rect -196 -33753 -184 -33719
rect 184 -33753 196 -33719
rect -196 -33759 196 -33753
rect -196 -33827 196 -33821
rect -196 -33861 -184 -33827
rect 184 -33861 196 -33827
rect -196 -33867 196 -33861
rect -252 -33920 -206 -33908
rect -252 -34096 -246 -33920
rect -212 -34096 -206 -33920
rect -252 -34108 -206 -34096
rect 206 -33920 252 -33908
rect 206 -34096 212 -33920
rect 246 -34096 252 -33920
rect 206 -34108 252 -34096
rect -196 -34155 196 -34149
rect -196 -34189 -184 -34155
rect 184 -34189 196 -34155
rect -196 -34195 196 -34189
rect -196 -34263 196 -34257
rect -196 -34297 -184 -34263
rect 184 -34297 196 -34263
rect -196 -34303 196 -34297
rect -252 -34356 -206 -34344
rect -252 -34532 -246 -34356
rect -212 -34532 -206 -34356
rect -252 -34544 -206 -34532
rect 206 -34356 252 -34344
rect 206 -34532 212 -34356
rect 246 -34532 252 -34356
rect 206 -34544 252 -34532
rect -196 -34591 196 -34585
rect -196 -34625 -184 -34591
rect 184 -34625 196 -34591
rect -196 -34631 196 -34625
rect -196 -34699 196 -34693
rect -196 -34733 -184 -34699
rect 184 -34733 196 -34699
rect -196 -34739 196 -34733
rect -252 -34792 -206 -34780
rect -252 -34968 -246 -34792
rect -212 -34968 -206 -34792
rect -252 -34980 -206 -34968
rect 206 -34792 252 -34780
rect 206 -34968 212 -34792
rect 246 -34968 252 -34792
rect 206 -34980 252 -34968
rect -196 -35027 196 -35021
rect -196 -35061 -184 -35027
rect 184 -35061 196 -35027
rect -196 -35067 196 -35061
rect -196 -35135 196 -35129
rect -196 -35169 -184 -35135
rect 184 -35169 196 -35135
rect -196 -35175 196 -35169
rect -252 -35228 -206 -35216
rect -252 -35404 -246 -35228
rect -212 -35404 -206 -35228
rect -252 -35416 -206 -35404
rect 206 -35228 252 -35216
rect 206 -35404 212 -35228
rect 246 -35404 252 -35228
rect 206 -35416 252 -35404
rect -196 -35463 196 -35457
rect -196 -35497 -184 -35463
rect 184 -35497 196 -35463
rect -196 -35503 196 -35497
rect -196 -35571 196 -35565
rect -196 -35605 -184 -35571
rect 184 -35605 196 -35571
rect -196 -35611 196 -35605
rect -252 -35664 -206 -35652
rect -252 -35840 -246 -35664
rect -212 -35840 -206 -35664
rect -252 -35852 -206 -35840
rect 206 -35664 252 -35652
rect 206 -35840 212 -35664
rect 246 -35840 252 -35664
rect 206 -35852 252 -35840
rect -196 -35899 196 -35893
rect -196 -35933 -184 -35899
rect 184 -35933 196 -35899
rect -196 -35939 196 -35933
rect -196 -36007 196 -36001
rect -196 -36041 -184 -36007
rect 184 -36041 196 -36007
rect -196 -36047 196 -36041
rect -252 -36100 -206 -36088
rect -252 -36276 -246 -36100
rect -212 -36276 -206 -36100
rect -252 -36288 -206 -36276
rect 206 -36100 252 -36088
rect 206 -36276 212 -36100
rect 246 -36276 252 -36100
rect 206 -36288 252 -36276
rect -196 -36335 196 -36329
rect -196 -36369 -184 -36335
rect 184 -36369 196 -36335
rect -196 -36375 196 -36369
rect -196 -36443 196 -36437
rect -196 -36477 -184 -36443
rect 184 -36477 196 -36443
rect -196 -36483 196 -36477
rect -252 -36536 -206 -36524
rect -252 -36712 -246 -36536
rect -212 -36712 -206 -36536
rect -252 -36724 -206 -36712
rect 206 -36536 252 -36524
rect 206 -36712 212 -36536
rect 246 -36712 252 -36536
rect 206 -36724 252 -36712
rect -196 -36771 196 -36765
rect -196 -36805 -184 -36771
rect 184 -36805 196 -36771
rect -196 -36811 196 -36805
rect -196 -36879 196 -36873
rect -196 -36913 -184 -36879
rect 184 -36913 196 -36879
rect -196 -36919 196 -36913
rect -252 -36972 -206 -36960
rect -252 -37148 -246 -36972
rect -212 -37148 -206 -36972
rect -252 -37160 -206 -37148
rect 206 -36972 252 -36960
rect 206 -37148 212 -36972
rect 246 -37148 252 -36972
rect 206 -37160 252 -37148
rect -196 -37207 196 -37201
rect -196 -37241 -184 -37207
rect 184 -37241 196 -37207
rect -196 -37247 196 -37241
rect -196 -37315 196 -37309
rect -196 -37349 -184 -37315
rect 184 -37349 196 -37315
rect -196 -37355 196 -37349
rect -252 -37408 -206 -37396
rect -252 -37584 -246 -37408
rect -212 -37584 -206 -37408
rect -252 -37596 -206 -37584
rect 206 -37408 252 -37396
rect 206 -37584 212 -37408
rect 246 -37584 252 -37408
rect 206 -37596 252 -37584
rect -196 -37643 196 -37637
rect -196 -37677 -184 -37643
rect 184 -37677 196 -37643
rect -196 -37683 196 -37677
rect -196 -37751 196 -37745
rect -196 -37785 -184 -37751
rect 184 -37785 196 -37751
rect -196 -37791 196 -37785
rect -252 -37844 -206 -37832
rect -252 -38020 -246 -37844
rect -212 -38020 -206 -37844
rect -252 -38032 -206 -38020
rect 206 -37844 252 -37832
rect 206 -38020 212 -37844
rect 246 -38020 252 -37844
rect 206 -38032 252 -38020
rect -196 -38079 196 -38073
rect -196 -38113 -184 -38079
rect 184 -38113 196 -38079
rect -196 -38119 196 -38113
rect -196 -38187 196 -38181
rect -196 -38221 -184 -38187
rect 184 -38221 196 -38187
rect -196 -38227 196 -38221
rect -252 -38280 -206 -38268
rect -252 -38456 -246 -38280
rect -212 -38456 -206 -38280
rect -252 -38468 -206 -38456
rect 206 -38280 252 -38268
rect 206 -38456 212 -38280
rect 246 -38456 252 -38280
rect 206 -38468 252 -38456
rect -196 -38515 196 -38509
rect -196 -38549 -184 -38515
rect 184 -38549 196 -38515
rect -196 -38555 196 -38549
rect -196 -38623 196 -38617
rect -196 -38657 -184 -38623
rect 184 -38657 196 -38623
rect -196 -38663 196 -38657
rect -252 -38716 -206 -38704
rect -252 -38892 -246 -38716
rect -212 -38892 -206 -38716
rect -252 -38904 -206 -38892
rect 206 -38716 252 -38704
rect 206 -38892 212 -38716
rect 246 -38892 252 -38716
rect 206 -38904 252 -38892
rect -196 -38951 196 -38945
rect -196 -38985 -184 -38951
rect 184 -38985 196 -38951
rect -196 -38991 196 -38985
rect -196 -39059 196 -39053
rect -196 -39093 -184 -39059
rect 184 -39093 196 -39059
rect -196 -39099 196 -39093
rect -252 -39152 -206 -39140
rect -252 -39328 -246 -39152
rect -212 -39328 -206 -39152
rect -252 -39340 -206 -39328
rect 206 -39152 252 -39140
rect 206 -39328 212 -39152
rect 246 -39328 252 -39152
rect 206 -39340 252 -39328
rect -196 -39387 196 -39381
rect -196 -39421 -184 -39387
rect 184 -39421 196 -39387
rect -196 -39427 196 -39421
rect -196 -39495 196 -39489
rect -196 -39529 -184 -39495
rect 184 -39529 196 -39495
rect -196 -39535 196 -39529
rect -252 -39588 -206 -39576
rect -252 -39764 -246 -39588
rect -212 -39764 -206 -39588
rect -252 -39776 -206 -39764
rect 206 -39588 252 -39576
rect 206 -39764 212 -39588
rect 246 -39764 252 -39588
rect 206 -39776 252 -39764
rect -196 -39823 196 -39817
rect -196 -39857 -184 -39823
rect 184 -39857 196 -39823
rect -196 -39863 196 -39857
rect -196 -39931 196 -39925
rect -196 -39965 -184 -39931
rect 184 -39965 196 -39931
rect -196 -39971 196 -39965
rect -252 -40024 -206 -40012
rect -252 -40200 -246 -40024
rect -212 -40200 -206 -40024
rect -252 -40212 -206 -40200
rect 206 -40024 252 -40012
rect 206 -40200 212 -40024
rect 246 -40200 252 -40024
rect 206 -40212 252 -40200
rect -196 -40259 196 -40253
rect -196 -40293 -184 -40259
rect 184 -40293 196 -40259
rect -196 -40299 196 -40293
rect -196 -40367 196 -40361
rect -196 -40401 -184 -40367
rect 184 -40401 196 -40367
rect -196 -40407 196 -40401
rect -252 -40460 -206 -40448
rect -252 -40636 -246 -40460
rect -212 -40636 -206 -40460
rect -252 -40648 -206 -40636
rect 206 -40460 252 -40448
rect 206 -40636 212 -40460
rect 246 -40636 252 -40460
rect 206 -40648 252 -40636
rect -196 -40695 196 -40689
rect -196 -40729 -184 -40695
rect 184 -40729 196 -40695
rect -196 -40735 196 -40729
rect -196 -40803 196 -40797
rect -196 -40837 -184 -40803
rect 184 -40837 196 -40803
rect -196 -40843 196 -40837
rect -252 -40896 -206 -40884
rect -252 -41072 -246 -40896
rect -212 -41072 -206 -40896
rect -252 -41084 -206 -41072
rect 206 -40896 252 -40884
rect 206 -41072 212 -40896
rect 246 -41072 252 -40896
rect 206 -41084 252 -41072
rect -196 -41131 196 -41125
rect -196 -41165 -184 -41131
rect 184 -41165 196 -41131
rect -196 -41171 196 -41165
rect -196 -41239 196 -41233
rect -196 -41273 -184 -41239
rect 184 -41273 196 -41239
rect -196 -41279 196 -41273
rect -252 -41332 -206 -41320
rect -252 -41508 -246 -41332
rect -212 -41508 -206 -41332
rect -252 -41520 -206 -41508
rect 206 -41332 252 -41320
rect 206 -41508 212 -41332
rect 246 -41508 252 -41332
rect 206 -41520 252 -41508
rect -196 -41567 196 -41561
rect -196 -41601 -184 -41567
rect 184 -41601 196 -41567
rect -196 -41607 196 -41601
rect -196 -41675 196 -41669
rect -196 -41709 -184 -41675
rect 184 -41709 196 -41675
rect -196 -41715 196 -41709
rect -252 -41768 -206 -41756
rect -252 -41944 -246 -41768
rect -212 -41944 -206 -41768
rect -252 -41956 -206 -41944
rect 206 -41768 252 -41756
rect 206 -41944 212 -41768
rect 246 -41944 252 -41768
rect 206 -41956 252 -41944
rect -196 -42003 196 -41997
rect -196 -42037 -184 -42003
rect 184 -42037 196 -42003
rect -196 -42043 196 -42037
rect -196 -42111 196 -42105
rect -196 -42145 -184 -42111
rect 184 -42145 196 -42111
rect -196 -42151 196 -42145
rect -252 -42204 -206 -42192
rect -252 -42380 -246 -42204
rect -212 -42380 -206 -42204
rect -252 -42392 -206 -42380
rect 206 -42204 252 -42192
rect 206 -42380 212 -42204
rect 246 -42380 252 -42204
rect 206 -42392 252 -42380
rect -196 -42439 196 -42433
rect -196 -42473 -184 -42439
rect 184 -42473 196 -42439
rect -196 -42479 196 -42473
rect -196 -42547 196 -42541
rect -196 -42581 -184 -42547
rect 184 -42581 196 -42547
rect -196 -42587 196 -42581
rect -252 -42640 -206 -42628
rect -252 -42816 -246 -42640
rect -212 -42816 -206 -42640
rect -252 -42828 -206 -42816
rect 206 -42640 252 -42628
rect 206 -42816 212 -42640
rect 246 -42816 252 -42640
rect 206 -42828 252 -42816
rect -196 -42875 196 -42869
rect -196 -42909 -184 -42875
rect 184 -42909 196 -42875
rect -196 -42915 196 -42909
rect -196 -42983 196 -42977
rect -196 -43017 -184 -42983
rect 184 -43017 196 -42983
rect -196 -43023 196 -43017
rect -252 -43076 -206 -43064
rect -252 -43252 -246 -43076
rect -212 -43252 -206 -43076
rect -252 -43264 -206 -43252
rect 206 -43076 252 -43064
rect 206 -43252 212 -43076
rect 246 -43252 252 -43076
rect 206 -43264 252 -43252
rect -196 -43311 196 -43305
rect -196 -43345 -184 -43311
rect 184 -43345 196 -43311
rect -196 -43351 196 -43345
rect -196 -43419 196 -43413
rect -196 -43453 -184 -43419
rect 184 -43453 196 -43419
rect -196 -43459 196 -43453
rect -252 -43512 -206 -43500
rect -252 -43688 -246 -43512
rect -212 -43688 -206 -43512
rect -252 -43700 -206 -43688
rect 206 -43512 252 -43500
rect 206 -43688 212 -43512
rect 246 -43688 252 -43512
rect 206 -43700 252 -43688
rect -196 -43747 196 -43741
rect -196 -43781 -184 -43747
rect 184 -43781 196 -43747
rect -196 -43787 196 -43781
rect -196 -43855 196 -43849
rect -196 -43889 -184 -43855
rect 184 -43889 196 -43855
rect -196 -43895 196 -43889
rect -252 -43948 -206 -43936
rect -252 -44124 -246 -43948
rect -212 -44124 -206 -43948
rect -252 -44136 -206 -44124
rect 206 -43948 252 -43936
rect 206 -44124 212 -43948
rect 246 -44124 252 -43948
rect 206 -44136 252 -44124
rect -196 -44183 196 -44177
rect -196 -44217 -184 -44183
rect 184 -44217 196 -44183
rect -196 -44223 196 -44217
rect -196 -44291 196 -44285
rect -196 -44325 -184 -44291
rect 184 -44325 196 -44291
rect -196 -44331 196 -44325
rect -252 -44384 -206 -44372
rect -252 -44560 -246 -44384
rect -212 -44560 -206 -44384
rect -252 -44572 -206 -44560
rect 206 -44384 252 -44372
rect 206 -44560 212 -44384
rect 246 -44560 252 -44384
rect 206 -44572 252 -44560
rect -196 -44619 196 -44613
rect -196 -44653 -184 -44619
rect 184 -44653 196 -44619
rect -196 -44659 196 -44653
rect -196 -44727 196 -44721
rect -196 -44761 -184 -44727
rect 184 -44761 196 -44727
rect -196 -44767 196 -44761
rect -252 -44820 -206 -44808
rect -252 -44996 -246 -44820
rect -212 -44996 -206 -44820
rect -252 -45008 -206 -44996
rect 206 -44820 252 -44808
rect 206 -44996 212 -44820
rect 246 -44996 252 -44820
rect 206 -45008 252 -44996
rect -196 -45055 196 -45049
rect -196 -45089 -184 -45055
rect 184 -45089 196 -45055
rect -196 -45095 196 -45089
rect -196 -45163 196 -45157
rect -196 -45197 -184 -45163
rect 184 -45197 196 -45163
rect -196 -45203 196 -45197
rect -252 -45256 -206 -45244
rect -252 -45432 -246 -45256
rect -212 -45432 -206 -45256
rect -252 -45444 -206 -45432
rect 206 -45256 252 -45244
rect 206 -45432 212 -45256
rect 246 -45432 252 -45256
rect 206 -45444 252 -45432
rect -196 -45491 196 -45485
rect -196 -45525 -184 -45491
rect 184 -45525 196 -45491
rect -196 -45531 196 -45525
rect -196 -45599 196 -45593
rect -196 -45633 -184 -45599
rect 184 -45633 196 -45599
rect -196 -45639 196 -45633
rect -252 -45692 -206 -45680
rect -252 -45868 -246 -45692
rect -212 -45868 -206 -45692
rect -252 -45880 -206 -45868
rect 206 -45692 252 -45680
rect 206 -45868 212 -45692
rect 246 -45868 252 -45692
rect 206 -45880 252 -45868
rect -196 -45927 196 -45921
rect -196 -45961 -184 -45927
rect 184 -45961 196 -45927
rect -196 -45967 196 -45961
rect -196 -46035 196 -46029
rect -196 -46069 -184 -46035
rect 184 -46069 196 -46035
rect -196 -46075 196 -46069
rect -252 -46128 -206 -46116
rect -252 -46304 -246 -46128
rect -212 -46304 -206 -46128
rect -252 -46316 -206 -46304
rect 206 -46128 252 -46116
rect 206 -46304 212 -46128
rect 246 -46304 252 -46128
rect 206 -46316 252 -46304
rect -196 -46363 196 -46357
rect -196 -46397 -184 -46363
rect 184 -46397 196 -46363
rect -196 -46403 196 -46397
rect -196 -46471 196 -46465
rect -196 -46505 -184 -46471
rect 184 -46505 196 -46471
rect -196 -46511 196 -46505
rect -252 -46564 -206 -46552
rect -252 -46740 -246 -46564
rect -212 -46740 -206 -46564
rect -252 -46752 -206 -46740
rect 206 -46564 252 -46552
rect 206 -46740 212 -46564
rect 246 -46740 252 -46564
rect 206 -46752 252 -46740
rect -196 -46799 196 -46793
rect -196 -46833 -184 -46799
rect 184 -46833 196 -46799
rect -196 -46839 196 -46833
rect -196 -46907 196 -46901
rect -196 -46941 -184 -46907
rect 184 -46941 196 -46907
rect -196 -46947 196 -46941
rect -252 -47000 -206 -46988
rect -252 -47176 -246 -47000
rect -212 -47176 -206 -47000
rect -252 -47188 -206 -47176
rect 206 -47000 252 -46988
rect 206 -47176 212 -47000
rect 246 -47176 252 -47000
rect 206 -47188 252 -47176
rect -196 -47235 196 -47229
rect -196 -47269 -184 -47235
rect 184 -47269 196 -47235
rect -196 -47275 196 -47269
rect -196 -47343 196 -47337
rect -196 -47377 -184 -47343
rect 184 -47377 196 -47343
rect -196 -47383 196 -47377
rect -252 -47436 -206 -47424
rect -252 -47612 -246 -47436
rect -212 -47612 -206 -47436
rect -252 -47624 -206 -47612
rect 206 -47436 252 -47424
rect 206 -47612 212 -47436
rect 246 -47612 252 -47436
rect 206 -47624 252 -47612
rect -196 -47671 196 -47665
rect -196 -47705 -184 -47671
rect 184 -47705 196 -47671
rect -196 -47711 196 -47705
rect -196 -47779 196 -47773
rect -196 -47813 -184 -47779
rect 184 -47813 196 -47779
rect -196 -47819 196 -47813
rect -252 -47872 -206 -47860
rect -252 -48048 -246 -47872
rect -212 -48048 -206 -47872
rect -252 -48060 -206 -48048
rect 206 -47872 252 -47860
rect 206 -48048 212 -47872
rect 246 -48048 252 -47872
rect 206 -48060 252 -48048
rect -196 -48107 196 -48101
rect -196 -48141 -184 -48107
rect 184 -48141 196 -48107
rect -196 -48147 196 -48141
rect -196 -48215 196 -48209
rect -196 -48249 -184 -48215
rect 184 -48249 196 -48215
rect -196 -48255 196 -48249
rect -252 -48308 -206 -48296
rect -252 -48484 -246 -48308
rect -212 -48484 -206 -48308
rect -252 -48496 -206 -48484
rect 206 -48308 252 -48296
rect 206 -48484 212 -48308
rect 246 -48484 252 -48308
rect 206 -48496 252 -48484
rect -196 -48543 196 -48537
rect -196 -48577 -184 -48543
rect 184 -48577 196 -48543
rect -196 -48583 196 -48577
rect -196 -48651 196 -48645
rect -196 -48685 -184 -48651
rect 184 -48685 196 -48651
rect -196 -48691 196 -48685
rect -252 -48744 -206 -48732
rect -252 -48920 -246 -48744
rect -212 -48920 -206 -48744
rect -252 -48932 -206 -48920
rect 206 -48744 252 -48732
rect 206 -48920 212 -48744
rect 246 -48920 252 -48744
rect 206 -48932 252 -48920
rect -196 -48979 196 -48973
rect -196 -49013 -184 -48979
rect 184 -49013 196 -48979
rect -196 -49019 196 -49013
rect -196 -49087 196 -49081
rect -196 -49121 -184 -49087
rect 184 -49121 196 -49087
rect -196 -49127 196 -49121
rect -252 -49180 -206 -49168
rect -252 -49356 -246 -49180
rect -212 -49356 -206 -49180
rect -252 -49368 -206 -49356
rect 206 -49180 252 -49168
rect 206 -49356 212 -49180
rect 246 -49356 252 -49180
rect 206 -49368 252 -49356
rect -196 -49415 196 -49409
rect -196 -49449 -184 -49415
rect 184 -49449 196 -49415
rect -196 -49455 196 -49449
rect -196 -49523 196 -49517
rect -196 -49557 -184 -49523
rect 184 -49557 196 -49523
rect -196 -49563 196 -49557
rect -252 -49616 -206 -49604
rect -252 -49792 -246 -49616
rect -212 -49792 -206 -49616
rect -252 -49804 -206 -49792
rect 206 -49616 252 -49604
rect 206 -49792 212 -49616
rect 246 -49792 252 -49616
rect 206 -49804 252 -49792
rect -196 -49851 196 -49845
rect -196 -49885 -184 -49851
rect 184 -49885 196 -49851
rect -196 -49891 196 -49885
rect -196 -49959 196 -49953
rect -196 -49993 -184 -49959
rect 184 -49993 196 -49959
rect -196 -49999 196 -49993
rect -252 -50052 -206 -50040
rect -252 -50228 -246 -50052
rect -212 -50228 -206 -50052
rect -252 -50240 -206 -50228
rect 206 -50052 252 -50040
rect 206 -50228 212 -50052
rect 246 -50228 252 -50052
rect 206 -50240 252 -50228
rect -196 -50287 196 -50281
rect -196 -50321 -184 -50287
rect 184 -50321 196 -50287
rect -196 -50327 196 -50321
rect -196 -50395 196 -50389
rect -196 -50429 -184 -50395
rect 184 -50429 196 -50395
rect -196 -50435 196 -50429
rect -252 -50488 -206 -50476
rect -252 -50664 -246 -50488
rect -212 -50664 -206 -50488
rect -252 -50676 -206 -50664
rect 206 -50488 252 -50476
rect 206 -50664 212 -50488
rect 246 -50664 252 -50488
rect 206 -50676 252 -50664
rect -196 -50723 196 -50717
rect -196 -50757 -184 -50723
rect 184 -50757 196 -50723
rect -196 -50763 196 -50757
rect -196 -50831 196 -50825
rect -196 -50865 -184 -50831
rect 184 -50865 196 -50831
rect -196 -50871 196 -50865
rect -252 -50924 -206 -50912
rect -252 -51100 -246 -50924
rect -212 -51100 -206 -50924
rect -252 -51112 -206 -51100
rect 206 -50924 252 -50912
rect 206 -51100 212 -50924
rect 246 -51100 252 -50924
rect 206 -51112 252 -51100
rect -196 -51159 196 -51153
rect -196 -51193 -184 -51159
rect 184 -51193 196 -51159
rect -196 -51199 196 -51193
rect -196 -51267 196 -51261
rect -196 -51301 -184 -51267
rect 184 -51301 196 -51267
rect -196 -51307 196 -51301
rect -252 -51360 -206 -51348
rect -252 -51536 -246 -51360
rect -212 -51536 -206 -51360
rect -252 -51548 -206 -51536
rect 206 -51360 252 -51348
rect 206 -51536 212 -51360
rect 246 -51536 252 -51360
rect 206 -51548 252 -51536
rect -196 -51595 196 -51589
rect -196 -51629 -184 -51595
rect 184 -51629 196 -51595
rect -196 -51635 196 -51629
rect -196 -51703 196 -51697
rect -196 -51737 -184 -51703
rect 184 -51737 196 -51703
rect -196 -51743 196 -51737
rect -252 -51796 -206 -51784
rect -252 -51972 -246 -51796
rect -212 -51972 -206 -51796
rect -252 -51984 -206 -51972
rect 206 -51796 252 -51784
rect 206 -51972 212 -51796
rect 246 -51972 252 -51796
rect 206 -51984 252 -51972
rect -196 -52031 196 -52025
rect -196 -52065 -184 -52031
rect 184 -52065 196 -52031
rect -196 -52071 196 -52065
rect -196 -52139 196 -52133
rect -196 -52173 -184 -52139
rect 184 -52173 196 -52139
rect -196 -52179 196 -52173
rect -252 -52232 -206 -52220
rect -252 -52408 -246 -52232
rect -212 -52408 -206 -52232
rect -252 -52420 -206 -52408
rect 206 -52232 252 -52220
rect 206 -52408 212 -52232
rect 246 -52408 252 -52232
rect 206 -52420 252 -52408
rect -196 -52467 196 -52461
rect -196 -52501 -184 -52467
rect 184 -52501 196 -52467
rect -196 -52507 196 -52501
rect -196 -52575 196 -52569
rect -196 -52609 -184 -52575
rect 184 -52609 196 -52575
rect -196 -52615 196 -52609
rect -252 -52668 -206 -52656
rect -252 -52844 -246 -52668
rect -212 -52844 -206 -52668
rect -252 -52856 -206 -52844
rect 206 -52668 252 -52656
rect 206 -52844 212 -52668
rect 246 -52844 252 -52668
rect 206 -52856 252 -52844
rect -196 -52903 196 -52897
rect -196 -52937 -184 -52903
rect 184 -52937 196 -52903
rect -196 -52943 196 -52937
rect -196 -53011 196 -53005
rect -196 -53045 -184 -53011
rect 184 -53045 196 -53011
rect -196 -53051 196 -53045
rect -252 -53104 -206 -53092
rect -252 -53280 -246 -53104
rect -212 -53280 -206 -53104
rect -252 -53292 -206 -53280
rect 206 -53104 252 -53092
rect 206 -53280 212 -53104
rect 246 -53280 252 -53104
rect 206 -53292 252 -53280
rect -196 -53339 196 -53333
rect -196 -53373 -184 -53339
rect 184 -53373 196 -53339
rect -196 -53379 196 -53373
rect -196 -53447 196 -53441
rect -196 -53481 -184 -53447
rect 184 -53481 196 -53447
rect -196 -53487 196 -53481
rect -252 -53540 -206 -53528
rect -252 -53716 -246 -53540
rect -212 -53716 -206 -53540
rect -252 -53728 -206 -53716
rect 206 -53540 252 -53528
rect 206 -53716 212 -53540
rect 246 -53716 252 -53540
rect 206 -53728 252 -53716
rect -196 -53775 196 -53769
rect -196 -53809 -184 -53775
rect 184 -53809 196 -53775
rect -196 -53815 196 -53809
rect -196 -53883 196 -53877
rect -196 -53917 -184 -53883
rect 184 -53917 196 -53883
rect -196 -53923 196 -53917
rect -252 -53976 -206 -53964
rect -252 -54152 -246 -53976
rect -212 -54152 -206 -53976
rect -252 -54164 -206 -54152
rect 206 -53976 252 -53964
rect 206 -54152 212 -53976
rect 246 -54152 252 -53976
rect 206 -54164 252 -54152
rect -196 -54211 196 -54205
rect -196 -54245 -184 -54211
rect 184 -54245 196 -54211
rect -196 -54251 196 -54245
rect -196 -54319 196 -54313
rect -196 -54353 -184 -54319
rect 184 -54353 196 -54319
rect -196 -54359 196 -54353
rect -252 -54412 -206 -54400
rect -252 -54588 -246 -54412
rect -212 -54588 -206 -54412
rect -252 -54600 -206 -54588
rect 206 -54412 252 -54400
rect 206 -54588 212 -54412
rect 246 -54588 252 -54412
rect 206 -54600 252 -54588
rect -196 -54647 196 -54641
rect -196 -54681 -184 -54647
rect 184 -54681 196 -54647
rect -196 -54687 196 -54681
rect -196 -54755 196 -54749
rect -196 -54789 -184 -54755
rect 184 -54789 196 -54755
rect -196 -54795 196 -54789
rect -252 -54848 -206 -54836
rect -252 -55024 -246 -54848
rect -212 -55024 -206 -54848
rect -252 -55036 -206 -55024
rect 206 -54848 252 -54836
rect 206 -55024 212 -54848
rect 246 -55024 252 -54848
rect 206 -55036 252 -55024
rect -196 -55083 196 -55077
rect -196 -55117 -184 -55083
rect 184 -55117 196 -55083
rect -196 -55123 196 -55117
rect -196 -55191 196 -55185
rect -196 -55225 -184 -55191
rect 184 -55225 196 -55191
rect -196 -55231 196 -55225
rect -252 -55284 -206 -55272
rect -252 -55460 -246 -55284
rect -212 -55460 -206 -55284
rect -252 -55472 -206 -55460
rect 206 -55284 252 -55272
rect 206 -55460 212 -55284
rect 246 -55460 252 -55284
rect 206 -55472 252 -55460
rect -196 -55519 196 -55513
rect -196 -55553 -184 -55519
rect 184 -55553 196 -55519
rect -196 -55559 196 -55553
rect -196 -55627 196 -55621
rect -196 -55661 -184 -55627
rect 184 -55661 196 -55627
rect -196 -55667 196 -55661
rect -252 -55720 -206 -55708
rect -252 -55896 -246 -55720
rect -212 -55896 -206 -55720
rect -252 -55908 -206 -55896
rect 206 -55720 252 -55708
rect 206 -55896 212 -55720
rect 246 -55896 252 -55720
rect 206 -55908 252 -55896
rect -196 -55955 196 -55949
rect -196 -55989 -184 -55955
rect 184 -55989 196 -55955
rect -196 -55995 196 -55989
rect -196 -56063 196 -56057
rect -196 -56097 -184 -56063
rect 184 -56097 196 -56063
rect -196 -56103 196 -56097
rect -252 -56156 -206 -56144
rect -252 -56332 -246 -56156
rect -212 -56332 -206 -56156
rect -252 -56344 -206 -56332
rect 206 -56156 252 -56144
rect 206 -56332 212 -56156
rect 246 -56332 252 -56156
rect 206 -56344 252 -56332
rect -196 -56391 196 -56385
rect -196 -56425 -184 -56391
rect 184 -56425 196 -56391
rect -196 -56431 196 -56425
rect -196 -56499 196 -56493
rect -196 -56533 -184 -56499
rect 184 -56533 196 -56499
rect -196 -56539 196 -56533
rect -252 -56592 -206 -56580
rect -252 -56768 -246 -56592
rect -212 -56768 -206 -56592
rect -252 -56780 -206 -56768
rect 206 -56592 252 -56580
rect 206 -56768 212 -56592
rect 246 -56768 252 -56592
rect 206 -56780 252 -56768
rect -196 -56827 196 -56821
rect -196 -56861 -184 -56827
rect 184 -56861 196 -56827
rect -196 -56867 196 -56861
rect -196 -56935 196 -56929
rect -196 -56969 -184 -56935
rect 184 -56969 196 -56935
rect -196 -56975 196 -56969
rect -252 -57028 -206 -57016
rect -252 -57204 -246 -57028
rect -212 -57204 -206 -57028
rect -252 -57216 -206 -57204
rect 206 -57028 252 -57016
rect 206 -57204 212 -57028
rect 246 -57204 252 -57028
rect 206 -57216 252 -57204
rect -196 -57263 196 -57257
rect -196 -57297 -184 -57263
rect 184 -57297 196 -57263
rect -196 -57303 196 -57297
rect -196 -57371 196 -57365
rect -196 -57405 -184 -57371
rect 184 -57405 196 -57371
rect -196 -57411 196 -57405
rect -252 -57464 -206 -57452
rect -252 -57640 -246 -57464
rect -212 -57640 -206 -57464
rect -252 -57652 -206 -57640
rect 206 -57464 252 -57452
rect 206 -57640 212 -57464
rect 246 -57640 252 -57464
rect 206 -57652 252 -57640
rect -196 -57699 196 -57693
rect -196 -57733 -184 -57699
rect 184 -57733 196 -57699
rect -196 -57739 196 -57733
rect -196 -57807 196 -57801
rect -196 -57841 -184 -57807
rect 184 -57841 196 -57807
rect -196 -57847 196 -57841
rect -252 -57900 -206 -57888
rect -252 -58076 -246 -57900
rect -212 -58076 -206 -57900
rect -252 -58088 -206 -58076
rect 206 -57900 252 -57888
rect 206 -58076 212 -57900
rect 246 -58076 252 -57900
rect 206 -58088 252 -58076
rect -196 -58135 196 -58129
rect -196 -58169 -184 -58135
rect 184 -58169 196 -58135
rect -196 -58175 196 -58169
rect -196 -58243 196 -58237
rect -196 -58277 -184 -58243
rect 184 -58277 196 -58243
rect -196 -58283 196 -58277
rect -252 -58336 -206 -58324
rect -252 -58512 -246 -58336
rect -212 -58512 -206 -58336
rect -252 -58524 -206 -58512
rect 206 -58336 252 -58324
rect 206 -58512 212 -58336
rect 246 -58512 252 -58336
rect 206 -58524 252 -58512
rect -196 -58571 196 -58565
rect -196 -58605 -184 -58571
rect 184 -58605 196 -58571
rect -196 -58611 196 -58605
rect -196 -58679 196 -58673
rect -196 -58713 -184 -58679
rect 184 -58713 196 -58679
rect -196 -58719 196 -58713
rect -252 -58772 -206 -58760
rect -252 -58948 -246 -58772
rect -212 -58948 -206 -58772
rect -252 -58960 -206 -58948
rect 206 -58772 252 -58760
rect 206 -58948 212 -58772
rect 246 -58948 252 -58772
rect 206 -58960 252 -58948
rect -196 -59007 196 -59001
rect -196 -59041 -184 -59007
rect 184 -59041 196 -59007
rect -196 -59047 196 -59041
rect -196 -59115 196 -59109
rect -196 -59149 -184 -59115
rect 184 -59149 196 -59115
rect -196 -59155 196 -59149
rect -252 -59208 -206 -59196
rect -252 -59384 -246 -59208
rect -212 -59384 -206 -59208
rect -252 -59396 -206 -59384
rect 206 -59208 252 -59196
rect 206 -59384 212 -59208
rect 246 -59384 252 -59208
rect 206 -59396 252 -59384
rect -196 -59443 196 -59437
rect -196 -59477 -184 -59443
rect 184 -59477 196 -59443
rect -196 -59483 196 -59477
rect -196 -59551 196 -59545
rect -196 -59585 -184 -59551
rect 184 -59585 196 -59551
rect -196 -59591 196 -59585
rect -252 -59644 -206 -59632
rect -252 -59820 -246 -59644
rect -212 -59820 -206 -59644
rect -252 -59832 -206 -59820
rect 206 -59644 252 -59632
rect 206 -59820 212 -59644
rect 246 -59820 252 -59644
rect 206 -59832 252 -59820
rect -196 -59879 196 -59873
rect -196 -59913 -184 -59879
rect 184 -59913 196 -59879
rect -196 -59919 196 -59913
rect -196 -59987 196 -59981
rect -196 -60021 -184 -59987
rect 184 -60021 196 -59987
rect -196 -60027 196 -60021
rect -252 -60080 -206 -60068
rect -252 -60256 -246 -60080
rect -212 -60256 -206 -60080
rect -252 -60268 -206 -60256
rect 206 -60080 252 -60068
rect 206 -60256 212 -60080
rect 246 -60256 252 -60080
rect 206 -60268 252 -60256
rect -196 -60315 196 -60309
rect -196 -60349 -184 -60315
rect 184 -60349 196 -60315
rect -196 -60355 196 -60349
rect -196 -60423 196 -60417
rect -196 -60457 -184 -60423
rect 184 -60457 196 -60423
rect -196 -60463 196 -60457
rect -252 -60516 -206 -60504
rect -252 -60692 -246 -60516
rect -212 -60692 -206 -60516
rect -252 -60704 -206 -60692
rect 206 -60516 252 -60504
rect 206 -60692 212 -60516
rect 246 -60692 252 -60516
rect 206 -60704 252 -60692
rect -196 -60751 196 -60745
rect -196 -60785 -184 -60751
rect 184 -60785 196 -60751
rect -196 -60791 196 -60785
rect -196 -60859 196 -60853
rect -196 -60893 -184 -60859
rect 184 -60893 196 -60859
rect -196 -60899 196 -60893
rect -252 -60952 -206 -60940
rect -252 -61128 -246 -60952
rect -212 -61128 -206 -60952
rect -252 -61140 -206 -61128
rect 206 -60952 252 -60940
rect 206 -61128 212 -60952
rect 246 -61128 252 -60952
rect 206 -61140 252 -61128
rect -196 -61187 196 -61181
rect -196 -61221 -184 -61187
rect 184 -61221 196 -61187
rect -196 -61227 196 -61221
rect -196 -61295 196 -61289
rect -196 -61329 -184 -61295
rect 184 -61329 196 -61295
rect -196 -61335 196 -61329
rect -252 -61388 -206 -61376
rect -252 -61564 -246 -61388
rect -212 -61564 -206 -61388
rect -252 -61576 -206 -61564
rect 206 -61388 252 -61376
rect 206 -61564 212 -61388
rect 246 -61564 252 -61388
rect 206 -61576 252 -61564
rect -196 -61623 196 -61617
rect -196 -61657 -184 -61623
rect 184 -61657 196 -61623
rect -196 -61663 196 -61657
rect -196 -61731 196 -61725
rect -196 -61765 -184 -61731
rect 184 -61765 196 -61731
rect -196 -61771 196 -61765
rect -252 -61824 -206 -61812
rect -252 -62000 -246 -61824
rect -212 -62000 -206 -61824
rect -252 -62012 -206 -62000
rect 206 -61824 252 -61812
rect 206 -62000 212 -61824
rect 246 -62000 252 -61824
rect 206 -62012 252 -62000
rect -196 -62059 196 -62053
rect -196 -62093 -184 -62059
rect 184 -62093 196 -62059
rect -196 -62099 196 -62093
rect -196 -62167 196 -62161
rect -196 -62201 -184 -62167
rect 184 -62201 196 -62167
rect -196 -62207 196 -62201
rect -252 -62260 -206 -62248
rect -252 -62436 -246 -62260
rect -212 -62436 -206 -62260
rect -252 -62448 -206 -62436
rect 206 -62260 252 -62248
rect 206 -62436 212 -62260
rect 246 -62436 252 -62260
rect 206 -62448 252 -62436
rect -196 -62495 196 -62489
rect -196 -62529 -184 -62495
rect 184 -62529 196 -62495
rect -196 -62535 196 -62529
rect -196 -62603 196 -62597
rect -196 -62637 -184 -62603
rect 184 -62637 196 -62603
rect -196 -62643 196 -62637
rect -252 -62696 -206 -62684
rect -252 -62872 -246 -62696
rect -212 -62872 -206 -62696
rect -252 -62884 -206 -62872
rect 206 -62696 252 -62684
rect 206 -62872 212 -62696
rect 246 -62872 252 -62696
rect 206 -62884 252 -62872
rect -196 -62931 196 -62925
rect -196 -62965 -184 -62931
rect 184 -62965 196 -62931
rect -196 -62971 196 -62965
rect -196 -63039 196 -63033
rect -196 -63073 -184 -63039
rect 184 -63073 196 -63039
rect -196 -63079 196 -63073
rect -252 -63132 -206 -63120
rect -252 -63308 -246 -63132
rect -212 -63308 -206 -63132
rect -252 -63320 -206 -63308
rect 206 -63132 252 -63120
rect 206 -63308 212 -63132
rect 246 -63308 252 -63132
rect 206 -63320 252 -63308
rect -196 -63367 196 -63361
rect -196 -63401 -184 -63367
rect 184 -63401 196 -63367
rect -196 -63407 196 -63401
rect -196 -63475 196 -63469
rect -196 -63509 -184 -63475
rect 184 -63509 196 -63475
rect -196 -63515 196 -63509
rect -252 -63568 -206 -63556
rect -252 -63744 -246 -63568
rect -212 -63744 -206 -63568
rect -252 -63756 -206 -63744
rect 206 -63568 252 -63556
rect 206 -63744 212 -63568
rect 246 -63744 252 -63568
rect 206 -63756 252 -63744
rect -196 -63803 196 -63797
rect -196 -63837 -184 -63803
rect 184 -63837 196 -63803
rect -196 -63843 196 -63837
rect -196 -63911 196 -63905
rect -196 -63945 -184 -63911
rect 184 -63945 196 -63911
rect -196 -63951 196 -63945
rect -252 -64004 -206 -63992
rect -252 -64180 -246 -64004
rect -212 -64180 -206 -64004
rect -252 -64192 -206 -64180
rect 206 -64004 252 -63992
rect 206 -64180 212 -64004
rect 246 -64180 252 -64004
rect 206 -64192 252 -64180
rect -196 -64239 196 -64233
rect -196 -64273 -184 -64239
rect 184 -64273 196 -64239
rect -196 -64279 196 -64273
rect -196 -64347 196 -64341
rect -196 -64381 -184 -64347
rect 184 -64381 196 -64347
rect -196 -64387 196 -64381
rect -252 -64440 -206 -64428
rect -252 -64616 -246 -64440
rect -212 -64616 -206 -64440
rect -252 -64628 -206 -64616
rect 206 -64440 252 -64428
rect 206 -64616 212 -64440
rect 246 -64616 252 -64440
rect 206 -64628 252 -64616
rect -196 -64675 196 -64669
rect -196 -64709 -184 -64675
rect 184 -64709 196 -64675
rect -196 -64715 196 -64709
rect -196 -64783 196 -64777
rect -196 -64817 -184 -64783
rect 184 -64817 196 -64783
rect -196 -64823 196 -64817
rect -252 -64876 -206 -64864
rect -252 -65052 -246 -64876
rect -212 -65052 -206 -64876
rect -252 -65064 -206 -65052
rect 206 -64876 252 -64864
rect 206 -65052 212 -64876
rect 246 -65052 252 -64876
rect 206 -65064 252 -65052
rect -196 -65111 196 -65105
rect -196 -65145 -184 -65111
rect 184 -65145 196 -65111
rect -196 -65151 196 -65145
rect -196 -65219 196 -65213
rect -196 -65253 -184 -65219
rect 184 -65253 196 -65219
rect -196 -65259 196 -65253
rect -252 -65312 -206 -65300
rect -252 -65488 -246 -65312
rect -212 -65488 -206 -65312
rect -252 -65500 -206 -65488
rect 206 -65312 252 -65300
rect 206 -65488 212 -65312
rect 246 -65488 252 -65312
rect 206 -65500 252 -65488
rect -196 -65547 196 -65541
rect -196 -65581 -184 -65547
rect 184 -65581 196 -65547
rect -196 -65587 196 -65581
rect -196 -65655 196 -65649
rect -196 -65689 -184 -65655
rect 184 -65689 196 -65655
rect -196 -65695 196 -65689
rect -252 -65748 -206 -65736
rect -252 -65924 -246 -65748
rect -212 -65924 -206 -65748
rect -252 -65936 -206 -65924
rect 206 -65748 252 -65736
rect 206 -65924 212 -65748
rect 246 -65924 252 -65748
rect 206 -65936 252 -65924
rect -196 -65983 196 -65977
rect -196 -66017 -184 -65983
rect 184 -66017 196 -65983
rect -196 -66023 196 -66017
rect -196 -66091 196 -66085
rect -196 -66125 -184 -66091
rect 184 -66125 196 -66091
rect -196 -66131 196 -66125
rect -252 -66184 -206 -66172
rect -252 -66360 -246 -66184
rect -212 -66360 -206 -66184
rect -252 -66372 -206 -66360
rect 206 -66184 252 -66172
rect 206 -66360 212 -66184
rect 246 -66360 252 -66184
rect 206 -66372 252 -66360
rect -196 -66419 196 -66413
rect -196 -66453 -184 -66419
rect 184 -66453 196 -66419
rect -196 -66459 196 -66453
rect -196 -66527 196 -66521
rect -196 -66561 -184 -66527
rect 184 -66561 196 -66527
rect -196 -66567 196 -66561
rect -252 -66620 -206 -66608
rect -252 -66796 -246 -66620
rect -212 -66796 -206 -66620
rect -252 -66808 -206 -66796
rect 206 -66620 252 -66608
rect 206 -66796 212 -66620
rect 246 -66796 252 -66620
rect 206 -66808 252 -66796
rect -196 -66855 196 -66849
rect -196 -66889 -184 -66855
rect 184 -66889 196 -66855
rect -196 -66895 196 -66889
rect -196 -66963 196 -66957
rect -196 -66997 -184 -66963
rect 184 -66997 196 -66963
rect -196 -67003 196 -66997
rect -252 -67056 -206 -67044
rect -252 -67232 -246 -67056
rect -212 -67232 -206 -67056
rect -252 -67244 -206 -67232
rect 206 -67056 252 -67044
rect 206 -67232 212 -67056
rect 246 -67232 252 -67056
rect 206 -67244 252 -67232
rect -196 -67291 196 -67285
rect -196 -67325 -184 -67291
rect 184 -67325 196 -67291
rect -196 -67331 196 -67325
rect -196 -67399 196 -67393
rect -196 -67433 -184 -67399
rect 184 -67433 196 -67399
rect -196 -67439 196 -67433
rect -252 -67492 -206 -67480
rect -252 -67668 -246 -67492
rect -212 -67668 -206 -67492
rect -252 -67680 -206 -67668
rect 206 -67492 252 -67480
rect 206 -67668 212 -67492
rect 246 -67668 252 -67492
rect 206 -67680 252 -67668
rect -196 -67727 196 -67721
rect -196 -67761 -184 -67727
rect 184 -67761 196 -67727
rect -196 -67767 196 -67761
rect -196 -67835 196 -67829
rect -196 -67869 -184 -67835
rect 184 -67869 196 -67835
rect -196 -67875 196 -67869
rect -252 -67928 -206 -67916
rect -252 -68104 -246 -67928
rect -212 -68104 -206 -67928
rect -252 -68116 -206 -68104
rect 206 -67928 252 -67916
rect 206 -68104 212 -67928
rect 246 -68104 252 -67928
rect 206 -68116 252 -68104
rect -196 -68163 196 -68157
rect -196 -68197 -184 -68163
rect 184 -68197 196 -68163
rect -196 -68203 196 -68197
rect -196 -68271 196 -68265
rect -196 -68305 -184 -68271
rect 184 -68305 196 -68271
rect -196 -68311 196 -68305
rect -252 -68364 -206 -68352
rect -252 -68540 -246 -68364
rect -212 -68540 -206 -68364
rect -252 -68552 -206 -68540
rect 206 -68364 252 -68352
rect 206 -68540 212 -68364
rect 246 -68540 252 -68364
rect 206 -68552 252 -68540
rect -196 -68599 196 -68593
rect -196 -68633 -184 -68599
rect 184 -68633 196 -68599
rect -196 -68639 196 -68633
rect -196 -68707 196 -68701
rect -196 -68741 -184 -68707
rect 184 -68741 196 -68707
rect -196 -68747 196 -68741
rect -252 -68800 -206 -68788
rect -252 -68976 -246 -68800
rect -212 -68976 -206 -68800
rect -252 -68988 -206 -68976
rect 206 -68800 252 -68788
rect 206 -68976 212 -68800
rect 246 -68976 252 -68800
rect 206 -68988 252 -68976
rect -196 -69035 196 -69029
rect -196 -69069 -184 -69035
rect 184 -69069 196 -69035
rect -196 -69075 196 -69069
rect -196 -69143 196 -69137
rect -196 -69177 -184 -69143
rect 184 -69177 196 -69143
rect -196 -69183 196 -69177
rect -252 -69236 -206 -69224
rect -252 -69412 -246 -69236
rect -212 -69412 -206 -69236
rect -252 -69424 -206 -69412
rect 206 -69236 252 -69224
rect 206 -69412 212 -69236
rect 246 -69412 252 -69236
rect 206 -69424 252 -69412
rect -196 -69471 196 -69465
rect -196 -69505 -184 -69471
rect 184 -69505 196 -69471
rect -196 -69511 196 -69505
rect -196 -69579 196 -69573
rect -196 -69613 -184 -69579
rect 184 -69613 196 -69579
rect -196 -69619 196 -69613
rect -252 -69672 -206 -69660
rect -252 -69848 -246 -69672
rect -212 -69848 -206 -69672
rect -252 -69860 -206 -69848
rect 206 -69672 252 -69660
rect 206 -69848 212 -69672
rect 246 -69848 252 -69672
rect 206 -69860 252 -69848
rect -196 -69907 196 -69901
rect -196 -69941 -184 -69907
rect 184 -69941 196 -69907
rect -196 -69947 196 -69941
rect -196 -70015 196 -70009
rect -196 -70049 -184 -70015
rect 184 -70049 196 -70015
rect -196 -70055 196 -70049
rect -252 -70108 -206 -70096
rect -252 -70284 -246 -70108
rect -212 -70284 -206 -70108
rect -252 -70296 -206 -70284
rect 206 -70108 252 -70096
rect 206 -70284 212 -70108
rect 246 -70284 252 -70108
rect 206 -70296 252 -70284
rect -196 -70343 196 -70337
rect -196 -70377 -184 -70343
rect 184 -70377 196 -70343
rect -196 -70383 196 -70377
rect -196 -70451 196 -70445
rect -196 -70485 -184 -70451
rect 184 -70485 196 -70451
rect -196 -70491 196 -70485
rect -252 -70544 -206 -70532
rect -252 -70720 -246 -70544
rect -212 -70720 -206 -70544
rect -252 -70732 -206 -70720
rect 206 -70544 252 -70532
rect 206 -70720 212 -70544
rect 246 -70720 252 -70544
rect 206 -70732 252 -70720
rect -196 -70779 196 -70773
rect -196 -70813 -184 -70779
rect 184 -70813 196 -70779
rect -196 -70819 196 -70813
rect -196 -70887 196 -70881
rect -196 -70921 -184 -70887
rect 184 -70921 196 -70887
rect -196 -70927 196 -70921
rect -252 -70980 -206 -70968
rect -252 -71156 -246 -70980
rect -212 -71156 -206 -70980
rect -252 -71168 -206 -71156
rect 206 -70980 252 -70968
rect 206 -71156 212 -70980
rect 246 -71156 252 -70980
rect 206 -71168 252 -71156
rect -196 -71215 196 -71209
rect -196 -71249 -184 -71215
rect 184 -71249 196 -71215
rect -196 -71255 196 -71249
rect -196 -71323 196 -71317
rect -196 -71357 -184 -71323
rect 184 -71357 196 -71323
rect -196 -71363 196 -71357
rect -252 -71416 -206 -71404
rect -252 -71592 -246 -71416
rect -212 -71592 -206 -71416
rect -252 -71604 -206 -71592
rect 206 -71416 252 -71404
rect 206 -71592 212 -71416
rect 246 -71592 252 -71416
rect 206 -71604 252 -71592
rect -196 -71651 196 -71645
rect -196 -71685 -184 -71651
rect 184 -71685 196 -71651
rect -196 -71691 196 -71685
rect -196 -71759 196 -71753
rect -196 -71793 -184 -71759
rect 184 -71793 196 -71759
rect -196 -71799 196 -71793
rect -252 -71852 -206 -71840
rect -252 -72028 -246 -71852
rect -212 -72028 -206 -71852
rect -252 -72040 -206 -72028
rect 206 -71852 252 -71840
rect 206 -72028 212 -71852
rect 246 -72028 252 -71852
rect 206 -72040 252 -72028
rect -196 -72087 196 -72081
rect -196 -72121 -184 -72087
rect 184 -72121 196 -72087
rect -196 -72127 196 -72121
rect -196 -72195 196 -72189
rect -196 -72229 -184 -72195
rect 184 -72229 196 -72195
rect -196 -72235 196 -72229
rect -252 -72288 -206 -72276
rect -252 -72464 -246 -72288
rect -212 -72464 -206 -72288
rect -252 -72476 -206 -72464
rect 206 -72288 252 -72276
rect 206 -72464 212 -72288
rect 246 -72464 252 -72288
rect 206 -72476 252 -72464
rect -196 -72523 196 -72517
rect -196 -72557 -184 -72523
rect 184 -72557 196 -72523
rect -196 -72563 196 -72557
rect -196 -72631 196 -72625
rect -196 -72665 -184 -72631
rect 184 -72665 196 -72631
rect -196 -72671 196 -72665
rect -252 -72724 -206 -72712
rect -252 -72900 -246 -72724
rect -212 -72900 -206 -72724
rect -252 -72912 -206 -72900
rect 206 -72724 252 -72712
rect 206 -72900 212 -72724
rect 246 -72900 252 -72724
rect 206 -72912 252 -72900
rect -196 -72959 196 -72953
rect -196 -72993 -184 -72959
rect 184 -72993 196 -72959
rect -196 -72999 196 -72993
rect -196 -73067 196 -73061
rect -196 -73101 -184 -73067
rect 184 -73101 196 -73067
rect -196 -73107 196 -73101
rect -252 -73160 -206 -73148
rect -252 -73336 -246 -73160
rect -212 -73336 -206 -73160
rect -252 -73348 -206 -73336
rect 206 -73160 252 -73148
rect 206 -73336 212 -73160
rect 246 -73336 252 -73160
rect 206 -73348 252 -73336
rect -196 -73395 196 -73389
rect -196 -73429 -184 -73395
rect 184 -73429 196 -73395
rect -196 -73435 196 -73429
rect -196 -73503 196 -73497
rect -196 -73537 -184 -73503
rect 184 -73537 196 -73503
rect -196 -73543 196 -73537
rect -252 -73596 -206 -73584
rect -252 -73772 -246 -73596
rect -212 -73772 -206 -73596
rect -252 -73784 -206 -73772
rect 206 -73596 252 -73584
rect 206 -73772 212 -73596
rect 246 -73772 252 -73596
rect 206 -73784 252 -73772
rect -196 -73831 196 -73825
rect -196 -73865 -184 -73831
rect 184 -73865 196 -73831
rect -196 -73871 196 -73865
rect -196 -73939 196 -73933
rect -196 -73973 -184 -73939
rect 184 -73973 196 -73939
rect -196 -73979 196 -73973
rect -252 -74032 -206 -74020
rect -252 -74208 -246 -74032
rect -212 -74208 -206 -74032
rect -252 -74220 -206 -74208
rect 206 -74032 252 -74020
rect 206 -74208 212 -74032
rect 246 -74208 252 -74032
rect 206 -74220 252 -74208
rect -196 -74267 196 -74261
rect -196 -74301 -184 -74267
rect 184 -74301 196 -74267
rect -196 -74307 196 -74301
rect -196 -74375 196 -74369
rect -196 -74409 -184 -74375
rect 184 -74409 196 -74375
rect -196 -74415 196 -74409
rect -252 -74468 -206 -74456
rect -252 -74644 -246 -74468
rect -212 -74644 -206 -74468
rect -252 -74656 -206 -74644
rect 206 -74468 252 -74456
rect 206 -74644 212 -74468
rect 246 -74644 252 -74468
rect 206 -74656 252 -74644
rect -196 -74703 196 -74697
rect -196 -74737 -184 -74703
rect 184 -74737 196 -74703
rect -196 -74743 196 -74737
rect -196 -74811 196 -74805
rect -196 -74845 -184 -74811
rect 184 -74845 196 -74811
rect -196 -74851 196 -74845
rect -252 -74904 -206 -74892
rect -252 -75080 -246 -74904
rect -212 -75080 -206 -74904
rect -252 -75092 -206 -75080
rect 206 -74904 252 -74892
rect 206 -75080 212 -74904
rect 246 -75080 252 -74904
rect 206 -75092 252 -75080
rect -196 -75139 196 -75133
rect -196 -75173 -184 -75139
rect 184 -75173 196 -75139
rect -196 -75179 196 -75173
rect -196 -75247 196 -75241
rect -196 -75281 -184 -75247
rect 184 -75281 196 -75247
rect -196 -75287 196 -75281
rect -252 -75340 -206 -75328
rect -252 -75516 -246 -75340
rect -212 -75516 -206 -75340
rect -252 -75528 -206 -75516
rect 206 -75340 252 -75328
rect 206 -75516 212 -75340
rect 246 -75516 252 -75340
rect 206 -75528 252 -75516
rect -196 -75575 196 -75569
rect -196 -75609 -184 -75575
rect 184 -75609 196 -75575
rect -196 -75615 196 -75609
rect -196 -75683 196 -75677
rect -196 -75717 -184 -75683
rect 184 -75717 196 -75683
rect -196 -75723 196 -75717
rect -252 -75776 -206 -75764
rect -252 -75952 -246 -75776
rect -212 -75952 -206 -75776
rect -252 -75964 -206 -75952
rect 206 -75776 252 -75764
rect 206 -75952 212 -75776
rect 246 -75952 252 -75776
rect 206 -75964 252 -75952
rect -196 -76011 196 -76005
rect -196 -76045 -184 -76011
rect 184 -76045 196 -76011
rect -196 -76051 196 -76045
rect -196 -76119 196 -76113
rect -196 -76153 -184 -76119
rect 184 -76153 196 -76119
rect -196 -76159 196 -76153
rect -252 -76212 -206 -76200
rect -252 -76388 -246 -76212
rect -212 -76388 -206 -76212
rect -252 -76400 -206 -76388
rect 206 -76212 252 -76200
rect 206 -76388 212 -76212
rect 246 -76388 252 -76212
rect 206 -76400 252 -76388
rect -196 -76447 196 -76441
rect -196 -76481 -184 -76447
rect 184 -76481 196 -76447
rect -196 -76487 196 -76481
rect -196 -76555 196 -76549
rect -196 -76589 -184 -76555
rect 184 -76589 196 -76555
rect -196 -76595 196 -76589
rect -252 -76648 -206 -76636
rect -252 -76824 -246 -76648
rect -212 -76824 -206 -76648
rect -252 -76836 -206 -76824
rect 206 -76648 252 -76636
rect 206 -76824 212 -76648
rect 246 -76824 252 -76648
rect 206 -76836 252 -76824
rect -196 -76883 196 -76877
rect -196 -76917 -184 -76883
rect 184 -76917 196 -76883
rect -196 -76923 196 -76917
rect -196 -76991 196 -76985
rect -196 -77025 -184 -76991
rect 184 -77025 196 -76991
rect -196 -77031 196 -77025
rect -252 -77084 -206 -77072
rect -252 -77260 -246 -77084
rect -212 -77260 -206 -77084
rect -252 -77272 -206 -77260
rect 206 -77084 252 -77072
rect 206 -77260 212 -77084
rect 246 -77260 252 -77084
rect 206 -77272 252 -77260
rect -196 -77319 196 -77313
rect -196 -77353 -184 -77319
rect 184 -77353 196 -77319
rect -196 -77359 196 -77353
rect -196 -77427 196 -77421
rect -196 -77461 -184 -77427
rect 184 -77461 196 -77427
rect -196 -77467 196 -77461
rect -252 -77520 -206 -77508
rect -252 -77696 -246 -77520
rect -212 -77696 -206 -77520
rect -252 -77708 -206 -77696
rect 206 -77520 252 -77508
rect 206 -77696 212 -77520
rect 246 -77696 252 -77520
rect 206 -77708 252 -77696
rect -196 -77755 196 -77749
rect -196 -77789 -184 -77755
rect 184 -77789 196 -77755
rect -196 -77795 196 -77789
rect -196 -77863 196 -77857
rect -196 -77897 -184 -77863
rect 184 -77897 196 -77863
rect -196 -77903 196 -77897
rect -252 -77956 -206 -77944
rect -252 -78132 -246 -77956
rect -212 -78132 -206 -77956
rect -252 -78144 -206 -78132
rect 206 -77956 252 -77944
rect 206 -78132 212 -77956
rect 246 -78132 252 -77956
rect 206 -78144 252 -78132
rect -196 -78191 196 -78185
rect -196 -78225 -184 -78191
rect 184 -78225 196 -78191
rect -196 -78231 196 -78225
rect -196 -78299 196 -78293
rect -196 -78333 -184 -78299
rect 184 -78333 196 -78299
rect -196 -78339 196 -78333
rect -252 -78392 -206 -78380
rect -252 -78568 -246 -78392
rect -212 -78568 -206 -78392
rect -252 -78580 -206 -78568
rect 206 -78392 252 -78380
rect 206 -78568 212 -78392
rect 246 -78568 252 -78392
rect 206 -78580 252 -78568
rect -196 -78627 196 -78621
rect -196 -78661 -184 -78627
rect 184 -78661 196 -78627
rect -196 -78667 196 -78661
rect -196 -78735 196 -78729
rect -196 -78769 -184 -78735
rect 184 -78769 196 -78735
rect -196 -78775 196 -78769
rect -252 -78828 -206 -78816
rect -252 -79004 -246 -78828
rect -212 -79004 -206 -78828
rect -252 -79016 -206 -79004
rect 206 -78828 252 -78816
rect 206 -79004 212 -78828
rect 246 -79004 252 -78828
rect 206 -79016 252 -79004
rect -196 -79063 196 -79057
rect -196 -79097 -184 -79063
rect 184 -79097 196 -79063
rect -196 -79103 196 -79097
rect -196 -79171 196 -79165
rect -196 -79205 -184 -79171
rect 184 -79205 196 -79171
rect -196 -79211 196 -79205
rect -252 -79264 -206 -79252
rect -252 -79440 -246 -79264
rect -212 -79440 -206 -79264
rect -252 -79452 -206 -79440
rect 206 -79264 252 -79252
rect 206 -79440 212 -79264
rect 246 -79440 252 -79264
rect 206 -79452 252 -79440
rect -196 -79499 196 -79493
rect -196 -79533 -184 -79499
rect 184 -79533 196 -79499
rect -196 -79539 196 -79533
rect -196 -79607 196 -79601
rect -196 -79641 -184 -79607
rect 184 -79641 196 -79607
rect -196 -79647 196 -79641
rect -252 -79700 -206 -79688
rect -252 -79876 -246 -79700
rect -212 -79876 -206 -79700
rect -252 -79888 -206 -79876
rect 206 -79700 252 -79688
rect 206 -79876 212 -79700
rect 246 -79876 252 -79700
rect 206 -79888 252 -79876
rect -196 -79935 196 -79929
rect -196 -79969 -184 -79935
rect 184 -79969 196 -79935
rect -196 -79975 196 -79969
rect -196 -80043 196 -80037
rect -196 -80077 -184 -80043
rect 184 -80077 196 -80043
rect -196 -80083 196 -80077
rect -252 -80136 -206 -80124
rect -252 -80312 -246 -80136
rect -212 -80312 -206 -80136
rect -252 -80324 -206 -80312
rect 206 -80136 252 -80124
rect 206 -80312 212 -80136
rect 246 -80312 252 -80136
rect 206 -80324 252 -80312
rect -196 -80371 196 -80365
rect -196 -80405 -184 -80371
rect 184 -80405 196 -80371
rect -196 -80411 196 -80405
rect -196 -80479 196 -80473
rect -196 -80513 -184 -80479
rect 184 -80513 196 -80479
rect -196 -80519 196 -80513
rect -252 -80572 -206 -80560
rect -252 -80748 -246 -80572
rect -212 -80748 -206 -80572
rect -252 -80760 -206 -80748
rect 206 -80572 252 -80560
rect 206 -80748 212 -80572
rect 246 -80748 252 -80572
rect 206 -80760 252 -80748
rect -196 -80807 196 -80801
rect -196 -80841 -184 -80807
rect 184 -80841 196 -80807
rect -196 -80847 196 -80841
rect -196 -80915 196 -80909
rect -196 -80949 -184 -80915
rect 184 -80949 196 -80915
rect -196 -80955 196 -80949
rect -252 -81008 -206 -80996
rect -252 -81184 -246 -81008
rect -212 -81184 -206 -81008
rect -252 -81196 -206 -81184
rect 206 -81008 252 -80996
rect 206 -81184 212 -81008
rect 246 -81184 252 -81008
rect 206 -81196 252 -81184
rect -196 -81243 196 -81237
rect -196 -81277 -184 -81243
rect 184 -81277 196 -81243
rect -196 -81283 196 -81277
rect -196 -81351 196 -81345
rect -196 -81385 -184 -81351
rect 184 -81385 196 -81351
rect -196 -81391 196 -81385
rect -252 -81444 -206 -81432
rect -252 -81620 -246 -81444
rect -212 -81620 -206 -81444
rect -252 -81632 -206 -81620
rect 206 -81444 252 -81432
rect 206 -81620 212 -81444
rect 246 -81620 252 -81444
rect 206 -81632 252 -81620
rect -196 -81679 196 -81673
rect -196 -81713 -184 -81679
rect 184 -81713 196 -81679
rect -196 -81719 196 -81713
rect -196 -81787 196 -81781
rect -196 -81821 -184 -81787
rect 184 -81821 196 -81787
rect -196 -81827 196 -81821
rect -252 -81880 -206 -81868
rect -252 -82056 -246 -81880
rect -212 -82056 -206 -81880
rect -252 -82068 -206 -82056
rect 206 -81880 252 -81868
rect 206 -82056 212 -81880
rect 246 -82056 252 -81880
rect 206 -82068 252 -82056
rect -196 -82115 196 -82109
rect -196 -82149 -184 -82115
rect 184 -82149 196 -82115
rect -196 -82155 196 -82149
rect -196 -82223 196 -82217
rect -196 -82257 -184 -82223
rect 184 -82257 196 -82223
rect -196 -82263 196 -82257
rect -252 -82316 -206 -82304
rect -252 -82492 -246 -82316
rect -212 -82492 -206 -82316
rect -252 -82504 -206 -82492
rect 206 -82316 252 -82304
rect 206 -82492 212 -82316
rect 246 -82492 252 -82316
rect 206 -82504 252 -82492
rect -196 -82551 196 -82545
rect -196 -82585 -184 -82551
rect 184 -82585 196 -82551
rect -196 -82591 196 -82585
rect -196 -82659 196 -82653
rect -196 -82693 -184 -82659
rect 184 -82693 196 -82659
rect -196 -82699 196 -82693
rect -252 -82752 -206 -82740
rect -252 -82928 -246 -82752
rect -212 -82928 -206 -82752
rect -252 -82940 -206 -82928
rect 206 -82752 252 -82740
rect 206 -82928 212 -82752
rect 246 -82928 252 -82752
rect 206 -82940 252 -82928
rect -196 -82987 196 -82981
rect -196 -83021 -184 -82987
rect 184 -83021 196 -82987
rect -196 -83027 196 -83021
rect -196 -83095 196 -83089
rect -196 -83129 -184 -83095
rect 184 -83129 196 -83095
rect -196 -83135 196 -83129
rect -252 -83188 -206 -83176
rect -252 -83364 -246 -83188
rect -212 -83364 -206 -83188
rect -252 -83376 -206 -83364
rect 206 -83188 252 -83176
rect 206 -83364 212 -83188
rect 246 -83364 252 -83188
rect 206 -83376 252 -83364
rect -196 -83423 196 -83417
rect -196 -83457 -184 -83423
rect 184 -83457 196 -83423
rect -196 -83463 196 -83457
rect -196 -83531 196 -83525
rect -196 -83565 -184 -83531
rect 184 -83565 196 -83531
rect -196 -83571 196 -83565
rect -252 -83624 -206 -83612
rect -252 -83800 -246 -83624
rect -212 -83800 -206 -83624
rect -252 -83812 -206 -83800
rect 206 -83624 252 -83612
rect 206 -83800 212 -83624
rect 246 -83800 252 -83624
rect 206 -83812 252 -83800
rect -196 -83859 196 -83853
rect -196 -83893 -184 -83859
rect 184 -83893 196 -83859
rect -196 -83899 196 -83893
rect -196 -83967 196 -83961
rect -196 -84001 -184 -83967
rect 184 -84001 196 -83967
rect -196 -84007 196 -84001
rect -252 -84060 -206 -84048
rect -252 -84236 -246 -84060
rect -212 -84236 -206 -84060
rect -252 -84248 -206 -84236
rect 206 -84060 252 -84048
rect 206 -84236 212 -84060
rect 246 -84236 252 -84060
rect 206 -84248 252 -84236
rect -196 -84295 196 -84289
rect -196 -84329 -184 -84295
rect 184 -84329 196 -84295
rect -196 -84335 196 -84329
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -343 -84414 343 84414
string parameters w 1 l 2 m 387 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
