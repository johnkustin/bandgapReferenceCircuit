magic
tech sky130A
magscale 1 2
timestamp 1622081478
<< nwell >>
rect -1101 -497 1101 497
<< mvpmos >>
rect -843 -200 -683 200
rect -625 -200 -465 200
rect -407 -200 -247 200
rect -189 -200 -29 200
rect 29 -200 189 200
rect 247 -200 407 200
rect 465 -200 625 200
rect 683 -200 843 200
<< mvpdiff >>
rect -901 187 -843 200
rect -901 153 -889 187
rect -855 153 -843 187
rect -901 119 -843 153
rect -901 85 -889 119
rect -855 85 -843 119
rect -901 51 -843 85
rect -901 17 -889 51
rect -855 17 -843 51
rect -901 -17 -843 17
rect -901 -51 -889 -17
rect -855 -51 -843 -17
rect -901 -85 -843 -51
rect -901 -119 -889 -85
rect -855 -119 -843 -85
rect -901 -153 -843 -119
rect -901 -187 -889 -153
rect -855 -187 -843 -153
rect -901 -200 -843 -187
rect -683 187 -625 200
rect -683 153 -671 187
rect -637 153 -625 187
rect -683 119 -625 153
rect -683 85 -671 119
rect -637 85 -625 119
rect -683 51 -625 85
rect -683 17 -671 51
rect -637 17 -625 51
rect -683 -17 -625 17
rect -683 -51 -671 -17
rect -637 -51 -625 -17
rect -683 -85 -625 -51
rect -683 -119 -671 -85
rect -637 -119 -625 -85
rect -683 -153 -625 -119
rect -683 -187 -671 -153
rect -637 -187 -625 -153
rect -683 -200 -625 -187
rect -465 187 -407 200
rect -465 153 -453 187
rect -419 153 -407 187
rect -465 119 -407 153
rect -465 85 -453 119
rect -419 85 -407 119
rect -465 51 -407 85
rect -465 17 -453 51
rect -419 17 -407 51
rect -465 -17 -407 17
rect -465 -51 -453 -17
rect -419 -51 -407 -17
rect -465 -85 -407 -51
rect -465 -119 -453 -85
rect -419 -119 -407 -85
rect -465 -153 -407 -119
rect -465 -187 -453 -153
rect -419 -187 -407 -153
rect -465 -200 -407 -187
rect -247 187 -189 200
rect -247 153 -235 187
rect -201 153 -189 187
rect -247 119 -189 153
rect -247 85 -235 119
rect -201 85 -189 119
rect -247 51 -189 85
rect -247 17 -235 51
rect -201 17 -189 51
rect -247 -17 -189 17
rect -247 -51 -235 -17
rect -201 -51 -189 -17
rect -247 -85 -189 -51
rect -247 -119 -235 -85
rect -201 -119 -189 -85
rect -247 -153 -189 -119
rect -247 -187 -235 -153
rect -201 -187 -189 -153
rect -247 -200 -189 -187
rect -29 187 29 200
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -200 29 -187
rect 189 187 247 200
rect 189 153 201 187
rect 235 153 247 187
rect 189 119 247 153
rect 189 85 201 119
rect 235 85 247 119
rect 189 51 247 85
rect 189 17 201 51
rect 235 17 247 51
rect 189 -17 247 17
rect 189 -51 201 -17
rect 235 -51 247 -17
rect 189 -85 247 -51
rect 189 -119 201 -85
rect 235 -119 247 -85
rect 189 -153 247 -119
rect 189 -187 201 -153
rect 235 -187 247 -153
rect 189 -200 247 -187
rect 407 187 465 200
rect 407 153 419 187
rect 453 153 465 187
rect 407 119 465 153
rect 407 85 419 119
rect 453 85 465 119
rect 407 51 465 85
rect 407 17 419 51
rect 453 17 465 51
rect 407 -17 465 17
rect 407 -51 419 -17
rect 453 -51 465 -17
rect 407 -85 465 -51
rect 407 -119 419 -85
rect 453 -119 465 -85
rect 407 -153 465 -119
rect 407 -187 419 -153
rect 453 -187 465 -153
rect 407 -200 465 -187
rect 625 187 683 200
rect 625 153 637 187
rect 671 153 683 187
rect 625 119 683 153
rect 625 85 637 119
rect 671 85 683 119
rect 625 51 683 85
rect 625 17 637 51
rect 671 17 683 51
rect 625 -17 683 17
rect 625 -51 637 -17
rect 671 -51 683 -17
rect 625 -85 683 -51
rect 625 -119 637 -85
rect 671 -119 683 -85
rect 625 -153 683 -119
rect 625 -187 637 -153
rect 671 -187 683 -153
rect 625 -200 683 -187
rect 843 187 901 200
rect 843 153 855 187
rect 889 153 901 187
rect 843 119 901 153
rect 843 85 855 119
rect 889 85 901 119
rect 843 51 901 85
rect 843 17 855 51
rect 889 17 901 51
rect 843 -17 901 17
rect 843 -51 855 -17
rect 889 -51 901 -17
rect 843 -85 901 -51
rect 843 -119 855 -85
rect 889 -119 901 -85
rect 843 -153 901 -119
rect 843 -187 855 -153
rect 889 -187 901 -153
rect 843 -200 901 -187
<< mvpdiffc >>
rect -889 153 -855 187
rect -889 85 -855 119
rect -889 17 -855 51
rect -889 -51 -855 -17
rect -889 -119 -855 -85
rect -889 -187 -855 -153
rect -671 153 -637 187
rect -671 85 -637 119
rect -671 17 -637 51
rect -671 -51 -637 -17
rect -671 -119 -637 -85
rect -671 -187 -637 -153
rect -453 153 -419 187
rect -453 85 -419 119
rect -453 17 -419 51
rect -453 -51 -419 -17
rect -453 -119 -419 -85
rect -453 -187 -419 -153
rect -235 153 -201 187
rect -235 85 -201 119
rect -235 17 -201 51
rect -235 -51 -201 -17
rect -235 -119 -201 -85
rect -235 -187 -201 -153
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect 201 153 235 187
rect 201 85 235 119
rect 201 17 235 51
rect 201 -51 235 -17
rect 201 -119 235 -85
rect 201 -187 235 -153
rect 419 153 453 187
rect 419 85 453 119
rect 419 17 453 51
rect 419 -51 453 -17
rect 419 -119 453 -85
rect 419 -187 453 -153
rect 637 153 671 187
rect 637 85 671 119
rect 637 17 671 51
rect 637 -51 671 -17
rect 637 -119 671 -85
rect 637 -187 671 -153
rect 855 153 889 187
rect 855 85 889 119
rect 855 17 889 51
rect 855 -51 889 -17
rect 855 -119 889 -85
rect 855 -187 889 -153
<< mvnsubdiff >>
rect -1035 419 1035 431
rect -1035 385 -901 419
rect -867 385 -833 419
rect -799 385 -765 419
rect -731 385 -697 419
rect -663 385 -629 419
rect -595 385 -561 419
rect -527 385 -493 419
rect -459 385 -425 419
rect -391 385 -357 419
rect -323 385 -289 419
rect -255 385 -221 419
rect -187 385 -153 419
rect -119 385 -85 419
rect -51 385 -17 419
rect 17 385 51 419
rect 85 385 119 419
rect 153 385 187 419
rect 221 385 255 419
rect 289 385 323 419
rect 357 385 391 419
rect 425 385 459 419
rect 493 385 527 419
rect 561 385 595 419
rect 629 385 663 419
rect 697 385 731 419
rect 765 385 799 419
rect 833 385 867 419
rect 901 385 1035 419
rect -1035 373 1035 385
rect -1035 323 -977 373
rect -1035 289 -1023 323
rect -989 289 -977 323
rect 977 323 1035 373
rect -1035 255 -977 289
rect -1035 221 -1023 255
rect -989 221 -977 255
rect -1035 187 -977 221
rect 977 289 989 323
rect 1023 289 1035 323
rect 977 255 1035 289
rect 977 221 989 255
rect 1023 221 1035 255
rect -1035 153 -1023 187
rect -989 153 -977 187
rect -1035 119 -977 153
rect -1035 85 -1023 119
rect -989 85 -977 119
rect -1035 51 -977 85
rect -1035 17 -1023 51
rect -989 17 -977 51
rect -1035 -17 -977 17
rect -1035 -51 -1023 -17
rect -989 -51 -977 -17
rect -1035 -85 -977 -51
rect -1035 -119 -1023 -85
rect -989 -119 -977 -85
rect -1035 -153 -977 -119
rect -1035 -187 -1023 -153
rect -989 -187 -977 -153
rect -1035 -221 -977 -187
rect 977 187 1035 221
rect 977 153 989 187
rect 1023 153 1035 187
rect 977 119 1035 153
rect 977 85 989 119
rect 1023 85 1035 119
rect 977 51 1035 85
rect 977 17 989 51
rect 1023 17 1035 51
rect 977 -17 1035 17
rect 977 -51 989 -17
rect 1023 -51 1035 -17
rect 977 -85 1035 -51
rect 977 -119 989 -85
rect 1023 -119 1035 -85
rect 977 -153 1035 -119
rect 977 -187 989 -153
rect 1023 -187 1035 -153
rect -1035 -255 -1023 -221
rect -989 -255 -977 -221
rect -1035 -289 -977 -255
rect -1035 -323 -1023 -289
rect -989 -323 -977 -289
rect 977 -221 1035 -187
rect 977 -255 989 -221
rect 1023 -255 1035 -221
rect 977 -289 1035 -255
rect -1035 -373 -977 -323
rect 977 -323 989 -289
rect 1023 -323 1035 -289
rect 977 -373 1035 -323
rect -1035 -385 1035 -373
rect -1035 -419 -901 -385
rect -867 -419 -833 -385
rect -799 -419 -765 -385
rect -731 -419 -697 -385
rect -663 -419 -629 -385
rect -595 -419 -561 -385
rect -527 -419 -493 -385
rect -459 -419 -425 -385
rect -391 -419 -357 -385
rect -323 -419 -289 -385
rect -255 -419 -221 -385
rect -187 -419 -153 -385
rect -119 -419 -85 -385
rect -51 -419 -17 -385
rect 17 -419 51 -385
rect 85 -419 119 -385
rect 153 -419 187 -385
rect 221 -419 255 -385
rect 289 -419 323 -385
rect 357 -419 391 -385
rect 425 -419 459 -385
rect 493 -419 527 -385
rect 561 -419 595 -385
rect 629 -419 663 -385
rect 697 -419 731 -385
rect 765 -419 799 -385
rect 833 -419 867 -385
rect 901 -419 1035 -385
rect -1035 -431 1035 -419
<< mvnsubdiffcont >>
rect -901 385 -867 419
rect -833 385 -799 419
rect -765 385 -731 419
rect -697 385 -663 419
rect -629 385 -595 419
rect -561 385 -527 419
rect -493 385 -459 419
rect -425 385 -391 419
rect -357 385 -323 419
rect -289 385 -255 419
rect -221 385 -187 419
rect -153 385 -119 419
rect -85 385 -51 419
rect -17 385 17 419
rect 51 385 85 419
rect 119 385 153 419
rect 187 385 221 419
rect 255 385 289 419
rect 323 385 357 419
rect 391 385 425 419
rect 459 385 493 419
rect 527 385 561 419
rect 595 385 629 419
rect 663 385 697 419
rect 731 385 765 419
rect 799 385 833 419
rect 867 385 901 419
rect -1023 289 -989 323
rect -1023 221 -989 255
rect 989 289 1023 323
rect 989 221 1023 255
rect -1023 153 -989 187
rect -1023 85 -989 119
rect -1023 17 -989 51
rect -1023 -51 -989 -17
rect -1023 -119 -989 -85
rect -1023 -187 -989 -153
rect 989 153 1023 187
rect 989 85 1023 119
rect 989 17 1023 51
rect 989 -51 1023 -17
rect 989 -119 1023 -85
rect 989 -187 1023 -153
rect -1023 -255 -989 -221
rect -1023 -323 -989 -289
rect 989 -255 1023 -221
rect 989 -323 1023 -289
rect -901 -419 -867 -385
rect -833 -419 -799 -385
rect -765 -419 -731 -385
rect -697 -419 -663 -385
rect -629 -419 -595 -385
rect -561 -419 -527 -385
rect -493 -419 -459 -385
rect -425 -419 -391 -385
rect -357 -419 -323 -385
rect -289 -419 -255 -385
rect -221 -419 -187 -385
rect -153 -419 -119 -385
rect -85 -419 -51 -385
rect -17 -419 17 -385
rect 51 -419 85 -385
rect 119 -419 153 -385
rect 187 -419 221 -385
rect 255 -419 289 -385
rect 323 -419 357 -385
rect 391 -419 425 -385
rect 459 -419 493 -385
rect 527 -419 561 -385
rect 595 -419 629 -385
rect 663 -419 697 -385
rect 731 -419 765 -385
rect 799 -419 833 -385
rect 867 -419 901 -385
<< poly >>
rect -843 281 -683 297
rect -843 247 -814 281
rect -780 247 -746 281
rect -712 247 -683 281
rect -843 200 -683 247
rect -625 281 -465 297
rect -625 247 -596 281
rect -562 247 -528 281
rect -494 247 -465 281
rect -625 200 -465 247
rect -407 281 -247 297
rect -407 247 -378 281
rect -344 247 -310 281
rect -276 247 -247 281
rect -407 200 -247 247
rect -189 281 -29 297
rect -189 247 -160 281
rect -126 247 -92 281
rect -58 247 -29 281
rect -189 200 -29 247
rect 29 281 189 297
rect 29 247 58 281
rect 92 247 126 281
rect 160 247 189 281
rect 29 200 189 247
rect 247 281 407 297
rect 247 247 276 281
rect 310 247 344 281
rect 378 247 407 281
rect 247 200 407 247
rect 465 281 625 297
rect 465 247 494 281
rect 528 247 562 281
rect 596 247 625 281
rect 465 200 625 247
rect 683 281 843 297
rect 683 247 712 281
rect 746 247 780 281
rect 814 247 843 281
rect 683 200 843 247
rect -843 -247 -683 -200
rect -843 -281 -814 -247
rect -780 -281 -746 -247
rect -712 -281 -683 -247
rect -843 -297 -683 -281
rect -625 -247 -465 -200
rect -625 -281 -596 -247
rect -562 -281 -528 -247
rect -494 -281 -465 -247
rect -625 -297 -465 -281
rect -407 -247 -247 -200
rect -407 -281 -378 -247
rect -344 -281 -310 -247
rect -276 -281 -247 -247
rect -407 -297 -247 -281
rect -189 -247 -29 -200
rect -189 -281 -160 -247
rect -126 -281 -92 -247
rect -58 -281 -29 -247
rect -189 -297 -29 -281
rect 29 -247 189 -200
rect 29 -281 58 -247
rect 92 -281 126 -247
rect 160 -281 189 -247
rect 29 -297 189 -281
rect 247 -247 407 -200
rect 247 -281 276 -247
rect 310 -281 344 -247
rect 378 -281 407 -247
rect 247 -297 407 -281
rect 465 -247 625 -200
rect 465 -281 494 -247
rect 528 -281 562 -247
rect 596 -281 625 -247
rect 465 -297 625 -281
rect 683 -247 843 -200
rect 683 -281 712 -247
rect 746 -281 780 -247
rect 814 -281 843 -247
rect 683 -297 843 -281
<< polycont >>
rect -814 247 -780 281
rect -746 247 -712 281
rect -596 247 -562 281
rect -528 247 -494 281
rect -378 247 -344 281
rect -310 247 -276 281
rect -160 247 -126 281
rect -92 247 -58 281
rect 58 247 92 281
rect 126 247 160 281
rect 276 247 310 281
rect 344 247 378 281
rect 494 247 528 281
rect 562 247 596 281
rect 712 247 746 281
rect 780 247 814 281
rect -814 -281 -780 -247
rect -746 -281 -712 -247
rect -596 -281 -562 -247
rect -528 -281 -494 -247
rect -378 -281 -344 -247
rect -310 -281 -276 -247
rect -160 -281 -126 -247
rect -92 -281 -58 -247
rect 58 -281 92 -247
rect 126 -281 160 -247
rect 276 -281 310 -247
rect 344 -281 378 -247
rect 494 -281 528 -247
rect 562 -281 596 -247
rect 712 -281 746 -247
rect 780 -281 814 -247
<< locali >>
rect -1023 385 -901 419
rect -847 385 -833 419
rect -775 385 -765 419
rect -703 385 -697 419
rect -631 385 -629 419
rect -595 385 -593 419
rect -527 385 -521 419
rect -459 385 -449 419
rect -391 385 -377 419
rect -323 385 -305 419
rect -255 385 -233 419
rect -187 385 -161 419
rect -119 385 -89 419
rect -51 385 -17 419
rect 17 385 51 419
rect 89 385 119 419
rect 161 385 187 419
rect 233 385 255 419
rect 305 385 323 419
rect 377 385 391 419
rect 449 385 459 419
rect 521 385 527 419
rect 593 385 595 419
rect 629 385 631 419
rect 697 385 703 419
rect 765 385 775 419
rect 833 385 847 419
rect 901 385 1023 419
rect -1023 353 -989 385
rect -1023 281 -989 289
rect 989 323 1023 385
rect -843 247 -816 281
rect -780 247 -746 281
rect -710 247 -683 281
rect -625 247 -598 281
rect -562 247 -528 281
rect -492 247 -465 281
rect -407 247 -380 281
rect -344 247 -310 281
rect -274 247 -247 281
rect -189 247 -162 281
rect -126 247 -92 281
rect -56 247 -29 281
rect 29 247 56 281
rect 92 247 126 281
rect 162 247 189 281
rect 247 247 274 281
rect 310 247 344 281
rect 380 247 407 281
rect 465 247 492 281
rect 528 247 562 281
rect 598 247 625 281
rect 683 247 710 281
rect 746 247 780 281
rect 816 247 843 281
rect 989 255 1023 289
rect -1023 209 -989 221
rect -1023 137 -989 153
rect -1023 65 -989 85
rect -1023 -17 -989 17
rect -1023 -85 -989 -51
rect -1023 -153 -989 -119
rect -1023 -221 -989 -187
rect -889 187 -855 204
rect -889 149 -855 153
rect -889 77 -855 85
rect -889 -17 -855 17
rect -889 -85 -855 -51
rect -889 -153 -855 -119
rect -889 -204 -855 -187
rect -671 187 -637 204
rect -671 119 -637 153
rect -671 51 -637 85
rect -671 -17 -637 17
rect -671 -85 -637 -77
rect -671 -153 -637 -149
rect -671 -204 -637 -187
rect -453 187 -419 204
rect -453 149 -419 153
rect -453 77 -419 85
rect -453 -17 -419 17
rect -453 -85 -419 -51
rect -453 -153 -419 -119
rect -453 -204 -419 -187
rect -235 187 -201 204
rect -235 119 -201 153
rect -235 51 -201 85
rect -235 -17 -201 17
rect -235 -85 -201 -77
rect -235 -153 -201 -149
rect -235 -204 -201 -187
rect -17 187 17 204
rect -17 149 17 153
rect -17 77 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -204 17 -187
rect 201 187 235 204
rect 201 119 235 153
rect 201 51 235 85
rect 201 -17 235 17
rect 201 -85 235 -77
rect 201 -153 235 -149
rect 201 -204 235 -187
rect 419 187 453 204
rect 419 149 453 153
rect 419 77 453 85
rect 419 -17 453 17
rect 419 -85 453 -51
rect 419 -153 453 -119
rect 419 -204 453 -187
rect 637 187 671 204
rect 637 119 671 153
rect 637 51 671 85
rect 637 -17 671 17
rect 637 -85 671 -77
rect 637 -153 671 -149
rect 637 -204 671 -187
rect 855 187 889 204
rect 855 149 889 153
rect 855 77 889 85
rect 855 -17 889 17
rect 855 -85 889 -51
rect 855 -153 889 -119
rect 855 -204 889 -187
rect 989 187 1023 221
rect 989 119 1023 153
rect 989 51 1023 85
rect 989 -17 1023 17
rect 989 -85 1023 -51
rect 989 -153 1023 -119
rect 989 -221 1023 -187
rect -1023 -289 -989 -255
rect -843 -281 -816 -247
rect -780 -281 -746 -247
rect -710 -281 -683 -247
rect -625 -281 -598 -247
rect -562 -281 -528 -247
rect -492 -281 -465 -247
rect -407 -281 -380 -247
rect -344 -281 -310 -247
rect -274 -281 -247 -247
rect -189 -281 -162 -247
rect -126 -281 -92 -247
rect -56 -281 -29 -247
rect 29 -281 56 -247
rect 92 -281 126 -247
rect 162 -281 189 -247
rect 247 -281 274 -247
rect 310 -281 344 -247
rect 380 -281 407 -247
rect 465 -281 492 -247
rect 528 -281 562 -247
rect 598 -281 625 -247
rect 683 -281 710 -247
rect 746 -281 780 -247
rect 816 -281 843 -247
rect -1023 -385 -989 -323
rect 989 -289 1023 -255
rect 989 -385 1023 -323
rect -1023 -419 -901 -385
rect -867 -419 -833 -385
rect -799 -419 -765 -385
rect -731 -419 -697 -385
rect -663 -419 -629 -385
rect -595 -419 -561 -385
rect -527 -419 -493 -385
rect -459 -419 -425 -385
rect -391 -419 -357 -385
rect -323 -419 -289 -385
rect -255 -419 -221 -385
rect -187 -419 -153 -385
rect -119 -419 -85 -385
rect -51 -419 -17 -385
rect 17 -419 51 -385
rect 85 -419 119 -385
rect 153 -419 187 -385
rect 221 -419 255 -385
rect 289 -419 323 -385
rect 357 -419 391 -385
rect 425 -419 459 -385
rect 493 -419 527 -385
rect 561 -419 595 -385
rect 629 -419 663 -385
rect 697 -419 731 -385
rect 765 -419 799 -385
rect 833 -419 867 -385
rect 901 -419 1023 -385
<< viali >>
rect -881 385 -867 419
rect -867 385 -847 419
rect -809 385 -799 419
rect -799 385 -775 419
rect -737 385 -731 419
rect -731 385 -703 419
rect -665 385 -663 419
rect -663 385 -631 419
rect -593 385 -561 419
rect -561 385 -559 419
rect -521 385 -493 419
rect -493 385 -487 419
rect -449 385 -425 419
rect -425 385 -415 419
rect -377 385 -357 419
rect -357 385 -343 419
rect -305 385 -289 419
rect -289 385 -271 419
rect -233 385 -221 419
rect -221 385 -199 419
rect -161 385 -153 419
rect -153 385 -127 419
rect -89 385 -85 419
rect -85 385 -55 419
rect -17 385 17 419
rect 55 385 85 419
rect 85 385 89 419
rect 127 385 153 419
rect 153 385 161 419
rect 199 385 221 419
rect 221 385 233 419
rect 271 385 289 419
rect 289 385 305 419
rect 343 385 357 419
rect 357 385 377 419
rect 415 385 425 419
rect 425 385 449 419
rect 487 385 493 419
rect 493 385 521 419
rect 559 385 561 419
rect 561 385 593 419
rect 631 385 663 419
rect 663 385 665 419
rect 703 385 731 419
rect 731 385 737 419
rect 775 385 799 419
rect 799 385 809 419
rect 847 385 867 419
rect 867 385 881 419
rect -1023 323 -989 353
rect -1023 319 -989 323
rect -1023 255 -989 281
rect -1023 247 -989 255
rect -816 247 -814 281
rect -814 247 -782 281
rect -744 247 -712 281
rect -712 247 -710 281
rect -598 247 -596 281
rect -596 247 -564 281
rect -526 247 -494 281
rect -494 247 -492 281
rect -380 247 -378 281
rect -378 247 -346 281
rect -308 247 -276 281
rect -276 247 -274 281
rect -162 247 -160 281
rect -160 247 -128 281
rect -90 247 -58 281
rect -58 247 -56 281
rect 56 247 58 281
rect 58 247 90 281
rect 128 247 160 281
rect 160 247 162 281
rect 274 247 276 281
rect 276 247 308 281
rect 346 247 378 281
rect 378 247 380 281
rect 492 247 494 281
rect 494 247 526 281
rect 564 247 596 281
rect 596 247 598 281
rect 710 247 712 281
rect 712 247 744 281
rect 782 247 814 281
rect 814 247 816 281
rect -1023 187 -989 209
rect -1023 175 -989 187
rect -1023 119 -989 137
rect -1023 103 -989 119
rect -1023 51 -989 65
rect -1023 31 -989 51
rect -889 119 -855 149
rect -889 115 -855 119
rect -889 51 -855 77
rect -889 43 -855 51
rect -671 -51 -637 -43
rect -671 -77 -637 -51
rect -671 -119 -637 -115
rect -671 -149 -637 -119
rect -453 119 -419 149
rect -453 115 -419 119
rect -453 51 -419 77
rect -453 43 -419 51
rect -235 -51 -201 -43
rect -235 -77 -201 -51
rect -235 -119 -201 -115
rect -235 -149 -201 -119
rect -17 119 17 149
rect -17 115 17 119
rect -17 51 17 77
rect -17 43 17 51
rect 201 -51 235 -43
rect 201 -77 235 -51
rect 201 -119 235 -115
rect 201 -149 235 -119
rect 419 119 453 149
rect 419 115 453 119
rect 419 51 453 77
rect 419 43 453 51
rect 637 -51 671 -43
rect 637 -77 671 -51
rect 637 -119 671 -115
rect 637 -149 671 -119
rect 855 119 889 149
rect 855 115 889 119
rect 855 51 889 77
rect 855 43 889 51
rect -816 -281 -814 -247
rect -814 -281 -782 -247
rect -744 -281 -712 -247
rect -712 -281 -710 -247
rect -598 -281 -596 -247
rect -596 -281 -564 -247
rect -526 -281 -494 -247
rect -494 -281 -492 -247
rect -380 -281 -378 -247
rect -378 -281 -346 -247
rect -308 -281 -276 -247
rect -276 -281 -274 -247
rect -162 -281 -160 -247
rect -160 -281 -128 -247
rect -90 -281 -58 -247
rect -58 -281 -56 -247
rect 56 -281 58 -247
rect 58 -281 90 -247
rect 128 -281 160 -247
rect 160 -281 162 -247
rect 274 -281 276 -247
rect 276 -281 308 -247
rect 346 -281 378 -247
rect 378 -281 380 -247
rect 492 -281 494 -247
rect 494 -281 526 -247
rect 564 -281 596 -247
rect 596 -281 598 -247
rect 710 -281 712 -247
rect 712 -281 744 -247
rect 782 -281 814 -247
rect 814 -281 816 -247
<< metal1 >>
rect -902 419 902 425
rect -1029 353 -983 397
rect -902 385 -881 419
rect -847 385 -809 419
rect -775 385 -737 419
rect -703 385 -665 419
rect -631 385 -593 419
rect -559 385 -521 419
rect -487 385 -449 419
rect -415 385 -377 419
rect -343 385 -305 419
rect -271 385 -233 419
rect -199 385 -161 419
rect -127 385 -89 419
rect -55 385 -17 419
rect 17 385 55 419
rect 89 385 127 419
rect 161 385 199 419
rect 233 385 271 419
rect 305 385 343 419
rect 377 385 415 419
rect 449 385 487 419
rect 521 385 559 419
rect 593 385 631 419
rect 665 385 703 419
rect 737 385 775 419
rect 809 385 847 419
rect 881 385 902 419
rect -902 379 902 385
rect -1029 319 -1023 353
rect -989 319 -983 353
rect -1029 281 -983 319
rect -1029 247 -1023 281
rect -989 247 -983 281
rect -1029 209 -983 247
rect -839 281 -687 287
rect -839 247 -816 281
rect -782 247 -744 281
rect -710 247 -687 281
rect -839 241 -687 247
rect -621 281 -469 287
rect -621 247 -598 281
rect -564 247 -526 281
rect -492 247 -469 281
rect -621 241 -469 247
rect -403 281 -251 287
rect -403 247 -380 281
rect -346 247 -308 281
rect -274 247 -251 281
rect -403 241 -251 247
rect -185 281 -33 287
rect -185 247 -162 281
rect -128 247 -90 281
rect -56 247 -33 281
rect -185 241 -33 247
rect 33 281 185 287
rect 33 247 56 281
rect 90 247 128 281
rect 162 247 185 281
rect 33 241 185 247
rect 251 281 403 287
rect 251 247 274 281
rect 308 247 346 281
rect 380 247 403 281
rect 251 241 403 247
rect 469 281 621 287
rect 469 247 492 281
rect 526 247 564 281
rect 598 247 621 281
rect 469 241 621 247
rect 687 281 839 287
rect 687 247 710 281
rect 744 247 782 281
rect 816 247 839 281
rect 687 241 839 247
rect -1029 175 -1023 209
rect -989 175 -983 209
rect -1029 137 -983 175
rect -1029 103 -1023 137
rect -989 103 -983 137
rect -1029 65 -983 103
rect -1029 31 -1023 65
rect -989 31 -983 65
rect -1029 -12 -983 31
rect -895 149 -849 183
rect -895 115 -889 149
rect -855 115 -849 149
rect -895 77 -849 115
rect -895 43 -889 77
rect -855 43 -849 77
rect -895 9 -849 43
rect -459 149 -413 183
rect -459 115 -453 149
rect -419 115 -413 149
rect -459 77 -413 115
rect -459 43 -453 77
rect -419 43 -413 77
rect -459 9 -413 43
rect -23 149 23 183
rect -23 115 -17 149
rect 17 115 23 149
rect -23 77 23 115
rect -23 43 -17 77
rect 17 43 23 77
rect -23 9 23 43
rect 413 149 459 183
rect 413 115 419 149
rect 453 115 459 149
rect 413 77 459 115
rect 413 43 419 77
rect 453 43 459 77
rect 413 9 459 43
rect 849 149 895 183
rect 849 115 855 149
rect 889 115 895 149
rect 849 77 895 115
rect 849 43 855 77
rect 889 43 895 77
rect 849 9 895 43
rect -677 -43 -631 -9
rect -677 -77 -671 -43
rect -637 -77 -631 -43
rect -677 -115 -631 -77
rect -677 -149 -671 -115
rect -637 -149 -631 -115
rect -677 -183 -631 -149
rect -241 -43 -195 -9
rect -241 -77 -235 -43
rect -201 -77 -195 -43
rect -241 -115 -195 -77
rect -241 -149 -235 -115
rect -201 -149 -195 -115
rect -241 -183 -195 -149
rect 195 -43 241 -9
rect 195 -77 201 -43
rect 235 -77 241 -43
rect 195 -115 241 -77
rect 195 -149 201 -115
rect 235 -149 241 -115
rect 195 -183 241 -149
rect 631 -43 677 -9
rect 631 -77 637 -43
rect 671 -77 677 -43
rect 631 -115 677 -77
rect 631 -149 637 -115
rect 671 -149 677 -115
rect 631 -183 677 -149
rect -839 -247 -687 -241
rect -839 -281 -816 -247
rect -782 -281 -744 -247
rect -710 -281 -687 -247
rect -839 -287 -687 -281
rect -621 -247 -469 -241
rect -621 -281 -598 -247
rect -564 -281 -526 -247
rect -492 -281 -469 -247
rect -621 -287 -469 -281
rect -403 -247 -251 -241
rect -403 -281 -380 -247
rect -346 -281 -308 -247
rect -274 -281 -251 -247
rect -403 -287 -251 -281
rect -185 -247 -33 -241
rect -185 -281 -162 -247
rect -128 -281 -90 -247
rect -56 -281 -33 -247
rect -185 -287 -33 -281
rect 33 -247 185 -241
rect 33 -281 56 -247
rect 90 -281 128 -247
rect 162 -281 185 -247
rect 33 -287 185 -281
rect 251 -247 403 -241
rect 251 -281 274 -247
rect 308 -281 346 -247
rect 380 -281 403 -247
rect 251 -287 403 -281
rect 469 -247 621 -241
rect 469 -281 492 -247
rect 526 -281 564 -247
rect 598 -281 621 -247
rect 469 -287 621 -281
rect 687 -247 839 -241
rect 687 -281 710 -247
rect 744 -281 782 -247
rect 816 -281 839 -247
rect 687 -287 839 -281
<< properties >>
string FIXED_BBOX -1006 -402 1006 402
<< end >>
