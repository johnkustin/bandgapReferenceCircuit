magic
tech sky130A
magscale 1 2
timestamp 1620324069
<< nwell >>
rect -12306 -2798 12306 2764
<< pmoslvt >>
rect -12212 -2736 -11812 2664
rect -11640 -2736 -11240 2664
rect -11068 -2736 -10668 2664
rect -10496 -2736 -10096 2664
rect -9924 -2736 -9524 2664
rect -9352 -2736 -8952 2664
rect -8780 -2736 -8380 2664
rect -8208 -2736 -7808 2664
rect -7636 -2736 -7236 2664
rect -7064 -2736 -6664 2664
rect -6492 -2736 -6092 2664
rect -5920 -2736 -5520 2664
rect -5348 -2736 -4948 2664
rect -4776 -2736 -4376 2664
rect -4204 -2736 -3804 2664
rect -3632 -2736 -3232 2664
rect -3060 -2736 -2660 2664
rect -2488 -2736 -2088 2664
rect -1916 -2736 -1516 2664
rect -1344 -2736 -944 2664
rect -772 -2736 -372 2664
rect -200 -2736 200 2664
rect 372 -2736 772 2664
rect 944 -2736 1344 2664
rect 1516 -2736 1916 2664
rect 2088 -2736 2488 2664
rect 2660 -2736 3060 2664
rect 3232 -2736 3632 2664
rect 3804 -2736 4204 2664
rect 4376 -2736 4776 2664
rect 4948 -2736 5348 2664
rect 5520 -2736 5920 2664
rect 6092 -2736 6492 2664
rect 6664 -2736 7064 2664
rect 7236 -2736 7636 2664
rect 7808 -2736 8208 2664
rect 8380 -2736 8780 2664
rect 8952 -2736 9352 2664
rect 9524 -2736 9924 2664
rect 10096 -2736 10496 2664
rect 10668 -2736 11068 2664
rect 11240 -2736 11640 2664
rect 11812 -2736 12212 2664
<< pdiff >>
rect -12270 2652 -12212 2664
rect -12270 -2724 -12258 2652
rect -12224 -2724 -12212 2652
rect -12270 -2736 -12212 -2724
rect -11812 2652 -11754 2664
rect -11812 -2724 -11800 2652
rect -11766 -2724 -11754 2652
rect -11812 -2736 -11754 -2724
rect -11698 2652 -11640 2664
rect -11698 -2724 -11686 2652
rect -11652 -2724 -11640 2652
rect -11698 -2736 -11640 -2724
rect -11240 2652 -11182 2664
rect -11240 -2724 -11228 2652
rect -11194 -2724 -11182 2652
rect -11240 -2736 -11182 -2724
rect -11126 2652 -11068 2664
rect -11126 -2724 -11114 2652
rect -11080 -2724 -11068 2652
rect -11126 -2736 -11068 -2724
rect -10668 2652 -10610 2664
rect -10668 -2724 -10656 2652
rect -10622 -2724 -10610 2652
rect -10668 -2736 -10610 -2724
rect -10554 2652 -10496 2664
rect -10554 -2724 -10542 2652
rect -10508 -2724 -10496 2652
rect -10554 -2736 -10496 -2724
rect -10096 2652 -10038 2664
rect -10096 -2724 -10084 2652
rect -10050 -2724 -10038 2652
rect -10096 -2736 -10038 -2724
rect -9982 2652 -9924 2664
rect -9982 -2724 -9970 2652
rect -9936 -2724 -9924 2652
rect -9982 -2736 -9924 -2724
rect -9524 2652 -9466 2664
rect -9524 -2724 -9512 2652
rect -9478 -2724 -9466 2652
rect -9524 -2736 -9466 -2724
rect -9410 2652 -9352 2664
rect -9410 -2724 -9398 2652
rect -9364 -2724 -9352 2652
rect -9410 -2736 -9352 -2724
rect -8952 2652 -8894 2664
rect -8952 -2724 -8940 2652
rect -8906 -2724 -8894 2652
rect -8952 -2736 -8894 -2724
rect -8838 2652 -8780 2664
rect -8838 -2724 -8826 2652
rect -8792 -2724 -8780 2652
rect -8838 -2736 -8780 -2724
rect -8380 2652 -8322 2664
rect -8380 -2724 -8368 2652
rect -8334 -2724 -8322 2652
rect -8380 -2736 -8322 -2724
rect -8266 2652 -8208 2664
rect -8266 -2724 -8254 2652
rect -8220 -2724 -8208 2652
rect -8266 -2736 -8208 -2724
rect -7808 2652 -7750 2664
rect -7808 -2724 -7796 2652
rect -7762 -2724 -7750 2652
rect -7808 -2736 -7750 -2724
rect -7694 2652 -7636 2664
rect -7694 -2724 -7682 2652
rect -7648 -2724 -7636 2652
rect -7694 -2736 -7636 -2724
rect -7236 2652 -7178 2664
rect -7236 -2724 -7224 2652
rect -7190 -2724 -7178 2652
rect -7236 -2736 -7178 -2724
rect -7122 2652 -7064 2664
rect -7122 -2724 -7110 2652
rect -7076 -2724 -7064 2652
rect -7122 -2736 -7064 -2724
rect -6664 2652 -6606 2664
rect -6664 -2724 -6652 2652
rect -6618 -2724 -6606 2652
rect -6664 -2736 -6606 -2724
rect -6550 2652 -6492 2664
rect -6550 -2724 -6538 2652
rect -6504 -2724 -6492 2652
rect -6550 -2736 -6492 -2724
rect -6092 2652 -6034 2664
rect -6092 -2724 -6080 2652
rect -6046 -2724 -6034 2652
rect -6092 -2736 -6034 -2724
rect -5978 2652 -5920 2664
rect -5978 -2724 -5966 2652
rect -5932 -2724 -5920 2652
rect -5978 -2736 -5920 -2724
rect -5520 2652 -5462 2664
rect -5520 -2724 -5508 2652
rect -5474 -2724 -5462 2652
rect -5520 -2736 -5462 -2724
rect -5406 2652 -5348 2664
rect -5406 -2724 -5394 2652
rect -5360 -2724 -5348 2652
rect -5406 -2736 -5348 -2724
rect -4948 2652 -4890 2664
rect -4948 -2724 -4936 2652
rect -4902 -2724 -4890 2652
rect -4948 -2736 -4890 -2724
rect -4834 2652 -4776 2664
rect -4834 -2724 -4822 2652
rect -4788 -2724 -4776 2652
rect -4834 -2736 -4776 -2724
rect -4376 2652 -4318 2664
rect -4376 -2724 -4364 2652
rect -4330 -2724 -4318 2652
rect -4376 -2736 -4318 -2724
rect -4262 2652 -4204 2664
rect -4262 -2724 -4250 2652
rect -4216 -2724 -4204 2652
rect -4262 -2736 -4204 -2724
rect -3804 2652 -3746 2664
rect -3804 -2724 -3792 2652
rect -3758 -2724 -3746 2652
rect -3804 -2736 -3746 -2724
rect -3690 2652 -3632 2664
rect -3690 -2724 -3678 2652
rect -3644 -2724 -3632 2652
rect -3690 -2736 -3632 -2724
rect -3232 2652 -3174 2664
rect -3232 -2724 -3220 2652
rect -3186 -2724 -3174 2652
rect -3232 -2736 -3174 -2724
rect -3118 2652 -3060 2664
rect -3118 -2724 -3106 2652
rect -3072 -2724 -3060 2652
rect -3118 -2736 -3060 -2724
rect -2660 2652 -2602 2664
rect -2660 -2724 -2648 2652
rect -2614 -2724 -2602 2652
rect -2660 -2736 -2602 -2724
rect -2546 2652 -2488 2664
rect -2546 -2724 -2534 2652
rect -2500 -2724 -2488 2652
rect -2546 -2736 -2488 -2724
rect -2088 2652 -2030 2664
rect -2088 -2724 -2076 2652
rect -2042 -2724 -2030 2652
rect -2088 -2736 -2030 -2724
rect -1974 2652 -1916 2664
rect -1974 -2724 -1962 2652
rect -1928 -2724 -1916 2652
rect -1974 -2736 -1916 -2724
rect -1516 2652 -1458 2664
rect -1516 -2724 -1504 2652
rect -1470 -2724 -1458 2652
rect -1516 -2736 -1458 -2724
rect -1402 2652 -1344 2664
rect -1402 -2724 -1390 2652
rect -1356 -2724 -1344 2652
rect -1402 -2736 -1344 -2724
rect -944 2652 -886 2664
rect -944 -2724 -932 2652
rect -898 -2724 -886 2652
rect -944 -2736 -886 -2724
rect -830 2652 -772 2664
rect -830 -2724 -818 2652
rect -784 -2724 -772 2652
rect -830 -2736 -772 -2724
rect -372 2652 -314 2664
rect -372 -2724 -360 2652
rect -326 -2724 -314 2652
rect -372 -2736 -314 -2724
rect -258 2652 -200 2664
rect -258 -2724 -246 2652
rect -212 -2724 -200 2652
rect -258 -2736 -200 -2724
rect 200 2652 258 2664
rect 200 -2724 212 2652
rect 246 -2724 258 2652
rect 200 -2736 258 -2724
rect 314 2652 372 2664
rect 314 -2724 326 2652
rect 360 -2724 372 2652
rect 314 -2736 372 -2724
rect 772 2652 830 2664
rect 772 -2724 784 2652
rect 818 -2724 830 2652
rect 772 -2736 830 -2724
rect 886 2652 944 2664
rect 886 -2724 898 2652
rect 932 -2724 944 2652
rect 886 -2736 944 -2724
rect 1344 2652 1402 2664
rect 1344 -2724 1356 2652
rect 1390 -2724 1402 2652
rect 1344 -2736 1402 -2724
rect 1458 2652 1516 2664
rect 1458 -2724 1470 2652
rect 1504 -2724 1516 2652
rect 1458 -2736 1516 -2724
rect 1916 2652 1974 2664
rect 1916 -2724 1928 2652
rect 1962 -2724 1974 2652
rect 1916 -2736 1974 -2724
rect 2030 2652 2088 2664
rect 2030 -2724 2042 2652
rect 2076 -2724 2088 2652
rect 2030 -2736 2088 -2724
rect 2488 2652 2546 2664
rect 2488 -2724 2500 2652
rect 2534 -2724 2546 2652
rect 2488 -2736 2546 -2724
rect 2602 2652 2660 2664
rect 2602 -2724 2614 2652
rect 2648 -2724 2660 2652
rect 2602 -2736 2660 -2724
rect 3060 2652 3118 2664
rect 3060 -2724 3072 2652
rect 3106 -2724 3118 2652
rect 3060 -2736 3118 -2724
rect 3174 2652 3232 2664
rect 3174 -2724 3186 2652
rect 3220 -2724 3232 2652
rect 3174 -2736 3232 -2724
rect 3632 2652 3690 2664
rect 3632 -2724 3644 2652
rect 3678 -2724 3690 2652
rect 3632 -2736 3690 -2724
rect 3746 2652 3804 2664
rect 3746 -2724 3758 2652
rect 3792 -2724 3804 2652
rect 3746 -2736 3804 -2724
rect 4204 2652 4262 2664
rect 4204 -2724 4216 2652
rect 4250 -2724 4262 2652
rect 4204 -2736 4262 -2724
rect 4318 2652 4376 2664
rect 4318 -2724 4330 2652
rect 4364 -2724 4376 2652
rect 4318 -2736 4376 -2724
rect 4776 2652 4834 2664
rect 4776 -2724 4788 2652
rect 4822 -2724 4834 2652
rect 4776 -2736 4834 -2724
rect 4890 2652 4948 2664
rect 4890 -2724 4902 2652
rect 4936 -2724 4948 2652
rect 4890 -2736 4948 -2724
rect 5348 2652 5406 2664
rect 5348 -2724 5360 2652
rect 5394 -2724 5406 2652
rect 5348 -2736 5406 -2724
rect 5462 2652 5520 2664
rect 5462 -2724 5474 2652
rect 5508 -2724 5520 2652
rect 5462 -2736 5520 -2724
rect 5920 2652 5978 2664
rect 5920 -2724 5932 2652
rect 5966 -2724 5978 2652
rect 5920 -2736 5978 -2724
rect 6034 2652 6092 2664
rect 6034 -2724 6046 2652
rect 6080 -2724 6092 2652
rect 6034 -2736 6092 -2724
rect 6492 2652 6550 2664
rect 6492 -2724 6504 2652
rect 6538 -2724 6550 2652
rect 6492 -2736 6550 -2724
rect 6606 2652 6664 2664
rect 6606 -2724 6618 2652
rect 6652 -2724 6664 2652
rect 6606 -2736 6664 -2724
rect 7064 2652 7122 2664
rect 7064 -2724 7076 2652
rect 7110 -2724 7122 2652
rect 7064 -2736 7122 -2724
rect 7178 2652 7236 2664
rect 7178 -2724 7190 2652
rect 7224 -2724 7236 2652
rect 7178 -2736 7236 -2724
rect 7636 2652 7694 2664
rect 7636 -2724 7648 2652
rect 7682 -2724 7694 2652
rect 7636 -2736 7694 -2724
rect 7750 2652 7808 2664
rect 7750 -2724 7762 2652
rect 7796 -2724 7808 2652
rect 7750 -2736 7808 -2724
rect 8208 2652 8266 2664
rect 8208 -2724 8220 2652
rect 8254 -2724 8266 2652
rect 8208 -2736 8266 -2724
rect 8322 2652 8380 2664
rect 8322 -2724 8334 2652
rect 8368 -2724 8380 2652
rect 8322 -2736 8380 -2724
rect 8780 2652 8838 2664
rect 8780 -2724 8792 2652
rect 8826 -2724 8838 2652
rect 8780 -2736 8838 -2724
rect 8894 2652 8952 2664
rect 8894 -2724 8906 2652
rect 8940 -2724 8952 2652
rect 8894 -2736 8952 -2724
rect 9352 2652 9410 2664
rect 9352 -2724 9364 2652
rect 9398 -2724 9410 2652
rect 9352 -2736 9410 -2724
rect 9466 2652 9524 2664
rect 9466 -2724 9478 2652
rect 9512 -2724 9524 2652
rect 9466 -2736 9524 -2724
rect 9924 2652 9982 2664
rect 9924 -2724 9936 2652
rect 9970 -2724 9982 2652
rect 9924 -2736 9982 -2724
rect 10038 2652 10096 2664
rect 10038 -2724 10050 2652
rect 10084 -2724 10096 2652
rect 10038 -2736 10096 -2724
rect 10496 2652 10554 2664
rect 10496 -2724 10508 2652
rect 10542 -2724 10554 2652
rect 10496 -2736 10554 -2724
rect 10610 2652 10668 2664
rect 10610 -2724 10622 2652
rect 10656 -2724 10668 2652
rect 10610 -2736 10668 -2724
rect 11068 2652 11126 2664
rect 11068 -2724 11080 2652
rect 11114 -2724 11126 2652
rect 11068 -2736 11126 -2724
rect 11182 2652 11240 2664
rect 11182 -2724 11194 2652
rect 11228 -2724 11240 2652
rect 11182 -2736 11240 -2724
rect 11640 2652 11698 2664
rect 11640 -2724 11652 2652
rect 11686 -2724 11698 2652
rect 11640 -2736 11698 -2724
rect 11754 2652 11812 2664
rect 11754 -2724 11766 2652
rect 11800 -2724 11812 2652
rect 11754 -2736 11812 -2724
rect 12212 2652 12270 2664
rect 12212 -2724 12224 2652
rect 12258 -2724 12270 2652
rect 12212 -2736 12270 -2724
<< pdiffc >>
rect -12258 -2724 -12224 2652
rect -11800 -2724 -11766 2652
rect -11686 -2724 -11652 2652
rect -11228 -2724 -11194 2652
rect -11114 -2724 -11080 2652
rect -10656 -2724 -10622 2652
rect -10542 -2724 -10508 2652
rect -10084 -2724 -10050 2652
rect -9970 -2724 -9936 2652
rect -9512 -2724 -9478 2652
rect -9398 -2724 -9364 2652
rect -8940 -2724 -8906 2652
rect -8826 -2724 -8792 2652
rect -8368 -2724 -8334 2652
rect -8254 -2724 -8220 2652
rect -7796 -2724 -7762 2652
rect -7682 -2724 -7648 2652
rect -7224 -2724 -7190 2652
rect -7110 -2724 -7076 2652
rect -6652 -2724 -6618 2652
rect -6538 -2724 -6504 2652
rect -6080 -2724 -6046 2652
rect -5966 -2724 -5932 2652
rect -5508 -2724 -5474 2652
rect -5394 -2724 -5360 2652
rect -4936 -2724 -4902 2652
rect -4822 -2724 -4788 2652
rect -4364 -2724 -4330 2652
rect -4250 -2724 -4216 2652
rect -3792 -2724 -3758 2652
rect -3678 -2724 -3644 2652
rect -3220 -2724 -3186 2652
rect -3106 -2724 -3072 2652
rect -2648 -2724 -2614 2652
rect -2534 -2724 -2500 2652
rect -2076 -2724 -2042 2652
rect -1962 -2724 -1928 2652
rect -1504 -2724 -1470 2652
rect -1390 -2724 -1356 2652
rect -932 -2724 -898 2652
rect -818 -2724 -784 2652
rect -360 -2724 -326 2652
rect -246 -2724 -212 2652
rect 212 -2724 246 2652
rect 326 -2724 360 2652
rect 784 -2724 818 2652
rect 898 -2724 932 2652
rect 1356 -2724 1390 2652
rect 1470 -2724 1504 2652
rect 1928 -2724 1962 2652
rect 2042 -2724 2076 2652
rect 2500 -2724 2534 2652
rect 2614 -2724 2648 2652
rect 3072 -2724 3106 2652
rect 3186 -2724 3220 2652
rect 3644 -2724 3678 2652
rect 3758 -2724 3792 2652
rect 4216 -2724 4250 2652
rect 4330 -2724 4364 2652
rect 4788 -2724 4822 2652
rect 4902 -2724 4936 2652
rect 5360 -2724 5394 2652
rect 5474 -2724 5508 2652
rect 5932 -2724 5966 2652
rect 6046 -2724 6080 2652
rect 6504 -2724 6538 2652
rect 6618 -2724 6652 2652
rect 7076 -2724 7110 2652
rect 7190 -2724 7224 2652
rect 7648 -2724 7682 2652
rect 7762 -2724 7796 2652
rect 8220 -2724 8254 2652
rect 8334 -2724 8368 2652
rect 8792 -2724 8826 2652
rect 8906 -2724 8940 2652
rect 9364 -2724 9398 2652
rect 9478 -2724 9512 2652
rect 9936 -2724 9970 2652
rect 10050 -2724 10084 2652
rect 10508 -2724 10542 2652
rect 10622 -2724 10656 2652
rect 11080 -2724 11114 2652
rect 11194 -2724 11228 2652
rect 11652 -2724 11686 2652
rect 11766 -2724 11800 2652
rect 12224 -2724 12258 2652
<< poly >>
rect -12212 2745 -11812 2761
rect -12212 2711 -12196 2745
rect -11828 2711 -11812 2745
rect -12212 2664 -11812 2711
rect -11640 2745 -11240 2761
rect -11640 2711 -11624 2745
rect -11256 2711 -11240 2745
rect -11640 2664 -11240 2711
rect -11068 2745 -10668 2761
rect -11068 2711 -11052 2745
rect -10684 2711 -10668 2745
rect -11068 2664 -10668 2711
rect -10496 2745 -10096 2761
rect -10496 2711 -10480 2745
rect -10112 2711 -10096 2745
rect -10496 2664 -10096 2711
rect -9924 2745 -9524 2761
rect -9924 2711 -9908 2745
rect -9540 2711 -9524 2745
rect -9924 2664 -9524 2711
rect -9352 2745 -8952 2761
rect -9352 2711 -9336 2745
rect -8968 2711 -8952 2745
rect -9352 2664 -8952 2711
rect -8780 2745 -8380 2761
rect -8780 2711 -8764 2745
rect -8396 2711 -8380 2745
rect -8780 2664 -8380 2711
rect -8208 2745 -7808 2761
rect -8208 2711 -8192 2745
rect -7824 2711 -7808 2745
rect -8208 2664 -7808 2711
rect -7636 2745 -7236 2761
rect -7636 2711 -7620 2745
rect -7252 2711 -7236 2745
rect -7636 2664 -7236 2711
rect -7064 2745 -6664 2761
rect -7064 2711 -7048 2745
rect -6680 2711 -6664 2745
rect -7064 2664 -6664 2711
rect -6492 2745 -6092 2761
rect -6492 2711 -6476 2745
rect -6108 2711 -6092 2745
rect -6492 2664 -6092 2711
rect -5920 2745 -5520 2761
rect -5920 2711 -5904 2745
rect -5536 2711 -5520 2745
rect -5920 2664 -5520 2711
rect -5348 2745 -4948 2761
rect -5348 2711 -5332 2745
rect -4964 2711 -4948 2745
rect -5348 2664 -4948 2711
rect -4776 2745 -4376 2761
rect -4776 2711 -4760 2745
rect -4392 2711 -4376 2745
rect -4776 2664 -4376 2711
rect -4204 2745 -3804 2761
rect -4204 2711 -4188 2745
rect -3820 2711 -3804 2745
rect -4204 2664 -3804 2711
rect -3632 2745 -3232 2761
rect -3632 2711 -3616 2745
rect -3248 2711 -3232 2745
rect -3632 2664 -3232 2711
rect -3060 2745 -2660 2761
rect -3060 2711 -3044 2745
rect -2676 2711 -2660 2745
rect -3060 2664 -2660 2711
rect -2488 2745 -2088 2761
rect -2488 2711 -2472 2745
rect -2104 2711 -2088 2745
rect -2488 2664 -2088 2711
rect -1916 2745 -1516 2761
rect -1916 2711 -1900 2745
rect -1532 2711 -1516 2745
rect -1916 2664 -1516 2711
rect -1344 2745 -944 2761
rect -1344 2711 -1328 2745
rect -960 2711 -944 2745
rect -1344 2664 -944 2711
rect -772 2745 -372 2761
rect -772 2711 -756 2745
rect -388 2711 -372 2745
rect -772 2664 -372 2711
rect -200 2745 200 2761
rect -200 2711 -184 2745
rect 184 2711 200 2745
rect -200 2664 200 2711
rect 372 2745 772 2761
rect 372 2711 388 2745
rect 756 2711 772 2745
rect 372 2664 772 2711
rect 944 2745 1344 2761
rect 944 2711 960 2745
rect 1328 2711 1344 2745
rect 944 2664 1344 2711
rect 1516 2745 1916 2761
rect 1516 2711 1532 2745
rect 1900 2711 1916 2745
rect 1516 2664 1916 2711
rect 2088 2745 2488 2761
rect 2088 2711 2104 2745
rect 2472 2711 2488 2745
rect 2088 2664 2488 2711
rect 2660 2745 3060 2761
rect 2660 2711 2676 2745
rect 3044 2711 3060 2745
rect 2660 2664 3060 2711
rect 3232 2745 3632 2761
rect 3232 2711 3248 2745
rect 3616 2711 3632 2745
rect 3232 2664 3632 2711
rect 3804 2745 4204 2761
rect 3804 2711 3820 2745
rect 4188 2711 4204 2745
rect 3804 2664 4204 2711
rect 4376 2745 4776 2761
rect 4376 2711 4392 2745
rect 4760 2711 4776 2745
rect 4376 2664 4776 2711
rect 4948 2745 5348 2761
rect 4948 2711 4964 2745
rect 5332 2711 5348 2745
rect 4948 2664 5348 2711
rect 5520 2745 5920 2761
rect 5520 2711 5536 2745
rect 5904 2711 5920 2745
rect 5520 2664 5920 2711
rect 6092 2745 6492 2761
rect 6092 2711 6108 2745
rect 6476 2711 6492 2745
rect 6092 2664 6492 2711
rect 6664 2745 7064 2761
rect 6664 2711 6680 2745
rect 7048 2711 7064 2745
rect 6664 2664 7064 2711
rect 7236 2745 7636 2761
rect 7236 2711 7252 2745
rect 7620 2711 7636 2745
rect 7236 2664 7636 2711
rect 7808 2745 8208 2761
rect 7808 2711 7824 2745
rect 8192 2711 8208 2745
rect 7808 2664 8208 2711
rect 8380 2745 8780 2761
rect 8380 2711 8396 2745
rect 8764 2711 8780 2745
rect 8380 2664 8780 2711
rect 8952 2745 9352 2761
rect 8952 2711 8968 2745
rect 9336 2711 9352 2745
rect 8952 2664 9352 2711
rect 9524 2745 9924 2761
rect 9524 2711 9540 2745
rect 9908 2711 9924 2745
rect 9524 2664 9924 2711
rect 10096 2745 10496 2761
rect 10096 2711 10112 2745
rect 10480 2711 10496 2745
rect 10096 2664 10496 2711
rect 10668 2745 11068 2761
rect 10668 2711 10684 2745
rect 11052 2711 11068 2745
rect 10668 2664 11068 2711
rect 11240 2745 11640 2761
rect 11240 2711 11256 2745
rect 11624 2711 11640 2745
rect 11240 2664 11640 2711
rect 11812 2745 12212 2761
rect 11812 2711 11828 2745
rect 12196 2711 12212 2745
rect 11812 2664 12212 2711
rect -12212 -2762 -11812 -2736
rect -11640 -2762 -11240 -2736
rect -11068 -2762 -10668 -2736
rect -10496 -2762 -10096 -2736
rect -9924 -2762 -9524 -2736
rect -9352 -2762 -8952 -2736
rect -8780 -2762 -8380 -2736
rect -8208 -2762 -7808 -2736
rect -7636 -2762 -7236 -2736
rect -7064 -2762 -6664 -2736
rect -6492 -2762 -6092 -2736
rect -5920 -2762 -5520 -2736
rect -5348 -2762 -4948 -2736
rect -4776 -2762 -4376 -2736
rect -4204 -2762 -3804 -2736
rect -3632 -2762 -3232 -2736
rect -3060 -2762 -2660 -2736
rect -2488 -2762 -2088 -2736
rect -1916 -2762 -1516 -2736
rect -1344 -2762 -944 -2736
rect -772 -2762 -372 -2736
rect -200 -2762 200 -2736
rect 372 -2762 772 -2736
rect 944 -2762 1344 -2736
rect 1516 -2762 1916 -2736
rect 2088 -2762 2488 -2736
rect 2660 -2762 3060 -2736
rect 3232 -2762 3632 -2736
rect 3804 -2762 4204 -2736
rect 4376 -2762 4776 -2736
rect 4948 -2762 5348 -2736
rect 5520 -2762 5920 -2736
rect 6092 -2762 6492 -2736
rect 6664 -2762 7064 -2736
rect 7236 -2762 7636 -2736
rect 7808 -2762 8208 -2736
rect 8380 -2762 8780 -2736
rect 8952 -2762 9352 -2736
rect 9524 -2762 9924 -2736
rect 10096 -2762 10496 -2736
rect 10668 -2762 11068 -2736
rect 11240 -2762 11640 -2736
rect 11812 -2762 12212 -2736
<< polycont >>
rect -12196 2711 -11828 2745
rect -11624 2711 -11256 2745
rect -11052 2711 -10684 2745
rect -10480 2711 -10112 2745
rect -9908 2711 -9540 2745
rect -9336 2711 -8968 2745
rect -8764 2711 -8396 2745
rect -8192 2711 -7824 2745
rect -7620 2711 -7252 2745
rect -7048 2711 -6680 2745
rect -6476 2711 -6108 2745
rect -5904 2711 -5536 2745
rect -5332 2711 -4964 2745
rect -4760 2711 -4392 2745
rect -4188 2711 -3820 2745
rect -3616 2711 -3248 2745
rect -3044 2711 -2676 2745
rect -2472 2711 -2104 2745
rect -1900 2711 -1532 2745
rect -1328 2711 -960 2745
rect -756 2711 -388 2745
rect -184 2711 184 2745
rect 388 2711 756 2745
rect 960 2711 1328 2745
rect 1532 2711 1900 2745
rect 2104 2711 2472 2745
rect 2676 2711 3044 2745
rect 3248 2711 3616 2745
rect 3820 2711 4188 2745
rect 4392 2711 4760 2745
rect 4964 2711 5332 2745
rect 5536 2711 5904 2745
rect 6108 2711 6476 2745
rect 6680 2711 7048 2745
rect 7252 2711 7620 2745
rect 7824 2711 8192 2745
rect 8396 2711 8764 2745
rect 8968 2711 9336 2745
rect 9540 2711 9908 2745
rect 10112 2711 10480 2745
rect 10684 2711 11052 2745
rect 11256 2711 11624 2745
rect 11828 2711 12196 2745
<< locali >>
rect -12212 2711 -12196 2745
rect -11828 2711 -11812 2745
rect -11640 2711 -11624 2745
rect -11256 2711 -11240 2745
rect -11068 2711 -11052 2745
rect -10684 2711 -10668 2745
rect -10496 2711 -10480 2745
rect -10112 2711 -10096 2745
rect -9924 2711 -9908 2745
rect -9540 2711 -9524 2745
rect -9352 2711 -9336 2745
rect -8968 2711 -8952 2745
rect -8780 2711 -8764 2745
rect -8396 2711 -8380 2745
rect -8208 2711 -8192 2745
rect -7824 2711 -7808 2745
rect -7636 2711 -7620 2745
rect -7252 2711 -7236 2745
rect -7064 2711 -7048 2745
rect -6680 2711 -6664 2745
rect -6492 2711 -6476 2745
rect -6108 2711 -6092 2745
rect -5920 2711 -5904 2745
rect -5536 2711 -5520 2745
rect -5348 2711 -5332 2745
rect -4964 2711 -4948 2745
rect -4776 2711 -4760 2745
rect -4392 2711 -4376 2745
rect -4204 2711 -4188 2745
rect -3820 2711 -3804 2745
rect -3632 2711 -3616 2745
rect -3248 2711 -3232 2745
rect -3060 2711 -3044 2745
rect -2676 2711 -2660 2745
rect -2488 2711 -2472 2745
rect -2104 2711 -2088 2745
rect -1916 2711 -1900 2745
rect -1532 2711 -1516 2745
rect -1344 2711 -1328 2745
rect -960 2711 -944 2745
rect -772 2711 -756 2745
rect -388 2711 -372 2745
rect -200 2711 -184 2745
rect 184 2711 200 2745
rect 372 2711 388 2745
rect 756 2711 772 2745
rect 944 2711 960 2745
rect 1328 2711 1344 2745
rect 1516 2711 1532 2745
rect 1900 2711 1916 2745
rect 2088 2711 2104 2745
rect 2472 2711 2488 2745
rect 2660 2711 2676 2745
rect 3044 2711 3060 2745
rect 3232 2711 3248 2745
rect 3616 2711 3632 2745
rect 3804 2711 3820 2745
rect 4188 2711 4204 2745
rect 4376 2711 4392 2745
rect 4760 2711 4776 2745
rect 4948 2711 4964 2745
rect 5332 2711 5348 2745
rect 5520 2711 5536 2745
rect 5904 2711 5920 2745
rect 6092 2711 6108 2745
rect 6476 2711 6492 2745
rect 6664 2711 6680 2745
rect 7048 2711 7064 2745
rect 7236 2711 7252 2745
rect 7620 2711 7636 2745
rect 7808 2711 7824 2745
rect 8192 2711 8208 2745
rect 8380 2711 8396 2745
rect 8764 2711 8780 2745
rect 8952 2711 8968 2745
rect 9336 2711 9352 2745
rect 9524 2711 9540 2745
rect 9908 2711 9924 2745
rect 10096 2711 10112 2745
rect 10480 2711 10496 2745
rect 10668 2711 10684 2745
rect 11052 2711 11068 2745
rect 11240 2711 11256 2745
rect 11624 2711 11640 2745
rect 11812 2711 11828 2745
rect 12196 2711 12212 2745
rect -12258 2652 -12224 2668
rect -12258 -2740 -12224 -2724
rect -11800 2652 -11766 2668
rect -11800 -2740 -11766 -2724
rect -11686 2652 -11652 2668
rect -11686 -2740 -11652 -2724
rect -11228 2652 -11194 2668
rect -11228 -2740 -11194 -2724
rect -11114 2652 -11080 2668
rect -11114 -2740 -11080 -2724
rect -10656 2652 -10622 2668
rect -10656 -2740 -10622 -2724
rect -10542 2652 -10508 2668
rect -10542 -2740 -10508 -2724
rect -10084 2652 -10050 2668
rect -10084 -2740 -10050 -2724
rect -9970 2652 -9936 2668
rect -9970 -2740 -9936 -2724
rect -9512 2652 -9478 2668
rect -9512 -2740 -9478 -2724
rect -9398 2652 -9364 2668
rect -9398 -2740 -9364 -2724
rect -8940 2652 -8906 2668
rect -8940 -2740 -8906 -2724
rect -8826 2652 -8792 2668
rect -8826 -2740 -8792 -2724
rect -8368 2652 -8334 2668
rect -8368 -2740 -8334 -2724
rect -8254 2652 -8220 2668
rect -8254 -2740 -8220 -2724
rect -7796 2652 -7762 2668
rect -7796 -2740 -7762 -2724
rect -7682 2652 -7648 2668
rect -7682 -2740 -7648 -2724
rect -7224 2652 -7190 2668
rect -7224 -2740 -7190 -2724
rect -7110 2652 -7076 2668
rect -7110 -2740 -7076 -2724
rect -6652 2652 -6618 2668
rect -6652 -2740 -6618 -2724
rect -6538 2652 -6504 2668
rect -6538 -2740 -6504 -2724
rect -6080 2652 -6046 2668
rect -6080 -2740 -6046 -2724
rect -5966 2652 -5932 2668
rect -5966 -2740 -5932 -2724
rect -5508 2652 -5474 2668
rect -5508 -2740 -5474 -2724
rect -5394 2652 -5360 2668
rect -5394 -2740 -5360 -2724
rect -4936 2652 -4902 2668
rect -4936 -2740 -4902 -2724
rect -4822 2652 -4788 2668
rect -4822 -2740 -4788 -2724
rect -4364 2652 -4330 2668
rect -4364 -2740 -4330 -2724
rect -4250 2652 -4216 2668
rect -4250 -2740 -4216 -2724
rect -3792 2652 -3758 2668
rect -3792 -2740 -3758 -2724
rect -3678 2652 -3644 2668
rect -3678 -2740 -3644 -2724
rect -3220 2652 -3186 2668
rect -3220 -2740 -3186 -2724
rect -3106 2652 -3072 2668
rect -3106 -2740 -3072 -2724
rect -2648 2652 -2614 2668
rect -2648 -2740 -2614 -2724
rect -2534 2652 -2500 2668
rect -2534 -2740 -2500 -2724
rect -2076 2652 -2042 2668
rect -2076 -2740 -2042 -2724
rect -1962 2652 -1928 2668
rect -1962 -2740 -1928 -2724
rect -1504 2652 -1470 2668
rect -1504 -2740 -1470 -2724
rect -1390 2652 -1356 2668
rect -1390 -2740 -1356 -2724
rect -932 2652 -898 2668
rect -932 -2740 -898 -2724
rect -818 2652 -784 2668
rect -818 -2740 -784 -2724
rect -360 2652 -326 2668
rect -360 -2740 -326 -2724
rect -246 2652 -212 2668
rect -246 -2740 -212 -2724
rect 212 2652 246 2668
rect 212 -2740 246 -2724
rect 326 2652 360 2668
rect 326 -2740 360 -2724
rect 784 2652 818 2668
rect 784 -2740 818 -2724
rect 898 2652 932 2668
rect 898 -2740 932 -2724
rect 1356 2652 1390 2668
rect 1356 -2740 1390 -2724
rect 1470 2652 1504 2668
rect 1470 -2740 1504 -2724
rect 1928 2652 1962 2668
rect 1928 -2740 1962 -2724
rect 2042 2652 2076 2668
rect 2042 -2740 2076 -2724
rect 2500 2652 2534 2668
rect 2500 -2740 2534 -2724
rect 2614 2652 2648 2668
rect 2614 -2740 2648 -2724
rect 3072 2652 3106 2668
rect 3072 -2740 3106 -2724
rect 3186 2652 3220 2668
rect 3186 -2740 3220 -2724
rect 3644 2652 3678 2668
rect 3644 -2740 3678 -2724
rect 3758 2652 3792 2668
rect 3758 -2740 3792 -2724
rect 4216 2652 4250 2668
rect 4216 -2740 4250 -2724
rect 4330 2652 4364 2668
rect 4330 -2740 4364 -2724
rect 4788 2652 4822 2668
rect 4788 -2740 4822 -2724
rect 4902 2652 4936 2668
rect 4902 -2740 4936 -2724
rect 5360 2652 5394 2668
rect 5360 -2740 5394 -2724
rect 5474 2652 5508 2668
rect 5474 -2740 5508 -2724
rect 5932 2652 5966 2668
rect 5932 -2740 5966 -2724
rect 6046 2652 6080 2668
rect 6046 -2740 6080 -2724
rect 6504 2652 6538 2668
rect 6504 -2740 6538 -2724
rect 6618 2652 6652 2668
rect 6618 -2740 6652 -2724
rect 7076 2652 7110 2668
rect 7076 -2740 7110 -2724
rect 7190 2652 7224 2668
rect 7190 -2740 7224 -2724
rect 7648 2652 7682 2668
rect 7648 -2740 7682 -2724
rect 7762 2652 7796 2668
rect 7762 -2740 7796 -2724
rect 8220 2652 8254 2668
rect 8220 -2740 8254 -2724
rect 8334 2652 8368 2668
rect 8334 -2740 8368 -2724
rect 8792 2652 8826 2668
rect 8792 -2740 8826 -2724
rect 8906 2652 8940 2668
rect 8906 -2740 8940 -2724
rect 9364 2652 9398 2668
rect 9364 -2740 9398 -2724
rect 9478 2652 9512 2668
rect 9478 -2740 9512 -2724
rect 9936 2652 9970 2668
rect 9936 -2740 9970 -2724
rect 10050 2652 10084 2668
rect 10050 -2740 10084 -2724
rect 10508 2652 10542 2668
rect 10508 -2740 10542 -2724
rect 10622 2652 10656 2668
rect 10622 -2740 10656 -2724
rect 11080 2652 11114 2668
rect 11080 -2740 11114 -2724
rect 11194 2652 11228 2668
rect 11194 -2740 11228 -2724
rect 11652 2652 11686 2668
rect 11652 -2740 11686 -2724
rect 11766 2652 11800 2668
rect 11766 -2740 11800 -2724
rect 12224 2652 12258 2668
rect 12224 -2740 12258 -2724
<< viali >>
rect -12196 2711 -11828 2745
rect -11624 2711 -11256 2745
rect -11052 2711 -10684 2745
rect -10480 2711 -10112 2745
rect -9908 2711 -9540 2745
rect -9336 2711 -8968 2745
rect -8764 2711 -8396 2745
rect -8192 2711 -7824 2745
rect -7620 2711 -7252 2745
rect -7048 2711 -6680 2745
rect -6476 2711 -6108 2745
rect -5904 2711 -5536 2745
rect -5332 2711 -4964 2745
rect -4760 2711 -4392 2745
rect -4188 2711 -3820 2745
rect -3616 2711 -3248 2745
rect -3044 2711 -2676 2745
rect -2472 2711 -2104 2745
rect -1900 2711 -1532 2745
rect -1328 2711 -960 2745
rect -756 2711 -388 2745
rect -184 2711 184 2745
rect 388 2711 756 2745
rect 960 2711 1328 2745
rect 1532 2711 1900 2745
rect 2104 2711 2472 2745
rect 2676 2711 3044 2745
rect 3248 2711 3616 2745
rect 3820 2711 4188 2745
rect 4392 2711 4760 2745
rect 4964 2711 5332 2745
rect 5536 2711 5904 2745
rect 6108 2711 6476 2745
rect 6680 2711 7048 2745
rect 7252 2711 7620 2745
rect 7824 2711 8192 2745
rect 8396 2711 8764 2745
rect 8968 2711 9336 2745
rect 9540 2711 9908 2745
rect 10112 2711 10480 2745
rect 10684 2711 11052 2745
rect 11256 2711 11624 2745
rect 11828 2711 12196 2745
rect -12258 -2724 -12224 2652
rect -11800 -2724 -11766 2652
rect -11686 -2724 -11652 2652
rect -11228 -2724 -11194 2652
rect -11114 -2724 -11080 2652
rect -10656 -2724 -10622 2652
rect -10542 -2724 -10508 2652
rect -10084 -2724 -10050 2652
rect -9970 -2724 -9936 2652
rect -9512 -2724 -9478 2652
rect -9398 -2724 -9364 2652
rect -8940 -2724 -8906 2652
rect -8826 -2724 -8792 2652
rect -8368 -2724 -8334 2652
rect -8254 -2724 -8220 2652
rect -7796 -2724 -7762 2652
rect -7682 -2724 -7648 2652
rect -7224 -2724 -7190 2652
rect -7110 -2724 -7076 2652
rect -6652 -2724 -6618 2652
rect -6538 -2724 -6504 2652
rect -6080 -2724 -6046 2652
rect -5966 -2724 -5932 2652
rect -5508 -2724 -5474 2652
rect -5394 -2724 -5360 2652
rect -4936 -2724 -4902 2652
rect -4822 -2724 -4788 2652
rect -4364 -2724 -4330 2652
rect -4250 -2724 -4216 2652
rect -3792 -2724 -3758 2652
rect -3678 -2724 -3644 2652
rect -3220 -2724 -3186 2652
rect -3106 -2724 -3072 2652
rect -2648 -2724 -2614 2652
rect -2534 -2724 -2500 2652
rect -2076 -2724 -2042 2652
rect -1962 -2724 -1928 2652
rect -1504 -2724 -1470 2652
rect -1390 -2724 -1356 2652
rect -932 -2724 -898 2652
rect -818 -2724 -784 2652
rect -360 -2724 -326 2652
rect -246 -2724 -212 2652
rect 212 -2724 246 2652
rect 326 -2724 360 2652
rect 784 -2724 818 2652
rect 898 -2724 932 2652
rect 1356 -2724 1390 2652
rect 1470 -2724 1504 2652
rect 1928 -2724 1962 2652
rect 2042 -2724 2076 2652
rect 2500 -2724 2534 2652
rect 2614 -2724 2648 2652
rect 3072 -2724 3106 2652
rect 3186 -2724 3220 2652
rect 3644 -2724 3678 2652
rect 3758 -2724 3792 2652
rect 4216 -2724 4250 2652
rect 4330 -2724 4364 2652
rect 4788 -2724 4822 2652
rect 4902 -2724 4936 2652
rect 5360 -2724 5394 2652
rect 5474 -2724 5508 2652
rect 5932 -2724 5966 2652
rect 6046 -2724 6080 2652
rect 6504 -2724 6538 2652
rect 6618 -2724 6652 2652
rect 7076 -2724 7110 2652
rect 7190 -2724 7224 2652
rect 7648 -2724 7682 2652
rect 7762 -2724 7796 2652
rect 8220 -2724 8254 2652
rect 8334 -2724 8368 2652
rect 8792 -2724 8826 2652
rect 8906 -2724 8940 2652
rect 9364 -2724 9398 2652
rect 9478 -2724 9512 2652
rect 9936 -2724 9970 2652
rect 10050 -2724 10084 2652
rect 10508 -2724 10542 2652
rect 10622 -2724 10656 2652
rect 11080 -2724 11114 2652
rect 11194 -2724 11228 2652
rect 11652 -2724 11686 2652
rect 11766 -2724 11800 2652
rect 12224 -2724 12258 2652
<< metal1 >>
rect -12208 2745 -11816 2751
rect -12208 2711 -12196 2745
rect -11828 2711 -11816 2745
rect -12208 2705 -11816 2711
rect -11636 2745 -11244 2751
rect -11636 2711 -11624 2745
rect -11256 2711 -11244 2745
rect -11636 2705 -11244 2711
rect -11064 2745 -10672 2751
rect -11064 2711 -11052 2745
rect -10684 2711 -10672 2745
rect -11064 2705 -10672 2711
rect -10492 2745 -10100 2751
rect -10492 2711 -10480 2745
rect -10112 2711 -10100 2745
rect -10492 2705 -10100 2711
rect -9920 2745 -9528 2751
rect -9920 2711 -9908 2745
rect -9540 2711 -9528 2745
rect -9920 2705 -9528 2711
rect -9348 2745 -8956 2751
rect -9348 2711 -9336 2745
rect -8968 2711 -8956 2745
rect -9348 2705 -8956 2711
rect -8776 2745 -8384 2751
rect -8776 2711 -8764 2745
rect -8396 2711 -8384 2745
rect -8776 2705 -8384 2711
rect -8204 2745 -7812 2751
rect -8204 2711 -8192 2745
rect -7824 2711 -7812 2745
rect -8204 2705 -7812 2711
rect -7632 2745 -7240 2751
rect -7632 2711 -7620 2745
rect -7252 2711 -7240 2745
rect -7632 2705 -7240 2711
rect -7060 2745 -6668 2751
rect -7060 2711 -7048 2745
rect -6680 2711 -6668 2745
rect -7060 2705 -6668 2711
rect -6488 2745 -6096 2751
rect -6488 2711 -6476 2745
rect -6108 2711 -6096 2745
rect -6488 2705 -6096 2711
rect -5916 2745 -5524 2751
rect -5916 2711 -5904 2745
rect -5536 2711 -5524 2745
rect -5916 2705 -5524 2711
rect -5344 2745 -4952 2751
rect -5344 2711 -5332 2745
rect -4964 2711 -4952 2745
rect -5344 2705 -4952 2711
rect -4772 2745 -4380 2751
rect -4772 2711 -4760 2745
rect -4392 2711 -4380 2745
rect -4772 2705 -4380 2711
rect -4200 2745 -3808 2751
rect -4200 2711 -4188 2745
rect -3820 2711 -3808 2745
rect -4200 2705 -3808 2711
rect -3628 2745 -3236 2751
rect -3628 2711 -3616 2745
rect -3248 2711 -3236 2745
rect -3628 2705 -3236 2711
rect -3056 2745 -2664 2751
rect -3056 2711 -3044 2745
rect -2676 2711 -2664 2745
rect -3056 2705 -2664 2711
rect -2484 2745 -2092 2751
rect -2484 2711 -2472 2745
rect -2104 2711 -2092 2745
rect -2484 2705 -2092 2711
rect -1912 2745 -1520 2751
rect -1912 2711 -1900 2745
rect -1532 2711 -1520 2745
rect -1912 2705 -1520 2711
rect -1340 2745 -948 2751
rect -1340 2711 -1328 2745
rect -960 2711 -948 2745
rect -1340 2705 -948 2711
rect -768 2745 -376 2751
rect -768 2711 -756 2745
rect -388 2711 -376 2745
rect -768 2705 -376 2711
rect -196 2745 196 2751
rect -196 2711 -184 2745
rect 184 2711 196 2745
rect -196 2705 196 2711
rect 376 2745 768 2751
rect 376 2711 388 2745
rect 756 2711 768 2745
rect 376 2705 768 2711
rect 948 2745 1340 2751
rect 948 2711 960 2745
rect 1328 2711 1340 2745
rect 948 2705 1340 2711
rect 1520 2745 1912 2751
rect 1520 2711 1532 2745
rect 1900 2711 1912 2745
rect 1520 2705 1912 2711
rect 2092 2745 2484 2751
rect 2092 2711 2104 2745
rect 2472 2711 2484 2745
rect 2092 2705 2484 2711
rect 2664 2745 3056 2751
rect 2664 2711 2676 2745
rect 3044 2711 3056 2745
rect 2664 2705 3056 2711
rect 3236 2745 3628 2751
rect 3236 2711 3248 2745
rect 3616 2711 3628 2745
rect 3236 2705 3628 2711
rect 3808 2745 4200 2751
rect 3808 2711 3820 2745
rect 4188 2711 4200 2745
rect 3808 2705 4200 2711
rect 4380 2745 4772 2751
rect 4380 2711 4392 2745
rect 4760 2711 4772 2745
rect 4380 2705 4772 2711
rect 4952 2745 5344 2751
rect 4952 2711 4964 2745
rect 5332 2711 5344 2745
rect 4952 2705 5344 2711
rect 5524 2745 5916 2751
rect 5524 2711 5536 2745
rect 5904 2711 5916 2745
rect 5524 2705 5916 2711
rect 6096 2745 6488 2751
rect 6096 2711 6108 2745
rect 6476 2711 6488 2745
rect 6096 2705 6488 2711
rect 6668 2745 7060 2751
rect 6668 2711 6680 2745
rect 7048 2711 7060 2745
rect 6668 2705 7060 2711
rect 7240 2745 7632 2751
rect 7240 2711 7252 2745
rect 7620 2711 7632 2745
rect 7240 2705 7632 2711
rect 7812 2745 8204 2751
rect 7812 2711 7824 2745
rect 8192 2711 8204 2745
rect 7812 2705 8204 2711
rect 8384 2745 8776 2751
rect 8384 2711 8396 2745
rect 8764 2711 8776 2745
rect 8384 2705 8776 2711
rect 8956 2745 9348 2751
rect 8956 2711 8968 2745
rect 9336 2711 9348 2745
rect 8956 2705 9348 2711
rect 9528 2745 9920 2751
rect 9528 2711 9540 2745
rect 9908 2711 9920 2745
rect 9528 2705 9920 2711
rect 10100 2745 10492 2751
rect 10100 2711 10112 2745
rect 10480 2711 10492 2745
rect 10100 2705 10492 2711
rect 10672 2745 11064 2751
rect 10672 2711 10684 2745
rect 11052 2711 11064 2745
rect 10672 2705 11064 2711
rect 11244 2745 11636 2751
rect 11244 2711 11256 2745
rect 11624 2711 11636 2745
rect 11244 2705 11636 2711
rect 11816 2745 12208 2751
rect 11816 2711 11828 2745
rect 12196 2711 12208 2745
rect 11816 2705 12208 2711
rect -12264 2652 -12218 2664
rect -12264 -2724 -12258 2652
rect -12224 -2724 -12218 2652
rect -12264 -2736 -12218 -2724
rect -11806 2652 -11760 2664
rect -11806 -2724 -11800 2652
rect -11766 -2724 -11760 2652
rect -11806 -2736 -11760 -2724
rect -11692 2652 -11646 2664
rect -11692 -2724 -11686 2652
rect -11652 -2724 -11646 2652
rect -11692 -2736 -11646 -2724
rect -11234 2652 -11188 2664
rect -11234 -2724 -11228 2652
rect -11194 -2724 -11188 2652
rect -11234 -2736 -11188 -2724
rect -11120 2652 -11074 2664
rect -11120 -2724 -11114 2652
rect -11080 -2724 -11074 2652
rect -11120 -2736 -11074 -2724
rect -10662 2652 -10616 2664
rect -10662 -2724 -10656 2652
rect -10622 -2724 -10616 2652
rect -10662 -2736 -10616 -2724
rect -10548 2652 -10502 2664
rect -10548 -2724 -10542 2652
rect -10508 -2724 -10502 2652
rect -10548 -2736 -10502 -2724
rect -10090 2652 -10044 2664
rect -10090 -2724 -10084 2652
rect -10050 -2724 -10044 2652
rect -10090 -2736 -10044 -2724
rect -9976 2652 -9930 2664
rect -9976 -2724 -9970 2652
rect -9936 -2724 -9930 2652
rect -9976 -2736 -9930 -2724
rect -9518 2652 -9472 2664
rect -9518 -2724 -9512 2652
rect -9478 -2724 -9472 2652
rect -9518 -2736 -9472 -2724
rect -9404 2652 -9358 2664
rect -9404 -2724 -9398 2652
rect -9364 -2724 -9358 2652
rect -9404 -2736 -9358 -2724
rect -8946 2652 -8900 2664
rect -8946 -2724 -8940 2652
rect -8906 -2724 -8900 2652
rect -8946 -2736 -8900 -2724
rect -8832 2652 -8786 2664
rect -8832 -2724 -8826 2652
rect -8792 -2724 -8786 2652
rect -8832 -2736 -8786 -2724
rect -8374 2652 -8328 2664
rect -8374 -2724 -8368 2652
rect -8334 -2724 -8328 2652
rect -8374 -2736 -8328 -2724
rect -8260 2652 -8214 2664
rect -8260 -2724 -8254 2652
rect -8220 -2724 -8214 2652
rect -8260 -2736 -8214 -2724
rect -7802 2652 -7756 2664
rect -7802 -2724 -7796 2652
rect -7762 -2724 -7756 2652
rect -7802 -2736 -7756 -2724
rect -7688 2652 -7642 2664
rect -7688 -2724 -7682 2652
rect -7648 -2724 -7642 2652
rect -7688 -2736 -7642 -2724
rect -7230 2652 -7184 2664
rect -7230 -2724 -7224 2652
rect -7190 -2724 -7184 2652
rect -7230 -2736 -7184 -2724
rect -7116 2652 -7070 2664
rect -7116 -2724 -7110 2652
rect -7076 -2724 -7070 2652
rect -7116 -2736 -7070 -2724
rect -6658 2652 -6612 2664
rect -6658 -2724 -6652 2652
rect -6618 -2724 -6612 2652
rect -6658 -2736 -6612 -2724
rect -6544 2652 -6498 2664
rect -6544 -2724 -6538 2652
rect -6504 -2724 -6498 2652
rect -6544 -2736 -6498 -2724
rect -6086 2652 -6040 2664
rect -6086 -2724 -6080 2652
rect -6046 -2724 -6040 2652
rect -6086 -2736 -6040 -2724
rect -5972 2652 -5926 2664
rect -5972 -2724 -5966 2652
rect -5932 -2724 -5926 2652
rect -5972 -2736 -5926 -2724
rect -5514 2652 -5468 2664
rect -5514 -2724 -5508 2652
rect -5474 -2724 -5468 2652
rect -5514 -2736 -5468 -2724
rect -5400 2652 -5354 2664
rect -5400 -2724 -5394 2652
rect -5360 -2724 -5354 2652
rect -5400 -2736 -5354 -2724
rect -4942 2652 -4896 2664
rect -4942 -2724 -4936 2652
rect -4902 -2724 -4896 2652
rect -4942 -2736 -4896 -2724
rect -4828 2652 -4782 2664
rect -4828 -2724 -4822 2652
rect -4788 -2724 -4782 2652
rect -4828 -2736 -4782 -2724
rect -4370 2652 -4324 2664
rect -4370 -2724 -4364 2652
rect -4330 -2724 -4324 2652
rect -4370 -2736 -4324 -2724
rect -4256 2652 -4210 2664
rect -4256 -2724 -4250 2652
rect -4216 -2724 -4210 2652
rect -4256 -2736 -4210 -2724
rect -3798 2652 -3752 2664
rect -3798 -2724 -3792 2652
rect -3758 -2724 -3752 2652
rect -3798 -2736 -3752 -2724
rect -3684 2652 -3638 2664
rect -3684 -2724 -3678 2652
rect -3644 -2724 -3638 2652
rect -3684 -2736 -3638 -2724
rect -3226 2652 -3180 2664
rect -3226 -2724 -3220 2652
rect -3186 -2724 -3180 2652
rect -3226 -2736 -3180 -2724
rect -3112 2652 -3066 2664
rect -3112 -2724 -3106 2652
rect -3072 -2724 -3066 2652
rect -3112 -2736 -3066 -2724
rect -2654 2652 -2608 2664
rect -2654 -2724 -2648 2652
rect -2614 -2724 -2608 2652
rect -2654 -2736 -2608 -2724
rect -2540 2652 -2494 2664
rect -2540 -2724 -2534 2652
rect -2500 -2724 -2494 2652
rect -2540 -2736 -2494 -2724
rect -2082 2652 -2036 2664
rect -2082 -2724 -2076 2652
rect -2042 -2724 -2036 2652
rect -2082 -2736 -2036 -2724
rect -1968 2652 -1922 2664
rect -1968 -2724 -1962 2652
rect -1928 -2724 -1922 2652
rect -1968 -2736 -1922 -2724
rect -1510 2652 -1464 2664
rect -1510 -2724 -1504 2652
rect -1470 -2724 -1464 2652
rect -1510 -2736 -1464 -2724
rect -1396 2652 -1350 2664
rect -1396 -2724 -1390 2652
rect -1356 -2724 -1350 2652
rect -1396 -2736 -1350 -2724
rect -938 2652 -892 2664
rect -938 -2724 -932 2652
rect -898 -2724 -892 2652
rect -938 -2736 -892 -2724
rect -824 2652 -778 2664
rect -824 -2724 -818 2652
rect -784 -2724 -778 2652
rect -824 -2736 -778 -2724
rect -366 2652 -320 2664
rect -366 -2724 -360 2652
rect -326 -2724 -320 2652
rect -366 -2736 -320 -2724
rect -252 2652 -206 2664
rect -252 -2724 -246 2652
rect -212 -2724 -206 2652
rect -252 -2736 -206 -2724
rect 206 2652 252 2664
rect 206 -2724 212 2652
rect 246 -2724 252 2652
rect 206 -2736 252 -2724
rect 320 2652 366 2664
rect 320 -2724 326 2652
rect 360 -2724 366 2652
rect 320 -2736 366 -2724
rect 778 2652 824 2664
rect 778 -2724 784 2652
rect 818 -2724 824 2652
rect 778 -2736 824 -2724
rect 892 2652 938 2664
rect 892 -2724 898 2652
rect 932 -2724 938 2652
rect 892 -2736 938 -2724
rect 1350 2652 1396 2664
rect 1350 -2724 1356 2652
rect 1390 -2724 1396 2652
rect 1350 -2736 1396 -2724
rect 1464 2652 1510 2664
rect 1464 -2724 1470 2652
rect 1504 -2724 1510 2652
rect 1464 -2736 1510 -2724
rect 1922 2652 1968 2664
rect 1922 -2724 1928 2652
rect 1962 -2724 1968 2652
rect 1922 -2736 1968 -2724
rect 2036 2652 2082 2664
rect 2036 -2724 2042 2652
rect 2076 -2724 2082 2652
rect 2036 -2736 2082 -2724
rect 2494 2652 2540 2664
rect 2494 -2724 2500 2652
rect 2534 -2724 2540 2652
rect 2494 -2736 2540 -2724
rect 2608 2652 2654 2664
rect 2608 -2724 2614 2652
rect 2648 -2724 2654 2652
rect 2608 -2736 2654 -2724
rect 3066 2652 3112 2664
rect 3066 -2724 3072 2652
rect 3106 -2724 3112 2652
rect 3066 -2736 3112 -2724
rect 3180 2652 3226 2664
rect 3180 -2724 3186 2652
rect 3220 -2724 3226 2652
rect 3180 -2736 3226 -2724
rect 3638 2652 3684 2664
rect 3638 -2724 3644 2652
rect 3678 -2724 3684 2652
rect 3638 -2736 3684 -2724
rect 3752 2652 3798 2664
rect 3752 -2724 3758 2652
rect 3792 -2724 3798 2652
rect 3752 -2736 3798 -2724
rect 4210 2652 4256 2664
rect 4210 -2724 4216 2652
rect 4250 -2724 4256 2652
rect 4210 -2736 4256 -2724
rect 4324 2652 4370 2664
rect 4324 -2724 4330 2652
rect 4364 -2724 4370 2652
rect 4324 -2736 4370 -2724
rect 4782 2652 4828 2664
rect 4782 -2724 4788 2652
rect 4822 -2724 4828 2652
rect 4782 -2736 4828 -2724
rect 4896 2652 4942 2664
rect 4896 -2724 4902 2652
rect 4936 -2724 4942 2652
rect 4896 -2736 4942 -2724
rect 5354 2652 5400 2664
rect 5354 -2724 5360 2652
rect 5394 -2724 5400 2652
rect 5354 -2736 5400 -2724
rect 5468 2652 5514 2664
rect 5468 -2724 5474 2652
rect 5508 -2724 5514 2652
rect 5468 -2736 5514 -2724
rect 5926 2652 5972 2664
rect 5926 -2724 5932 2652
rect 5966 -2724 5972 2652
rect 5926 -2736 5972 -2724
rect 6040 2652 6086 2664
rect 6040 -2724 6046 2652
rect 6080 -2724 6086 2652
rect 6040 -2736 6086 -2724
rect 6498 2652 6544 2664
rect 6498 -2724 6504 2652
rect 6538 -2724 6544 2652
rect 6498 -2736 6544 -2724
rect 6612 2652 6658 2664
rect 6612 -2724 6618 2652
rect 6652 -2724 6658 2652
rect 6612 -2736 6658 -2724
rect 7070 2652 7116 2664
rect 7070 -2724 7076 2652
rect 7110 -2724 7116 2652
rect 7070 -2736 7116 -2724
rect 7184 2652 7230 2664
rect 7184 -2724 7190 2652
rect 7224 -2724 7230 2652
rect 7184 -2736 7230 -2724
rect 7642 2652 7688 2664
rect 7642 -2724 7648 2652
rect 7682 -2724 7688 2652
rect 7642 -2736 7688 -2724
rect 7756 2652 7802 2664
rect 7756 -2724 7762 2652
rect 7796 -2724 7802 2652
rect 7756 -2736 7802 -2724
rect 8214 2652 8260 2664
rect 8214 -2724 8220 2652
rect 8254 -2724 8260 2652
rect 8214 -2736 8260 -2724
rect 8328 2652 8374 2664
rect 8328 -2724 8334 2652
rect 8368 -2724 8374 2652
rect 8328 -2736 8374 -2724
rect 8786 2652 8832 2664
rect 8786 -2724 8792 2652
rect 8826 -2724 8832 2652
rect 8786 -2736 8832 -2724
rect 8900 2652 8946 2664
rect 8900 -2724 8906 2652
rect 8940 -2724 8946 2652
rect 8900 -2736 8946 -2724
rect 9358 2652 9404 2664
rect 9358 -2724 9364 2652
rect 9398 -2724 9404 2652
rect 9358 -2736 9404 -2724
rect 9472 2652 9518 2664
rect 9472 -2724 9478 2652
rect 9512 -2724 9518 2652
rect 9472 -2736 9518 -2724
rect 9930 2652 9976 2664
rect 9930 -2724 9936 2652
rect 9970 -2724 9976 2652
rect 9930 -2736 9976 -2724
rect 10044 2652 10090 2664
rect 10044 -2724 10050 2652
rect 10084 -2724 10090 2652
rect 10044 -2736 10090 -2724
rect 10502 2652 10548 2664
rect 10502 -2724 10508 2652
rect 10542 -2724 10548 2652
rect 10502 -2736 10548 -2724
rect 10616 2652 10662 2664
rect 10616 -2724 10622 2652
rect 10656 -2724 10662 2652
rect 10616 -2736 10662 -2724
rect 11074 2652 11120 2664
rect 11074 -2724 11080 2652
rect 11114 -2724 11120 2652
rect 11074 -2736 11120 -2724
rect 11188 2652 11234 2664
rect 11188 -2724 11194 2652
rect 11228 -2724 11234 2652
rect 11188 -2736 11234 -2724
rect 11646 2652 11692 2664
rect 11646 -2724 11652 2652
rect 11686 -2724 11692 2652
rect 11646 -2736 11692 -2724
rect 11760 2652 11806 2664
rect 11760 -2724 11766 2652
rect 11800 -2724 11806 2652
rect 11760 -2736 11806 -2724
rect 12218 2652 12264 2664
rect 12218 -2724 12224 2652
rect 12258 -2724 12264 2652
rect 12218 -2736 12264 -2724
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 27 l 2 m 1 nf 43 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
