magic
tech sky130A
magscale 1 2
timestamp 1620318829
<< nwell >>
rect -812 -419 812 419
<< pmos >>
rect -616 -200 -416 200
rect -358 -200 -158 200
rect -100 -200 100 200
rect 158 -200 358 200
rect 416 -200 616 200
<< pdiff >>
rect -674 188 -616 200
rect -674 -188 -662 188
rect -628 -188 -616 188
rect -674 -200 -616 -188
rect -416 188 -358 200
rect -416 -188 -404 188
rect -370 -188 -358 188
rect -416 -200 -358 -188
rect -158 188 -100 200
rect -158 -188 -146 188
rect -112 -188 -100 188
rect -158 -200 -100 -188
rect 100 188 158 200
rect 100 -188 112 188
rect 146 -188 158 188
rect 100 -200 158 -188
rect 358 188 416 200
rect 358 -188 370 188
rect 404 -188 416 188
rect 358 -200 416 -188
rect 616 188 674 200
rect 616 -188 628 188
rect 662 -188 674 188
rect 616 -200 674 -188
<< pdiffc >>
rect -662 -188 -628 188
rect -404 -188 -370 188
rect -146 -188 -112 188
rect 112 -188 146 188
rect 370 -188 404 188
rect 628 -188 662 188
<< nsubdiff >>
rect -776 349 -680 383
rect 680 349 776 383
rect -776 287 -742 349
rect 742 287 776 349
rect -776 -349 -742 -287
rect 742 -349 776 -287
rect -776 -383 -680 -349
rect 680 -383 776 -349
<< nsubdiffcont >>
rect -680 349 680 383
rect -776 -287 -742 287
rect 742 -287 776 287
rect -680 -383 680 -349
<< poly >>
rect -616 281 -416 297
rect -616 247 -600 281
rect -432 247 -416 281
rect -616 200 -416 247
rect -358 281 -158 297
rect -358 247 -342 281
rect -174 247 -158 281
rect -358 200 -158 247
rect -100 281 100 297
rect -100 247 -84 281
rect 84 247 100 281
rect -100 200 100 247
rect 158 281 358 297
rect 158 247 174 281
rect 342 247 358 281
rect 158 200 358 247
rect 416 281 616 297
rect 416 247 432 281
rect 600 247 616 281
rect 416 200 616 247
rect -616 -247 -416 -200
rect -616 -281 -600 -247
rect -432 -281 -416 -247
rect -616 -297 -416 -281
rect -358 -247 -158 -200
rect -358 -281 -342 -247
rect -174 -281 -158 -247
rect -358 -297 -158 -281
rect -100 -247 100 -200
rect -100 -281 -84 -247
rect 84 -281 100 -247
rect -100 -297 100 -281
rect 158 -247 358 -200
rect 158 -281 174 -247
rect 342 -281 358 -247
rect 158 -297 358 -281
rect 416 -247 616 -200
rect 416 -281 432 -247
rect 600 -281 616 -247
rect 416 -297 616 -281
<< polycont >>
rect -600 247 -432 281
rect -342 247 -174 281
rect -84 247 84 281
rect 174 247 342 281
rect 432 247 600 281
rect -600 -281 -432 -247
rect -342 -281 -174 -247
rect -84 -281 84 -247
rect 174 -281 342 -247
rect 432 -281 600 -247
<< locali >>
rect -776 349 -680 383
rect 680 349 776 383
rect -776 287 -742 349
rect 742 287 776 349
rect -616 247 -600 281
rect -432 247 -416 281
rect -358 247 -342 281
rect -174 247 -158 281
rect -100 247 -84 281
rect 84 247 100 281
rect 158 247 174 281
rect 342 247 358 281
rect 416 247 432 281
rect 600 247 616 281
rect -662 188 -628 204
rect -662 -204 -628 -188
rect -404 188 -370 204
rect -404 -204 -370 -188
rect -146 188 -112 204
rect -146 -204 -112 -188
rect 112 188 146 204
rect 112 -204 146 -188
rect 370 188 404 204
rect 370 -204 404 -188
rect 628 188 662 204
rect 628 -204 662 -188
rect -616 -281 -600 -247
rect -432 -281 -416 -247
rect -358 -281 -342 -247
rect -174 -281 -158 -247
rect -100 -281 -84 -247
rect 84 -281 100 -247
rect 158 -281 174 -247
rect 342 -281 358 -247
rect 416 -281 432 -247
rect 600 -281 616 -247
rect -776 -349 -742 -287
rect 742 -349 776 -287
rect -776 -383 -680 -349
rect 680 -383 776 -349
<< viali >>
rect -600 247 -432 281
rect -342 247 -174 281
rect -84 247 84 281
rect 174 247 342 281
rect 432 247 600 281
rect -662 -188 -628 188
rect -404 -188 -370 188
rect -146 -188 -112 188
rect 112 -188 146 188
rect 370 -188 404 188
rect 628 -188 662 188
rect -600 -281 -432 -247
rect -342 -281 -174 -247
rect -84 -281 84 -247
rect 174 -281 342 -247
rect 432 -281 600 -247
<< metal1 >>
rect -612 281 -420 287
rect -612 247 -600 281
rect -432 247 -420 281
rect -612 241 -420 247
rect -354 281 -162 287
rect -354 247 -342 281
rect -174 247 -162 281
rect -354 241 -162 247
rect -96 281 96 287
rect -96 247 -84 281
rect 84 247 96 281
rect -96 241 96 247
rect 162 281 354 287
rect 162 247 174 281
rect 342 247 354 281
rect 162 241 354 247
rect 420 281 612 287
rect 420 247 432 281
rect 600 247 612 281
rect 420 241 612 247
rect -668 188 -622 200
rect -668 -188 -662 188
rect -628 -188 -622 188
rect -668 -200 -622 -188
rect -410 188 -364 200
rect -410 -188 -404 188
rect -370 -188 -364 188
rect -410 -200 -364 -188
rect -152 188 -106 200
rect -152 -188 -146 188
rect -112 -188 -106 188
rect -152 -200 -106 -188
rect 106 188 152 200
rect 106 -188 112 188
rect 146 -188 152 188
rect 106 -200 152 -188
rect 364 188 410 200
rect 364 -188 370 188
rect 404 -188 410 188
rect 364 -200 410 -188
rect 622 188 668 200
rect 622 -188 628 188
rect 662 -188 668 188
rect 622 -200 668 -188
rect -612 -247 -420 -241
rect -612 -281 -600 -247
rect -432 -281 -420 -247
rect -612 -287 -420 -281
rect -354 -247 -162 -241
rect -354 -281 -342 -247
rect -174 -281 -162 -247
rect -354 -287 -162 -281
rect -96 -247 96 -241
rect -96 -281 -84 -247
rect 84 -281 96 -247
rect -96 -287 96 -281
rect 162 -247 354 -241
rect 162 -281 174 -247
rect 342 -281 354 -247
rect 162 -287 354 -281
rect 420 -247 612 -241
rect 420 -281 432 -247
rect 600 -281 612 -247
rect 420 -287 612 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -759 -366 759 366
string parameters w 2 l 1 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
