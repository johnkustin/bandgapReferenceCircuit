magic
tech sky130A
magscale 1 2
timestamp 1620926822
<< error_p >>
rect -487 -231 -429 169
rect -29 -231 29 169
rect 429 -231 487 169
<< nmoslvt >>
rect -429 -231 -29 169
rect 29 -231 429 169
<< ndiff >>
rect -487 157 -429 169
rect -487 -219 -475 157
rect -441 -219 -429 157
rect -487 -231 -429 -219
rect -29 157 29 169
rect -29 -219 -17 157
rect 17 -219 29 157
rect -29 -231 29 -219
rect 429 157 487 169
rect 429 -219 441 157
rect 475 -219 487 157
rect 429 -231 487 -219
<< ndiffc >>
rect -475 -219 -441 157
rect -17 -219 17 157
rect 441 -219 475 157
<< poly >>
rect -429 241 -29 257
rect -429 207 -413 241
rect -45 207 -29 241
rect -429 169 -29 207
rect 29 241 429 257
rect 29 207 45 241
rect 413 207 429 241
rect 29 169 429 207
rect -429 -257 -29 -231
rect 29 -257 429 -231
<< polycont >>
rect -413 207 -45 241
rect 45 207 413 241
<< locali >>
rect -429 207 -413 241
rect -45 207 -29 241
rect 29 207 45 241
rect 413 207 429 241
rect -475 157 -441 173
rect -475 -235 -441 -219
rect -17 157 17 173
rect -17 -235 17 -219
rect 441 157 475 173
rect 441 -235 475 -219
<< viali >>
rect -413 207 -45 241
rect 45 207 413 241
rect -475 -219 -441 157
rect -17 -219 17 157
rect 441 -219 475 157
<< metal1 >>
rect -425 241 -33 247
rect -425 207 -413 241
rect -45 207 -33 241
rect -425 201 -33 207
rect 33 241 425 247
rect 33 207 45 241
rect 413 207 425 241
rect 33 201 425 207
rect -481 157 -435 169
rect -481 -219 -475 157
rect -441 -219 -435 157
rect -481 -231 -435 -219
rect -23 157 23 169
rect -23 -219 -17 157
rect 17 -219 23 157
rect -23 -231 23 -219
rect 435 157 481 169
rect 435 -219 441 157
rect 475 -219 481 157
rect 435 -231 481 -219
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 2 l 2 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
