magic
tech sky130A
magscale 1 2
timestamp 1622081478
<< nwell >>
rect -992 -497 992 497
<< mvpmos >>
rect -734 -200 -574 200
rect -516 -200 -356 200
rect -298 -200 -138 200
rect -80 -200 80 200
rect 138 -200 298 200
rect 356 -200 516 200
rect 574 -200 734 200
<< mvpdiff >>
rect -792 187 -734 200
rect -792 153 -780 187
rect -746 153 -734 187
rect -792 119 -734 153
rect -792 85 -780 119
rect -746 85 -734 119
rect -792 51 -734 85
rect -792 17 -780 51
rect -746 17 -734 51
rect -792 -17 -734 17
rect -792 -51 -780 -17
rect -746 -51 -734 -17
rect -792 -85 -734 -51
rect -792 -119 -780 -85
rect -746 -119 -734 -85
rect -792 -153 -734 -119
rect -792 -187 -780 -153
rect -746 -187 -734 -153
rect -792 -200 -734 -187
rect -574 187 -516 200
rect -574 153 -562 187
rect -528 153 -516 187
rect -574 119 -516 153
rect -574 85 -562 119
rect -528 85 -516 119
rect -574 51 -516 85
rect -574 17 -562 51
rect -528 17 -516 51
rect -574 -17 -516 17
rect -574 -51 -562 -17
rect -528 -51 -516 -17
rect -574 -85 -516 -51
rect -574 -119 -562 -85
rect -528 -119 -516 -85
rect -574 -153 -516 -119
rect -574 -187 -562 -153
rect -528 -187 -516 -153
rect -574 -200 -516 -187
rect -356 187 -298 200
rect -356 153 -344 187
rect -310 153 -298 187
rect -356 119 -298 153
rect -356 85 -344 119
rect -310 85 -298 119
rect -356 51 -298 85
rect -356 17 -344 51
rect -310 17 -298 51
rect -356 -17 -298 17
rect -356 -51 -344 -17
rect -310 -51 -298 -17
rect -356 -85 -298 -51
rect -356 -119 -344 -85
rect -310 -119 -298 -85
rect -356 -153 -298 -119
rect -356 -187 -344 -153
rect -310 -187 -298 -153
rect -356 -200 -298 -187
rect -138 187 -80 200
rect -138 153 -126 187
rect -92 153 -80 187
rect -138 119 -80 153
rect -138 85 -126 119
rect -92 85 -80 119
rect -138 51 -80 85
rect -138 17 -126 51
rect -92 17 -80 51
rect -138 -17 -80 17
rect -138 -51 -126 -17
rect -92 -51 -80 -17
rect -138 -85 -80 -51
rect -138 -119 -126 -85
rect -92 -119 -80 -85
rect -138 -153 -80 -119
rect -138 -187 -126 -153
rect -92 -187 -80 -153
rect -138 -200 -80 -187
rect 80 187 138 200
rect 80 153 92 187
rect 126 153 138 187
rect 80 119 138 153
rect 80 85 92 119
rect 126 85 138 119
rect 80 51 138 85
rect 80 17 92 51
rect 126 17 138 51
rect 80 -17 138 17
rect 80 -51 92 -17
rect 126 -51 138 -17
rect 80 -85 138 -51
rect 80 -119 92 -85
rect 126 -119 138 -85
rect 80 -153 138 -119
rect 80 -187 92 -153
rect 126 -187 138 -153
rect 80 -200 138 -187
rect 298 187 356 200
rect 298 153 310 187
rect 344 153 356 187
rect 298 119 356 153
rect 298 85 310 119
rect 344 85 356 119
rect 298 51 356 85
rect 298 17 310 51
rect 344 17 356 51
rect 298 -17 356 17
rect 298 -51 310 -17
rect 344 -51 356 -17
rect 298 -85 356 -51
rect 298 -119 310 -85
rect 344 -119 356 -85
rect 298 -153 356 -119
rect 298 -187 310 -153
rect 344 -187 356 -153
rect 298 -200 356 -187
rect 516 187 574 200
rect 516 153 528 187
rect 562 153 574 187
rect 516 119 574 153
rect 516 85 528 119
rect 562 85 574 119
rect 516 51 574 85
rect 516 17 528 51
rect 562 17 574 51
rect 516 -17 574 17
rect 516 -51 528 -17
rect 562 -51 574 -17
rect 516 -85 574 -51
rect 516 -119 528 -85
rect 562 -119 574 -85
rect 516 -153 574 -119
rect 516 -187 528 -153
rect 562 -187 574 -153
rect 516 -200 574 -187
rect 734 187 792 200
rect 734 153 746 187
rect 780 153 792 187
rect 734 119 792 153
rect 734 85 746 119
rect 780 85 792 119
rect 734 51 792 85
rect 734 17 746 51
rect 780 17 792 51
rect 734 -17 792 17
rect 734 -51 746 -17
rect 780 -51 792 -17
rect 734 -85 792 -51
rect 734 -119 746 -85
rect 780 -119 792 -85
rect 734 -153 792 -119
rect 734 -187 746 -153
rect 780 -187 792 -153
rect 734 -200 792 -187
<< mvpdiffc >>
rect -780 153 -746 187
rect -780 85 -746 119
rect -780 17 -746 51
rect -780 -51 -746 -17
rect -780 -119 -746 -85
rect -780 -187 -746 -153
rect -562 153 -528 187
rect -562 85 -528 119
rect -562 17 -528 51
rect -562 -51 -528 -17
rect -562 -119 -528 -85
rect -562 -187 -528 -153
rect -344 153 -310 187
rect -344 85 -310 119
rect -344 17 -310 51
rect -344 -51 -310 -17
rect -344 -119 -310 -85
rect -344 -187 -310 -153
rect -126 153 -92 187
rect -126 85 -92 119
rect -126 17 -92 51
rect -126 -51 -92 -17
rect -126 -119 -92 -85
rect -126 -187 -92 -153
rect 92 153 126 187
rect 92 85 126 119
rect 92 17 126 51
rect 92 -51 126 -17
rect 92 -119 126 -85
rect 92 -187 126 -153
rect 310 153 344 187
rect 310 85 344 119
rect 310 17 344 51
rect 310 -51 344 -17
rect 310 -119 344 -85
rect 310 -187 344 -153
rect 528 153 562 187
rect 528 85 562 119
rect 528 17 562 51
rect 528 -51 562 -17
rect 528 -119 562 -85
rect 528 -187 562 -153
rect 746 153 780 187
rect 746 85 780 119
rect 746 17 780 51
rect 746 -51 780 -17
rect 746 -119 780 -85
rect 746 -187 780 -153
<< mvnsubdiff >>
rect -926 419 926 431
rect -926 385 -799 419
rect -765 385 -731 419
rect -697 385 -663 419
rect -629 385 -595 419
rect -561 385 -527 419
rect -493 385 -459 419
rect -425 385 -391 419
rect -357 385 -323 419
rect -289 385 -255 419
rect -221 385 -187 419
rect -153 385 -119 419
rect -85 385 -51 419
rect -17 385 17 419
rect 51 385 85 419
rect 119 385 153 419
rect 187 385 221 419
rect 255 385 289 419
rect 323 385 357 419
rect 391 385 425 419
rect 459 385 493 419
rect 527 385 561 419
rect 595 385 629 419
rect 663 385 697 419
rect 731 385 765 419
rect 799 385 926 419
rect -926 373 926 385
rect -926 323 -868 373
rect -926 289 -914 323
rect -880 289 -868 323
rect 868 323 926 373
rect -926 255 -868 289
rect -926 221 -914 255
rect -880 221 -868 255
rect -926 187 -868 221
rect 868 289 880 323
rect 914 289 926 323
rect 868 255 926 289
rect 868 221 880 255
rect 914 221 926 255
rect -926 153 -914 187
rect -880 153 -868 187
rect -926 119 -868 153
rect -926 85 -914 119
rect -880 85 -868 119
rect -926 51 -868 85
rect -926 17 -914 51
rect -880 17 -868 51
rect -926 -17 -868 17
rect -926 -51 -914 -17
rect -880 -51 -868 -17
rect -926 -85 -868 -51
rect -926 -119 -914 -85
rect -880 -119 -868 -85
rect -926 -153 -868 -119
rect -926 -187 -914 -153
rect -880 -187 -868 -153
rect -926 -221 -868 -187
rect 868 187 926 221
rect 868 153 880 187
rect 914 153 926 187
rect 868 119 926 153
rect 868 85 880 119
rect 914 85 926 119
rect 868 51 926 85
rect 868 17 880 51
rect 914 17 926 51
rect 868 -17 926 17
rect 868 -51 880 -17
rect 914 -51 926 -17
rect 868 -85 926 -51
rect 868 -119 880 -85
rect 914 -119 926 -85
rect 868 -153 926 -119
rect 868 -187 880 -153
rect 914 -187 926 -153
rect -926 -255 -914 -221
rect -880 -255 -868 -221
rect -926 -289 -868 -255
rect -926 -323 -914 -289
rect -880 -323 -868 -289
rect 868 -221 926 -187
rect 868 -255 880 -221
rect 914 -255 926 -221
rect 868 -289 926 -255
rect -926 -373 -868 -323
rect 868 -323 880 -289
rect 914 -323 926 -289
rect 868 -373 926 -323
rect -926 -385 926 -373
rect -926 -419 -799 -385
rect -765 -419 -731 -385
rect -697 -419 -663 -385
rect -629 -419 -595 -385
rect -561 -419 -527 -385
rect -493 -419 -459 -385
rect -425 -419 -391 -385
rect -357 -419 -323 -385
rect -289 -419 -255 -385
rect -221 -419 -187 -385
rect -153 -419 -119 -385
rect -85 -419 -51 -385
rect -17 -419 17 -385
rect 51 -419 85 -385
rect 119 -419 153 -385
rect 187 -419 221 -385
rect 255 -419 289 -385
rect 323 -419 357 -385
rect 391 -419 425 -385
rect 459 -419 493 -385
rect 527 -419 561 -385
rect 595 -419 629 -385
rect 663 -419 697 -385
rect 731 -419 765 -385
rect 799 -419 926 -385
rect -926 -431 926 -419
<< mvnsubdiffcont >>
rect -799 385 -765 419
rect -731 385 -697 419
rect -663 385 -629 419
rect -595 385 -561 419
rect -527 385 -493 419
rect -459 385 -425 419
rect -391 385 -357 419
rect -323 385 -289 419
rect -255 385 -221 419
rect -187 385 -153 419
rect -119 385 -85 419
rect -51 385 -17 419
rect 17 385 51 419
rect 85 385 119 419
rect 153 385 187 419
rect 221 385 255 419
rect 289 385 323 419
rect 357 385 391 419
rect 425 385 459 419
rect 493 385 527 419
rect 561 385 595 419
rect 629 385 663 419
rect 697 385 731 419
rect 765 385 799 419
rect -914 289 -880 323
rect -914 221 -880 255
rect 880 289 914 323
rect 880 221 914 255
rect -914 153 -880 187
rect -914 85 -880 119
rect -914 17 -880 51
rect -914 -51 -880 -17
rect -914 -119 -880 -85
rect -914 -187 -880 -153
rect 880 153 914 187
rect 880 85 914 119
rect 880 17 914 51
rect 880 -51 914 -17
rect 880 -119 914 -85
rect 880 -187 914 -153
rect -914 -255 -880 -221
rect -914 -323 -880 -289
rect 880 -255 914 -221
rect 880 -323 914 -289
rect -799 -419 -765 -385
rect -731 -419 -697 -385
rect -663 -419 -629 -385
rect -595 -419 -561 -385
rect -527 -419 -493 -385
rect -459 -419 -425 -385
rect -391 -419 -357 -385
rect -323 -419 -289 -385
rect -255 -419 -221 -385
rect -187 -419 -153 -385
rect -119 -419 -85 -385
rect -51 -419 -17 -385
rect 17 -419 51 -385
rect 85 -419 119 -385
rect 153 -419 187 -385
rect 221 -419 255 -385
rect 289 -419 323 -385
rect 357 -419 391 -385
rect 425 -419 459 -385
rect 493 -419 527 -385
rect 561 -419 595 -385
rect 629 -419 663 -385
rect 697 -419 731 -385
rect 765 -419 799 -385
<< poly >>
rect -734 281 -574 297
rect -734 247 -705 281
rect -671 247 -637 281
rect -603 247 -574 281
rect -734 200 -574 247
rect -516 281 -356 297
rect -516 247 -487 281
rect -453 247 -419 281
rect -385 247 -356 281
rect -516 200 -356 247
rect -298 281 -138 297
rect -298 247 -269 281
rect -235 247 -201 281
rect -167 247 -138 281
rect -298 200 -138 247
rect -80 281 80 297
rect -80 247 -51 281
rect -17 247 17 281
rect 51 247 80 281
rect -80 200 80 247
rect 138 281 298 297
rect 138 247 167 281
rect 201 247 235 281
rect 269 247 298 281
rect 138 200 298 247
rect 356 281 516 297
rect 356 247 385 281
rect 419 247 453 281
rect 487 247 516 281
rect 356 200 516 247
rect 574 281 734 297
rect 574 247 603 281
rect 637 247 671 281
rect 705 247 734 281
rect 574 200 734 247
rect -734 -247 -574 -200
rect -734 -281 -705 -247
rect -671 -281 -637 -247
rect -603 -281 -574 -247
rect -734 -297 -574 -281
rect -516 -247 -356 -200
rect -516 -281 -487 -247
rect -453 -281 -419 -247
rect -385 -281 -356 -247
rect -516 -297 -356 -281
rect -298 -247 -138 -200
rect -298 -281 -269 -247
rect -235 -281 -201 -247
rect -167 -281 -138 -247
rect -298 -297 -138 -281
rect -80 -247 80 -200
rect -80 -281 -51 -247
rect -17 -281 17 -247
rect 51 -281 80 -247
rect -80 -297 80 -281
rect 138 -247 298 -200
rect 138 -281 167 -247
rect 201 -281 235 -247
rect 269 -281 298 -247
rect 138 -297 298 -281
rect 356 -247 516 -200
rect 356 -281 385 -247
rect 419 -281 453 -247
rect 487 -281 516 -247
rect 356 -297 516 -281
rect 574 -247 734 -200
rect 574 -281 603 -247
rect 637 -281 671 -247
rect 705 -281 734 -247
rect 574 -297 734 -281
<< polycont >>
rect -705 247 -671 281
rect -637 247 -603 281
rect -487 247 -453 281
rect -419 247 -385 281
rect -269 247 -235 281
rect -201 247 -167 281
rect -51 247 -17 281
rect 17 247 51 281
rect 167 247 201 281
rect 235 247 269 281
rect 385 247 419 281
rect 453 247 487 281
rect 603 247 637 281
rect 671 247 705 281
rect -705 -281 -671 -247
rect -637 -281 -603 -247
rect -487 -281 -453 -247
rect -419 -281 -385 -247
rect -269 -281 -235 -247
rect -201 -281 -167 -247
rect -51 -281 -17 -247
rect 17 -281 51 -247
rect 167 -281 201 -247
rect 235 -281 269 -247
rect 385 -281 419 -247
rect 453 -281 487 -247
rect 603 -281 637 -247
rect 671 -281 705 -247
<< locali >>
rect -914 385 -799 419
rect -739 385 -731 419
rect -667 385 -663 419
rect -561 385 -557 419
rect -493 385 -485 419
rect -425 385 -413 419
rect -357 385 -341 419
rect -289 385 -269 419
rect -221 385 -197 419
rect -153 385 -125 419
rect -85 385 -53 419
rect -17 385 17 419
rect 53 385 85 419
rect 125 385 153 419
rect 197 385 221 419
rect 269 385 289 419
rect 341 385 357 419
rect 413 385 425 419
rect 485 385 493 419
rect 557 385 561 419
rect 663 385 667 419
rect 731 385 739 419
rect 799 385 914 419
rect -914 372 -880 385
rect -914 323 -880 338
rect 880 323 914 385
rect -914 255 -880 266
rect -734 247 -707 281
rect -671 247 -637 281
rect -601 247 -574 281
rect -516 247 -489 281
rect -453 247 -419 281
rect -383 247 -356 281
rect -298 247 -271 281
rect -235 247 -201 281
rect -165 247 -138 281
rect -80 247 -53 281
rect -17 247 17 281
rect 53 247 80 281
rect 138 247 165 281
rect 201 247 235 281
rect 271 247 298 281
rect 356 247 383 281
rect 419 247 453 281
rect 489 247 516 281
rect 574 247 601 281
rect 637 247 671 281
rect 707 247 734 281
rect 880 255 914 289
rect -914 187 -880 194
rect -914 119 -880 122
rect -914 84 -880 85
rect -914 -17 -880 17
rect -914 -85 -880 -51
rect -914 -153 -880 -119
rect -914 -221 -880 -187
rect -780 187 -746 204
rect -780 149 -746 153
rect -780 77 -746 85
rect -780 -17 -746 17
rect -780 -85 -746 -51
rect -780 -153 -746 -119
rect -780 -204 -746 -187
rect -562 187 -528 204
rect -562 119 -528 153
rect -562 51 -528 85
rect -562 -17 -528 17
rect -562 -85 -528 -77
rect -562 -153 -528 -149
rect -562 -204 -528 -187
rect -344 187 -310 204
rect -344 149 -310 153
rect -344 77 -310 85
rect -344 -17 -310 17
rect -344 -85 -310 -51
rect -344 -153 -310 -119
rect -344 -204 -310 -187
rect -126 187 -92 204
rect -126 119 -92 153
rect -126 51 -92 85
rect -126 -17 -92 17
rect -126 -85 -92 -77
rect -126 -153 -92 -149
rect -126 -204 -92 -187
rect 92 187 126 204
rect 92 149 126 153
rect 92 77 126 85
rect 92 -17 126 17
rect 92 -85 126 -51
rect 92 -153 126 -119
rect 92 -204 126 -187
rect 310 187 344 204
rect 310 119 344 153
rect 310 51 344 85
rect 310 -17 344 17
rect 310 -85 344 -77
rect 310 -153 344 -149
rect 310 -204 344 -187
rect 528 187 562 204
rect 528 149 562 153
rect 528 77 562 85
rect 528 -17 562 17
rect 528 -85 562 -51
rect 528 -153 562 -119
rect 528 -204 562 -187
rect 746 187 780 204
rect 746 119 780 153
rect 746 51 780 85
rect 746 -17 780 17
rect 746 -85 780 -77
rect 746 -153 780 -149
rect 746 -204 780 -187
rect 880 187 914 221
rect 880 119 914 153
rect 880 51 914 85
rect 880 -17 914 17
rect 880 -85 914 -51
rect 880 -153 914 -119
rect 880 -221 914 -187
rect -914 -289 -880 -255
rect -734 -281 -707 -247
rect -671 -281 -637 -247
rect -601 -281 -574 -247
rect -516 -281 -489 -247
rect -453 -281 -419 -247
rect -383 -281 -356 -247
rect -298 -281 -271 -247
rect -235 -281 -201 -247
rect -165 -281 -138 -247
rect -80 -281 -53 -247
rect -17 -281 17 -247
rect 53 -281 80 -247
rect 138 -281 165 -247
rect 201 -281 235 -247
rect 271 -281 298 -247
rect 356 -281 383 -247
rect 419 -281 453 -247
rect 489 -281 516 -247
rect 574 -281 601 -247
rect 637 -281 671 -247
rect 707 -281 734 -247
rect -914 -385 -880 -323
rect 880 -289 914 -255
rect 880 -385 914 -323
rect -914 -419 -799 -385
rect -765 -419 -731 -385
rect -697 -419 -663 -385
rect -629 -419 -595 -385
rect -561 -419 -527 -385
rect -493 -419 -459 -385
rect -425 -419 -391 -385
rect -357 -419 -323 -385
rect -289 -419 -255 -385
rect -221 -419 -187 -385
rect -153 -419 -119 -385
rect -85 -419 -51 -385
rect -17 -419 17 -385
rect 51 -419 85 -385
rect 119 -419 153 -385
rect 187 -419 221 -385
rect 255 -419 289 -385
rect 323 -419 357 -385
rect 391 -419 425 -385
rect 459 -419 493 -385
rect 527 -419 561 -385
rect 595 -419 629 -385
rect 663 -419 697 -385
rect 731 -419 765 -385
rect 799 -419 914 -385
<< viali >>
rect -773 385 -765 419
rect -765 385 -739 419
rect -701 385 -697 419
rect -697 385 -667 419
rect -629 385 -595 419
rect -557 385 -527 419
rect -527 385 -523 419
rect -485 385 -459 419
rect -459 385 -451 419
rect -413 385 -391 419
rect -391 385 -379 419
rect -341 385 -323 419
rect -323 385 -307 419
rect -269 385 -255 419
rect -255 385 -235 419
rect -197 385 -187 419
rect -187 385 -163 419
rect -125 385 -119 419
rect -119 385 -91 419
rect -53 385 -51 419
rect -51 385 -19 419
rect 19 385 51 419
rect 51 385 53 419
rect 91 385 119 419
rect 119 385 125 419
rect 163 385 187 419
rect 187 385 197 419
rect 235 385 255 419
rect 255 385 269 419
rect 307 385 323 419
rect 323 385 341 419
rect 379 385 391 419
rect 391 385 413 419
rect 451 385 459 419
rect 459 385 485 419
rect 523 385 527 419
rect 527 385 557 419
rect 595 385 629 419
rect 667 385 697 419
rect 697 385 701 419
rect 739 385 765 419
rect 765 385 773 419
rect -914 338 -880 372
rect -914 289 -880 300
rect -914 266 -880 289
rect -707 247 -705 281
rect -705 247 -673 281
rect -635 247 -603 281
rect -603 247 -601 281
rect -489 247 -487 281
rect -487 247 -455 281
rect -417 247 -385 281
rect -385 247 -383 281
rect -271 247 -269 281
rect -269 247 -237 281
rect -199 247 -167 281
rect -167 247 -165 281
rect -53 247 -51 281
rect -51 247 -19 281
rect 19 247 51 281
rect 51 247 53 281
rect 165 247 167 281
rect 167 247 199 281
rect 237 247 269 281
rect 269 247 271 281
rect 383 247 385 281
rect 385 247 417 281
rect 455 247 487 281
rect 487 247 489 281
rect 601 247 603 281
rect 603 247 635 281
rect 673 247 705 281
rect 705 247 707 281
rect -914 221 -880 228
rect -914 194 -880 221
rect -914 153 -880 156
rect -914 122 -880 153
rect -914 51 -880 84
rect -914 50 -880 51
rect -780 119 -746 149
rect -780 115 -746 119
rect -780 51 -746 77
rect -780 43 -746 51
rect -562 -51 -528 -43
rect -562 -77 -528 -51
rect -562 -119 -528 -115
rect -562 -149 -528 -119
rect -344 119 -310 149
rect -344 115 -310 119
rect -344 51 -310 77
rect -344 43 -310 51
rect -126 -51 -92 -43
rect -126 -77 -92 -51
rect -126 -119 -92 -115
rect -126 -149 -92 -119
rect 92 119 126 149
rect 92 115 126 119
rect 92 51 126 77
rect 92 43 126 51
rect 310 -51 344 -43
rect 310 -77 344 -51
rect 310 -119 344 -115
rect 310 -149 344 -119
rect 528 119 562 149
rect 528 115 562 119
rect 528 51 562 77
rect 528 43 562 51
rect 746 -51 780 -43
rect 746 -77 780 -51
rect 746 -119 780 -115
rect 746 -149 780 -119
rect -707 -281 -705 -247
rect -705 -281 -673 -247
rect -635 -281 -603 -247
rect -603 -281 -601 -247
rect -489 -281 -487 -247
rect -487 -281 -455 -247
rect -417 -281 -385 -247
rect -385 -281 -383 -247
rect -271 -281 -269 -247
rect -269 -281 -237 -247
rect -199 -281 -167 -247
rect -167 -281 -165 -247
rect -53 -281 -51 -247
rect -51 -281 -19 -247
rect 19 -281 51 -247
rect 51 -281 53 -247
rect 165 -281 167 -247
rect 167 -281 199 -247
rect 237 -281 269 -247
rect 269 -281 271 -247
rect 383 -281 385 -247
rect 385 -281 417 -247
rect 455 -281 487 -247
rect 487 -281 489 -247
rect 601 -281 603 -247
rect 603 -281 635 -247
rect 673 -281 705 -247
rect 705 -281 707 -247
<< metal1 >>
rect -804 419 804 425
rect -920 372 -874 397
rect -804 385 -773 419
rect -739 385 -701 419
rect -667 385 -629 419
rect -595 385 -557 419
rect -523 385 -485 419
rect -451 385 -413 419
rect -379 385 -341 419
rect -307 385 -269 419
rect -235 385 -197 419
rect -163 385 -125 419
rect -91 385 -53 419
rect -19 385 19 419
rect 53 385 91 419
rect 125 385 163 419
rect 197 385 235 419
rect 269 385 307 419
rect 341 385 379 419
rect 413 385 451 419
rect 485 385 523 419
rect 557 385 595 419
rect 629 385 667 419
rect 701 385 739 419
rect 773 385 804 419
rect -804 379 804 385
rect -920 338 -914 372
rect -880 338 -874 372
rect -920 300 -874 338
rect -920 266 -914 300
rect -880 266 -874 300
rect -920 228 -874 266
rect -730 281 -578 287
rect -730 247 -707 281
rect -673 247 -635 281
rect -601 247 -578 281
rect -730 241 -578 247
rect -512 281 -360 287
rect -512 247 -489 281
rect -455 247 -417 281
rect -383 247 -360 281
rect -512 241 -360 247
rect -294 281 -142 287
rect -294 247 -271 281
rect -237 247 -199 281
rect -165 247 -142 281
rect -294 241 -142 247
rect -76 281 76 287
rect -76 247 -53 281
rect -19 247 19 281
rect 53 247 76 281
rect -76 241 76 247
rect 142 281 294 287
rect 142 247 165 281
rect 199 247 237 281
rect 271 247 294 281
rect 142 241 294 247
rect 360 281 512 287
rect 360 247 383 281
rect 417 247 455 281
rect 489 247 512 281
rect 360 241 512 247
rect 578 281 730 287
rect 578 247 601 281
rect 635 247 673 281
rect 707 247 730 281
rect 578 241 730 247
rect -920 194 -914 228
rect -880 194 -874 228
rect -920 156 -874 194
rect -920 122 -914 156
rect -880 122 -874 156
rect -920 84 -874 122
rect -920 50 -914 84
rect -880 50 -874 84
rect -920 26 -874 50
rect -786 149 -740 183
rect -786 115 -780 149
rect -746 115 -740 149
rect -786 77 -740 115
rect -786 43 -780 77
rect -746 43 -740 77
rect -786 9 -740 43
rect -350 149 -304 183
rect -350 115 -344 149
rect -310 115 -304 149
rect -350 77 -304 115
rect -350 43 -344 77
rect -310 43 -304 77
rect -350 9 -304 43
rect 86 149 132 183
rect 86 115 92 149
rect 126 115 132 149
rect 86 77 132 115
rect 86 43 92 77
rect 126 43 132 77
rect 86 9 132 43
rect 522 149 568 183
rect 522 115 528 149
rect 562 115 568 149
rect 522 77 568 115
rect 522 43 528 77
rect 562 43 568 77
rect 522 9 568 43
rect -568 -43 -522 -9
rect -568 -77 -562 -43
rect -528 -77 -522 -43
rect -568 -115 -522 -77
rect -568 -149 -562 -115
rect -528 -149 -522 -115
rect -568 -183 -522 -149
rect -132 -43 -86 -9
rect -132 -77 -126 -43
rect -92 -77 -86 -43
rect -132 -115 -86 -77
rect -132 -149 -126 -115
rect -92 -149 -86 -115
rect -132 -183 -86 -149
rect 304 -43 350 -9
rect 304 -77 310 -43
rect 344 -77 350 -43
rect 304 -115 350 -77
rect 304 -149 310 -115
rect 344 -149 350 -115
rect 304 -183 350 -149
rect 740 -43 786 -9
rect 740 -77 746 -43
rect 780 -77 786 -43
rect 740 -115 786 -77
rect 740 -149 746 -115
rect 780 -149 786 -115
rect 740 -183 786 -149
rect -730 -247 -578 -241
rect -730 -281 -707 -247
rect -673 -281 -635 -247
rect -601 -281 -578 -247
rect -730 -287 -578 -281
rect -512 -247 -360 -241
rect -512 -281 -489 -247
rect -455 -281 -417 -247
rect -383 -281 -360 -247
rect -512 -287 -360 -281
rect -294 -247 -142 -241
rect -294 -281 -271 -247
rect -237 -281 -199 -247
rect -165 -281 -142 -247
rect -294 -287 -142 -281
rect -76 -247 76 -241
rect -76 -281 -53 -247
rect -19 -281 19 -247
rect 53 -281 76 -247
rect -76 -287 76 -281
rect 142 -247 294 -241
rect 142 -281 165 -247
rect 199 -281 237 -247
rect 271 -281 294 -247
rect 142 -287 294 -281
rect 360 -247 512 -241
rect 360 -281 383 -247
rect 417 -281 455 -247
rect 489 -281 512 -247
rect 360 -287 512 -281
rect 578 -247 730 -241
rect 578 -281 601 -247
rect 635 -281 673 -247
rect 707 -281 730 -247
rect 578 -287 730 -281
<< properties >>
string FIXED_BBOX -897 -402 897 402
<< end >>
