magic
tech sky130A
magscale 1 2
timestamp 1622081478
<< pwell >>
rect -298 -448 298 448
<< mvnmos >>
rect -80 -200 80 200
<< mvndiff >>
rect -138 187 -80 200
rect -138 153 -126 187
rect -92 153 -80 187
rect -138 119 -80 153
rect -138 85 -126 119
rect -92 85 -80 119
rect -138 51 -80 85
rect -138 17 -126 51
rect -92 17 -80 51
rect -138 -17 -80 17
rect -138 -51 -126 -17
rect -92 -51 -80 -17
rect -138 -85 -80 -51
rect -138 -119 -126 -85
rect -92 -119 -80 -85
rect -138 -153 -80 -119
rect -138 -187 -126 -153
rect -92 -187 -80 -153
rect -138 -200 -80 -187
rect 80 187 138 200
rect 80 153 92 187
rect 126 153 138 187
rect 80 119 138 153
rect 80 85 92 119
rect 126 85 138 119
rect 80 51 138 85
rect 80 17 92 51
rect 126 17 138 51
rect 80 -17 138 17
rect 80 -51 92 -17
rect 126 -51 138 -17
rect 80 -85 138 -51
rect 80 -119 92 -85
rect 126 -119 138 -85
rect 80 -153 138 -119
rect 80 -187 92 -153
rect 126 -187 138 -153
rect 80 -200 138 -187
<< mvndiffc >>
rect -126 153 -92 187
rect -126 85 -92 119
rect -126 17 -92 51
rect -126 -51 -92 -17
rect -126 -119 -92 -85
rect -126 -187 -92 -153
rect 92 153 126 187
rect 92 85 126 119
rect 92 17 126 51
rect 92 -51 126 -17
rect 92 -119 126 -85
rect 92 -187 126 -153
<< mvpsubdiff >>
rect -272 410 272 422
rect -272 376 -153 410
rect -119 376 -85 410
rect -51 376 -17 410
rect 17 376 51 410
rect 85 376 119 410
rect 153 376 272 410
rect -272 364 272 376
rect -272 -364 -214 364
rect 214 289 272 364
rect 214 255 226 289
rect 260 255 272 289
rect 214 221 272 255
rect 214 187 226 221
rect 260 187 272 221
rect 214 153 272 187
rect 214 119 226 153
rect 260 119 272 153
rect 214 85 272 119
rect 214 51 226 85
rect 260 51 272 85
rect 214 17 272 51
rect 214 -17 226 17
rect 260 -17 272 17
rect 214 -51 272 -17
rect 214 -85 226 -51
rect 260 -85 272 -51
rect 214 -119 272 -85
rect 214 -153 226 -119
rect 260 -153 272 -119
rect 214 -187 272 -153
rect 214 -221 226 -187
rect 260 -221 272 -187
rect 214 -255 272 -221
rect 214 -289 226 -255
rect 260 -289 272 -255
rect 214 -364 272 -289
rect -272 -376 272 -364
rect -272 -410 -153 -376
rect -119 -410 -85 -376
rect -51 -410 -17 -376
rect 17 -410 51 -376
rect 85 -410 119 -376
rect 153 -410 272 -376
rect -272 -422 272 -410
<< mvpsubdiffcont >>
rect -153 376 -119 410
rect -85 376 -51 410
rect -17 376 17 410
rect 51 376 85 410
rect 119 376 153 410
rect 226 255 260 289
rect 226 187 260 221
rect 226 119 260 153
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect 226 -153 260 -119
rect 226 -221 260 -187
rect 226 -289 260 -255
rect -153 -410 -119 -376
rect -85 -410 -51 -376
rect -17 -410 17 -376
rect 51 -410 85 -376
rect 119 -410 153 -376
<< poly >>
rect -80 272 80 288
rect -80 238 -51 272
rect -17 238 17 272
rect 51 238 80 272
rect -80 200 80 238
rect -80 -238 80 -200
rect -80 -272 -51 -238
rect -17 -272 17 -238
rect 51 -272 80 -238
rect -80 -288 80 -272
<< polycont >>
rect -51 238 -17 272
rect 17 238 51 272
rect -51 -272 -17 -238
rect 17 -272 51 -238
<< locali >>
rect -260 376 -153 410
rect -119 376 -85 410
rect -51 376 -17 410
rect 17 376 51 410
rect 85 376 119 410
rect 153 376 260 410
rect -260 -46 -226 376
rect 226 289 260 376
rect -80 238 -53 272
rect -17 238 17 272
rect 53 238 80 272
rect 226 221 260 255
rect -260 -118 -226 -80
rect -260 -190 -226 -152
rect -126 187 -92 204
rect -126 119 -92 127
rect -126 51 -92 55
rect -126 -55 -92 -51
rect -126 -127 -92 -119
rect -126 -204 -92 -187
rect 92 187 126 204
rect 92 119 126 127
rect 92 51 126 55
rect 92 -55 126 -51
rect 92 -127 126 -119
rect 92 -204 126 -187
rect 226 153 260 187
rect 226 85 260 119
rect 226 17 260 51
rect 226 -51 260 -17
rect 226 -119 260 -85
rect 226 -187 260 -153
rect -260 -262 -226 -224
rect -80 -272 -53 -238
rect -17 -272 17 -238
rect 53 -272 80 -238
rect 226 -255 260 -221
rect -260 -334 -226 -296
rect -260 -376 -226 -368
rect 226 -376 260 -289
rect -260 -410 -153 -376
rect -119 -410 -85 -376
rect -51 -410 -17 -376
rect 17 -410 51 -376
rect 85 -410 119 -376
rect 153 -410 260 -376
<< viali >>
rect -53 238 -51 272
rect -51 238 -19 272
rect 19 238 51 272
rect 51 238 53 272
rect -260 -80 -226 -46
rect -260 -152 -226 -118
rect -260 -224 -226 -190
rect -126 153 -92 161
rect -126 127 -92 153
rect -126 85 -92 89
rect -126 55 -92 85
rect -126 -17 -92 17
rect -126 -85 -92 -55
rect -126 -89 -92 -85
rect -126 -153 -92 -127
rect -126 -161 -92 -153
rect 92 153 126 161
rect 92 127 126 153
rect 92 85 126 89
rect 92 55 126 85
rect 92 -17 126 17
rect 92 -85 126 -55
rect 92 -89 126 -85
rect 92 -153 126 -127
rect 92 -161 126 -153
rect -260 -296 -226 -262
rect -53 -272 -51 -238
rect -51 -272 -19 -238
rect 19 -272 51 -238
rect 51 -272 53 -238
rect -260 -368 -226 -334
<< metal1 >>
rect -76 272 76 278
rect -76 238 -53 272
rect -19 238 19 272
rect 53 238 76 272
rect -76 232 76 238
rect -132 161 -86 200
rect -132 127 -126 161
rect -92 127 -86 161
rect -132 89 -86 127
rect -132 55 -126 89
rect -92 55 -86 89
rect -132 17 -86 55
rect -132 -17 -126 17
rect -92 -17 -86 17
rect -266 -46 -220 -26
rect -266 -80 -260 -46
rect -226 -80 -220 -46
rect -266 -118 -220 -80
rect -266 -152 -260 -118
rect -226 -152 -220 -118
rect -266 -190 -220 -152
rect -266 -224 -260 -190
rect -226 -224 -220 -190
rect -132 -55 -86 -17
rect -132 -89 -126 -55
rect -92 -89 -86 -55
rect -132 -127 -86 -89
rect -132 -161 -126 -127
rect -92 -161 -86 -127
rect -132 -200 -86 -161
rect 86 161 132 200
rect 86 127 92 161
rect 126 127 132 161
rect 86 89 132 127
rect 86 55 92 89
rect 126 55 132 89
rect 86 17 132 55
rect 86 -17 92 17
rect 126 -17 132 17
rect 86 -55 132 -17
rect 86 -89 92 -55
rect 126 -89 132 -55
rect 86 -127 132 -89
rect 86 -161 92 -127
rect 126 -161 132 -127
rect 86 -200 132 -161
rect -266 -262 -220 -224
rect -266 -296 -260 -262
rect -226 -296 -220 -262
rect -76 -238 76 -232
rect -76 -272 -53 -238
rect -19 -272 19 -238
rect 53 -272 76 -238
rect -76 -278 76 -272
rect -266 -334 -220 -296
rect -266 -368 -260 -334
rect -226 -368 -220 -334
rect -266 -388 -220 -368
<< properties >>
string FIXED_BBOX -242 -392 242 392
<< end >>
