magic
tech sky130A
magscale 1 2
timestamp 1620244706
<< error_p >>
rect -989 912 -919 1056
rect -671 912 -601 1056
rect -353 912 -283 1056
rect -35 912 35 1056
rect 283 912 353 1056
rect 601 912 671 1056
rect 919 912 989 1056
rect -989 -808 -919 -664
rect -671 -808 -601 -664
rect -353 -808 -283 -664
rect -35 -808 35 -664
rect 283 -808 353 -664
rect 601 -808 671 -664
rect 919 -808 989 -664
<< pwell >>
rect -1155 -2694 1155 2694
<< psubdiff >>
rect -1119 2624 -1023 2658
rect 1023 2624 1119 2658
rect -1119 2562 -1085 2624
rect 1085 2562 1119 2624
rect -1119 -2624 -1085 -2562
rect 1085 -2624 1119 -2562
rect -1119 -2658 -1023 -2624
rect 1023 -2658 1119 -2624
<< psubdiffcont >>
rect -1023 2624 1023 2658
rect -1119 -2562 -1085 2562
rect 1085 -2562 1119 2562
rect -1023 -2658 1023 -2624
<< xpolycontact >>
rect -989 2096 -919 2528
rect -989 912 -919 1344
rect -671 2096 -601 2528
rect -671 912 -601 1344
rect -353 2096 -283 2528
rect -353 912 -283 1344
rect -35 2096 35 2528
rect -35 912 35 1344
rect 283 2096 353 2528
rect 283 912 353 1344
rect 601 2096 671 2528
rect 601 912 671 1344
rect 919 2096 989 2528
rect 919 912 989 1344
rect -989 376 -919 808
rect -989 -808 -919 -376
rect -671 376 -601 808
rect -671 -808 -601 -376
rect -353 376 -283 808
rect -353 -808 -283 -376
rect -35 376 35 808
rect -35 -808 35 -376
rect 283 376 353 808
rect 283 -808 353 -376
rect 601 376 671 808
rect 601 -808 671 -376
rect 919 376 989 808
rect 919 -808 989 -376
rect -989 -1344 -919 -912
rect -989 -2528 -919 -2096
rect -671 -1344 -601 -912
rect -671 -2528 -601 -2096
rect -353 -1344 -283 -912
rect -353 -2528 -283 -2096
rect -35 -1344 35 -912
rect -35 -2528 35 -2096
rect 283 -1344 353 -912
rect 283 -2528 353 -2096
rect 601 -1344 671 -912
rect 601 -2528 671 -2096
rect 919 -1344 989 -912
rect 919 -2528 989 -2096
<< xpolyres >>
rect -989 1344 -919 2096
rect -671 1344 -601 2096
rect -353 1344 -283 2096
rect -35 1344 35 2096
rect 283 1344 353 2096
rect 601 1344 671 2096
rect 919 1344 989 2096
rect -989 -376 -919 376
rect -671 -376 -601 376
rect -353 -376 -283 376
rect -35 -376 35 376
rect 283 -376 353 376
rect 601 -376 671 376
rect 919 -376 989 376
rect -989 -2096 -919 -1344
rect -671 -2096 -601 -1344
rect -353 -2096 -283 -1344
rect -35 -2096 35 -1344
rect 283 -2096 353 -1344
rect 601 -2096 671 -1344
rect 919 -2096 989 -1344
<< locali >>
rect -1119 2624 -1023 2658
rect 1023 2624 1119 2658
rect -1119 2562 -1085 2624
rect 1085 2562 1119 2624
rect -1119 -2624 -1085 -2562
rect 1085 -2624 1119 -2562
rect -1119 -2658 -1023 -2624
rect 1023 -2658 1119 -2624
<< viali >>
rect -973 2113 -935 2510
rect -655 2113 -617 2510
rect -337 2113 -299 2510
rect -19 2113 19 2510
rect 299 2113 337 2510
rect 617 2113 655 2510
rect 935 2113 973 2510
rect -973 930 -935 1327
rect -655 930 -617 1327
rect -337 930 -299 1327
rect -19 930 19 1327
rect 299 930 337 1327
rect 617 930 655 1327
rect 935 930 973 1327
rect -973 393 -935 790
rect -655 393 -617 790
rect -337 393 -299 790
rect -19 393 19 790
rect 299 393 337 790
rect 617 393 655 790
rect 935 393 973 790
rect -973 -790 -935 -393
rect -655 -790 -617 -393
rect -337 -790 -299 -393
rect -19 -790 19 -393
rect 299 -790 337 -393
rect 617 -790 655 -393
rect 935 -790 973 -393
rect -973 -1327 -935 -930
rect -655 -1327 -617 -930
rect -337 -1327 -299 -930
rect -19 -1327 19 -930
rect 299 -1327 337 -930
rect 617 -1327 655 -930
rect 935 -1327 973 -930
rect -973 -2510 -935 -2113
rect -655 -2510 -617 -2113
rect -337 -2510 -299 -2113
rect -19 -2510 19 -2113
rect 299 -2510 337 -2113
rect 617 -2510 655 -2113
rect 935 -2510 973 -2113
<< metal1 >>
rect -979 2510 -929 2522
rect -979 2113 -973 2510
rect -935 2113 -929 2510
rect -979 2101 -929 2113
rect -661 2510 -611 2522
rect -661 2113 -655 2510
rect -617 2113 -611 2510
rect -661 2101 -611 2113
rect -343 2510 -293 2522
rect -343 2113 -337 2510
rect -299 2113 -293 2510
rect -343 2101 -293 2113
rect -25 2510 25 2522
rect -25 2113 -19 2510
rect 19 2113 25 2510
rect -25 2101 25 2113
rect 293 2510 343 2522
rect 293 2113 299 2510
rect 337 2113 343 2510
rect 293 2101 343 2113
rect 611 2510 661 2522
rect 611 2113 617 2510
rect 655 2113 661 2510
rect 611 2101 661 2113
rect 929 2510 979 2522
rect 929 2113 935 2510
rect 973 2113 979 2510
rect 929 2101 979 2113
rect -979 1327 -929 1339
rect -979 930 -973 1327
rect -935 930 -929 1327
rect -979 918 -929 930
rect -661 1327 -611 1339
rect -661 930 -655 1327
rect -617 930 -611 1327
rect -661 918 -611 930
rect -343 1327 -293 1339
rect -343 930 -337 1327
rect -299 930 -293 1327
rect -343 918 -293 930
rect -25 1327 25 1339
rect -25 930 -19 1327
rect 19 930 25 1327
rect -25 918 25 930
rect 293 1327 343 1339
rect 293 930 299 1327
rect 337 930 343 1327
rect 293 918 343 930
rect 611 1327 661 1339
rect 611 930 617 1327
rect 655 930 661 1327
rect 611 918 661 930
rect 929 1327 979 1339
rect 929 930 935 1327
rect 973 930 979 1327
rect 929 918 979 930
rect -979 790 -929 802
rect -979 393 -973 790
rect -935 393 -929 790
rect -979 381 -929 393
rect -661 790 -611 802
rect -661 393 -655 790
rect -617 393 -611 790
rect -661 381 -611 393
rect -343 790 -293 802
rect -343 393 -337 790
rect -299 393 -293 790
rect -343 381 -293 393
rect -25 790 25 802
rect -25 393 -19 790
rect 19 393 25 790
rect -25 381 25 393
rect 293 790 343 802
rect 293 393 299 790
rect 337 393 343 790
rect 293 381 343 393
rect 611 790 661 802
rect 611 393 617 790
rect 655 393 661 790
rect 611 381 661 393
rect 929 790 979 802
rect 929 393 935 790
rect 973 393 979 790
rect 929 381 979 393
rect -979 -393 -929 -381
rect -979 -790 -973 -393
rect -935 -790 -929 -393
rect -979 -802 -929 -790
rect -661 -393 -611 -381
rect -661 -790 -655 -393
rect -617 -790 -611 -393
rect -661 -802 -611 -790
rect -343 -393 -293 -381
rect -343 -790 -337 -393
rect -299 -790 -293 -393
rect -343 -802 -293 -790
rect -25 -393 25 -381
rect -25 -790 -19 -393
rect 19 -790 25 -393
rect -25 -802 25 -790
rect 293 -393 343 -381
rect 293 -790 299 -393
rect 337 -790 343 -393
rect 293 -802 343 -790
rect 611 -393 661 -381
rect 611 -790 617 -393
rect 655 -790 661 -393
rect 611 -802 661 -790
rect 929 -393 979 -381
rect 929 -790 935 -393
rect 973 -790 979 -393
rect 929 -802 979 -790
rect -979 -930 -929 -918
rect -979 -1327 -973 -930
rect -935 -1327 -929 -930
rect -979 -1339 -929 -1327
rect -661 -930 -611 -918
rect -661 -1327 -655 -930
rect -617 -1327 -611 -930
rect -661 -1339 -611 -1327
rect -343 -930 -293 -918
rect -343 -1327 -337 -930
rect -299 -1327 -293 -930
rect -343 -1339 -293 -1327
rect -25 -930 25 -918
rect -25 -1327 -19 -930
rect 19 -1327 25 -930
rect -25 -1339 25 -1327
rect 293 -930 343 -918
rect 293 -1327 299 -930
rect 337 -1327 343 -930
rect 293 -1339 343 -1327
rect 611 -930 661 -918
rect 611 -1327 617 -930
rect 655 -1327 661 -930
rect 611 -1339 661 -1327
rect 929 -930 979 -918
rect 929 -1327 935 -930
rect 973 -1327 979 -930
rect 929 -1339 979 -1327
rect -979 -2113 -929 -2101
rect -979 -2510 -973 -2113
rect -935 -2510 -929 -2113
rect -979 -2522 -929 -2510
rect -661 -2113 -611 -2101
rect -661 -2510 -655 -2113
rect -617 -2510 -611 -2113
rect -661 -2522 -611 -2510
rect -343 -2113 -293 -2101
rect -343 -2510 -337 -2113
rect -299 -2510 -293 -2113
rect -343 -2522 -293 -2510
rect -25 -2113 25 -2101
rect -25 -2510 -19 -2113
rect 19 -2510 25 -2113
rect -25 -2522 25 -2510
rect 293 -2113 343 -2101
rect 293 -2510 299 -2113
rect 337 -2510 343 -2113
rect 293 -2522 343 -2510
rect 611 -2113 661 -2101
rect 611 -2510 617 -2113
rect 655 -2510 661 -2113
rect 611 -2522 661 -2510
rect 929 -2113 979 -2101
rect 929 -2510 935 -2113
rect 973 -2510 979 -2113
rect 929 -2522 979 -2510
<< res0p35 >>
rect -991 1342 -917 2098
rect -673 1342 -599 2098
rect -355 1342 -281 2098
rect -37 1342 37 2098
rect 281 1342 355 2098
rect 599 1342 673 2098
rect 917 1342 991 2098
rect -991 -378 -917 378
rect -673 -378 -599 378
rect -355 -378 -281 378
rect -37 -378 37 378
rect 281 -378 355 378
rect 599 -378 673 378
rect 917 -378 991 378
rect -991 -2098 -917 -1342
rect -673 -2098 -599 -1342
rect -355 -2098 -281 -1342
rect -37 -2098 37 -1342
rect 281 -2098 355 -1342
rect 599 -2098 673 -1342
rect 917 -2098 991 -1342
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string FIXED_BBOX -1102 -2641 1102 2641
string parameters w 0.350 l 3.763 m 3 nx 7 wmin 0.350 lmin 0.50 rho 2000 val 22.188k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
