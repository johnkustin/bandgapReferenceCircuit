magic
tech sky130A
magscale 1 2
timestamp 1620324069
<< nwell >>
rect -9912 -2798 9912 2764
<< pmoslvt >>
rect -9818 -2736 -9418 2664
rect -9360 -2736 -8960 2664
rect -8902 -2736 -8502 2664
rect -8444 -2736 -8044 2664
rect -7986 -2736 -7586 2664
rect -7528 -2736 -7128 2664
rect -7070 -2736 -6670 2664
rect -6612 -2736 -6212 2664
rect -6154 -2736 -5754 2664
rect -5696 -2736 -5296 2664
rect -5238 -2736 -4838 2664
rect -4780 -2736 -4380 2664
rect -4322 -2736 -3922 2664
rect -3864 -2736 -3464 2664
rect -3406 -2736 -3006 2664
rect -2948 -2736 -2548 2664
rect -2490 -2736 -2090 2664
rect -2032 -2736 -1632 2664
rect -1574 -2736 -1174 2664
rect -1116 -2736 -716 2664
rect -658 -2736 -258 2664
rect -200 -2736 200 2664
rect 258 -2736 658 2664
rect 716 -2736 1116 2664
rect 1174 -2736 1574 2664
rect 1632 -2736 2032 2664
rect 2090 -2736 2490 2664
rect 2548 -2736 2948 2664
rect 3006 -2736 3406 2664
rect 3464 -2736 3864 2664
rect 3922 -2736 4322 2664
rect 4380 -2736 4780 2664
rect 4838 -2736 5238 2664
rect 5296 -2736 5696 2664
rect 5754 -2736 6154 2664
rect 6212 -2736 6612 2664
rect 6670 -2736 7070 2664
rect 7128 -2736 7528 2664
rect 7586 -2736 7986 2664
rect 8044 -2736 8444 2664
rect 8502 -2736 8902 2664
rect 8960 -2736 9360 2664
rect 9418 -2736 9818 2664
<< pdiff >>
rect -9876 2652 -9818 2664
rect -9876 -2724 -9864 2652
rect -9830 -2724 -9818 2652
rect -9876 -2736 -9818 -2724
rect -9418 2652 -9360 2664
rect -9418 -2724 -9406 2652
rect -9372 -2724 -9360 2652
rect -9418 -2736 -9360 -2724
rect -8960 2652 -8902 2664
rect -8960 -2724 -8948 2652
rect -8914 -2724 -8902 2652
rect -8960 -2736 -8902 -2724
rect -8502 2652 -8444 2664
rect -8502 -2724 -8490 2652
rect -8456 -2724 -8444 2652
rect -8502 -2736 -8444 -2724
rect -8044 2652 -7986 2664
rect -8044 -2724 -8032 2652
rect -7998 -2724 -7986 2652
rect -8044 -2736 -7986 -2724
rect -7586 2652 -7528 2664
rect -7586 -2724 -7574 2652
rect -7540 -2724 -7528 2652
rect -7586 -2736 -7528 -2724
rect -7128 2652 -7070 2664
rect -7128 -2724 -7116 2652
rect -7082 -2724 -7070 2652
rect -7128 -2736 -7070 -2724
rect -6670 2652 -6612 2664
rect -6670 -2724 -6658 2652
rect -6624 -2724 -6612 2652
rect -6670 -2736 -6612 -2724
rect -6212 2652 -6154 2664
rect -6212 -2724 -6200 2652
rect -6166 -2724 -6154 2652
rect -6212 -2736 -6154 -2724
rect -5754 2652 -5696 2664
rect -5754 -2724 -5742 2652
rect -5708 -2724 -5696 2652
rect -5754 -2736 -5696 -2724
rect -5296 2652 -5238 2664
rect -5296 -2724 -5284 2652
rect -5250 -2724 -5238 2652
rect -5296 -2736 -5238 -2724
rect -4838 2652 -4780 2664
rect -4838 -2724 -4826 2652
rect -4792 -2724 -4780 2652
rect -4838 -2736 -4780 -2724
rect -4380 2652 -4322 2664
rect -4380 -2724 -4368 2652
rect -4334 -2724 -4322 2652
rect -4380 -2736 -4322 -2724
rect -3922 2652 -3864 2664
rect -3922 -2724 -3910 2652
rect -3876 -2724 -3864 2652
rect -3922 -2736 -3864 -2724
rect -3464 2652 -3406 2664
rect -3464 -2724 -3452 2652
rect -3418 -2724 -3406 2652
rect -3464 -2736 -3406 -2724
rect -3006 2652 -2948 2664
rect -3006 -2724 -2994 2652
rect -2960 -2724 -2948 2652
rect -3006 -2736 -2948 -2724
rect -2548 2652 -2490 2664
rect -2548 -2724 -2536 2652
rect -2502 -2724 -2490 2652
rect -2548 -2736 -2490 -2724
rect -2090 2652 -2032 2664
rect -2090 -2724 -2078 2652
rect -2044 -2724 -2032 2652
rect -2090 -2736 -2032 -2724
rect -1632 2652 -1574 2664
rect -1632 -2724 -1620 2652
rect -1586 -2724 -1574 2652
rect -1632 -2736 -1574 -2724
rect -1174 2652 -1116 2664
rect -1174 -2724 -1162 2652
rect -1128 -2724 -1116 2652
rect -1174 -2736 -1116 -2724
rect -716 2652 -658 2664
rect -716 -2724 -704 2652
rect -670 -2724 -658 2652
rect -716 -2736 -658 -2724
rect -258 2652 -200 2664
rect -258 -2724 -246 2652
rect -212 -2724 -200 2652
rect -258 -2736 -200 -2724
rect 200 2652 258 2664
rect 200 -2724 212 2652
rect 246 -2724 258 2652
rect 200 -2736 258 -2724
rect 658 2652 716 2664
rect 658 -2724 670 2652
rect 704 -2724 716 2652
rect 658 -2736 716 -2724
rect 1116 2652 1174 2664
rect 1116 -2724 1128 2652
rect 1162 -2724 1174 2652
rect 1116 -2736 1174 -2724
rect 1574 2652 1632 2664
rect 1574 -2724 1586 2652
rect 1620 -2724 1632 2652
rect 1574 -2736 1632 -2724
rect 2032 2652 2090 2664
rect 2032 -2724 2044 2652
rect 2078 -2724 2090 2652
rect 2032 -2736 2090 -2724
rect 2490 2652 2548 2664
rect 2490 -2724 2502 2652
rect 2536 -2724 2548 2652
rect 2490 -2736 2548 -2724
rect 2948 2652 3006 2664
rect 2948 -2724 2960 2652
rect 2994 -2724 3006 2652
rect 2948 -2736 3006 -2724
rect 3406 2652 3464 2664
rect 3406 -2724 3418 2652
rect 3452 -2724 3464 2652
rect 3406 -2736 3464 -2724
rect 3864 2652 3922 2664
rect 3864 -2724 3876 2652
rect 3910 -2724 3922 2652
rect 3864 -2736 3922 -2724
rect 4322 2652 4380 2664
rect 4322 -2724 4334 2652
rect 4368 -2724 4380 2652
rect 4322 -2736 4380 -2724
rect 4780 2652 4838 2664
rect 4780 -2724 4792 2652
rect 4826 -2724 4838 2652
rect 4780 -2736 4838 -2724
rect 5238 2652 5296 2664
rect 5238 -2724 5250 2652
rect 5284 -2724 5296 2652
rect 5238 -2736 5296 -2724
rect 5696 2652 5754 2664
rect 5696 -2724 5708 2652
rect 5742 -2724 5754 2652
rect 5696 -2736 5754 -2724
rect 6154 2652 6212 2664
rect 6154 -2724 6166 2652
rect 6200 -2724 6212 2652
rect 6154 -2736 6212 -2724
rect 6612 2652 6670 2664
rect 6612 -2724 6624 2652
rect 6658 -2724 6670 2652
rect 6612 -2736 6670 -2724
rect 7070 2652 7128 2664
rect 7070 -2724 7082 2652
rect 7116 -2724 7128 2652
rect 7070 -2736 7128 -2724
rect 7528 2652 7586 2664
rect 7528 -2724 7540 2652
rect 7574 -2724 7586 2652
rect 7528 -2736 7586 -2724
rect 7986 2652 8044 2664
rect 7986 -2724 7998 2652
rect 8032 -2724 8044 2652
rect 7986 -2736 8044 -2724
rect 8444 2652 8502 2664
rect 8444 -2724 8456 2652
rect 8490 -2724 8502 2652
rect 8444 -2736 8502 -2724
rect 8902 2652 8960 2664
rect 8902 -2724 8914 2652
rect 8948 -2724 8960 2652
rect 8902 -2736 8960 -2724
rect 9360 2652 9418 2664
rect 9360 -2724 9372 2652
rect 9406 -2724 9418 2652
rect 9360 -2736 9418 -2724
rect 9818 2652 9876 2664
rect 9818 -2724 9830 2652
rect 9864 -2724 9876 2652
rect 9818 -2736 9876 -2724
<< pdiffc >>
rect -9864 -2724 -9830 2652
rect -9406 -2724 -9372 2652
rect -8948 -2724 -8914 2652
rect -8490 -2724 -8456 2652
rect -8032 -2724 -7998 2652
rect -7574 -2724 -7540 2652
rect -7116 -2724 -7082 2652
rect -6658 -2724 -6624 2652
rect -6200 -2724 -6166 2652
rect -5742 -2724 -5708 2652
rect -5284 -2724 -5250 2652
rect -4826 -2724 -4792 2652
rect -4368 -2724 -4334 2652
rect -3910 -2724 -3876 2652
rect -3452 -2724 -3418 2652
rect -2994 -2724 -2960 2652
rect -2536 -2724 -2502 2652
rect -2078 -2724 -2044 2652
rect -1620 -2724 -1586 2652
rect -1162 -2724 -1128 2652
rect -704 -2724 -670 2652
rect -246 -2724 -212 2652
rect 212 -2724 246 2652
rect 670 -2724 704 2652
rect 1128 -2724 1162 2652
rect 1586 -2724 1620 2652
rect 2044 -2724 2078 2652
rect 2502 -2724 2536 2652
rect 2960 -2724 2994 2652
rect 3418 -2724 3452 2652
rect 3876 -2724 3910 2652
rect 4334 -2724 4368 2652
rect 4792 -2724 4826 2652
rect 5250 -2724 5284 2652
rect 5708 -2724 5742 2652
rect 6166 -2724 6200 2652
rect 6624 -2724 6658 2652
rect 7082 -2724 7116 2652
rect 7540 -2724 7574 2652
rect 7998 -2724 8032 2652
rect 8456 -2724 8490 2652
rect 8914 -2724 8948 2652
rect 9372 -2724 9406 2652
rect 9830 -2724 9864 2652
<< poly >>
rect -9818 2745 -9418 2761
rect -9818 2711 -9802 2745
rect -9434 2711 -9418 2745
rect -9818 2664 -9418 2711
rect -9360 2745 -8960 2761
rect -9360 2711 -9344 2745
rect -8976 2711 -8960 2745
rect -9360 2664 -8960 2711
rect -8902 2745 -8502 2761
rect -8902 2711 -8886 2745
rect -8518 2711 -8502 2745
rect -8902 2664 -8502 2711
rect -8444 2745 -8044 2761
rect -8444 2711 -8428 2745
rect -8060 2711 -8044 2745
rect -8444 2664 -8044 2711
rect -7986 2745 -7586 2761
rect -7986 2711 -7970 2745
rect -7602 2711 -7586 2745
rect -7986 2664 -7586 2711
rect -7528 2745 -7128 2761
rect -7528 2711 -7512 2745
rect -7144 2711 -7128 2745
rect -7528 2664 -7128 2711
rect -7070 2745 -6670 2761
rect -7070 2711 -7054 2745
rect -6686 2711 -6670 2745
rect -7070 2664 -6670 2711
rect -6612 2745 -6212 2761
rect -6612 2711 -6596 2745
rect -6228 2711 -6212 2745
rect -6612 2664 -6212 2711
rect -6154 2745 -5754 2761
rect -6154 2711 -6138 2745
rect -5770 2711 -5754 2745
rect -6154 2664 -5754 2711
rect -5696 2745 -5296 2761
rect -5696 2711 -5680 2745
rect -5312 2711 -5296 2745
rect -5696 2664 -5296 2711
rect -5238 2745 -4838 2761
rect -5238 2711 -5222 2745
rect -4854 2711 -4838 2745
rect -5238 2664 -4838 2711
rect -4780 2745 -4380 2761
rect -4780 2711 -4764 2745
rect -4396 2711 -4380 2745
rect -4780 2664 -4380 2711
rect -4322 2745 -3922 2761
rect -4322 2711 -4306 2745
rect -3938 2711 -3922 2745
rect -4322 2664 -3922 2711
rect -3864 2745 -3464 2761
rect -3864 2711 -3848 2745
rect -3480 2711 -3464 2745
rect -3864 2664 -3464 2711
rect -3406 2745 -3006 2761
rect -3406 2711 -3390 2745
rect -3022 2711 -3006 2745
rect -3406 2664 -3006 2711
rect -2948 2745 -2548 2761
rect -2948 2711 -2932 2745
rect -2564 2711 -2548 2745
rect -2948 2664 -2548 2711
rect -2490 2745 -2090 2761
rect -2490 2711 -2474 2745
rect -2106 2711 -2090 2745
rect -2490 2664 -2090 2711
rect -2032 2745 -1632 2761
rect -2032 2711 -2016 2745
rect -1648 2711 -1632 2745
rect -2032 2664 -1632 2711
rect -1574 2745 -1174 2761
rect -1574 2711 -1558 2745
rect -1190 2711 -1174 2745
rect -1574 2664 -1174 2711
rect -1116 2745 -716 2761
rect -1116 2711 -1100 2745
rect -732 2711 -716 2745
rect -1116 2664 -716 2711
rect -658 2745 -258 2761
rect -658 2711 -642 2745
rect -274 2711 -258 2745
rect -658 2664 -258 2711
rect -200 2745 200 2761
rect -200 2711 -184 2745
rect 184 2711 200 2745
rect -200 2664 200 2711
rect 258 2745 658 2761
rect 258 2711 274 2745
rect 642 2711 658 2745
rect 258 2664 658 2711
rect 716 2745 1116 2761
rect 716 2711 732 2745
rect 1100 2711 1116 2745
rect 716 2664 1116 2711
rect 1174 2745 1574 2761
rect 1174 2711 1190 2745
rect 1558 2711 1574 2745
rect 1174 2664 1574 2711
rect 1632 2745 2032 2761
rect 1632 2711 1648 2745
rect 2016 2711 2032 2745
rect 1632 2664 2032 2711
rect 2090 2745 2490 2761
rect 2090 2711 2106 2745
rect 2474 2711 2490 2745
rect 2090 2664 2490 2711
rect 2548 2745 2948 2761
rect 2548 2711 2564 2745
rect 2932 2711 2948 2745
rect 2548 2664 2948 2711
rect 3006 2745 3406 2761
rect 3006 2711 3022 2745
rect 3390 2711 3406 2745
rect 3006 2664 3406 2711
rect 3464 2745 3864 2761
rect 3464 2711 3480 2745
rect 3848 2711 3864 2745
rect 3464 2664 3864 2711
rect 3922 2745 4322 2761
rect 3922 2711 3938 2745
rect 4306 2711 4322 2745
rect 3922 2664 4322 2711
rect 4380 2745 4780 2761
rect 4380 2711 4396 2745
rect 4764 2711 4780 2745
rect 4380 2664 4780 2711
rect 4838 2745 5238 2761
rect 4838 2711 4854 2745
rect 5222 2711 5238 2745
rect 4838 2664 5238 2711
rect 5296 2745 5696 2761
rect 5296 2711 5312 2745
rect 5680 2711 5696 2745
rect 5296 2664 5696 2711
rect 5754 2745 6154 2761
rect 5754 2711 5770 2745
rect 6138 2711 6154 2745
rect 5754 2664 6154 2711
rect 6212 2745 6612 2761
rect 6212 2711 6228 2745
rect 6596 2711 6612 2745
rect 6212 2664 6612 2711
rect 6670 2745 7070 2761
rect 6670 2711 6686 2745
rect 7054 2711 7070 2745
rect 6670 2664 7070 2711
rect 7128 2745 7528 2761
rect 7128 2711 7144 2745
rect 7512 2711 7528 2745
rect 7128 2664 7528 2711
rect 7586 2745 7986 2761
rect 7586 2711 7602 2745
rect 7970 2711 7986 2745
rect 7586 2664 7986 2711
rect 8044 2745 8444 2761
rect 8044 2711 8060 2745
rect 8428 2711 8444 2745
rect 8044 2664 8444 2711
rect 8502 2745 8902 2761
rect 8502 2711 8518 2745
rect 8886 2711 8902 2745
rect 8502 2664 8902 2711
rect 8960 2745 9360 2761
rect 8960 2711 8976 2745
rect 9344 2711 9360 2745
rect 8960 2664 9360 2711
rect 9418 2745 9818 2761
rect 9418 2711 9434 2745
rect 9802 2711 9818 2745
rect 9418 2664 9818 2711
rect -9818 -2762 -9418 -2736
rect -9360 -2762 -8960 -2736
rect -8902 -2762 -8502 -2736
rect -8444 -2762 -8044 -2736
rect -7986 -2762 -7586 -2736
rect -7528 -2762 -7128 -2736
rect -7070 -2762 -6670 -2736
rect -6612 -2762 -6212 -2736
rect -6154 -2762 -5754 -2736
rect -5696 -2762 -5296 -2736
rect -5238 -2762 -4838 -2736
rect -4780 -2762 -4380 -2736
rect -4322 -2762 -3922 -2736
rect -3864 -2762 -3464 -2736
rect -3406 -2762 -3006 -2736
rect -2948 -2762 -2548 -2736
rect -2490 -2762 -2090 -2736
rect -2032 -2762 -1632 -2736
rect -1574 -2762 -1174 -2736
rect -1116 -2762 -716 -2736
rect -658 -2762 -258 -2736
rect -200 -2762 200 -2736
rect 258 -2762 658 -2736
rect 716 -2762 1116 -2736
rect 1174 -2762 1574 -2736
rect 1632 -2762 2032 -2736
rect 2090 -2762 2490 -2736
rect 2548 -2762 2948 -2736
rect 3006 -2762 3406 -2736
rect 3464 -2762 3864 -2736
rect 3922 -2762 4322 -2736
rect 4380 -2762 4780 -2736
rect 4838 -2762 5238 -2736
rect 5296 -2762 5696 -2736
rect 5754 -2762 6154 -2736
rect 6212 -2762 6612 -2736
rect 6670 -2762 7070 -2736
rect 7128 -2762 7528 -2736
rect 7586 -2762 7986 -2736
rect 8044 -2762 8444 -2736
rect 8502 -2762 8902 -2736
rect 8960 -2762 9360 -2736
rect 9418 -2762 9818 -2736
<< polycont >>
rect -9802 2711 -9434 2745
rect -9344 2711 -8976 2745
rect -8886 2711 -8518 2745
rect -8428 2711 -8060 2745
rect -7970 2711 -7602 2745
rect -7512 2711 -7144 2745
rect -7054 2711 -6686 2745
rect -6596 2711 -6228 2745
rect -6138 2711 -5770 2745
rect -5680 2711 -5312 2745
rect -5222 2711 -4854 2745
rect -4764 2711 -4396 2745
rect -4306 2711 -3938 2745
rect -3848 2711 -3480 2745
rect -3390 2711 -3022 2745
rect -2932 2711 -2564 2745
rect -2474 2711 -2106 2745
rect -2016 2711 -1648 2745
rect -1558 2711 -1190 2745
rect -1100 2711 -732 2745
rect -642 2711 -274 2745
rect -184 2711 184 2745
rect 274 2711 642 2745
rect 732 2711 1100 2745
rect 1190 2711 1558 2745
rect 1648 2711 2016 2745
rect 2106 2711 2474 2745
rect 2564 2711 2932 2745
rect 3022 2711 3390 2745
rect 3480 2711 3848 2745
rect 3938 2711 4306 2745
rect 4396 2711 4764 2745
rect 4854 2711 5222 2745
rect 5312 2711 5680 2745
rect 5770 2711 6138 2745
rect 6228 2711 6596 2745
rect 6686 2711 7054 2745
rect 7144 2711 7512 2745
rect 7602 2711 7970 2745
rect 8060 2711 8428 2745
rect 8518 2711 8886 2745
rect 8976 2711 9344 2745
rect 9434 2711 9802 2745
<< locali >>
rect -9818 2711 -9802 2745
rect -9434 2711 -9418 2745
rect -9360 2711 -9344 2745
rect -8976 2711 -8960 2745
rect -8902 2711 -8886 2745
rect -8518 2711 -8502 2745
rect -8444 2711 -8428 2745
rect -8060 2711 -8044 2745
rect -7986 2711 -7970 2745
rect -7602 2711 -7586 2745
rect -7528 2711 -7512 2745
rect -7144 2711 -7128 2745
rect -7070 2711 -7054 2745
rect -6686 2711 -6670 2745
rect -6612 2711 -6596 2745
rect -6228 2711 -6212 2745
rect -6154 2711 -6138 2745
rect -5770 2711 -5754 2745
rect -5696 2711 -5680 2745
rect -5312 2711 -5296 2745
rect -5238 2711 -5222 2745
rect -4854 2711 -4838 2745
rect -4780 2711 -4764 2745
rect -4396 2711 -4380 2745
rect -4322 2711 -4306 2745
rect -3938 2711 -3922 2745
rect -3864 2711 -3848 2745
rect -3480 2711 -3464 2745
rect -3406 2711 -3390 2745
rect -3022 2711 -3006 2745
rect -2948 2711 -2932 2745
rect -2564 2711 -2548 2745
rect -2490 2711 -2474 2745
rect -2106 2711 -2090 2745
rect -2032 2711 -2016 2745
rect -1648 2711 -1632 2745
rect -1574 2711 -1558 2745
rect -1190 2711 -1174 2745
rect -1116 2711 -1100 2745
rect -732 2711 -716 2745
rect -658 2711 -642 2745
rect -274 2711 -258 2745
rect -200 2711 -184 2745
rect 184 2711 200 2745
rect 258 2711 274 2745
rect 642 2711 658 2745
rect 716 2711 732 2745
rect 1100 2711 1116 2745
rect 1174 2711 1190 2745
rect 1558 2711 1574 2745
rect 1632 2711 1648 2745
rect 2016 2711 2032 2745
rect 2090 2711 2106 2745
rect 2474 2711 2490 2745
rect 2548 2711 2564 2745
rect 2932 2711 2948 2745
rect 3006 2711 3022 2745
rect 3390 2711 3406 2745
rect 3464 2711 3480 2745
rect 3848 2711 3864 2745
rect 3922 2711 3938 2745
rect 4306 2711 4322 2745
rect 4380 2711 4396 2745
rect 4764 2711 4780 2745
rect 4838 2711 4854 2745
rect 5222 2711 5238 2745
rect 5296 2711 5312 2745
rect 5680 2711 5696 2745
rect 5754 2711 5770 2745
rect 6138 2711 6154 2745
rect 6212 2711 6228 2745
rect 6596 2711 6612 2745
rect 6670 2711 6686 2745
rect 7054 2711 7070 2745
rect 7128 2711 7144 2745
rect 7512 2711 7528 2745
rect 7586 2711 7602 2745
rect 7970 2711 7986 2745
rect 8044 2711 8060 2745
rect 8428 2711 8444 2745
rect 8502 2711 8518 2745
rect 8886 2711 8902 2745
rect 8960 2711 8976 2745
rect 9344 2711 9360 2745
rect 9418 2711 9434 2745
rect 9802 2711 9818 2745
rect -9864 2652 -9830 2668
rect -9864 -2740 -9830 -2724
rect -9406 2652 -9372 2668
rect -9406 -2740 -9372 -2724
rect -8948 2652 -8914 2668
rect -8948 -2740 -8914 -2724
rect -8490 2652 -8456 2668
rect -8490 -2740 -8456 -2724
rect -8032 2652 -7998 2668
rect -8032 -2740 -7998 -2724
rect -7574 2652 -7540 2668
rect -7574 -2740 -7540 -2724
rect -7116 2652 -7082 2668
rect -7116 -2740 -7082 -2724
rect -6658 2652 -6624 2668
rect -6658 -2740 -6624 -2724
rect -6200 2652 -6166 2668
rect -6200 -2740 -6166 -2724
rect -5742 2652 -5708 2668
rect -5742 -2740 -5708 -2724
rect -5284 2652 -5250 2668
rect -5284 -2740 -5250 -2724
rect -4826 2652 -4792 2668
rect -4826 -2740 -4792 -2724
rect -4368 2652 -4334 2668
rect -4368 -2740 -4334 -2724
rect -3910 2652 -3876 2668
rect -3910 -2740 -3876 -2724
rect -3452 2652 -3418 2668
rect -3452 -2740 -3418 -2724
rect -2994 2652 -2960 2668
rect -2994 -2740 -2960 -2724
rect -2536 2652 -2502 2668
rect -2536 -2740 -2502 -2724
rect -2078 2652 -2044 2668
rect -2078 -2740 -2044 -2724
rect -1620 2652 -1586 2668
rect -1620 -2740 -1586 -2724
rect -1162 2652 -1128 2668
rect -1162 -2740 -1128 -2724
rect -704 2652 -670 2668
rect -704 -2740 -670 -2724
rect -246 2652 -212 2668
rect -246 -2740 -212 -2724
rect 212 2652 246 2668
rect 212 -2740 246 -2724
rect 670 2652 704 2668
rect 670 -2740 704 -2724
rect 1128 2652 1162 2668
rect 1128 -2740 1162 -2724
rect 1586 2652 1620 2668
rect 1586 -2740 1620 -2724
rect 2044 2652 2078 2668
rect 2044 -2740 2078 -2724
rect 2502 2652 2536 2668
rect 2502 -2740 2536 -2724
rect 2960 2652 2994 2668
rect 2960 -2740 2994 -2724
rect 3418 2652 3452 2668
rect 3418 -2740 3452 -2724
rect 3876 2652 3910 2668
rect 3876 -2740 3910 -2724
rect 4334 2652 4368 2668
rect 4334 -2740 4368 -2724
rect 4792 2652 4826 2668
rect 4792 -2740 4826 -2724
rect 5250 2652 5284 2668
rect 5250 -2740 5284 -2724
rect 5708 2652 5742 2668
rect 5708 -2740 5742 -2724
rect 6166 2652 6200 2668
rect 6166 -2740 6200 -2724
rect 6624 2652 6658 2668
rect 6624 -2740 6658 -2724
rect 7082 2652 7116 2668
rect 7082 -2740 7116 -2724
rect 7540 2652 7574 2668
rect 7540 -2740 7574 -2724
rect 7998 2652 8032 2668
rect 7998 -2740 8032 -2724
rect 8456 2652 8490 2668
rect 8456 -2740 8490 -2724
rect 8914 2652 8948 2668
rect 8914 -2740 8948 -2724
rect 9372 2652 9406 2668
rect 9372 -2740 9406 -2724
rect 9830 2652 9864 2668
rect 9830 -2740 9864 -2724
<< viali >>
rect -9802 2711 -9434 2745
rect -9344 2711 -8976 2745
rect -8886 2711 -8518 2745
rect -8428 2711 -8060 2745
rect -7970 2711 -7602 2745
rect -7512 2711 -7144 2745
rect -7054 2711 -6686 2745
rect -6596 2711 -6228 2745
rect -6138 2711 -5770 2745
rect -5680 2711 -5312 2745
rect -5222 2711 -4854 2745
rect -4764 2711 -4396 2745
rect -4306 2711 -3938 2745
rect -3848 2711 -3480 2745
rect -3390 2711 -3022 2745
rect -2932 2711 -2564 2745
rect -2474 2711 -2106 2745
rect -2016 2711 -1648 2745
rect -1558 2711 -1190 2745
rect -1100 2711 -732 2745
rect -642 2711 -274 2745
rect -184 2711 184 2745
rect 274 2711 642 2745
rect 732 2711 1100 2745
rect 1190 2711 1558 2745
rect 1648 2711 2016 2745
rect 2106 2711 2474 2745
rect 2564 2711 2932 2745
rect 3022 2711 3390 2745
rect 3480 2711 3848 2745
rect 3938 2711 4306 2745
rect 4396 2711 4764 2745
rect 4854 2711 5222 2745
rect 5312 2711 5680 2745
rect 5770 2711 6138 2745
rect 6228 2711 6596 2745
rect 6686 2711 7054 2745
rect 7144 2711 7512 2745
rect 7602 2711 7970 2745
rect 8060 2711 8428 2745
rect 8518 2711 8886 2745
rect 8976 2711 9344 2745
rect 9434 2711 9802 2745
rect -9864 -2724 -9830 2652
rect -9406 -2724 -9372 2652
rect -8948 -2724 -8914 2652
rect -8490 -2724 -8456 2652
rect -8032 -2724 -7998 2652
rect -7574 -2724 -7540 2652
rect -7116 -2724 -7082 2652
rect -6658 -2724 -6624 2652
rect -6200 -2724 -6166 2652
rect -5742 -2724 -5708 2652
rect -5284 -2724 -5250 2652
rect -4826 -2724 -4792 2652
rect -4368 -2724 -4334 2652
rect -3910 -2724 -3876 2652
rect -3452 -2724 -3418 2652
rect -2994 -2724 -2960 2652
rect -2536 -2724 -2502 2652
rect -2078 -2724 -2044 2652
rect -1620 -2724 -1586 2652
rect -1162 -2724 -1128 2652
rect -704 -2724 -670 2652
rect -246 -2724 -212 2652
rect 212 -2724 246 2652
rect 670 -2724 704 2652
rect 1128 -2724 1162 2652
rect 1586 -2724 1620 2652
rect 2044 -2724 2078 2652
rect 2502 -2724 2536 2652
rect 2960 -2724 2994 2652
rect 3418 -2724 3452 2652
rect 3876 -2724 3910 2652
rect 4334 -2724 4368 2652
rect 4792 -2724 4826 2652
rect 5250 -2724 5284 2652
rect 5708 -2724 5742 2652
rect 6166 -2724 6200 2652
rect 6624 -2724 6658 2652
rect 7082 -2724 7116 2652
rect 7540 -2724 7574 2652
rect 7998 -2724 8032 2652
rect 8456 -2724 8490 2652
rect 8914 -2724 8948 2652
rect 9372 -2724 9406 2652
rect 9830 -2724 9864 2652
<< metal1 >>
rect -9814 2745 -9422 2751
rect -9814 2711 -9802 2745
rect -9434 2711 -9422 2745
rect -9814 2705 -9422 2711
rect -9356 2745 -8964 2751
rect -9356 2711 -9344 2745
rect -8976 2711 -8964 2745
rect -9356 2705 -8964 2711
rect -8898 2745 -8506 2751
rect -8898 2711 -8886 2745
rect -8518 2711 -8506 2745
rect -8898 2705 -8506 2711
rect -8440 2745 -8048 2751
rect -8440 2711 -8428 2745
rect -8060 2711 -8048 2745
rect -8440 2705 -8048 2711
rect -7982 2745 -7590 2751
rect -7982 2711 -7970 2745
rect -7602 2711 -7590 2745
rect -7982 2705 -7590 2711
rect -7524 2745 -7132 2751
rect -7524 2711 -7512 2745
rect -7144 2711 -7132 2745
rect -7524 2705 -7132 2711
rect -7066 2745 -6674 2751
rect -7066 2711 -7054 2745
rect -6686 2711 -6674 2745
rect -7066 2705 -6674 2711
rect -6608 2745 -6216 2751
rect -6608 2711 -6596 2745
rect -6228 2711 -6216 2745
rect -6608 2705 -6216 2711
rect -6150 2745 -5758 2751
rect -6150 2711 -6138 2745
rect -5770 2711 -5758 2745
rect -6150 2705 -5758 2711
rect -5692 2745 -5300 2751
rect -5692 2711 -5680 2745
rect -5312 2711 -5300 2745
rect -5692 2705 -5300 2711
rect -5234 2745 -4842 2751
rect -5234 2711 -5222 2745
rect -4854 2711 -4842 2745
rect -5234 2705 -4842 2711
rect -4776 2745 -4384 2751
rect -4776 2711 -4764 2745
rect -4396 2711 -4384 2745
rect -4776 2705 -4384 2711
rect -4318 2745 -3926 2751
rect -4318 2711 -4306 2745
rect -3938 2711 -3926 2745
rect -4318 2705 -3926 2711
rect -3860 2745 -3468 2751
rect -3860 2711 -3848 2745
rect -3480 2711 -3468 2745
rect -3860 2705 -3468 2711
rect -3402 2745 -3010 2751
rect -3402 2711 -3390 2745
rect -3022 2711 -3010 2745
rect -3402 2705 -3010 2711
rect -2944 2745 -2552 2751
rect -2944 2711 -2932 2745
rect -2564 2711 -2552 2745
rect -2944 2705 -2552 2711
rect -2486 2745 -2094 2751
rect -2486 2711 -2474 2745
rect -2106 2711 -2094 2745
rect -2486 2705 -2094 2711
rect -2028 2745 -1636 2751
rect -2028 2711 -2016 2745
rect -1648 2711 -1636 2745
rect -2028 2705 -1636 2711
rect -1570 2745 -1178 2751
rect -1570 2711 -1558 2745
rect -1190 2711 -1178 2745
rect -1570 2705 -1178 2711
rect -1112 2745 -720 2751
rect -1112 2711 -1100 2745
rect -732 2711 -720 2745
rect -1112 2705 -720 2711
rect -654 2745 -262 2751
rect -654 2711 -642 2745
rect -274 2711 -262 2745
rect -654 2705 -262 2711
rect -196 2745 196 2751
rect -196 2711 -184 2745
rect 184 2711 196 2745
rect -196 2705 196 2711
rect 262 2745 654 2751
rect 262 2711 274 2745
rect 642 2711 654 2745
rect 262 2705 654 2711
rect 720 2745 1112 2751
rect 720 2711 732 2745
rect 1100 2711 1112 2745
rect 720 2705 1112 2711
rect 1178 2745 1570 2751
rect 1178 2711 1190 2745
rect 1558 2711 1570 2745
rect 1178 2705 1570 2711
rect 1636 2745 2028 2751
rect 1636 2711 1648 2745
rect 2016 2711 2028 2745
rect 1636 2705 2028 2711
rect 2094 2745 2486 2751
rect 2094 2711 2106 2745
rect 2474 2711 2486 2745
rect 2094 2705 2486 2711
rect 2552 2745 2944 2751
rect 2552 2711 2564 2745
rect 2932 2711 2944 2745
rect 2552 2705 2944 2711
rect 3010 2745 3402 2751
rect 3010 2711 3022 2745
rect 3390 2711 3402 2745
rect 3010 2705 3402 2711
rect 3468 2745 3860 2751
rect 3468 2711 3480 2745
rect 3848 2711 3860 2745
rect 3468 2705 3860 2711
rect 3926 2745 4318 2751
rect 3926 2711 3938 2745
rect 4306 2711 4318 2745
rect 3926 2705 4318 2711
rect 4384 2745 4776 2751
rect 4384 2711 4396 2745
rect 4764 2711 4776 2745
rect 4384 2705 4776 2711
rect 4842 2745 5234 2751
rect 4842 2711 4854 2745
rect 5222 2711 5234 2745
rect 4842 2705 5234 2711
rect 5300 2745 5692 2751
rect 5300 2711 5312 2745
rect 5680 2711 5692 2745
rect 5300 2705 5692 2711
rect 5758 2745 6150 2751
rect 5758 2711 5770 2745
rect 6138 2711 6150 2745
rect 5758 2705 6150 2711
rect 6216 2745 6608 2751
rect 6216 2711 6228 2745
rect 6596 2711 6608 2745
rect 6216 2705 6608 2711
rect 6674 2745 7066 2751
rect 6674 2711 6686 2745
rect 7054 2711 7066 2745
rect 6674 2705 7066 2711
rect 7132 2745 7524 2751
rect 7132 2711 7144 2745
rect 7512 2711 7524 2745
rect 7132 2705 7524 2711
rect 7590 2745 7982 2751
rect 7590 2711 7602 2745
rect 7970 2711 7982 2745
rect 7590 2705 7982 2711
rect 8048 2745 8440 2751
rect 8048 2711 8060 2745
rect 8428 2711 8440 2745
rect 8048 2705 8440 2711
rect 8506 2745 8898 2751
rect 8506 2711 8518 2745
rect 8886 2711 8898 2745
rect 8506 2705 8898 2711
rect 8964 2745 9356 2751
rect 8964 2711 8976 2745
rect 9344 2711 9356 2745
rect 8964 2705 9356 2711
rect 9422 2745 9814 2751
rect 9422 2711 9434 2745
rect 9802 2711 9814 2745
rect 9422 2705 9814 2711
rect -9870 2652 -9824 2664
rect -9870 -2724 -9864 2652
rect -9830 -2724 -9824 2652
rect -9870 -2736 -9824 -2724
rect -9412 2652 -9366 2664
rect -9412 -2724 -9406 2652
rect -9372 -2724 -9366 2652
rect -9412 -2736 -9366 -2724
rect -8954 2652 -8908 2664
rect -8954 -2724 -8948 2652
rect -8914 -2724 -8908 2652
rect -8954 -2736 -8908 -2724
rect -8496 2652 -8450 2664
rect -8496 -2724 -8490 2652
rect -8456 -2724 -8450 2652
rect -8496 -2736 -8450 -2724
rect -8038 2652 -7992 2664
rect -8038 -2724 -8032 2652
rect -7998 -2724 -7992 2652
rect -8038 -2736 -7992 -2724
rect -7580 2652 -7534 2664
rect -7580 -2724 -7574 2652
rect -7540 -2724 -7534 2652
rect -7580 -2736 -7534 -2724
rect -7122 2652 -7076 2664
rect -7122 -2724 -7116 2652
rect -7082 -2724 -7076 2652
rect -7122 -2736 -7076 -2724
rect -6664 2652 -6618 2664
rect -6664 -2724 -6658 2652
rect -6624 -2724 -6618 2652
rect -6664 -2736 -6618 -2724
rect -6206 2652 -6160 2664
rect -6206 -2724 -6200 2652
rect -6166 -2724 -6160 2652
rect -6206 -2736 -6160 -2724
rect -5748 2652 -5702 2664
rect -5748 -2724 -5742 2652
rect -5708 -2724 -5702 2652
rect -5748 -2736 -5702 -2724
rect -5290 2652 -5244 2664
rect -5290 -2724 -5284 2652
rect -5250 -2724 -5244 2652
rect -5290 -2736 -5244 -2724
rect -4832 2652 -4786 2664
rect -4832 -2724 -4826 2652
rect -4792 -2724 -4786 2652
rect -4832 -2736 -4786 -2724
rect -4374 2652 -4328 2664
rect -4374 -2724 -4368 2652
rect -4334 -2724 -4328 2652
rect -4374 -2736 -4328 -2724
rect -3916 2652 -3870 2664
rect -3916 -2724 -3910 2652
rect -3876 -2724 -3870 2652
rect -3916 -2736 -3870 -2724
rect -3458 2652 -3412 2664
rect -3458 -2724 -3452 2652
rect -3418 -2724 -3412 2652
rect -3458 -2736 -3412 -2724
rect -3000 2652 -2954 2664
rect -3000 -2724 -2994 2652
rect -2960 -2724 -2954 2652
rect -3000 -2736 -2954 -2724
rect -2542 2652 -2496 2664
rect -2542 -2724 -2536 2652
rect -2502 -2724 -2496 2652
rect -2542 -2736 -2496 -2724
rect -2084 2652 -2038 2664
rect -2084 -2724 -2078 2652
rect -2044 -2724 -2038 2652
rect -2084 -2736 -2038 -2724
rect -1626 2652 -1580 2664
rect -1626 -2724 -1620 2652
rect -1586 -2724 -1580 2652
rect -1626 -2736 -1580 -2724
rect -1168 2652 -1122 2664
rect -1168 -2724 -1162 2652
rect -1128 -2724 -1122 2652
rect -1168 -2736 -1122 -2724
rect -710 2652 -664 2664
rect -710 -2724 -704 2652
rect -670 -2724 -664 2652
rect -710 -2736 -664 -2724
rect -252 2652 -206 2664
rect -252 -2724 -246 2652
rect -212 -2724 -206 2652
rect -252 -2736 -206 -2724
rect 206 2652 252 2664
rect 206 -2724 212 2652
rect 246 -2724 252 2652
rect 206 -2736 252 -2724
rect 664 2652 710 2664
rect 664 -2724 670 2652
rect 704 -2724 710 2652
rect 664 -2736 710 -2724
rect 1122 2652 1168 2664
rect 1122 -2724 1128 2652
rect 1162 -2724 1168 2652
rect 1122 -2736 1168 -2724
rect 1580 2652 1626 2664
rect 1580 -2724 1586 2652
rect 1620 -2724 1626 2652
rect 1580 -2736 1626 -2724
rect 2038 2652 2084 2664
rect 2038 -2724 2044 2652
rect 2078 -2724 2084 2652
rect 2038 -2736 2084 -2724
rect 2496 2652 2542 2664
rect 2496 -2724 2502 2652
rect 2536 -2724 2542 2652
rect 2496 -2736 2542 -2724
rect 2954 2652 3000 2664
rect 2954 -2724 2960 2652
rect 2994 -2724 3000 2652
rect 2954 -2736 3000 -2724
rect 3412 2652 3458 2664
rect 3412 -2724 3418 2652
rect 3452 -2724 3458 2652
rect 3412 -2736 3458 -2724
rect 3870 2652 3916 2664
rect 3870 -2724 3876 2652
rect 3910 -2724 3916 2652
rect 3870 -2736 3916 -2724
rect 4328 2652 4374 2664
rect 4328 -2724 4334 2652
rect 4368 -2724 4374 2652
rect 4328 -2736 4374 -2724
rect 4786 2652 4832 2664
rect 4786 -2724 4792 2652
rect 4826 -2724 4832 2652
rect 4786 -2736 4832 -2724
rect 5244 2652 5290 2664
rect 5244 -2724 5250 2652
rect 5284 -2724 5290 2652
rect 5244 -2736 5290 -2724
rect 5702 2652 5748 2664
rect 5702 -2724 5708 2652
rect 5742 -2724 5748 2652
rect 5702 -2736 5748 -2724
rect 6160 2652 6206 2664
rect 6160 -2724 6166 2652
rect 6200 -2724 6206 2652
rect 6160 -2736 6206 -2724
rect 6618 2652 6664 2664
rect 6618 -2724 6624 2652
rect 6658 -2724 6664 2652
rect 6618 -2736 6664 -2724
rect 7076 2652 7122 2664
rect 7076 -2724 7082 2652
rect 7116 -2724 7122 2652
rect 7076 -2736 7122 -2724
rect 7534 2652 7580 2664
rect 7534 -2724 7540 2652
rect 7574 -2724 7580 2652
rect 7534 -2736 7580 -2724
rect 7992 2652 8038 2664
rect 7992 -2724 7998 2652
rect 8032 -2724 8038 2652
rect 7992 -2736 8038 -2724
rect 8450 2652 8496 2664
rect 8450 -2724 8456 2652
rect 8490 -2724 8496 2652
rect 8450 -2736 8496 -2724
rect 8908 2652 8954 2664
rect 8908 -2724 8914 2652
rect 8948 -2724 8954 2652
rect 8908 -2736 8954 -2724
rect 9366 2652 9412 2664
rect 9366 -2724 9372 2652
rect 9406 -2724 9412 2652
rect 9366 -2736 9412 -2724
rect 9824 2652 9870 2664
rect 9824 -2724 9830 2652
rect 9864 -2724 9870 2652
rect 9824 -2736 9870 -2724
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 27 l 2 m 1 nf 43 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
