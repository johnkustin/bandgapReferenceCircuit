magic
tech sky130A
magscale 1 2
timestamp 1622081478
<< metal3 >>
rect -3136 3072 3136 3100
rect -3136 3008 3052 3072
rect 3116 3008 3136 3072
rect -3136 2992 3136 3008
rect -3136 2928 3052 2992
rect 3116 2928 3136 2992
rect -3136 2912 3136 2928
rect -3136 2848 3052 2912
rect 3116 2848 3136 2912
rect -3136 2832 3136 2848
rect -3136 2768 3052 2832
rect 3116 2768 3136 2832
rect -3136 2752 3136 2768
rect -3136 2688 3052 2752
rect 3116 2688 3136 2752
rect -3136 2672 3136 2688
rect -3136 2608 3052 2672
rect 3116 2608 3136 2672
rect -3136 2592 3136 2608
rect -3136 2528 3052 2592
rect 3116 2528 3136 2592
rect -3136 2512 3136 2528
rect -3136 2448 3052 2512
rect 3116 2448 3136 2512
rect -3136 2432 3136 2448
rect -3136 2368 3052 2432
rect 3116 2368 3136 2432
rect -3136 2352 3136 2368
rect -3136 2288 3052 2352
rect 3116 2288 3136 2352
rect -3136 2272 3136 2288
rect -3136 2208 3052 2272
rect 3116 2208 3136 2272
rect -3136 2192 3136 2208
rect -3136 2128 3052 2192
rect 3116 2128 3136 2192
rect -3136 2112 3136 2128
rect -3136 2048 3052 2112
rect 3116 2048 3136 2112
rect -3136 2032 3136 2048
rect -3136 1968 3052 2032
rect 3116 1968 3136 2032
rect -3136 1952 3136 1968
rect -3136 1888 3052 1952
rect 3116 1888 3136 1952
rect -3136 1872 3136 1888
rect -3136 1808 3052 1872
rect 3116 1808 3136 1872
rect -3136 1792 3136 1808
rect -3136 1728 3052 1792
rect 3116 1728 3136 1792
rect -3136 1712 3136 1728
rect -3136 1648 3052 1712
rect 3116 1648 3136 1712
rect -3136 1632 3136 1648
rect -3136 1568 3052 1632
rect 3116 1568 3136 1632
rect -3136 1552 3136 1568
rect -3136 1488 3052 1552
rect 3116 1488 3136 1552
rect -3136 1472 3136 1488
rect -3136 1408 3052 1472
rect 3116 1408 3136 1472
rect -3136 1392 3136 1408
rect -3136 1328 3052 1392
rect 3116 1328 3136 1392
rect -3136 1312 3136 1328
rect -3136 1248 3052 1312
rect 3116 1248 3136 1312
rect -3136 1232 3136 1248
rect -3136 1168 3052 1232
rect 3116 1168 3136 1232
rect -3136 1152 3136 1168
rect -3136 1088 3052 1152
rect 3116 1088 3136 1152
rect -3136 1072 3136 1088
rect -3136 1008 3052 1072
rect 3116 1008 3136 1072
rect -3136 992 3136 1008
rect -3136 928 3052 992
rect 3116 928 3136 992
rect -3136 912 3136 928
rect -3136 848 3052 912
rect 3116 848 3136 912
rect -3136 832 3136 848
rect -3136 768 3052 832
rect 3116 768 3136 832
rect -3136 752 3136 768
rect -3136 688 3052 752
rect 3116 688 3136 752
rect -3136 672 3136 688
rect -3136 608 3052 672
rect 3116 608 3136 672
rect -3136 592 3136 608
rect -3136 528 3052 592
rect 3116 528 3136 592
rect -3136 512 3136 528
rect -3136 448 3052 512
rect 3116 448 3136 512
rect -3136 432 3136 448
rect -3136 368 3052 432
rect 3116 368 3136 432
rect -3136 352 3136 368
rect -3136 288 3052 352
rect 3116 288 3136 352
rect -3136 272 3136 288
rect -3136 208 3052 272
rect 3116 208 3136 272
rect -3136 192 3136 208
rect -3136 128 3052 192
rect 3116 128 3136 192
rect -3136 112 3136 128
rect -3136 48 3052 112
rect 3116 48 3136 112
rect -3136 32 3136 48
rect -3136 -32 3052 32
rect 3116 -32 3136 32
rect -3136 -48 3136 -32
rect -3136 -112 3052 -48
rect 3116 -112 3136 -48
rect -3136 -128 3136 -112
rect -3136 -192 3052 -128
rect 3116 -192 3136 -128
rect -3136 -208 3136 -192
rect -3136 -272 3052 -208
rect 3116 -272 3136 -208
rect -3136 -288 3136 -272
rect -3136 -352 3052 -288
rect 3116 -352 3136 -288
rect -3136 -368 3136 -352
rect -3136 -432 3052 -368
rect 3116 -432 3136 -368
rect -3136 -448 3136 -432
rect -3136 -512 3052 -448
rect 3116 -512 3136 -448
rect -3136 -528 3136 -512
rect -3136 -592 3052 -528
rect 3116 -592 3136 -528
rect -3136 -608 3136 -592
rect -3136 -672 3052 -608
rect 3116 -672 3136 -608
rect -3136 -688 3136 -672
rect -3136 -752 3052 -688
rect 3116 -752 3136 -688
rect -3136 -768 3136 -752
rect -3136 -832 3052 -768
rect 3116 -832 3136 -768
rect -3136 -848 3136 -832
rect -3136 -912 3052 -848
rect 3116 -912 3136 -848
rect -3136 -928 3136 -912
rect -3136 -992 3052 -928
rect 3116 -992 3136 -928
rect -3136 -1008 3136 -992
rect -3136 -1072 3052 -1008
rect 3116 -1072 3136 -1008
rect -3136 -1088 3136 -1072
rect -3136 -1152 3052 -1088
rect 3116 -1152 3136 -1088
rect -3136 -1168 3136 -1152
rect -3136 -1232 3052 -1168
rect 3116 -1232 3136 -1168
rect -3136 -1248 3136 -1232
rect -3136 -1312 3052 -1248
rect 3116 -1312 3136 -1248
rect -3136 -1328 3136 -1312
rect -3136 -1392 3052 -1328
rect 3116 -1392 3136 -1328
rect -3136 -1408 3136 -1392
rect -3136 -1472 3052 -1408
rect 3116 -1472 3136 -1408
rect -3136 -1488 3136 -1472
rect -3136 -1552 3052 -1488
rect 3116 -1552 3136 -1488
rect -3136 -1568 3136 -1552
rect -3136 -1632 3052 -1568
rect 3116 -1632 3136 -1568
rect -3136 -1648 3136 -1632
rect -3136 -1712 3052 -1648
rect 3116 -1712 3136 -1648
rect -3136 -1728 3136 -1712
rect -3136 -1792 3052 -1728
rect 3116 -1792 3136 -1728
rect -3136 -1808 3136 -1792
rect -3136 -1872 3052 -1808
rect 3116 -1872 3136 -1808
rect -3136 -1888 3136 -1872
rect -3136 -1952 3052 -1888
rect 3116 -1952 3136 -1888
rect -3136 -1968 3136 -1952
rect -3136 -2032 3052 -1968
rect 3116 -2032 3136 -1968
rect -3136 -2048 3136 -2032
rect -3136 -2112 3052 -2048
rect 3116 -2112 3136 -2048
rect -3136 -2128 3136 -2112
rect -3136 -2192 3052 -2128
rect 3116 -2192 3136 -2128
rect -3136 -2208 3136 -2192
rect -3136 -2272 3052 -2208
rect 3116 -2272 3136 -2208
rect -3136 -2288 3136 -2272
rect -3136 -2352 3052 -2288
rect 3116 -2352 3136 -2288
rect -3136 -2368 3136 -2352
rect -3136 -2432 3052 -2368
rect 3116 -2432 3136 -2368
rect -3136 -2448 3136 -2432
rect -3136 -2512 3052 -2448
rect 3116 -2512 3136 -2448
rect -3136 -2528 3136 -2512
rect -3136 -2592 3052 -2528
rect 3116 -2592 3136 -2528
rect -3136 -2608 3136 -2592
rect -3136 -2672 3052 -2608
rect 3116 -2672 3136 -2608
rect -3136 -2688 3136 -2672
rect -3136 -2752 3052 -2688
rect 3116 -2752 3136 -2688
rect -3136 -2768 3136 -2752
rect -3136 -2832 3052 -2768
rect 3116 -2832 3136 -2768
rect -3136 -2848 3136 -2832
rect -3136 -2912 3052 -2848
rect 3116 -2912 3136 -2848
rect -3136 -2928 3136 -2912
rect -3136 -2992 3052 -2928
rect 3116 -2992 3136 -2928
rect -3136 -3008 3136 -2992
rect -3136 -3072 3052 -3008
rect 3116 -3072 3136 -3008
rect -3136 -3100 3136 -3072
<< via3 >>
rect 3052 3008 3116 3072
rect 3052 2928 3116 2992
rect 3052 2848 3116 2912
rect 3052 2768 3116 2832
rect 3052 2688 3116 2752
rect 3052 2608 3116 2672
rect 3052 2528 3116 2592
rect 3052 2448 3116 2512
rect 3052 2368 3116 2432
rect 3052 2288 3116 2352
rect 3052 2208 3116 2272
rect 3052 2128 3116 2192
rect 3052 2048 3116 2112
rect 3052 1968 3116 2032
rect 3052 1888 3116 1952
rect 3052 1808 3116 1872
rect 3052 1728 3116 1792
rect 3052 1648 3116 1712
rect 3052 1568 3116 1632
rect 3052 1488 3116 1552
rect 3052 1408 3116 1472
rect 3052 1328 3116 1392
rect 3052 1248 3116 1312
rect 3052 1168 3116 1232
rect 3052 1088 3116 1152
rect 3052 1008 3116 1072
rect 3052 928 3116 992
rect 3052 848 3116 912
rect 3052 768 3116 832
rect 3052 688 3116 752
rect 3052 608 3116 672
rect 3052 528 3116 592
rect 3052 448 3116 512
rect 3052 368 3116 432
rect 3052 288 3116 352
rect 3052 208 3116 272
rect 3052 128 3116 192
rect 3052 48 3116 112
rect 3052 -32 3116 32
rect 3052 -112 3116 -48
rect 3052 -192 3116 -128
rect 3052 -272 3116 -208
rect 3052 -352 3116 -288
rect 3052 -432 3116 -368
rect 3052 -512 3116 -448
rect 3052 -592 3116 -528
rect 3052 -672 3116 -608
rect 3052 -752 3116 -688
rect 3052 -832 3116 -768
rect 3052 -912 3116 -848
rect 3052 -992 3116 -928
rect 3052 -1072 3116 -1008
rect 3052 -1152 3116 -1088
rect 3052 -1232 3116 -1168
rect 3052 -1312 3116 -1248
rect 3052 -1392 3116 -1328
rect 3052 -1472 3116 -1408
rect 3052 -1552 3116 -1488
rect 3052 -1632 3116 -1568
rect 3052 -1712 3116 -1648
rect 3052 -1792 3116 -1728
rect 3052 -1872 3116 -1808
rect 3052 -1952 3116 -1888
rect 3052 -2032 3116 -1968
rect 3052 -2112 3116 -2048
rect 3052 -2192 3116 -2128
rect 3052 -2272 3116 -2208
rect 3052 -2352 3116 -2288
rect 3052 -2432 3116 -2368
rect 3052 -2512 3116 -2448
rect 3052 -2592 3116 -2528
rect 3052 -2672 3116 -2608
rect 3052 -2752 3116 -2688
rect 3052 -2832 3116 -2768
rect 3052 -2912 3116 -2848
rect 3052 -2992 3116 -2928
rect 3052 -3072 3116 -3008
<< mimcap >>
rect -3036 2952 2964 3000
rect -3036 -2952 2356 2952
rect 2900 -2952 2964 2952
rect -3036 -3000 2964 -2952
<< mimcapcontact >>
rect 2356 -2952 2900 2952
<< metal4 >>
rect 3036 3072 3132 3088
rect 3036 3008 3052 3072
rect 3116 3008 3132 3072
rect 3036 2992 3132 3008
rect 2331 2952 2925 2961
rect 2331 -2952 2356 2952
rect 2900 -2952 2925 2952
rect 2331 -2961 2925 -2952
rect 3036 2928 3052 2992
rect 3116 2928 3132 2992
rect 3036 2912 3132 2928
rect 3036 2848 3052 2912
rect 3116 2848 3132 2912
rect 3036 2832 3132 2848
rect 3036 2768 3052 2832
rect 3116 2768 3132 2832
rect 3036 2752 3132 2768
rect 3036 2688 3052 2752
rect 3116 2688 3132 2752
rect 3036 2672 3132 2688
rect 3036 2608 3052 2672
rect 3116 2608 3132 2672
rect 3036 2592 3132 2608
rect 3036 2528 3052 2592
rect 3116 2528 3132 2592
rect 3036 2512 3132 2528
rect 3036 2448 3052 2512
rect 3116 2448 3132 2512
rect 3036 2432 3132 2448
rect 3036 2368 3052 2432
rect 3116 2368 3132 2432
rect 3036 2352 3132 2368
rect 3036 2288 3052 2352
rect 3116 2288 3132 2352
rect 3036 2272 3132 2288
rect 3036 2208 3052 2272
rect 3116 2208 3132 2272
rect 3036 2192 3132 2208
rect 3036 2128 3052 2192
rect 3116 2128 3132 2192
rect 3036 2112 3132 2128
rect 3036 2048 3052 2112
rect 3116 2048 3132 2112
rect 3036 2032 3132 2048
rect 3036 1968 3052 2032
rect 3116 1968 3132 2032
rect 3036 1952 3132 1968
rect 3036 1888 3052 1952
rect 3116 1888 3132 1952
rect 3036 1872 3132 1888
rect 3036 1808 3052 1872
rect 3116 1808 3132 1872
rect 3036 1792 3132 1808
rect 3036 1728 3052 1792
rect 3116 1728 3132 1792
rect 3036 1712 3132 1728
rect 3036 1648 3052 1712
rect 3116 1648 3132 1712
rect 3036 1632 3132 1648
rect 3036 1568 3052 1632
rect 3116 1568 3132 1632
rect 3036 1552 3132 1568
rect 3036 1488 3052 1552
rect 3116 1488 3132 1552
rect 3036 1472 3132 1488
rect 3036 1408 3052 1472
rect 3116 1408 3132 1472
rect 3036 1392 3132 1408
rect 3036 1328 3052 1392
rect 3116 1328 3132 1392
rect 3036 1312 3132 1328
rect 3036 1248 3052 1312
rect 3116 1248 3132 1312
rect 3036 1232 3132 1248
rect 3036 1168 3052 1232
rect 3116 1168 3132 1232
rect 3036 1152 3132 1168
rect 3036 1088 3052 1152
rect 3116 1088 3132 1152
rect 3036 1072 3132 1088
rect 3036 1008 3052 1072
rect 3116 1008 3132 1072
rect 3036 992 3132 1008
rect 3036 928 3052 992
rect 3116 928 3132 992
rect 3036 912 3132 928
rect 3036 848 3052 912
rect 3116 848 3132 912
rect 3036 832 3132 848
rect 3036 768 3052 832
rect 3116 768 3132 832
rect 3036 752 3132 768
rect 3036 688 3052 752
rect 3116 688 3132 752
rect 3036 672 3132 688
rect 3036 608 3052 672
rect 3116 608 3132 672
rect 3036 592 3132 608
rect 3036 528 3052 592
rect 3116 528 3132 592
rect 3036 512 3132 528
rect 3036 448 3052 512
rect 3116 448 3132 512
rect 3036 432 3132 448
rect 3036 368 3052 432
rect 3116 368 3132 432
rect 3036 352 3132 368
rect 3036 288 3052 352
rect 3116 288 3132 352
rect 3036 272 3132 288
rect 3036 208 3052 272
rect 3116 208 3132 272
rect 3036 192 3132 208
rect 3036 128 3052 192
rect 3116 128 3132 192
rect 3036 112 3132 128
rect 3036 48 3052 112
rect 3116 48 3132 112
rect 3036 32 3132 48
rect 3036 -32 3052 32
rect 3116 -32 3132 32
rect 3036 -48 3132 -32
rect 3036 -112 3052 -48
rect 3116 -112 3132 -48
rect 3036 -128 3132 -112
rect 3036 -192 3052 -128
rect 3116 -192 3132 -128
rect 3036 -208 3132 -192
rect 3036 -272 3052 -208
rect 3116 -272 3132 -208
rect 3036 -288 3132 -272
rect 3036 -352 3052 -288
rect 3116 -352 3132 -288
rect 3036 -368 3132 -352
rect 3036 -432 3052 -368
rect 3116 -432 3132 -368
rect 3036 -448 3132 -432
rect 3036 -512 3052 -448
rect 3116 -512 3132 -448
rect 3036 -528 3132 -512
rect 3036 -592 3052 -528
rect 3116 -592 3132 -528
rect 3036 -608 3132 -592
rect 3036 -672 3052 -608
rect 3116 -672 3132 -608
rect 3036 -688 3132 -672
rect 3036 -752 3052 -688
rect 3116 -752 3132 -688
rect 3036 -768 3132 -752
rect 3036 -832 3052 -768
rect 3116 -832 3132 -768
rect 3036 -848 3132 -832
rect 3036 -912 3052 -848
rect 3116 -912 3132 -848
rect 3036 -928 3132 -912
rect 3036 -992 3052 -928
rect 3116 -992 3132 -928
rect 3036 -1008 3132 -992
rect 3036 -1072 3052 -1008
rect 3116 -1072 3132 -1008
rect 3036 -1088 3132 -1072
rect 3036 -1152 3052 -1088
rect 3116 -1152 3132 -1088
rect 3036 -1168 3132 -1152
rect 3036 -1232 3052 -1168
rect 3116 -1232 3132 -1168
rect 3036 -1248 3132 -1232
rect 3036 -1312 3052 -1248
rect 3116 -1312 3132 -1248
rect 3036 -1328 3132 -1312
rect 3036 -1392 3052 -1328
rect 3116 -1392 3132 -1328
rect 3036 -1408 3132 -1392
rect 3036 -1472 3052 -1408
rect 3116 -1472 3132 -1408
rect 3036 -1488 3132 -1472
rect 3036 -1552 3052 -1488
rect 3116 -1552 3132 -1488
rect 3036 -1568 3132 -1552
rect 3036 -1632 3052 -1568
rect 3116 -1632 3132 -1568
rect 3036 -1648 3132 -1632
rect 3036 -1712 3052 -1648
rect 3116 -1712 3132 -1648
rect 3036 -1728 3132 -1712
rect 3036 -1792 3052 -1728
rect 3116 -1792 3132 -1728
rect 3036 -1808 3132 -1792
rect 3036 -1872 3052 -1808
rect 3116 -1872 3132 -1808
rect 3036 -1888 3132 -1872
rect 3036 -1952 3052 -1888
rect 3116 -1952 3132 -1888
rect 3036 -1968 3132 -1952
rect 3036 -2032 3052 -1968
rect 3116 -2032 3132 -1968
rect 3036 -2048 3132 -2032
rect 3036 -2112 3052 -2048
rect 3116 -2112 3132 -2048
rect 3036 -2128 3132 -2112
rect 3036 -2192 3052 -2128
rect 3116 -2192 3132 -2128
rect 3036 -2208 3132 -2192
rect 3036 -2272 3052 -2208
rect 3116 -2272 3132 -2208
rect 3036 -2288 3132 -2272
rect 3036 -2352 3052 -2288
rect 3116 -2352 3132 -2288
rect 3036 -2368 3132 -2352
rect 3036 -2432 3052 -2368
rect 3116 -2432 3132 -2368
rect 3036 -2448 3132 -2432
rect 3036 -2512 3052 -2448
rect 3116 -2512 3132 -2448
rect 3036 -2528 3132 -2512
rect 3036 -2592 3052 -2528
rect 3116 -2592 3132 -2528
rect 3036 -2608 3132 -2592
rect 3036 -2672 3052 -2608
rect 3116 -2672 3132 -2608
rect 3036 -2688 3132 -2672
rect 3036 -2752 3052 -2688
rect 3116 -2752 3132 -2688
rect 3036 -2768 3132 -2752
rect 3036 -2832 3052 -2768
rect 3116 -2832 3132 -2768
rect 3036 -2848 3132 -2832
rect 3036 -2912 3052 -2848
rect 3116 -2912 3132 -2848
rect 3036 -2928 3132 -2912
rect 3036 -2992 3052 -2928
rect 3116 -2992 3132 -2928
rect 3036 -3008 3132 -2992
rect 3036 -3072 3052 -3008
rect 3116 -3072 3132 -3008
rect 3036 -3088 3132 -3072
<< properties >>
string FIXED_BBOX -3136 -3100 3064 3100
<< end >>
