magic
tech sky130A
magscale 1 2
timestamp 1620775510
<< xpolycontact >>
rect -35 2184 35 2616
rect -35 -2616 35 -2184
<< xpolyres >>
rect -35 -2184 35 2184
<< viali >>
rect -19 2201 19 2598
rect -19 -2598 19 -2201
<< metal1 >>
rect -25 2598 25 2610
rect -25 2201 -19 2598
rect 19 2201 25 2598
rect -25 2189 25 2201
rect -25 -2201 25 -2189
rect -25 -2598 -19 -2201
rect 19 -2598 25 -2201
rect -25 -2610 25 -2598
<< res0p35 >>
rect -37 -2186 37 2186
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 21.839 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 124.903k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
