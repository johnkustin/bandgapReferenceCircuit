magic
tech sky130A
magscale 1 2
timestamp 1620417585
<< xpolycontact >>
rect -1307 376 -1237 808
rect -1307 -808 -1237 -376
rect -989 376 -919 808
rect -989 -808 -919 -376
rect -671 376 -601 808
rect -671 -808 -601 -376
rect -353 376 -283 808
rect -353 -808 -283 -376
rect -35 376 35 808
rect -35 -808 35 -376
rect 283 376 353 808
rect 283 -808 353 -376
rect 601 376 671 808
rect 601 -808 671 -376
rect 919 376 989 808
rect 919 -808 989 -376
rect 1237 376 1307 808
rect 1237 -808 1307 -376
<< xpolyres >>
rect -1307 -376 -1237 376
rect -989 -376 -919 376
rect -671 -376 -601 376
rect -353 -376 -283 376
rect -35 -376 35 376
rect 283 -376 353 376
rect 601 -376 671 376
rect 919 -376 989 376
rect 1237 -376 1307 376
<< viali >>
rect -1291 393 -1253 790
rect -973 393 -935 790
rect -655 393 -617 790
rect -337 393 -299 790
rect -19 393 19 790
rect 299 393 337 790
rect 617 393 655 790
rect 935 393 973 790
rect 1253 393 1291 790
rect -1291 -790 -1253 -393
rect -973 -790 -935 -393
rect -655 -790 -617 -393
rect -337 -790 -299 -393
rect -19 -790 19 -393
rect 299 -790 337 -393
rect 617 -790 655 -393
rect 935 -790 973 -393
rect 1253 -790 1291 -393
<< metal1 >>
rect -1297 790 -1247 802
rect -1297 393 -1291 790
rect -1253 393 -1247 790
rect -1297 381 -1247 393
rect -979 790 -929 802
rect -979 393 -973 790
rect -935 393 -929 790
rect -979 381 -929 393
rect -661 790 -611 802
rect -661 393 -655 790
rect -617 393 -611 790
rect -661 381 -611 393
rect -343 790 -293 802
rect -343 393 -337 790
rect -299 393 -293 790
rect -343 381 -293 393
rect -25 790 25 802
rect -25 393 -19 790
rect 19 393 25 790
rect -25 381 25 393
rect 293 790 343 802
rect 293 393 299 790
rect 337 393 343 790
rect 293 381 343 393
rect 611 790 661 802
rect 611 393 617 790
rect 655 393 661 790
rect 611 381 661 393
rect 929 790 979 802
rect 929 393 935 790
rect 973 393 979 790
rect 929 381 979 393
rect 1247 790 1297 802
rect 1247 393 1253 790
rect 1291 393 1297 790
rect 1247 381 1297 393
rect -1297 -393 -1247 -381
rect -1297 -790 -1291 -393
rect -1253 -790 -1247 -393
rect -1297 -802 -1247 -790
rect -979 -393 -929 -381
rect -979 -790 -973 -393
rect -935 -790 -929 -393
rect -979 -802 -929 -790
rect -661 -393 -611 -381
rect -661 -790 -655 -393
rect -617 -790 -611 -393
rect -661 -802 -611 -790
rect -343 -393 -293 -381
rect -343 -790 -337 -393
rect -299 -790 -293 -393
rect -343 -802 -293 -790
rect -25 -393 25 -381
rect -25 -790 -19 -393
rect 19 -790 25 -393
rect -25 -802 25 -790
rect 293 -393 343 -381
rect 293 -790 299 -393
rect 337 -790 343 -393
rect 293 -802 343 -790
rect 611 -393 661 -381
rect 611 -790 617 -393
rect 655 -790 661 -393
rect 611 -802 661 -790
rect 929 -393 979 -381
rect 929 -790 935 -393
rect 973 -790 979 -393
rect 929 -802 979 -790
rect 1247 -393 1297 -381
rect 1247 -790 1253 -393
rect 1291 -790 1297 -393
rect 1247 -802 1297 -790
<< res0p35 >>
rect -1309 -378 -1235 378
rect -991 -378 -917 378
rect -673 -378 -599 378
rect -355 -378 -281 378
rect -37 -378 37 378
rect 281 -378 355 378
rect 599 -378 673 378
rect 917 -378 991 378
rect 1235 -378 1309 378
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 3.763 m 1 nx 9 wmin 0.350 lmin 0.50 rho 2000 val 22.188k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
