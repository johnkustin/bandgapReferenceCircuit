magic
tech sky130A
magscale 1 2
timestamp 1621196701
<< error_p >>
rect -8649 9500 -8589 15700
rect -8569 9500 -8509 15700
rect -2930 9500 -2870 15700
rect -2850 9500 -2790 15700
rect 2789 9500 2849 15700
rect 2869 9500 2929 15700
rect 8508 9500 8568 15700
rect 8588 9500 8648 15700
rect -8649 3200 -8589 9400
rect -8569 3200 -8509 9400
rect -2930 3200 -2870 9400
rect -2850 3200 -2790 9400
rect 2789 3200 2849 9400
rect 2869 3200 2929 9400
rect 8508 3200 8568 9400
rect 8588 3200 8648 9400
rect -8649 -3100 -8589 3100
rect -8569 -3100 -8509 3100
rect -2930 -3100 -2870 3100
rect -2850 -3100 -2790 3100
rect 2789 -3100 2849 3100
rect 2869 -3100 2929 3100
rect 8508 -3100 8568 3100
rect 8588 -3100 8648 3100
rect -8649 -9400 -8589 -3200
rect -8569 -9400 -8509 -3200
rect -2930 -9400 -2870 -3200
rect -2850 -9400 -2790 -3200
rect 2789 -9400 2849 -3200
rect 2869 -9400 2929 -3200
rect 8508 -9400 8568 -3200
rect 8588 -9400 8648 -3200
rect -8649 -15700 -8589 -9500
rect -8569 -15700 -8509 -9500
rect -2930 -15700 -2870 -9500
rect -2850 -15700 -2790 -9500
rect 2789 -15700 2849 -9500
rect 2869 -15700 2929 -9500
rect 8508 -15700 8568 -9500
rect 8588 -15700 8648 -9500
<< metal3 >>
rect -14288 15672 -8589 15700
rect -14288 9528 -8673 15672
rect -8609 9528 -8589 15672
rect -14288 9500 -8589 9528
rect -8569 15672 -2870 15700
rect -8569 9528 -2954 15672
rect -2890 9528 -2870 15672
rect -8569 9500 -2870 9528
rect -2850 15672 2849 15700
rect -2850 9528 2765 15672
rect 2829 9528 2849 15672
rect -2850 9500 2849 9528
rect 2869 15672 8568 15700
rect 2869 9528 8484 15672
rect 8548 9528 8568 15672
rect 2869 9500 8568 9528
rect 8588 15672 14287 15700
rect 8588 9528 14203 15672
rect 14267 9528 14287 15672
rect 8588 9500 14287 9528
rect -14288 9372 -8589 9400
rect -14288 3228 -8673 9372
rect -8609 3228 -8589 9372
rect -14288 3200 -8589 3228
rect -8569 9372 -2870 9400
rect -8569 3228 -2954 9372
rect -2890 3228 -2870 9372
rect -8569 3200 -2870 3228
rect -2850 9372 2849 9400
rect -2850 3228 2765 9372
rect 2829 3228 2849 9372
rect -2850 3200 2849 3228
rect 2869 9372 8568 9400
rect 2869 3228 8484 9372
rect 8548 3228 8568 9372
rect 2869 3200 8568 3228
rect 8588 9372 14287 9400
rect 8588 3228 14203 9372
rect 14267 3228 14287 9372
rect 8588 3200 14287 3228
rect -14288 3072 -8589 3100
rect -14288 -3072 -8673 3072
rect -8609 -3072 -8589 3072
rect -14288 -3100 -8589 -3072
rect -8569 3072 -2870 3100
rect -8569 -3072 -2954 3072
rect -2890 -3072 -2870 3072
rect -8569 -3100 -2870 -3072
rect -2850 3072 2849 3100
rect -2850 -3072 2765 3072
rect 2829 -3072 2849 3072
rect -2850 -3100 2849 -3072
rect 2869 3072 8568 3100
rect 2869 -3072 8484 3072
rect 8548 -3072 8568 3072
rect 2869 -3100 8568 -3072
rect 8588 3072 14287 3100
rect 8588 -3072 14203 3072
rect 14267 -3072 14287 3072
rect 8588 -3100 14287 -3072
rect -14288 -3228 -8589 -3200
rect -14288 -9372 -8673 -3228
rect -8609 -9372 -8589 -3228
rect -14288 -9400 -8589 -9372
rect -8569 -3228 -2870 -3200
rect -8569 -9372 -2954 -3228
rect -2890 -9372 -2870 -3228
rect -8569 -9400 -2870 -9372
rect -2850 -3228 2849 -3200
rect -2850 -9372 2765 -3228
rect 2829 -9372 2849 -3228
rect -2850 -9400 2849 -9372
rect 2869 -3228 8568 -3200
rect 2869 -9372 8484 -3228
rect 8548 -9372 8568 -3228
rect 2869 -9400 8568 -9372
rect 8588 -3228 14287 -3200
rect 8588 -9372 14203 -3228
rect 14267 -9372 14287 -3228
rect 8588 -9400 14287 -9372
rect -14288 -9528 -8589 -9500
rect -14288 -15672 -8673 -9528
rect -8609 -15672 -8589 -9528
rect -14288 -15700 -8589 -15672
rect -8569 -9528 -2870 -9500
rect -8569 -15672 -2954 -9528
rect -2890 -15672 -2870 -9528
rect -8569 -15700 -2870 -15672
rect -2850 -9528 2849 -9500
rect -2850 -15672 2765 -9528
rect 2829 -15672 2849 -9528
rect -2850 -15700 2849 -15672
rect 2869 -9528 8568 -9500
rect 2869 -15672 8484 -9528
rect 8548 -15672 8568 -9528
rect 2869 -15700 8568 -15672
rect 8588 -9528 14287 -9500
rect 8588 -15672 14203 -9528
rect 14267 -15672 14287 -9528
rect 8588 -15700 14287 -15672
<< via3 >>
rect -8673 9528 -8609 15672
rect -2954 9528 -2890 15672
rect 2765 9528 2829 15672
rect 8484 9528 8548 15672
rect 14203 9528 14267 15672
rect -8673 3228 -8609 9372
rect -2954 3228 -2890 9372
rect 2765 3228 2829 9372
rect 8484 3228 8548 9372
rect 14203 3228 14267 9372
rect -8673 -3072 -8609 3072
rect -2954 -3072 -2890 3072
rect 2765 -3072 2829 3072
rect 8484 -3072 8548 3072
rect 14203 -3072 14267 3072
rect -8673 -9372 -8609 -3228
rect -2954 -9372 -2890 -3228
rect 2765 -9372 2829 -3228
rect 8484 -9372 8548 -3228
rect 14203 -9372 14267 -3228
rect -8673 -15672 -8609 -9528
rect -2954 -15672 -2890 -9528
rect 2765 -15672 2829 -9528
rect 8484 -15672 8548 -9528
rect 14203 -15672 14267 -9528
<< mimcap >>
rect -14188 15560 -8788 15600
rect -14188 9640 -14148 15560
rect -8828 9640 -8788 15560
rect -14188 9600 -8788 9640
rect -8469 15560 -3069 15600
rect -8469 9640 -8429 15560
rect -3109 9640 -3069 15560
rect -8469 9600 -3069 9640
rect -2750 15560 2650 15600
rect -2750 9640 -2710 15560
rect 2610 9640 2650 15560
rect -2750 9600 2650 9640
rect 2969 15560 8369 15600
rect 2969 9640 3009 15560
rect 8329 9640 8369 15560
rect 2969 9600 8369 9640
rect 8688 15560 14088 15600
rect 8688 9640 8728 15560
rect 14048 9640 14088 15560
rect 8688 9600 14088 9640
rect -14188 9260 -8788 9300
rect -14188 3340 -14148 9260
rect -8828 3340 -8788 9260
rect -14188 3300 -8788 3340
rect -8469 9260 -3069 9300
rect -8469 3340 -8429 9260
rect -3109 3340 -3069 9260
rect -8469 3300 -3069 3340
rect -2750 9260 2650 9300
rect -2750 3340 -2710 9260
rect 2610 3340 2650 9260
rect -2750 3300 2650 3340
rect 2969 9260 8369 9300
rect 2969 3340 3009 9260
rect 8329 3340 8369 9260
rect 2969 3300 8369 3340
rect 8688 9260 14088 9300
rect 8688 3340 8728 9260
rect 14048 3340 14088 9260
rect 8688 3300 14088 3340
rect -14188 2960 -8788 3000
rect -14188 -2960 -14148 2960
rect -8828 -2960 -8788 2960
rect -14188 -3000 -8788 -2960
rect -8469 2960 -3069 3000
rect -8469 -2960 -8429 2960
rect -3109 -2960 -3069 2960
rect -8469 -3000 -3069 -2960
rect -2750 2960 2650 3000
rect -2750 -2960 -2710 2960
rect 2610 -2960 2650 2960
rect -2750 -3000 2650 -2960
rect 2969 2960 8369 3000
rect 2969 -2960 3009 2960
rect 8329 -2960 8369 2960
rect 2969 -3000 8369 -2960
rect 8688 2960 14088 3000
rect 8688 -2960 8728 2960
rect 14048 -2960 14088 2960
rect 8688 -3000 14088 -2960
rect -14188 -3340 -8788 -3300
rect -14188 -9260 -14148 -3340
rect -8828 -9260 -8788 -3340
rect -14188 -9300 -8788 -9260
rect -8469 -3340 -3069 -3300
rect -8469 -9260 -8429 -3340
rect -3109 -9260 -3069 -3340
rect -8469 -9300 -3069 -9260
rect -2750 -3340 2650 -3300
rect -2750 -9260 -2710 -3340
rect 2610 -9260 2650 -3340
rect -2750 -9300 2650 -9260
rect 2969 -3340 8369 -3300
rect 2969 -9260 3009 -3340
rect 8329 -9260 8369 -3340
rect 2969 -9300 8369 -9260
rect 8688 -3340 14088 -3300
rect 8688 -9260 8728 -3340
rect 14048 -9260 14088 -3340
rect 8688 -9300 14088 -9260
rect -14188 -9640 -8788 -9600
rect -14188 -15560 -14148 -9640
rect -8828 -15560 -8788 -9640
rect -14188 -15600 -8788 -15560
rect -8469 -9640 -3069 -9600
rect -8469 -15560 -8429 -9640
rect -3109 -15560 -3069 -9640
rect -8469 -15600 -3069 -15560
rect -2750 -9640 2650 -9600
rect -2750 -15560 -2710 -9640
rect 2610 -15560 2650 -9640
rect -2750 -15600 2650 -15560
rect 2969 -9640 8369 -9600
rect 2969 -15560 3009 -9640
rect 8329 -15560 8369 -9640
rect 2969 -15600 8369 -15560
rect 8688 -9640 14088 -9600
rect 8688 -15560 8728 -9640
rect 14048 -15560 14088 -9640
rect 8688 -15600 14088 -15560
<< mimcapcontact >>
rect -14148 9640 -8828 15560
rect -8429 9640 -3109 15560
rect -2710 9640 2610 15560
rect 3009 9640 8329 15560
rect 8728 9640 14048 15560
rect -14148 3340 -8828 9260
rect -8429 3340 -3109 9260
rect -2710 3340 2610 9260
rect 3009 3340 8329 9260
rect 8728 3340 14048 9260
rect -14148 -2960 -8828 2960
rect -8429 -2960 -3109 2960
rect -2710 -2960 2610 2960
rect 3009 -2960 8329 2960
rect 8728 -2960 14048 2960
rect -14148 -9260 -8828 -3340
rect -8429 -9260 -3109 -3340
rect -2710 -9260 2610 -3340
rect 3009 -9260 8329 -3340
rect 8728 -9260 14048 -3340
rect -14148 -15560 -8828 -9640
rect -8429 -15560 -3109 -9640
rect -2710 -15560 2610 -9640
rect 3009 -15560 8329 -9640
rect 8728 -15560 14048 -9640
<< metal4 >>
rect -11540 15561 -11436 15750
rect -8720 15688 -8616 15750
rect -8720 15672 -8593 15688
rect -14149 15560 -8827 15561
rect -14149 9640 -14148 15560
rect -8828 9640 -8827 15560
rect -14149 9639 -8827 9640
rect -11540 9261 -11436 9639
rect -8720 9528 -8673 15672
rect -8609 9528 -8593 15672
rect -5821 15561 -5717 15750
rect -3001 15688 -2897 15750
rect -3001 15672 -2874 15688
rect -8430 15560 -3108 15561
rect -8430 9640 -8429 15560
rect -3109 9640 -3108 15560
rect -8430 9639 -3108 9640
rect -8720 9512 -8593 9528
rect -8720 9388 -8616 9512
rect -8720 9372 -8593 9388
rect -14149 9260 -8827 9261
rect -14149 3340 -14148 9260
rect -8828 3340 -8827 9260
rect -14149 3339 -8827 3340
rect -11540 2961 -11436 3339
rect -8720 3228 -8673 9372
rect -8609 3228 -8593 9372
rect -5821 9261 -5717 9639
rect -3001 9528 -2954 15672
rect -2890 9528 -2874 15672
rect -102 15561 2 15750
rect 2718 15688 2822 15750
rect 2718 15672 2845 15688
rect -2711 15560 2611 15561
rect -2711 9640 -2710 15560
rect 2610 9640 2611 15560
rect -2711 9639 2611 9640
rect -3001 9512 -2874 9528
rect -3001 9388 -2897 9512
rect -3001 9372 -2874 9388
rect -8430 9260 -3108 9261
rect -8430 3340 -8429 9260
rect -3109 3340 -3108 9260
rect -8430 3339 -3108 3340
rect -8720 3212 -8593 3228
rect -8720 3088 -8616 3212
rect -8720 3072 -8593 3088
rect -14149 2960 -8827 2961
rect -14149 -2960 -14148 2960
rect -8828 -2960 -8827 2960
rect -14149 -2961 -8827 -2960
rect -11540 -3339 -11436 -2961
rect -8720 -3072 -8673 3072
rect -8609 -3072 -8593 3072
rect -5821 2961 -5717 3339
rect -3001 3228 -2954 9372
rect -2890 3228 -2874 9372
rect -102 9261 2 9639
rect 2718 9528 2765 15672
rect 2829 9528 2845 15672
rect 5617 15561 5721 15750
rect 8437 15688 8541 15750
rect 8437 15672 8564 15688
rect 3008 15560 8330 15561
rect 3008 9640 3009 15560
rect 8329 9640 8330 15560
rect 3008 9639 8330 9640
rect 2718 9512 2845 9528
rect 2718 9388 2822 9512
rect 2718 9372 2845 9388
rect -2711 9260 2611 9261
rect -2711 3340 -2710 9260
rect 2610 3340 2611 9260
rect -2711 3339 2611 3340
rect -3001 3212 -2874 3228
rect -3001 3088 -2897 3212
rect -3001 3072 -2874 3088
rect -8430 2960 -3108 2961
rect -8430 -2960 -8429 2960
rect -3109 -2960 -3108 2960
rect -8430 -2961 -3108 -2960
rect -8720 -3088 -8593 -3072
rect -8720 -3212 -8616 -3088
rect -8720 -3228 -8593 -3212
rect -14149 -3340 -8827 -3339
rect -14149 -9260 -14148 -3340
rect -8828 -9260 -8827 -3340
rect -14149 -9261 -8827 -9260
rect -11540 -9639 -11436 -9261
rect -8720 -9372 -8673 -3228
rect -8609 -9372 -8593 -3228
rect -5821 -3339 -5717 -2961
rect -3001 -3072 -2954 3072
rect -2890 -3072 -2874 3072
rect -102 2961 2 3339
rect 2718 3228 2765 9372
rect 2829 3228 2845 9372
rect 5617 9261 5721 9639
rect 8437 9528 8484 15672
rect 8548 9528 8564 15672
rect 11336 15561 11440 15750
rect 14156 15688 14260 15750
rect 14156 15672 14283 15688
rect 8727 15560 14049 15561
rect 8727 9640 8728 15560
rect 14048 9640 14049 15560
rect 8727 9639 14049 9640
rect 8437 9512 8564 9528
rect 8437 9388 8541 9512
rect 8437 9372 8564 9388
rect 3008 9260 8330 9261
rect 3008 3340 3009 9260
rect 8329 3340 8330 9260
rect 3008 3339 8330 3340
rect 2718 3212 2845 3228
rect 2718 3088 2822 3212
rect 2718 3072 2845 3088
rect -2711 2960 2611 2961
rect -2711 -2960 -2710 2960
rect 2610 -2960 2611 2960
rect -2711 -2961 2611 -2960
rect -3001 -3088 -2874 -3072
rect -3001 -3212 -2897 -3088
rect -3001 -3228 -2874 -3212
rect -8430 -3340 -3108 -3339
rect -8430 -9260 -8429 -3340
rect -3109 -9260 -3108 -3340
rect -8430 -9261 -3108 -9260
rect -8720 -9388 -8593 -9372
rect -8720 -9512 -8616 -9388
rect -8720 -9528 -8593 -9512
rect -14149 -9640 -8827 -9639
rect -14149 -15560 -14148 -9640
rect -8828 -15560 -8827 -9640
rect -14149 -15561 -8827 -15560
rect -11540 -15750 -11436 -15561
rect -8720 -15672 -8673 -9528
rect -8609 -15672 -8593 -9528
rect -5821 -9639 -5717 -9261
rect -3001 -9372 -2954 -3228
rect -2890 -9372 -2874 -3228
rect -102 -3339 2 -2961
rect 2718 -3072 2765 3072
rect 2829 -3072 2845 3072
rect 5617 2961 5721 3339
rect 8437 3228 8484 9372
rect 8548 3228 8564 9372
rect 11336 9261 11440 9639
rect 14156 9528 14203 15672
rect 14267 9528 14283 15672
rect 14156 9512 14283 9528
rect 14156 9388 14260 9512
rect 14156 9372 14283 9388
rect 8727 9260 14049 9261
rect 8727 3340 8728 9260
rect 14048 3340 14049 9260
rect 8727 3339 14049 3340
rect 8437 3212 8564 3228
rect 8437 3088 8541 3212
rect 8437 3072 8564 3088
rect 3008 2960 8330 2961
rect 3008 -2960 3009 2960
rect 8329 -2960 8330 2960
rect 3008 -2961 8330 -2960
rect 2718 -3088 2845 -3072
rect 2718 -3212 2822 -3088
rect 2718 -3228 2845 -3212
rect -2711 -3340 2611 -3339
rect -2711 -9260 -2710 -3340
rect 2610 -9260 2611 -3340
rect -2711 -9261 2611 -9260
rect -3001 -9388 -2874 -9372
rect -3001 -9512 -2897 -9388
rect -3001 -9528 -2874 -9512
rect -8430 -9640 -3108 -9639
rect -8430 -15560 -8429 -9640
rect -3109 -15560 -3108 -9640
rect -8430 -15561 -3108 -15560
rect -8720 -15688 -8593 -15672
rect -8720 -15750 -8616 -15688
rect -5821 -15750 -5717 -15561
rect -3001 -15672 -2954 -9528
rect -2890 -15672 -2874 -9528
rect -102 -9639 2 -9261
rect 2718 -9372 2765 -3228
rect 2829 -9372 2845 -3228
rect 5617 -3339 5721 -2961
rect 8437 -3072 8484 3072
rect 8548 -3072 8564 3072
rect 11336 2961 11440 3339
rect 14156 3228 14203 9372
rect 14267 3228 14283 9372
rect 14156 3212 14283 3228
rect 14156 3088 14260 3212
rect 14156 3072 14283 3088
rect 8727 2960 14049 2961
rect 8727 -2960 8728 2960
rect 14048 -2960 14049 2960
rect 8727 -2961 14049 -2960
rect 8437 -3088 8564 -3072
rect 8437 -3212 8541 -3088
rect 8437 -3228 8564 -3212
rect 3008 -3340 8330 -3339
rect 3008 -9260 3009 -3340
rect 8329 -9260 8330 -3340
rect 3008 -9261 8330 -9260
rect 2718 -9388 2845 -9372
rect 2718 -9512 2822 -9388
rect 2718 -9528 2845 -9512
rect -2711 -9640 2611 -9639
rect -2711 -15560 -2710 -9640
rect 2610 -15560 2611 -9640
rect -2711 -15561 2611 -15560
rect -3001 -15688 -2874 -15672
rect -3001 -15750 -2897 -15688
rect -102 -15750 2 -15561
rect 2718 -15672 2765 -9528
rect 2829 -15672 2845 -9528
rect 5617 -9639 5721 -9261
rect 8437 -9372 8484 -3228
rect 8548 -9372 8564 -3228
rect 11336 -3339 11440 -2961
rect 14156 -3072 14203 3072
rect 14267 -3072 14283 3072
rect 14156 -3088 14283 -3072
rect 14156 -3212 14260 -3088
rect 14156 -3228 14283 -3212
rect 8727 -3340 14049 -3339
rect 8727 -9260 8728 -3340
rect 14048 -9260 14049 -3340
rect 8727 -9261 14049 -9260
rect 8437 -9388 8564 -9372
rect 8437 -9512 8541 -9388
rect 8437 -9528 8564 -9512
rect 3008 -9640 8330 -9639
rect 3008 -15560 3009 -9640
rect 8329 -15560 8330 -9640
rect 3008 -15561 8330 -15560
rect 2718 -15688 2845 -15672
rect 2718 -15750 2822 -15688
rect 5617 -15750 5721 -15561
rect 8437 -15672 8484 -9528
rect 8548 -15672 8564 -9528
rect 11336 -9639 11440 -9261
rect 14156 -9372 14203 -3228
rect 14267 -9372 14283 -3228
rect 14156 -9388 14283 -9372
rect 14156 -9512 14260 -9388
rect 14156 -9528 14283 -9512
rect 8727 -9640 14049 -9639
rect 8727 -15560 8728 -9640
rect 14048 -15560 14049 -9640
rect 8727 -15561 14049 -15560
rect 8437 -15688 8564 -15672
rect 8437 -15750 8541 -15688
rect 11336 -15750 11440 -15561
rect 14156 -15672 14203 -9528
rect 14267 -15672 14283 -9528
rect 14156 -15688 14283 -15672
rect 14156 -15750 14260 -15688
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 8588 9500 14188 15700
string parameters w 27 l 30 val 829.38 carea 1.00 cperi 0.17 nx 5 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
