magic
tech sky130A
magscale 1 2
timestamp 1621229569
<< nmoslvt >>
rect -200 -2731 200 2669
<< ndiff >>
rect -258 2657 -200 2669
rect -258 -2719 -246 2657
rect -212 -2719 -200 2657
rect -258 -2731 -200 -2719
rect 200 2657 258 2669
rect 200 -2719 212 2657
rect 246 -2719 258 2657
rect 200 -2731 258 -2719
<< ndiffc >>
rect -246 -2719 -212 2657
rect 212 -2719 246 2657
<< poly >>
rect -200 2741 200 2757
rect -200 2707 -184 2741
rect 184 2707 200 2741
rect -200 2669 200 2707
rect -200 -2757 200 -2731
<< polycont >>
rect -184 2707 184 2741
<< locali >>
rect -200 2707 -184 2741
rect 184 2707 200 2741
rect -246 2657 -212 2673
rect -246 -2735 -212 -2719
rect 212 2657 246 2673
rect 212 -2735 246 -2719
<< viali >>
rect -184 2707 184 2741
rect -246 -2719 -212 2657
rect 212 -2719 246 2657
<< metal1 >>
rect -196 2741 196 2747
rect -196 2707 -184 2741
rect 184 2707 196 2741
rect -196 2701 196 2707
rect -252 2657 -206 2669
rect -252 -2719 -246 2657
rect -212 -2719 -206 2657
rect -252 -2731 -206 -2719
rect 206 2657 252 2669
rect 206 -2719 212 2657
rect 246 -2719 252 2657
rect 206 -2731 252 -2719
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 27 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
