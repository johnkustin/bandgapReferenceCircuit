magic
tech sky130A
magscale 1 2
timestamp 1620316209
<< nwell >>
rect -294 -4400 294 4400
<< pmoslvt >>
rect -200 -4300 200 4300
<< pdiff >>
rect -258 4288 -200 4300
rect -258 -4288 -246 4288
rect -212 -4288 -200 4288
rect -258 -4300 -200 -4288
rect 200 4288 258 4300
rect 200 -4288 212 4288
rect 246 -4288 258 4288
rect 200 -4300 258 -4288
<< pdiffc >>
rect -246 -4288 -212 4288
rect 212 -4288 246 4288
<< poly >>
rect -200 4381 200 4397
rect -200 4347 -184 4381
rect 184 4347 200 4381
rect -200 4300 200 4347
rect -200 -4347 200 -4300
rect -200 -4381 -184 -4347
rect 184 -4381 200 -4347
rect -200 -4397 200 -4381
<< polycont >>
rect -184 4347 184 4381
rect -184 -4381 184 -4347
<< locali >>
rect -200 4347 -184 4381
rect 184 4347 200 4381
rect -246 4288 -212 4304
rect -246 -4304 -212 -4288
rect 212 4288 246 4304
rect 212 -4304 246 -4288
rect -200 -4381 -184 -4347
rect 184 -4381 200 -4347
<< viali >>
rect -184 4347 184 4381
rect -246 -4288 -212 4288
rect 212 -4288 246 4288
rect -184 -4381 184 -4347
<< metal1 >>
rect -196 4381 196 4387
rect -196 4347 -184 4381
rect 184 4347 196 4381
rect -196 4341 196 4347
rect -252 4288 -206 4300
rect -252 -4288 -246 4288
rect -212 -4288 -206 4288
rect -252 -4300 -206 -4288
rect 206 4288 252 4300
rect 206 -4288 212 4288
rect 246 -4288 252 4288
rect 206 -4300 252 -4288
rect -196 -4347 196 -4341
rect -196 -4381 -184 -4347
rect 184 -4381 196 -4347
rect -196 -4387 196 -4381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 43 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
