magic
tech sky130A
magscale 1 2
timestamp 1621231152
<< error_p >>
rect -2926 2850 -2886 3450
rect -2866 2850 -2826 3450
rect -2207 2850 -2167 3450
rect -2147 2850 -2107 3450
rect -1488 2850 -1448 3450
rect -1428 2850 -1388 3450
rect -769 2850 -729 3450
rect -709 2850 -669 3450
rect -50 2850 -10 3450
rect 10 2850 50 3450
rect 669 2850 709 3450
rect 729 2850 769 3450
rect 1388 2850 1428 3450
rect 1448 2850 1488 3450
rect 2107 2850 2147 3450
rect 2167 2850 2207 3450
rect 2826 2850 2866 3450
rect 2886 2850 2926 3450
rect -2926 2150 -2886 2750
rect -2866 2150 -2826 2750
rect -2207 2150 -2167 2750
rect -2147 2150 -2107 2750
rect -1488 2150 -1448 2750
rect -1428 2150 -1388 2750
rect -769 2150 -729 2750
rect -709 2150 -669 2750
rect -50 2150 -10 2750
rect 10 2150 50 2750
rect 669 2150 709 2750
rect 729 2150 769 2750
rect 1388 2150 1428 2750
rect 1448 2150 1488 2750
rect 2107 2150 2147 2750
rect 2167 2150 2207 2750
rect 2826 2150 2866 2750
rect 2886 2150 2926 2750
rect -2926 1450 -2886 2050
rect -2866 1450 -2826 2050
rect -2207 1450 -2167 2050
rect -2147 1450 -2107 2050
rect -1488 1450 -1448 2050
rect -1428 1450 -1388 2050
rect -769 1450 -729 2050
rect -709 1450 -669 2050
rect -50 1450 -10 2050
rect 10 1450 50 2050
rect 669 1450 709 2050
rect 729 1450 769 2050
rect 1388 1450 1428 2050
rect 1448 1450 1488 2050
rect 2107 1450 2147 2050
rect 2167 1450 2207 2050
rect 2826 1450 2866 2050
rect 2886 1450 2926 2050
rect -2926 750 -2886 1350
rect -2866 750 -2826 1350
rect -2207 750 -2167 1350
rect -2147 750 -2107 1350
rect -1488 750 -1448 1350
rect -1428 750 -1388 1350
rect -769 750 -729 1350
rect -709 750 -669 1350
rect -50 750 -10 1350
rect 10 750 50 1350
rect 669 750 709 1350
rect 729 750 769 1350
rect 1388 750 1428 1350
rect 1448 750 1488 1350
rect 2107 750 2147 1350
rect 2167 750 2207 1350
rect 2826 750 2866 1350
rect 2886 750 2926 1350
rect -2926 50 -2886 650
rect -2866 50 -2826 650
rect -2207 50 -2167 650
rect -2147 50 -2107 650
rect -1488 50 -1448 650
rect -1428 50 -1388 650
rect -769 50 -729 650
rect -709 50 -669 650
rect -50 50 -10 650
rect 10 50 50 650
rect 669 50 709 650
rect 729 50 769 650
rect 1388 50 1428 650
rect 1448 50 1488 650
rect 2107 50 2147 650
rect 2167 50 2207 650
rect 2826 50 2866 650
rect 2886 50 2926 650
rect -2926 -650 -2886 -50
rect -2866 -650 -2826 -50
rect -2207 -650 -2167 -50
rect -2147 -650 -2107 -50
rect -1488 -650 -1448 -50
rect -1428 -650 -1388 -50
rect -769 -650 -729 -50
rect -709 -650 -669 -50
rect -50 -650 -10 -50
rect 10 -650 50 -50
rect 669 -650 709 -50
rect 729 -650 769 -50
rect 1388 -650 1428 -50
rect 1448 -650 1488 -50
rect 2107 -650 2147 -50
rect 2167 -650 2207 -50
rect 2826 -650 2866 -50
rect 2886 -650 2926 -50
rect -2926 -1350 -2886 -750
rect -2866 -1350 -2826 -750
rect -2207 -1350 -2167 -750
rect -2147 -1350 -2107 -750
rect -1488 -1350 -1448 -750
rect -1428 -1350 -1388 -750
rect -769 -1350 -729 -750
rect -709 -1350 -669 -750
rect -50 -1350 -10 -750
rect 10 -1350 50 -750
rect 669 -1350 709 -750
rect 729 -1350 769 -750
rect 1388 -1350 1428 -750
rect 1448 -1350 1488 -750
rect 2107 -1350 2147 -750
rect 2167 -1350 2207 -750
rect 2826 -1350 2866 -750
rect 2886 -1350 2926 -750
rect -2926 -2050 -2886 -1450
rect -2866 -2050 -2826 -1450
rect -2207 -2050 -2167 -1450
rect -2147 -2050 -2107 -1450
rect -1488 -2050 -1448 -1450
rect -1428 -2050 -1388 -1450
rect -769 -2050 -729 -1450
rect -709 -2050 -669 -1450
rect -50 -2050 -10 -1450
rect 10 -2050 50 -1450
rect 669 -2050 709 -1450
rect 729 -2050 769 -1450
rect 1388 -2050 1428 -1450
rect 1448 -2050 1488 -1450
rect 2107 -2050 2147 -1450
rect 2167 -2050 2207 -1450
rect 2826 -2050 2866 -1450
rect 2886 -2050 2926 -1450
rect -2926 -2750 -2886 -2150
rect -2866 -2750 -2826 -2150
rect -2207 -2750 -2167 -2150
rect -2147 -2750 -2107 -2150
rect -1488 -2750 -1448 -2150
rect -1428 -2750 -1388 -2150
rect -769 -2750 -729 -2150
rect -709 -2750 -669 -2150
rect -50 -2750 -10 -2150
rect 10 -2750 50 -2150
rect 669 -2750 709 -2150
rect 729 -2750 769 -2150
rect 1388 -2750 1428 -2150
rect 1448 -2750 1488 -2150
rect 2107 -2750 2147 -2150
rect 2167 -2750 2207 -2150
rect 2826 -2750 2866 -2150
rect 2886 -2750 2926 -2150
rect -2926 -3450 -2886 -2850
rect -2866 -3450 -2826 -2850
rect -2207 -3450 -2167 -2850
rect -2147 -3450 -2107 -2850
rect -1488 -3450 -1448 -2850
rect -1428 -3450 -1388 -2850
rect -769 -3450 -729 -2850
rect -709 -3450 -669 -2850
rect -50 -3450 -10 -2850
rect 10 -3450 50 -2850
rect 669 -3450 709 -2850
rect 729 -3450 769 -2850
rect 1388 -3450 1428 -2850
rect 1448 -3450 1488 -2850
rect 2107 -3450 2147 -2850
rect 2167 -3450 2207 -2850
rect 2826 -3450 2866 -2850
rect 2886 -3450 2926 -2850
<< metal3 >>
rect -3585 3422 -2886 3450
rect -3585 2878 -2970 3422
rect -2906 2878 -2886 3422
rect -3585 2850 -2886 2878
rect -2866 3422 -2167 3450
rect -2866 2878 -2251 3422
rect -2187 2878 -2167 3422
rect -2866 2850 -2167 2878
rect -2147 3422 -1448 3450
rect -2147 2878 -1532 3422
rect -1468 2878 -1448 3422
rect -2147 2850 -1448 2878
rect -1428 3422 -729 3450
rect -1428 2878 -813 3422
rect -749 2878 -729 3422
rect -1428 2850 -729 2878
rect -709 3422 -10 3450
rect -709 2878 -94 3422
rect -30 2878 -10 3422
rect -709 2850 -10 2878
rect 10 3422 709 3450
rect 10 2878 625 3422
rect 689 2878 709 3422
rect 10 2850 709 2878
rect 729 3422 1428 3450
rect 729 2878 1344 3422
rect 1408 2878 1428 3422
rect 729 2850 1428 2878
rect 1448 3422 2147 3450
rect 1448 2878 2063 3422
rect 2127 2878 2147 3422
rect 1448 2850 2147 2878
rect 2167 3422 2866 3450
rect 2167 2878 2782 3422
rect 2846 2878 2866 3422
rect 2167 2850 2866 2878
rect 2886 3422 3585 3450
rect 2886 2878 3501 3422
rect 3565 2878 3585 3422
rect 2886 2850 3585 2878
rect -3585 2722 -2886 2750
rect -3585 2178 -2970 2722
rect -2906 2178 -2886 2722
rect -3585 2150 -2886 2178
rect -2866 2722 -2167 2750
rect -2866 2178 -2251 2722
rect -2187 2178 -2167 2722
rect -2866 2150 -2167 2178
rect -2147 2722 -1448 2750
rect -2147 2178 -1532 2722
rect -1468 2178 -1448 2722
rect -2147 2150 -1448 2178
rect -1428 2722 -729 2750
rect -1428 2178 -813 2722
rect -749 2178 -729 2722
rect -1428 2150 -729 2178
rect -709 2722 -10 2750
rect -709 2178 -94 2722
rect -30 2178 -10 2722
rect -709 2150 -10 2178
rect 10 2722 709 2750
rect 10 2178 625 2722
rect 689 2178 709 2722
rect 10 2150 709 2178
rect 729 2722 1428 2750
rect 729 2178 1344 2722
rect 1408 2178 1428 2722
rect 729 2150 1428 2178
rect 1448 2722 2147 2750
rect 1448 2178 2063 2722
rect 2127 2178 2147 2722
rect 1448 2150 2147 2178
rect 2167 2722 2866 2750
rect 2167 2178 2782 2722
rect 2846 2178 2866 2722
rect 2167 2150 2866 2178
rect 2886 2722 3585 2750
rect 2886 2178 3501 2722
rect 3565 2178 3585 2722
rect 2886 2150 3585 2178
rect -3585 2022 -2886 2050
rect -3585 1478 -2970 2022
rect -2906 1478 -2886 2022
rect -3585 1450 -2886 1478
rect -2866 2022 -2167 2050
rect -2866 1478 -2251 2022
rect -2187 1478 -2167 2022
rect -2866 1450 -2167 1478
rect -2147 2022 -1448 2050
rect -2147 1478 -1532 2022
rect -1468 1478 -1448 2022
rect -2147 1450 -1448 1478
rect -1428 2022 -729 2050
rect -1428 1478 -813 2022
rect -749 1478 -729 2022
rect -1428 1450 -729 1478
rect -709 2022 -10 2050
rect -709 1478 -94 2022
rect -30 1478 -10 2022
rect -709 1450 -10 1478
rect 10 2022 709 2050
rect 10 1478 625 2022
rect 689 1478 709 2022
rect 10 1450 709 1478
rect 729 2022 1428 2050
rect 729 1478 1344 2022
rect 1408 1478 1428 2022
rect 729 1450 1428 1478
rect 1448 2022 2147 2050
rect 1448 1478 2063 2022
rect 2127 1478 2147 2022
rect 1448 1450 2147 1478
rect 2167 2022 2866 2050
rect 2167 1478 2782 2022
rect 2846 1478 2866 2022
rect 2167 1450 2866 1478
rect 2886 2022 3585 2050
rect 2886 1478 3501 2022
rect 3565 1478 3585 2022
rect 2886 1450 3585 1478
rect -3585 1322 -2886 1350
rect -3585 778 -2970 1322
rect -2906 778 -2886 1322
rect -3585 750 -2886 778
rect -2866 1322 -2167 1350
rect -2866 778 -2251 1322
rect -2187 778 -2167 1322
rect -2866 750 -2167 778
rect -2147 1322 -1448 1350
rect -2147 778 -1532 1322
rect -1468 778 -1448 1322
rect -2147 750 -1448 778
rect -1428 1322 -729 1350
rect -1428 778 -813 1322
rect -749 778 -729 1322
rect -1428 750 -729 778
rect -709 1322 -10 1350
rect -709 778 -94 1322
rect -30 778 -10 1322
rect -709 750 -10 778
rect 10 1322 709 1350
rect 10 778 625 1322
rect 689 778 709 1322
rect 10 750 709 778
rect 729 1322 1428 1350
rect 729 778 1344 1322
rect 1408 778 1428 1322
rect 729 750 1428 778
rect 1448 1322 2147 1350
rect 1448 778 2063 1322
rect 2127 778 2147 1322
rect 1448 750 2147 778
rect 2167 1322 2866 1350
rect 2167 778 2782 1322
rect 2846 778 2866 1322
rect 2167 750 2866 778
rect 2886 1322 3585 1350
rect 2886 778 3501 1322
rect 3565 778 3585 1322
rect 2886 750 3585 778
rect -3585 622 -2886 650
rect -3585 78 -2970 622
rect -2906 78 -2886 622
rect -3585 50 -2886 78
rect -2866 622 -2167 650
rect -2866 78 -2251 622
rect -2187 78 -2167 622
rect -2866 50 -2167 78
rect -2147 622 -1448 650
rect -2147 78 -1532 622
rect -1468 78 -1448 622
rect -2147 50 -1448 78
rect -1428 622 -729 650
rect -1428 78 -813 622
rect -749 78 -729 622
rect -1428 50 -729 78
rect -709 622 -10 650
rect -709 78 -94 622
rect -30 78 -10 622
rect -709 50 -10 78
rect 10 622 709 650
rect 10 78 625 622
rect 689 78 709 622
rect 10 50 709 78
rect 729 622 1428 650
rect 729 78 1344 622
rect 1408 78 1428 622
rect 729 50 1428 78
rect 1448 622 2147 650
rect 1448 78 2063 622
rect 2127 78 2147 622
rect 1448 50 2147 78
rect 2167 622 2866 650
rect 2167 78 2782 622
rect 2846 78 2866 622
rect 2167 50 2866 78
rect 2886 622 3585 650
rect 2886 78 3501 622
rect 3565 78 3585 622
rect 2886 50 3585 78
rect -3585 -78 -2886 -50
rect -3585 -622 -2970 -78
rect -2906 -622 -2886 -78
rect -3585 -650 -2886 -622
rect -2866 -78 -2167 -50
rect -2866 -622 -2251 -78
rect -2187 -622 -2167 -78
rect -2866 -650 -2167 -622
rect -2147 -78 -1448 -50
rect -2147 -622 -1532 -78
rect -1468 -622 -1448 -78
rect -2147 -650 -1448 -622
rect -1428 -78 -729 -50
rect -1428 -622 -813 -78
rect -749 -622 -729 -78
rect -1428 -650 -729 -622
rect -709 -78 -10 -50
rect -709 -622 -94 -78
rect -30 -622 -10 -78
rect -709 -650 -10 -622
rect 10 -78 709 -50
rect 10 -622 625 -78
rect 689 -622 709 -78
rect 10 -650 709 -622
rect 729 -78 1428 -50
rect 729 -622 1344 -78
rect 1408 -622 1428 -78
rect 729 -650 1428 -622
rect 1448 -78 2147 -50
rect 1448 -622 2063 -78
rect 2127 -622 2147 -78
rect 1448 -650 2147 -622
rect 2167 -78 2866 -50
rect 2167 -622 2782 -78
rect 2846 -622 2866 -78
rect 2167 -650 2866 -622
rect 2886 -78 3585 -50
rect 2886 -622 3501 -78
rect 3565 -622 3585 -78
rect 2886 -650 3585 -622
rect -3585 -778 -2886 -750
rect -3585 -1322 -2970 -778
rect -2906 -1322 -2886 -778
rect -3585 -1350 -2886 -1322
rect -2866 -778 -2167 -750
rect -2866 -1322 -2251 -778
rect -2187 -1322 -2167 -778
rect -2866 -1350 -2167 -1322
rect -2147 -778 -1448 -750
rect -2147 -1322 -1532 -778
rect -1468 -1322 -1448 -778
rect -2147 -1350 -1448 -1322
rect -1428 -778 -729 -750
rect -1428 -1322 -813 -778
rect -749 -1322 -729 -778
rect -1428 -1350 -729 -1322
rect -709 -778 -10 -750
rect -709 -1322 -94 -778
rect -30 -1322 -10 -778
rect -709 -1350 -10 -1322
rect 10 -778 709 -750
rect 10 -1322 625 -778
rect 689 -1322 709 -778
rect 10 -1350 709 -1322
rect 729 -778 1428 -750
rect 729 -1322 1344 -778
rect 1408 -1322 1428 -778
rect 729 -1350 1428 -1322
rect 1448 -778 2147 -750
rect 1448 -1322 2063 -778
rect 2127 -1322 2147 -778
rect 1448 -1350 2147 -1322
rect 2167 -778 2866 -750
rect 2167 -1322 2782 -778
rect 2846 -1322 2866 -778
rect 2167 -1350 2866 -1322
rect 2886 -778 3585 -750
rect 2886 -1322 3501 -778
rect 3565 -1322 3585 -778
rect 2886 -1350 3585 -1322
rect -3585 -1478 -2886 -1450
rect -3585 -2022 -2970 -1478
rect -2906 -2022 -2886 -1478
rect -3585 -2050 -2886 -2022
rect -2866 -1478 -2167 -1450
rect -2866 -2022 -2251 -1478
rect -2187 -2022 -2167 -1478
rect -2866 -2050 -2167 -2022
rect -2147 -1478 -1448 -1450
rect -2147 -2022 -1532 -1478
rect -1468 -2022 -1448 -1478
rect -2147 -2050 -1448 -2022
rect -1428 -1478 -729 -1450
rect -1428 -2022 -813 -1478
rect -749 -2022 -729 -1478
rect -1428 -2050 -729 -2022
rect -709 -1478 -10 -1450
rect -709 -2022 -94 -1478
rect -30 -2022 -10 -1478
rect -709 -2050 -10 -2022
rect 10 -1478 709 -1450
rect 10 -2022 625 -1478
rect 689 -2022 709 -1478
rect 10 -2050 709 -2022
rect 729 -1478 1428 -1450
rect 729 -2022 1344 -1478
rect 1408 -2022 1428 -1478
rect 729 -2050 1428 -2022
rect 1448 -1478 2147 -1450
rect 1448 -2022 2063 -1478
rect 2127 -2022 2147 -1478
rect 1448 -2050 2147 -2022
rect 2167 -1478 2866 -1450
rect 2167 -2022 2782 -1478
rect 2846 -2022 2866 -1478
rect 2167 -2050 2866 -2022
rect 2886 -1478 3585 -1450
rect 2886 -2022 3501 -1478
rect 3565 -2022 3585 -1478
rect 2886 -2050 3585 -2022
rect -3585 -2178 -2886 -2150
rect -3585 -2722 -2970 -2178
rect -2906 -2722 -2886 -2178
rect -3585 -2750 -2886 -2722
rect -2866 -2178 -2167 -2150
rect -2866 -2722 -2251 -2178
rect -2187 -2722 -2167 -2178
rect -2866 -2750 -2167 -2722
rect -2147 -2178 -1448 -2150
rect -2147 -2722 -1532 -2178
rect -1468 -2722 -1448 -2178
rect -2147 -2750 -1448 -2722
rect -1428 -2178 -729 -2150
rect -1428 -2722 -813 -2178
rect -749 -2722 -729 -2178
rect -1428 -2750 -729 -2722
rect -709 -2178 -10 -2150
rect -709 -2722 -94 -2178
rect -30 -2722 -10 -2178
rect -709 -2750 -10 -2722
rect 10 -2178 709 -2150
rect 10 -2722 625 -2178
rect 689 -2722 709 -2178
rect 10 -2750 709 -2722
rect 729 -2178 1428 -2150
rect 729 -2722 1344 -2178
rect 1408 -2722 1428 -2178
rect 729 -2750 1428 -2722
rect 1448 -2178 2147 -2150
rect 1448 -2722 2063 -2178
rect 2127 -2722 2147 -2178
rect 1448 -2750 2147 -2722
rect 2167 -2178 2866 -2150
rect 2167 -2722 2782 -2178
rect 2846 -2722 2866 -2178
rect 2167 -2750 2866 -2722
rect 2886 -2178 3585 -2150
rect 2886 -2722 3501 -2178
rect 3565 -2722 3585 -2178
rect 2886 -2750 3585 -2722
rect -3585 -2878 -2886 -2850
rect -3585 -3422 -2970 -2878
rect -2906 -3422 -2886 -2878
rect -3585 -3450 -2886 -3422
rect -2866 -2878 -2167 -2850
rect -2866 -3422 -2251 -2878
rect -2187 -3422 -2167 -2878
rect -2866 -3450 -2167 -3422
rect -2147 -2878 -1448 -2850
rect -2147 -3422 -1532 -2878
rect -1468 -3422 -1448 -2878
rect -2147 -3450 -1448 -3422
rect -1428 -2878 -729 -2850
rect -1428 -3422 -813 -2878
rect -749 -3422 -729 -2878
rect -1428 -3450 -729 -3422
rect -709 -2878 -10 -2850
rect -709 -3422 -94 -2878
rect -30 -3422 -10 -2878
rect -709 -3450 -10 -3422
rect 10 -2878 709 -2850
rect 10 -3422 625 -2878
rect 689 -3422 709 -2878
rect 10 -3450 709 -3422
rect 729 -2878 1428 -2850
rect 729 -3422 1344 -2878
rect 1408 -3422 1428 -2878
rect 729 -3450 1428 -3422
rect 1448 -2878 2147 -2850
rect 1448 -3422 2063 -2878
rect 2127 -3422 2147 -2878
rect 1448 -3450 2147 -3422
rect 2167 -2878 2866 -2850
rect 2167 -3422 2782 -2878
rect 2846 -3422 2866 -2878
rect 2167 -3450 2866 -3422
rect 2886 -2878 3585 -2850
rect 2886 -3422 3501 -2878
rect 3565 -3422 3585 -2878
rect 2886 -3450 3585 -3422
<< via3 >>
rect -2970 2878 -2906 3422
rect -2251 2878 -2187 3422
rect -1532 2878 -1468 3422
rect -813 2878 -749 3422
rect -94 2878 -30 3422
rect 625 2878 689 3422
rect 1344 2878 1408 3422
rect 2063 2878 2127 3422
rect 2782 2878 2846 3422
rect 3501 2878 3565 3422
rect -2970 2178 -2906 2722
rect -2251 2178 -2187 2722
rect -1532 2178 -1468 2722
rect -813 2178 -749 2722
rect -94 2178 -30 2722
rect 625 2178 689 2722
rect 1344 2178 1408 2722
rect 2063 2178 2127 2722
rect 2782 2178 2846 2722
rect 3501 2178 3565 2722
rect -2970 1478 -2906 2022
rect -2251 1478 -2187 2022
rect -1532 1478 -1468 2022
rect -813 1478 -749 2022
rect -94 1478 -30 2022
rect 625 1478 689 2022
rect 1344 1478 1408 2022
rect 2063 1478 2127 2022
rect 2782 1478 2846 2022
rect 3501 1478 3565 2022
rect -2970 778 -2906 1322
rect -2251 778 -2187 1322
rect -1532 778 -1468 1322
rect -813 778 -749 1322
rect -94 778 -30 1322
rect 625 778 689 1322
rect 1344 778 1408 1322
rect 2063 778 2127 1322
rect 2782 778 2846 1322
rect 3501 778 3565 1322
rect -2970 78 -2906 622
rect -2251 78 -2187 622
rect -1532 78 -1468 622
rect -813 78 -749 622
rect -94 78 -30 622
rect 625 78 689 622
rect 1344 78 1408 622
rect 2063 78 2127 622
rect 2782 78 2846 622
rect 3501 78 3565 622
rect -2970 -622 -2906 -78
rect -2251 -622 -2187 -78
rect -1532 -622 -1468 -78
rect -813 -622 -749 -78
rect -94 -622 -30 -78
rect 625 -622 689 -78
rect 1344 -622 1408 -78
rect 2063 -622 2127 -78
rect 2782 -622 2846 -78
rect 3501 -622 3565 -78
rect -2970 -1322 -2906 -778
rect -2251 -1322 -2187 -778
rect -1532 -1322 -1468 -778
rect -813 -1322 -749 -778
rect -94 -1322 -30 -778
rect 625 -1322 689 -778
rect 1344 -1322 1408 -778
rect 2063 -1322 2127 -778
rect 2782 -1322 2846 -778
rect 3501 -1322 3565 -778
rect -2970 -2022 -2906 -1478
rect -2251 -2022 -2187 -1478
rect -1532 -2022 -1468 -1478
rect -813 -2022 -749 -1478
rect -94 -2022 -30 -1478
rect 625 -2022 689 -1478
rect 1344 -2022 1408 -1478
rect 2063 -2022 2127 -1478
rect 2782 -2022 2846 -1478
rect 3501 -2022 3565 -1478
rect -2970 -2722 -2906 -2178
rect -2251 -2722 -2187 -2178
rect -1532 -2722 -1468 -2178
rect -813 -2722 -749 -2178
rect -94 -2722 -30 -2178
rect 625 -2722 689 -2178
rect 1344 -2722 1408 -2178
rect 2063 -2722 2127 -2178
rect 2782 -2722 2846 -2178
rect 3501 -2722 3565 -2178
rect -2970 -3422 -2906 -2878
rect -2251 -3422 -2187 -2878
rect -1532 -3422 -1468 -2878
rect -813 -3422 -749 -2878
rect -94 -3422 -30 -2878
rect 625 -3422 689 -2878
rect 1344 -3422 1408 -2878
rect 2063 -3422 2127 -2878
rect 2782 -3422 2846 -2878
rect 3501 -3422 3565 -2878
<< mimcap >>
rect -3485 3310 -3085 3350
rect -3485 2990 -3445 3310
rect -3125 2990 -3085 3310
rect -3485 2950 -3085 2990
rect -2766 3310 -2366 3350
rect -2766 2990 -2726 3310
rect -2406 2990 -2366 3310
rect -2766 2950 -2366 2990
rect -2047 3310 -1647 3350
rect -2047 2990 -2007 3310
rect -1687 2990 -1647 3310
rect -2047 2950 -1647 2990
rect -1328 3310 -928 3350
rect -1328 2990 -1288 3310
rect -968 2990 -928 3310
rect -1328 2950 -928 2990
rect -609 3310 -209 3350
rect -609 2990 -569 3310
rect -249 2990 -209 3310
rect -609 2950 -209 2990
rect 110 3310 510 3350
rect 110 2990 150 3310
rect 470 2990 510 3310
rect 110 2950 510 2990
rect 829 3310 1229 3350
rect 829 2990 869 3310
rect 1189 2990 1229 3310
rect 829 2950 1229 2990
rect 1548 3310 1948 3350
rect 1548 2990 1588 3310
rect 1908 2990 1948 3310
rect 1548 2950 1948 2990
rect 2267 3310 2667 3350
rect 2267 2990 2307 3310
rect 2627 2990 2667 3310
rect 2267 2950 2667 2990
rect 2986 3310 3386 3350
rect 2986 2990 3026 3310
rect 3346 2990 3386 3310
rect 2986 2950 3386 2990
rect -3485 2610 -3085 2650
rect -3485 2290 -3445 2610
rect -3125 2290 -3085 2610
rect -3485 2250 -3085 2290
rect -2766 2610 -2366 2650
rect -2766 2290 -2726 2610
rect -2406 2290 -2366 2610
rect -2766 2250 -2366 2290
rect -2047 2610 -1647 2650
rect -2047 2290 -2007 2610
rect -1687 2290 -1647 2610
rect -2047 2250 -1647 2290
rect -1328 2610 -928 2650
rect -1328 2290 -1288 2610
rect -968 2290 -928 2610
rect -1328 2250 -928 2290
rect -609 2610 -209 2650
rect -609 2290 -569 2610
rect -249 2290 -209 2610
rect -609 2250 -209 2290
rect 110 2610 510 2650
rect 110 2290 150 2610
rect 470 2290 510 2610
rect 110 2250 510 2290
rect 829 2610 1229 2650
rect 829 2290 869 2610
rect 1189 2290 1229 2610
rect 829 2250 1229 2290
rect 1548 2610 1948 2650
rect 1548 2290 1588 2610
rect 1908 2290 1948 2610
rect 1548 2250 1948 2290
rect 2267 2610 2667 2650
rect 2267 2290 2307 2610
rect 2627 2290 2667 2610
rect 2267 2250 2667 2290
rect 2986 2610 3386 2650
rect 2986 2290 3026 2610
rect 3346 2290 3386 2610
rect 2986 2250 3386 2290
rect -3485 1910 -3085 1950
rect -3485 1590 -3445 1910
rect -3125 1590 -3085 1910
rect -3485 1550 -3085 1590
rect -2766 1910 -2366 1950
rect -2766 1590 -2726 1910
rect -2406 1590 -2366 1910
rect -2766 1550 -2366 1590
rect -2047 1910 -1647 1950
rect -2047 1590 -2007 1910
rect -1687 1590 -1647 1910
rect -2047 1550 -1647 1590
rect -1328 1910 -928 1950
rect -1328 1590 -1288 1910
rect -968 1590 -928 1910
rect -1328 1550 -928 1590
rect -609 1910 -209 1950
rect -609 1590 -569 1910
rect -249 1590 -209 1910
rect -609 1550 -209 1590
rect 110 1910 510 1950
rect 110 1590 150 1910
rect 470 1590 510 1910
rect 110 1550 510 1590
rect 829 1910 1229 1950
rect 829 1590 869 1910
rect 1189 1590 1229 1910
rect 829 1550 1229 1590
rect 1548 1910 1948 1950
rect 1548 1590 1588 1910
rect 1908 1590 1948 1910
rect 1548 1550 1948 1590
rect 2267 1910 2667 1950
rect 2267 1590 2307 1910
rect 2627 1590 2667 1910
rect 2267 1550 2667 1590
rect 2986 1910 3386 1950
rect 2986 1590 3026 1910
rect 3346 1590 3386 1910
rect 2986 1550 3386 1590
rect -3485 1210 -3085 1250
rect -3485 890 -3445 1210
rect -3125 890 -3085 1210
rect -3485 850 -3085 890
rect -2766 1210 -2366 1250
rect -2766 890 -2726 1210
rect -2406 890 -2366 1210
rect -2766 850 -2366 890
rect -2047 1210 -1647 1250
rect -2047 890 -2007 1210
rect -1687 890 -1647 1210
rect -2047 850 -1647 890
rect -1328 1210 -928 1250
rect -1328 890 -1288 1210
rect -968 890 -928 1210
rect -1328 850 -928 890
rect -609 1210 -209 1250
rect -609 890 -569 1210
rect -249 890 -209 1210
rect -609 850 -209 890
rect 110 1210 510 1250
rect 110 890 150 1210
rect 470 890 510 1210
rect 110 850 510 890
rect 829 1210 1229 1250
rect 829 890 869 1210
rect 1189 890 1229 1210
rect 829 850 1229 890
rect 1548 1210 1948 1250
rect 1548 890 1588 1210
rect 1908 890 1948 1210
rect 1548 850 1948 890
rect 2267 1210 2667 1250
rect 2267 890 2307 1210
rect 2627 890 2667 1210
rect 2267 850 2667 890
rect 2986 1210 3386 1250
rect 2986 890 3026 1210
rect 3346 890 3386 1210
rect 2986 850 3386 890
rect -3485 510 -3085 550
rect -3485 190 -3445 510
rect -3125 190 -3085 510
rect -3485 150 -3085 190
rect -2766 510 -2366 550
rect -2766 190 -2726 510
rect -2406 190 -2366 510
rect -2766 150 -2366 190
rect -2047 510 -1647 550
rect -2047 190 -2007 510
rect -1687 190 -1647 510
rect -2047 150 -1647 190
rect -1328 510 -928 550
rect -1328 190 -1288 510
rect -968 190 -928 510
rect -1328 150 -928 190
rect -609 510 -209 550
rect -609 190 -569 510
rect -249 190 -209 510
rect -609 150 -209 190
rect 110 510 510 550
rect 110 190 150 510
rect 470 190 510 510
rect 110 150 510 190
rect 829 510 1229 550
rect 829 190 869 510
rect 1189 190 1229 510
rect 829 150 1229 190
rect 1548 510 1948 550
rect 1548 190 1588 510
rect 1908 190 1948 510
rect 1548 150 1948 190
rect 2267 510 2667 550
rect 2267 190 2307 510
rect 2627 190 2667 510
rect 2267 150 2667 190
rect 2986 510 3386 550
rect 2986 190 3026 510
rect 3346 190 3386 510
rect 2986 150 3386 190
rect -3485 -190 -3085 -150
rect -3485 -510 -3445 -190
rect -3125 -510 -3085 -190
rect -3485 -550 -3085 -510
rect -2766 -190 -2366 -150
rect -2766 -510 -2726 -190
rect -2406 -510 -2366 -190
rect -2766 -550 -2366 -510
rect -2047 -190 -1647 -150
rect -2047 -510 -2007 -190
rect -1687 -510 -1647 -190
rect -2047 -550 -1647 -510
rect -1328 -190 -928 -150
rect -1328 -510 -1288 -190
rect -968 -510 -928 -190
rect -1328 -550 -928 -510
rect -609 -190 -209 -150
rect -609 -510 -569 -190
rect -249 -510 -209 -190
rect -609 -550 -209 -510
rect 110 -190 510 -150
rect 110 -510 150 -190
rect 470 -510 510 -190
rect 110 -550 510 -510
rect 829 -190 1229 -150
rect 829 -510 869 -190
rect 1189 -510 1229 -190
rect 829 -550 1229 -510
rect 1548 -190 1948 -150
rect 1548 -510 1588 -190
rect 1908 -510 1948 -190
rect 1548 -550 1948 -510
rect 2267 -190 2667 -150
rect 2267 -510 2307 -190
rect 2627 -510 2667 -190
rect 2267 -550 2667 -510
rect 2986 -190 3386 -150
rect 2986 -510 3026 -190
rect 3346 -510 3386 -190
rect 2986 -550 3386 -510
rect -3485 -890 -3085 -850
rect -3485 -1210 -3445 -890
rect -3125 -1210 -3085 -890
rect -3485 -1250 -3085 -1210
rect -2766 -890 -2366 -850
rect -2766 -1210 -2726 -890
rect -2406 -1210 -2366 -890
rect -2766 -1250 -2366 -1210
rect -2047 -890 -1647 -850
rect -2047 -1210 -2007 -890
rect -1687 -1210 -1647 -890
rect -2047 -1250 -1647 -1210
rect -1328 -890 -928 -850
rect -1328 -1210 -1288 -890
rect -968 -1210 -928 -890
rect -1328 -1250 -928 -1210
rect -609 -890 -209 -850
rect -609 -1210 -569 -890
rect -249 -1210 -209 -890
rect -609 -1250 -209 -1210
rect 110 -890 510 -850
rect 110 -1210 150 -890
rect 470 -1210 510 -890
rect 110 -1250 510 -1210
rect 829 -890 1229 -850
rect 829 -1210 869 -890
rect 1189 -1210 1229 -890
rect 829 -1250 1229 -1210
rect 1548 -890 1948 -850
rect 1548 -1210 1588 -890
rect 1908 -1210 1948 -890
rect 1548 -1250 1948 -1210
rect 2267 -890 2667 -850
rect 2267 -1210 2307 -890
rect 2627 -1210 2667 -890
rect 2267 -1250 2667 -1210
rect 2986 -890 3386 -850
rect 2986 -1210 3026 -890
rect 3346 -1210 3386 -890
rect 2986 -1250 3386 -1210
rect -3485 -1590 -3085 -1550
rect -3485 -1910 -3445 -1590
rect -3125 -1910 -3085 -1590
rect -3485 -1950 -3085 -1910
rect -2766 -1590 -2366 -1550
rect -2766 -1910 -2726 -1590
rect -2406 -1910 -2366 -1590
rect -2766 -1950 -2366 -1910
rect -2047 -1590 -1647 -1550
rect -2047 -1910 -2007 -1590
rect -1687 -1910 -1647 -1590
rect -2047 -1950 -1647 -1910
rect -1328 -1590 -928 -1550
rect -1328 -1910 -1288 -1590
rect -968 -1910 -928 -1590
rect -1328 -1950 -928 -1910
rect -609 -1590 -209 -1550
rect -609 -1910 -569 -1590
rect -249 -1910 -209 -1590
rect -609 -1950 -209 -1910
rect 110 -1590 510 -1550
rect 110 -1910 150 -1590
rect 470 -1910 510 -1590
rect 110 -1950 510 -1910
rect 829 -1590 1229 -1550
rect 829 -1910 869 -1590
rect 1189 -1910 1229 -1590
rect 829 -1950 1229 -1910
rect 1548 -1590 1948 -1550
rect 1548 -1910 1588 -1590
rect 1908 -1910 1948 -1590
rect 1548 -1950 1948 -1910
rect 2267 -1590 2667 -1550
rect 2267 -1910 2307 -1590
rect 2627 -1910 2667 -1590
rect 2267 -1950 2667 -1910
rect 2986 -1590 3386 -1550
rect 2986 -1910 3026 -1590
rect 3346 -1910 3386 -1590
rect 2986 -1950 3386 -1910
rect -3485 -2290 -3085 -2250
rect -3485 -2610 -3445 -2290
rect -3125 -2610 -3085 -2290
rect -3485 -2650 -3085 -2610
rect -2766 -2290 -2366 -2250
rect -2766 -2610 -2726 -2290
rect -2406 -2610 -2366 -2290
rect -2766 -2650 -2366 -2610
rect -2047 -2290 -1647 -2250
rect -2047 -2610 -2007 -2290
rect -1687 -2610 -1647 -2290
rect -2047 -2650 -1647 -2610
rect -1328 -2290 -928 -2250
rect -1328 -2610 -1288 -2290
rect -968 -2610 -928 -2290
rect -1328 -2650 -928 -2610
rect -609 -2290 -209 -2250
rect -609 -2610 -569 -2290
rect -249 -2610 -209 -2290
rect -609 -2650 -209 -2610
rect 110 -2290 510 -2250
rect 110 -2610 150 -2290
rect 470 -2610 510 -2290
rect 110 -2650 510 -2610
rect 829 -2290 1229 -2250
rect 829 -2610 869 -2290
rect 1189 -2610 1229 -2290
rect 829 -2650 1229 -2610
rect 1548 -2290 1948 -2250
rect 1548 -2610 1588 -2290
rect 1908 -2610 1948 -2290
rect 1548 -2650 1948 -2610
rect 2267 -2290 2667 -2250
rect 2267 -2610 2307 -2290
rect 2627 -2610 2667 -2290
rect 2267 -2650 2667 -2610
rect 2986 -2290 3386 -2250
rect 2986 -2610 3026 -2290
rect 3346 -2610 3386 -2290
rect 2986 -2650 3386 -2610
rect -3485 -2990 -3085 -2950
rect -3485 -3310 -3445 -2990
rect -3125 -3310 -3085 -2990
rect -3485 -3350 -3085 -3310
rect -2766 -2990 -2366 -2950
rect -2766 -3310 -2726 -2990
rect -2406 -3310 -2366 -2990
rect -2766 -3350 -2366 -3310
rect -2047 -2990 -1647 -2950
rect -2047 -3310 -2007 -2990
rect -1687 -3310 -1647 -2990
rect -2047 -3350 -1647 -3310
rect -1328 -2990 -928 -2950
rect -1328 -3310 -1288 -2990
rect -968 -3310 -928 -2990
rect -1328 -3350 -928 -3310
rect -609 -2990 -209 -2950
rect -609 -3310 -569 -2990
rect -249 -3310 -209 -2990
rect -609 -3350 -209 -3310
rect 110 -2990 510 -2950
rect 110 -3310 150 -2990
rect 470 -3310 510 -2990
rect 110 -3350 510 -3310
rect 829 -2990 1229 -2950
rect 829 -3310 869 -2990
rect 1189 -3310 1229 -2990
rect 829 -3350 1229 -3310
rect 1548 -2990 1948 -2950
rect 1548 -3310 1588 -2990
rect 1908 -3310 1948 -2990
rect 1548 -3350 1948 -3310
rect 2267 -2990 2667 -2950
rect 2267 -3310 2307 -2990
rect 2627 -3310 2667 -2990
rect 2267 -3350 2667 -3310
rect 2986 -2990 3386 -2950
rect 2986 -3310 3026 -2990
rect 3346 -3310 3386 -2990
rect 2986 -3350 3386 -3310
<< mimcapcontact >>
rect -3445 2990 -3125 3310
rect -2726 2990 -2406 3310
rect -2007 2990 -1687 3310
rect -1288 2990 -968 3310
rect -569 2990 -249 3310
rect 150 2990 470 3310
rect 869 2990 1189 3310
rect 1588 2990 1908 3310
rect 2307 2990 2627 3310
rect 3026 2990 3346 3310
rect -3445 2290 -3125 2610
rect -2726 2290 -2406 2610
rect -2007 2290 -1687 2610
rect -1288 2290 -968 2610
rect -569 2290 -249 2610
rect 150 2290 470 2610
rect 869 2290 1189 2610
rect 1588 2290 1908 2610
rect 2307 2290 2627 2610
rect 3026 2290 3346 2610
rect -3445 1590 -3125 1910
rect -2726 1590 -2406 1910
rect -2007 1590 -1687 1910
rect -1288 1590 -968 1910
rect -569 1590 -249 1910
rect 150 1590 470 1910
rect 869 1590 1189 1910
rect 1588 1590 1908 1910
rect 2307 1590 2627 1910
rect 3026 1590 3346 1910
rect -3445 890 -3125 1210
rect -2726 890 -2406 1210
rect -2007 890 -1687 1210
rect -1288 890 -968 1210
rect -569 890 -249 1210
rect 150 890 470 1210
rect 869 890 1189 1210
rect 1588 890 1908 1210
rect 2307 890 2627 1210
rect 3026 890 3346 1210
rect -3445 190 -3125 510
rect -2726 190 -2406 510
rect -2007 190 -1687 510
rect -1288 190 -968 510
rect -569 190 -249 510
rect 150 190 470 510
rect 869 190 1189 510
rect 1588 190 1908 510
rect 2307 190 2627 510
rect 3026 190 3346 510
rect -3445 -510 -3125 -190
rect -2726 -510 -2406 -190
rect -2007 -510 -1687 -190
rect -1288 -510 -968 -190
rect -569 -510 -249 -190
rect 150 -510 470 -190
rect 869 -510 1189 -190
rect 1588 -510 1908 -190
rect 2307 -510 2627 -190
rect 3026 -510 3346 -190
rect -3445 -1210 -3125 -890
rect -2726 -1210 -2406 -890
rect -2007 -1210 -1687 -890
rect -1288 -1210 -968 -890
rect -569 -1210 -249 -890
rect 150 -1210 470 -890
rect 869 -1210 1189 -890
rect 1588 -1210 1908 -890
rect 2307 -1210 2627 -890
rect 3026 -1210 3346 -890
rect -3445 -1910 -3125 -1590
rect -2726 -1910 -2406 -1590
rect -2007 -1910 -1687 -1590
rect -1288 -1910 -968 -1590
rect -569 -1910 -249 -1590
rect 150 -1910 470 -1590
rect 869 -1910 1189 -1590
rect 1588 -1910 1908 -1590
rect 2307 -1910 2627 -1590
rect 3026 -1910 3346 -1590
rect -3445 -2610 -3125 -2290
rect -2726 -2610 -2406 -2290
rect -2007 -2610 -1687 -2290
rect -1288 -2610 -968 -2290
rect -569 -2610 -249 -2290
rect 150 -2610 470 -2290
rect 869 -2610 1189 -2290
rect 1588 -2610 1908 -2290
rect 2307 -2610 2627 -2290
rect 3026 -2610 3346 -2290
rect -3445 -3310 -3125 -2990
rect -2726 -3310 -2406 -2990
rect -2007 -3310 -1687 -2990
rect -1288 -3310 -968 -2990
rect -569 -3310 -249 -2990
rect 150 -3310 470 -2990
rect 869 -3310 1189 -2990
rect 1588 -3310 1908 -2990
rect 2307 -3310 2627 -2990
rect 3026 -3310 3346 -2990
<< metal4 >>
rect -3337 3311 -3233 3500
rect -3017 3438 -2913 3500
rect -3017 3422 -2890 3438
rect -3446 3310 -3124 3311
rect -3446 2990 -3445 3310
rect -3125 2990 -3124 3310
rect -3446 2989 -3124 2990
rect -3337 2611 -3233 2989
rect -3017 2878 -2970 3422
rect -2906 2878 -2890 3422
rect -2618 3311 -2514 3500
rect -2298 3438 -2194 3500
rect -2298 3422 -2171 3438
rect -2727 3310 -2405 3311
rect -2727 2990 -2726 3310
rect -2406 2990 -2405 3310
rect -2727 2989 -2405 2990
rect -3017 2862 -2890 2878
rect -3017 2738 -2913 2862
rect -3017 2722 -2890 2738
rect -3446 2610 -3124 2611
rect -3446 2290 -3445 2610
rect -3125 2290 -3124 2610
rect -3446 2289 -3124 2290
rect -3337 1911 -3233 2289
rect -3017 2178 -2970 2722
rect -2906 2178 -2890 2722
rect -2618 2611 -2514 2989
rect -2298 2878 -2251 3422
rect -2187 2878 -2171 3422
rect -1899 3311 -1795 3500
rect -1579 3438 -1475 3500
rect -1579 3422 -1452 3438
rect -2008 3310 -1686 3311
rect -2008 2990 -2007 3310
rect -1687 2990 -1686 3310
rect -2008 2989 -1686 2990
rect -2298 2862 -2171 2878
rect -2298 2738 -2194 2862
rect -2298 2722 -2171 2738
rect -2727 2610 -2405 2611
rect -2727 2290 -2726 2610
rect -2406 2290 -2405 2610
rect -2727 2289 -2405 2290
rect -3017 2162 -2890 2178
rect -3017 2038 -2913 2162
rect -3017 2022 -2890 2038
rect -3446 1910 -3124 1911
rect -3446 1590 -3445 1910
rect -3125 1590 -3124 1910
rect -3446 1589 -3124 1590
rect -3337 1211 -3233 1589
rect -3017 1478 -2970 2022
rect -2906 1478 -2890 2022
rect -2618 1911 -2514 2289
rect -2298 2178 -2251 2722
rect -2187 2178 -2171 2722
rect -1899 2611 -1795 2989
rect -1579 2878 -1532 3422
rect -1468 2878 -1452 3422
rect -1180 3311 -1076 3500
rect -860 3438 -756 3500
rect -860 3422 -733 3438
rect -1289 3310 -967 3311
rect -1289 2990 -1288 3310
rect -968 2990 -967 3310
rect -1289 2989 -967 2990
rect -1579 2862 -1452 2878
rect -1579 2738 -1475 2862
rect -1579 2722 -1452 2738
rect -2008 2610 -1686 2611
rect -2008 2290 -2007 2610
rect -1687 2290 -1686 2610
rect -2008 2289 -1686 2290
rect -2298 2162 -2171 2178
rect -2298 2038 -2194 2162
rect -2298 2022 -2171 2038
rect -2727 1910 -2405 1911
rect -2727 1590 -2726 1910
rect -2406 1590 -2405 1910
rect -2727 1589 -2405 1590
rect -3017 1462 -2890 1478
rect -3017 1338 -2913 1462
rect -3017 1322 -2890 1338
rect -3446 1210 -3124 1211
rect -3446 890 -3445 1210
rect -3125 890 -3124 1210
rect -3446 889 -3124 890
rect -3337 511 -3233 889
rect -3017 778 -2970 1322
rect -2906 778 -2890 1322
rect -2618 1211 -2514 1589
rect -2298 1478 -2251 2022
rect -2187 1478 -2171 2022
rect -1899 1911 -1795 2289
rect -1579 2178 -1532 2722
rect -1468 2178 -1452 2722
rect -1180 2611 -1076 2989
rect -860 2878 -813 3422
rect -749 2878 -733 3422
rect -461 3311 -357 3500
rect -141 3438 -37 3500
rect -141 3422 -14 3438
rect -570 3310 -248 3311
rect -570 2990 -569 3310
rect -249 2990 -248 3310
rect -570 2989 -248 2990
rect -860 2862 -733 2878
rect -860 2738 -756 2862
rect -860 2722 -733 2738
rect -1289 2610 -967 2611
rect -1289 2290 -1288 2610
rect -968 2290 -967 2610
rect -1289 2289 -967 2290
rect -1579 2162 -1452 2178
rect -1579 2038 -1475 2162
rect -1579 2022 -1452 2038
rect -2008 1910 -1686 1911
rect -2008 1590 -2007 1910
rect -1687 1590 -1686 1910
rect -2008 1589 -1686 1590
rect -2298 1462 -2171 1478
rect -2298 1338 -2194 1462
rect -2298 1322 -2171 1338
rect -2727 1210 -2405 1211
rect -2727 890 -2726 1210
rect -2406 890 -2405 1210
rect -2727 889 -2405 890
rect -3017 762 -2890 778
rect -3017 638 -2913 762
rect -3017 622 -2890 638
rect -3446 510 -3124 511
rect -3446 190 -3445 510
rect -3125 190 -3124 510
rect -3446 189 -3124 190
rect -3337 -189 -3233 189
rect -3017 78 -2970 622
rect -2906 78 -2890 622
rect -2618 511 -2514 889
rect -2298 778 -2251 1322
rect -2187 778 -2171 1322
rect -1899 1211 -1795 1589
rect -1579 1478 -1532 2022
rect -1468 1478 -1452 2022
rect -1180 1911 -1076 2289
rect -860 2178 -813 2722
rect -749 2178 -733 2722
rect -461 2611 -357 2989
rect -141 2878 -94 3422
rect -30 2878 -14 3422
rect 258 3311 362 3500
rect 578 3438 682 3500
rect 578 3422 705 3438
rect 149 3310 471 3311
rect 149 2990 150 3310
rect 470 2990 471 3310
rect 149 2989 471 2990
rect -141 2862 -14 2878
rect -141 2738 -37 2862
rect -141 2722 -14 2738
rect -570 2610 -248 2611
rect -570 2290 -569 2610
rect -249 2290 -248 2610
rect -570 2289 -248 2290
rect -860 2162 -733 2178
rect -860 2038 -756 2162
rect -860 2022 -733 2038
rect -1289 1910 -967 1911
rect -1289 1590 -1288 1910
rect -968 1590 -967 1910
rect -1289 1589 -967 1590
rect -1579 1462 -1452 1478
rect -1579 1338 -1475 1462
rect -1579 1322 -1452 1338
rect -2008 1210 -1686 1211
rect -2008 890 -2007 1210
rect -1687 890 -1686 1210
rect -2008 889 -1686 890
rect -2298 762 -2171 778
rect -2298 638 -2194 762
rect -2298 622 -2171 638
rect -2727 510 -2405 511
rect -2727 190 -2726 510
rect -2406 190 -2405 510
rect -2727 189 -2405 190
rect -3017 62 -2890 78
rect -3017 -62 -2913 62
rect -3017 -78 -2890 -62
rect -3446 -190 -3124 -189
rect -3446 -510 -3445 -190
rect -3125 -510 -3124 -190
rect -3446 -511 -3124 -510
rect -3337 -889 -3233 -511
rect -3017 -622 -2970 -78
rect -2906 -622 -2890 -78
rect -2618 -189 -2514 189
rect -2298 78 -2251 622
rect -2187 78 -2171 622
rect -1899 511 -1795 889
rect -1579 778 -1532 1322
rect -1468 778 -1452 1322
rect -1180 1211 -1076 1589
rect -860 1478 -813 2022
rect -749 1478 -733 2022
rect -461 1911 -357 2289
rect -141 2178 -94 2722
rect -30 2178 -14 2722
rect 258 2611 362 2989
rect 578 2878 625 3422
rect 689 2878 705 3422
rect 977 3311 1081 3500
rect 1297 3438 1401 3500
rect 1297 3422 1424 3438
rect 868 3310 1190 3311
rect 868 2990 869 3310
rect 1189 2990 1190 3310
rect 868 2989 1190 2990
rect 578 2862 705 2878
rect 578 2738 682 2862
rect 578 2722 705 2738
rect 149 2610 471 2611
rect 149 2290 150 2610
rect 470 2290 471 2610
rect 149 2289 471 2290
rect -141 2162 -14 2178
rect -141 2038 -37 2162
rect -141 2022 -14 2038
rect -570 1910 -248 1911
rect -570 1590 -569 1910
rect -249 1590 -248 1910
rect -570 1589 -248 1590
rect -860 1462 -733 1478
rect -860 1338 -756 1462
rect -860 1322 -733 1338
rect -1289 1210 -967 1211
rect -1289 890 -1288 1210
rect -968 890 -967 1210
rect -1289 889 -967 890
rect -1579 762 -1452 778
rect -1579 638 -1475 762
rect -1579 622 -1452 638
rect -2008 510 -1686 511
rect -2008 190 -2007 510
rect -1687 190 -1686 510
rect -2008 189 -1686 190
rect -2298 62 -2171 78
rect -2298 -62 -2194 62
rect -2298 -78 -2171 -62
rect -2727 -190 -2405 -189
rect -2727 -510 -2726 -190
rect -2406 -510 -2405 -190
rect -2727 -511 -2405 -510
rect -3017 -638 -2890 -622
rect -3017 -762 -2913 -638
rect -3017 -778 -2890 -762
rect -3446 -890 -3124 -889
rect -3446 -1210 -3445 -890
rect -3125 -1210 -3124 -890
rect -3446 -1211 -3124 -1210
rect -3337 -1589 -3233 -1211
rect -3017 -1322 -2970 -778
rect -2906 -1322 -2890 -778
rect -2618 -889 -2514 -511
rect -2298 -622 -2251 -78
rect -2187 -622 -2171 -78
rect -1899 -189 -1795 189
rect -1579 78 -1532 622
rect -1468 78 -1452 622
rect -1180 511 -1076 889
rect -860 778 -813 1322
rect -749 778 -733 1322
rect -461 1211 -357 1589
rect -141 1478 -94 2022
rect -30 1478 -14 2022
rect 258 1911 362 2289
rect 578 2178 625 2722
rect 689 2178 705 2722
rect 977 2611 1081 2989
rect 1297 2878 1344 3422
rect 1408 2878 1424 3422
rect 1696 3311 1800 3500
rect 2016 3438 2120 3500
rect 2016 3422 2143 3438
rect 1587 3310 1909 3311
rect 1587 2990 1588 3310
rect 1908 2990 1909 3310
rect 1587 2989 1909 2990
rect 1297 2862 1424 2878
rect 1297 2738 1401 2862
rect 1297 2722 1424 2738
rect 868 2610 1190 2611
rect 868 2290 869 2610
rect 1189 2290 1190 2610
rect 868 2289 1190 2290
rect 578 2162 705 2178
rect 578 2038 682 2162
rect 578 2022 705 2038
rect 149 1910 471 1911
rect 149 1590 150 1910
rect 470 1590 471 1910
rect 149 1589 471 1590
rect -141 1462 -14 1478
rect -141 1338 -37 1462
rect -141 1322 -14 1338
rect -570 1210 -248 1211
rect -570 890 -569 1210
rect -249 890 -248 1210
rect -570 889 -248 890
rect -860 762 -733 778
rect -860 638 -756 762
rect -860 622 -733 638
rect -1289 510 -967 511
rect -1289 190 -1288 510
rect -968 190 -967 510
rect -1289 189 -967 190
rect -1579 62 -1452 78
rect -1579 -62 -1475 62
rect -1579 -78 -1452 -62
rect -2008 -190 -1686 -189
rect -2008 -510 -2007 -190
rect -1687 -510 -1686 -190
rect -2008 -511 -1686 -510
rect -2298 -638 -2171 -622
rect -2298 -762 -2194 -638
rect -2298 -778 -2171 -762
rect -2727 -890 -2405 -889
rect -2727 -1210 -2726 -890
rect -2406 -1210 -2405 -890
rect -2727 -1211 -2405 -1210
rect -3017 -1338 -2890 -1322
rect -3017 -1462 -2913 -1338
rect -3017 -1478 -2890 -1462
rect -3446 -1590 -3124 -1589
rect -3446 -1910 -3445 -1590
rect -3125 -1910 -3124 -1590
rect -3446 -1911 -3124 -1910
rect -3337 -2289 -3233 -1911
rect -3017 -2022 -2970 -1478
rect -2906 -2022 -2890 -1478
rect -2618 -1589 -2514 -1211
rect -2298 -1322 -2251 -778
rect -2187 -1322 -2171 -778
rect -1899 -889 -1795 -511
rect -1579 -622 -1532 -78
rect -1468 -622 -1452 -78
rect -1180 -189 -1076 189
rect -860 78 -813 622
rect -749 78 -733 622
rect -461 511 -357 889
rect -141 778 -94 1322
rect -30 778 -14 1322
rect 258 1211 362 1589
rect 578 1478 625 2022
rect 689 1478 705 2022
rect 977 1911 1081 2289
rect 1297 2178 1344 2722
rect 1408 2178 1424 2722
rect 1696 2611 1800 2989
rect 2016 2878 2063 3422
rect 2127 2878 2143 3422
rect 2415 3311 2519 3500
rect 2735 3438 2839 3500
rect 2735 3422 2862 3438
rect 2306 3310 2628 3311
rect 2306 2990 2307 3310
rect 2627 2990 2628 3310
rect 2306 2989 2628 2990
rect 2016 2862 2143 2878
rect 2016 2738 2120 2862
rect 2016 2722 2143 2738
rect 1587 2610 1909 2611
rect 1587 2290 1588 2610
rect 1908 2290 1909 2610
rect 1587 2289 1909 2290
rect 1297 2162 1424 2178
rect 1297 2038 1401 2162
rect 1297 2022 1424 2038
rect 868 1910 1190 1911
rect 868 1590 869 1910
rect 1189 1590 1190 1910
rect 868 1589 1190 1590
rect 578 1462 705 1478
rect 578 1338 682 1462
rect 578 1322 705 1338
rect 149 1210 471 1211
rect 149 890 150 1210
rect 470 890 471 1210
rect 149 889 471 890
rect -141 762 -14 778
rect -141 638 -37 762
rect -141 622 -14 638
rect -570 510 -248 511
rect -570 190 -569 510
rect -249 190 -248 510
rect -570 189 -248 190
rect -860 62 -733 78
rect -860 -62 -756 62
rect -860 -78 -733 -62
rect -1289 -190 -967 -189
rect -1289 -510 -1288 -190
rect -968 -510 -967 -190
rect -1289 -511 -967 -510
rect -1579 -638 -1452 -622
rect -1579 -762 -1475 -638
rect -1579 -778 -1452 -762
rect -2008 -890 -1686 -889
rect -2008 -1210 -2007 -890
rect -1687 -1210 -1686 -890
rect -2008 -1211 -1686 -1210
rect -2298 -1338 -2171 -1322
rect -2298 -1462 -2194 -1338
rect -2298 -1478 -2171 -1462
rect -2727 -1590 -2405 -1589
rect -2727 -1910 -2726 -1590
rect -2406 -1910 -2405 -1590
rect -2727 -1911 -2405 -1910
rect -3017 -2038 -2890 -2022
rect -3017 -2162 -2913 -2038
rect -3017 -2178 -2890 -2162
rect -3446 -2290 -3124 -2289
rect -3446 -2610 -3445 -2290
rect -3125 -2610 -3124 -2290
rect -3446 -2611 -3124 -2610
rect -3337 -2989 -3233 -2611
rect -3017 -2722 -2970 -2178
rect -2906 -2722 -2890 -2178
rect -2618 -2289 -2514 -1911
rect -2298 -2022 -2251 -1478
rect -2187 -2022 -2171 -1478
rect -1899 -1589 -1795 -1211
rect -1579 -1322 -1532 -778
rect -1468 -1322 -1452 -778
rect -1180 -889 -1076 -511
rect -860 -622 -813 -78
rect -749 -622 -733 -78
rect -461 -189 -357 189
rect -141 78 -94 622
rect -30 78 -14 622
rect 258 511 362 889
rect 578 778 625 1322
rect 689 778 705 1322
rect 977 1211 1081 1589
rect 1297 1478 1344 2022
rect 1408 1478 1424 2022
rect 1696 1911 1800 2289
rect 2016 2178 2063 2722
rect 2127 2178 2143 2722
rect 2415 2611 2519 2989
rect 2735 2878 2782 3422
rect 2846 2878 2862 3422
rect 3134 3311 3238 3500
rect 3454 3438 3558 3500
rect 3454 3422 3581 3438
rect 3025 3310 3347 3311
rect 3025 2990 3026 3310
rect 3346 2990 3347 3310
rect 3025 2989 3347 2990
rect 2735 2862 2862 2878
rect 2735 2738 2839 2862
rect 2735 2722 2862 2738
rect 2306 2610 2628 2611
rect 2306 2290 2307 2610
rect 2627 2290 2628 2610
rect 2306 2289 2628 2290
rect 2016 2162 2143 2178
rect 2016 2038 2120 2162
rect 2016 2022 2143 2038
rect 1587 1910 1909 1911
rect 1587 1590 1588 1910
rect 1908 1590 1909 1910
rect 1587 1589 1909 1590
rect 1297 1462 1424 1478
rect 1297 1338 1401 1462
rect 1297 1322 1424 1338
rect 868 1210 1190 1211
rect 868 890 869 1210
rect 1189 890 1190 1210
rect 868 889 1190 890
rect 578 762 705 778
rect 578 638 682 762
rect 578 622 705 638
rect 149 510 471 511
rect 149 190 150 510
rect 470 190 471 510
rect 149 189 471 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -570 -190 -248 -189
rect -570 -510 -569 -190
rect -249 -510 -248 -190
rect -570 -511 -248 -510
rect -860 -638 -733 -622
rect -860 -762 -756 -638
rect -860 -778 -733 -762
rect -1289 -890 -967 -889
rect -1289 -1210 -1288 -890
rect -968 -1210 -967 -890
rect -1289 -1211 -967 -1210
rect -1579 -1338 -1452 -1322
rect -1579 -1462 -1475 -1338
rect -1579 -1478 -1452 -1462
rect -2008 -1590 -1686 -1589
rect -2008 -1910 -2007 -1590
rect -1687 -1910 -1686 -1590
rect -2008 -1911 -1686 -1910
rect -2298 -2038 -2171 -2022
rect -2298 -2162 -2194 -2038
rect -2298 -2178 -2171 -2162
rect -2727 -2290 -2405 -2289
rect -2727 -2610 -2726 -2290
rect -2406 -2610 -2405 -2290
rect -2727 -2611 -2405 -2610
rect -3017 -2738 -2890 -2722
rect -3017 -2862 -2913 -2738
rect -3017 -2878 -2890 -2862
rect -3446 -2990 -3124 -2989
rect -3446 -3310 -3445 -2990
rect -3125 -3310 -3124 -2990
rect -3446 -3311 -3124 -3310
rect -3337 -3500 -3233 -3311
rect -3017 -3422 -2970 -2878
rect -2906 -3422 -2890 -2878
rect -2618 -2989 -2514 -2611
rect -2298 -2722 -2251 -2178
rect -2187 -2722 -2171 -2178
rect -1899 -2289 -1795 -1911
rect -1579 -2022 -1532 -1478
rect -1468 -2022 -1452 -1478
rect -1180 -1589 -1076 -1211
rect -860 -1322 -813 -778
rect -749 -1322 -733 -778
rect -461 -889 -357 -511
rect -141 -622 -94 -78
rect -30 -622 -14 -78
rect 258 -189 362 189
rect 578 78 625 622
rect 689 78 705 622
rect 977 511 1081 889
rect 1297 778 1344 1322
rect 1408 778 1424 1322
rect 1696 1211 1800 1589
rect 2016 1478 2063 2022
rect 2127 1478 2143 2022
rect 2415 1911 2519 2289
rect 2735 2178 2782 2722
rect 2846 2178 2862 2722
rect 3134 2611 3238 2989
rect 3454 2878 3501 3422
rect 3565 2878 3581 3422
rect 3454 2862 3581 2878
rect 3454 2738 3558 2862
rect 3454 2722 3581 2738
rect 3025 2610 3347 2611
rect 3025 2290 3026 2610
rect 3346 2290 3347 2610
rect 3025 2289 3347 2290
rect 2735 2162 2862 2178
rect 2735 2038 2839 2162
rect 2735 2022 2862 2038
rect 2306 1910 2628 1911
rect 2306 1590 2307 1910
rect 2627 1590 2628 1910
rect 2306 1589 2628 1590
rect 2016 1462 2143 1478
rect 2016 1338 2120 1462
rect 2016 1322 2143 1338
rect 1587 1210 1909 1211
rect 1587 890 1588 1210
rect 1908 890 1909 1210
rect 1587 889 1909 890
rect 1297 762 1424 778
rect 1297 638 1401 762
rect 1297 622 1424 638
rect 868 510 1190 511
rect 868 190 869 510
rect 1189 190 1190 510
rect 868 189 1190 190
rect 578 62 705 78
rect 578 -62 682 62
rect 578 -78 705 -62
rect 149 -190 471 -189
rect 149 -510 150 -190
rect 470 -510 471 -190
rect 149 -511 471 -510
rect -141 -638 -14 -622
rect -141 -762 -37 -638
rect -141 -778 -14 -762
rect -570 -890 -248 -889
rect -570 -1210 -569 -890
rect -249 -1210 -248 -890
rect -570 -1211 -248 -1210
rect -860 -1338 -733 -1322
rect -860 -1462 -756 -1338
rect -860 -1478 -733 -1462
rect -1289 -1590 -967 -1589
rect -1289 -1910 -1288 -1590
rect -968 -1910 -967 -1590
rect -1289 -1911 -967 -1910
rect -1579 -2038 -1452 -2022
rect -1579 -2162 -1475 -2038
rect -1579 -2178 -1452 -2162
rect -2008 -2290 -1686 -2289
rect -2008 -2610 -2007 -2290
rect -1687 -2610 -1686 -2290
rect -2008 -2611 -1686 -2610
rect -2298 -2738 -2171 -2722
rect -2298 -2862 -2194 -2738
rect -2298 -2878 -2171 -2862
rect -2727 -2990 -2405 -2989
rect -2727 -3310 -2726 -2990
rect -2406 -3310 -2405 -2990
rect -2727 -3311 -2405 -3310
rect -3017 -3438 -2890 -3422
rect -3017 -3500 -2913 -3438
rect -2618 -3500 -2514 -3311
rect -2298 -3422 -2251 -2878
rect -2187 -3422 -2171 -2878
rect -1899 -2989 -1795 -2611
rect -1579 -2722 -1532 -2178
rect -1468 -2722 -1452 -2178
rect -1180 -2289 -1076 -1911
rect -860 -2022 -813 -1478
rect -749 -2022 -733 -1478
rect -461 -1589 -357 -1211
rect -141 -1322 -94 -778
rect -30 -1322 -14 -778
rect 258 -889 362 -511
rect 578 -622 625 -78
rect 689 -622 705 -78
rect 977 -189 1081 189
rect 1297 78 1344 622
rect 1408 78 1424 622
rect 1696 511 1800 889
rect 2016 778 2063 1322
rect 2127 778 2143 1322
rect 2415 1211 2519 1589
rect 2735 1478 2782 2022
rect 2846 1478 2862 2022
rect 3134 1911 3238 2289
rect 3454 2178 3501 2722
rect 3565 2178 3581 2722
rect 3454 2162 3581 2178
rect 3454 2038 3558 2162
rect 3454 2022 3581 2038
rect 3025 1910 3347 1911
rect 3025 1590 3026 1910
rect 3346 1590 3347 1910
rect 3025 1589 3347 1590
rect 2735 1462 2862 1478
rect 2735 1338 2839 1462
rect 2735 1322 2862 1338
rect 2306 1210 2628 1211
rect 2306 890 2307 1210
rect 2627 890 2628 1210
rect 2306 889 2628 890
rect 2016 762 2143 778
rect 2016 638 2120 762
rect 2016 622 2143 638
rect 1587 510 1909 511
rect 1587 190 1588 510
rect 1908 190 1909 510
rect 1587 189 1909 190
rect 1297 62 1424 78
rect 1297 -62 1401 62
rect 1297 -78 1424 -62
rect 868 -190 1190 -189
rect 868 -510 869 -190
rect 1189 -510 1190 -190
rect 868 -511 1190 -510
rect 578 -638 705 -622
rect 578 -762 682 -638
rect 578 -778 705 -762
rect 149 -890 471 -889
rect 149 -1210 150 -890
rect 470 -1210 471 -890
rect 149 -1211 471 -1210
rect -141 -1338 -14 -1322
rect -141 -1462 -37 -1338
rect -141 -1478 -14 -1462
rect -570 -1590 -248 -1589
rect -570 -1910 -569 -1590
rect -249 -1910 -248 -1590
rect -570 -1911 -248 -1910
rect -860 -2038 -733 -2022
rect -860 -2162 -756 -2038
rect -860 -2178 -733 -2162
rect -1289 -2290 -967 -2289
rect -1289 -2610 -1288 -2290
rect -968 -2610 -967 -2290
rect -1289 -2611 -967 -2610
rect -1579 -2738 -1452 -2722
rect -1579 -2862 -1475 -2738
rect -1579 -2878 -1452 -2862
rect -2008 -2990 -1686 -2989
rect -2008 -3310 -2007 -2990
rect -1687 -3310 -1686 -2990
rect -2008 -3311 -1686 -3310
rect -2298 -3438 -2171 -3422
rect -2298 -3500 -2194 -3438
rect -1899 -3500 -1795 -3311
rect -1579 -3422 -1532 -2878
rect -1468 -3422 -1452 -2878
rect -1180 -2989 -1076 -2611
rect -860 -2722 -813 -2178
rect -749 -2722 -733 -2178
rect -461 -2289 -357 -1911
rect -141 -2022 -94 -1478
rect -30 -2022 -14 -1478
rect 258 -1589 362 -1211
rect 578 -1322 625 -778
rect 689 -1322 705 -778
rect 977 -889 1081 -511
rect 1297 -622 1344 -78
rect 1408 -622 1424 -78
rect 1696 -189 1800 189
rect 2016 78 2063 622
rect 2127 78 2143 622
rect 2415 511 2519 889
rect 2735 778 2782 1322
rect 2846 778 2862 1322
rect 3134 1211 3238 1589
rect 3454 1478 3501 2022
rect 3565 1478 3581 2022
rect 3454 1462 3581 1478
rect 3454 1338 3558 1462
rect 3454 1322 3581 1338
rect 3025 1210 3347 1211
rect 3025 890 3026 1210
rect 3346 890 3347 1210
rect 3025 889 3347 890
rect 2735 762 2862 778
rect 2735 638 2839 762
rect 2735 622 2862 638
rect 2306 510 2628 511
rect 2306 190 2307 510
rect 2627 190 2628 510
rect 2306 189 2628 190
rect 2016 62 2143 78
rect 2016 -62 2120 62
rect 2016 -78 2143 -62
rect 1587 -190 1909 -189
rect 1587 -510 1588 -190
rect 1908 -510 1909 -190
rect 1587 -511 1909 -510
rect 1297 -638 1424 -622
rect 1297 -762 1401 -638
rect 1297 -778 1424 -762
rect 868 -890 1190 -889
rect 868 -1210 869 -890
rect 1189 -1210 1190 -890
rect 868 -1211 1190 -1210
rect 578 -1338 705 -1322
rect 578 -1462 682 -1338
rect 578 -1478 705 -1462
rect 149 -1590 471 -1589
rect 149 -1910 150 -1590
rect 470 -1910 471 -1590
rect 149 -1911 471 -1910
rect -141 -2038 -14 -2022
rect -141 -2162 -37 -2038
rect -141 -2178 -14 -2162
rect -570 -2290 -248 -2289
rect -570 -2610 -569 -2290
rect -249 -2610 -248 -2290
rect -570 -2611 -248 -2610
rect -860 -2738 -733 -2722
rect -860 -2862 -756 -2738
rect -860 -2878 -733 -2862
rect -1289 -2990 -967 -2989
rect -1289 -3310 -1288 -2990
rect -968 -3310 -967 -2990
rect -1289 -3311 -967 -3310
rect -1579 -3438 -1452 -3422
rect -1579 -3500 -1475 -3438
rect -1180 -3500 -1076 -3311
rect -860 -3422 -813 -2878
rect -749 -3422 -733 -2878
rect -461 -2989 -357 -2611
rect -141 -2722 -94 -2178
rect -30 -2722 -14 -2178
rect 258 -2289 362 -1911
rect 578 -2022 625 -1478
rect 689 -2022 705 -1478
rect 977 -1589 1081 -1211
rect 1297 -1322 1344 -778
rect 1408 -1322 1424 -778
rect 1696 -889 1800 -511
rect 2016 -622 2063 -78
rect 2127 -622 2143 -78
rect 2415 -189 2519 189
rect 2735 78 2782 622
rect 2846 78 2862 622
rect 3134 511 3238 889
rect 3454 778 3501 1322
rect 3565 778 3581 1322
rect 3454 762 3581 778
rect 3454 638 3558 762
rect 3454 622 3581 638
rect 3025 510 3347 511
rect 3025 190 3026 510
rect 3346 190 3347 510
rect 3025 189 3347 190
rect 2735 62 2862 78
rect 2735 -62 2839 62
rect 2735 -78 2862 -62
rect 2306 -190 2628 -189
rect 2306 -510 2307 -190
rect 2627 -510 2628 -190
rect 2306 -511 2628 -510
rect 2016 -638 2143 -622
rect 2016 -762 2120 -638
rect 2016 -778 2143 -762
rect 1587 -890 1909 -889
rect 1587 -1210 1588 -890
rect 1908 -1210 1909 -890
rect 1587 -1211 1909 -1210
rect 1297 -1338 1424 -1322
rect 1297 -1462 1401 -1338
rect 1297 -1478 1424 -1462
rect 868 -1590 1190 -1589
rect 868 -1910 869 -1590
rect 1189 -1910 1190 -1590
rect 868 -1911 1190 -1910
rect 578 -2038 705 -2022
rect 578 -2162 682 -2038
rect 578 -2178 705 -2162
rect 149 -2290 471 -2289
rect 149 -2610 150 -2290
rect 470 -2610 471 -2290
rect 149 -2611 471 -2610
rect -141 -2738 -14 -2722
rect -141 -2862 -37 -2738
rect -141 -2878 -14 -2862
rect -570 -2990 -248 -2989
rect -570 -3310 -569 -2990
rect -249 -3310 -248 -2990
rect -570 -3311 -248 -3310
rect -860 -3438 -733 -3422
rect -860 -3500 -756 -3438
rect -461 -3500 -357 -3311
rect -141 -3422 -94 -2878
rect -30 -3422 -14 -2878
rect 258 -2989 362 -2611
rect 578 -2722 625 -2178
rect 689 -2722 705 -2178
rect 977 -2289 1081 -1911
rect 1297 -2022 1344 -1478
rect 1408 -2022 1424 -1478
rect 1696 -1589 1800 -1211
rect 2016 -1322 2063 -778
rect 2127 -1322 2143 -778
rect 2415 -889 2519 -511
rect 2735 -622 2782 -78
rect 2846 -622 2862 -78
rect 3134 -189 3238 189
rect 3454 78 3501 622
rect 3565 78 3581 622
rect 3454 62 3581 78
rect 3454 -62 3558 62
rect 3454 -78 3581 -62
rect 3025 -190 3347 -189
rect 3025 -510 3026 -190
rect 3346 -510 3347 -190
rect 3025 -511 3347 -510
rect 2735 -638 2862 -622
rect 2735 -762 2839 -638
rect 2735 -778 2862 -762
rect 2306 -890 2628 -889
rect 2306 -1210 2307 -890
rect 2627 -1210 2628 -890
rect 2306 -1211 2628 -1210
rect 2016 -1338 2143 -1322
rect 2016 -1462 2120 -1338
rect 2016 -1478 2143 -1462
rect 1587 -1590 1909 -1589
rect 1587 -1910 1588 -1590
rect 1908 -1910 1909 -1590
rect 1587 -1911 1909 -1910
rect 1297 -2038 1424 -2022
rect 1297 -2162 1401 -2038
rect 1297 -2178 1424 -2162
rect 868 -2290 1190 -2289
rect 868 -2610 869 -2290
rect 1189 -2610 1190 -2290
rect 868 -2611 1190 -2610
rect 578 -2738 705 -2722
rect 578 -2862 682 -2738
rect 578 -2878 705 -2862
rect 149 -2990 471 -2989
rect 149 -3310 150 -2990
rect 470 -3310 471 -2990
rect 149 -3311 471 -3310
rect -141 -3438 -14 -3422
rect -141 -3500 -37 -3438
rect 258 -3500 362 -3311
rect 578 -3422 625 -2878
rect 689 -3422 705 -2878
rect 977 -2989 1081 -2611
rect 1297 -2722 1344 -2178
rect 1408 -2722 1424 -2178
rect 1696 -2289 1800 -1911
rect 2016 -2022 2063 -1478
rect 2127 -2022 2143 -1478
rect 2415 -1589 2519 -1211
rect 2735 -1322 2782 -778
rect 2846 -1322 2862 -778
rect 3134 -889 3238 -511
rect 3454 -622 3501 -78
rect 3565 -622 3581 -78
rect 3454 -638 3581 -622
rect 3454 -762 3558 -638
rect 3454 -778 3581 -762
rect 3025 -890 3347 -889
rect 3025 -1210 3026 -890
rect 3346 -1210 3347 -890
rect 3025 -1211 3347 -1210
rect 2735 -1338 2862 -1322
rect 2735 -1462 2839 -1338
rect 2735 -1478 2862 -1462
rect 2306 -1590 2628 -1589
rect 2306 -1910 2307 -1590
rect 2627 -1910 2628 -1590
rect 2306 -1911 2628 -1910
rect 2016 -2038 2143 -2022
rect 2016 -2162 2120 -2038
rect 2016 -2178 2143 -2162
rect 1587 -2290 1909 -2289
rect 1587 -2610 1588 -2290
rect 1908 -2610 1909 -2290
rect 1587 -2611 1909 -2610
rect 1297 -2738 1424 -2722
rect 1297 -2862 1401 -2738
rect 1297 -2878 1424 -2862
rect 868 -2990 1190 -2989
rect 868 -3310 869 -2990
rect 1189 -3310 1190 -2990
rect 868 -3311 1190 -3310
rect 578 -3438 705 -3422
rect 578 -3500 682 -3438
rect 977 -3500 1081 -3311
rect 1297 -3422 1344 -2878
rect 1408 -3422 1424 -2878
rect 1696 -2989 1800 -2611
rect 2016 -2722 2063 -2178
rect 2127 -2722 2143 -2178
rect 2415 -2289 2519 -1911
rect 2735 -2022 2782 -1478
rect 2846 -2022 2862 -1478
rect 3134 -1589 3238 -1211
rect 3454 -1322 3501 -778
rect 3565 -1322 3581 -778
rect 3454 -1338 3581 -1322
rect 3454 -1462 3558 -1338
rect 3454 -1478 3581 -1462
rect 3025 -1590 3347 -1589
rect 3025 -1910 3026 -1590
rect 3346 -1910 3347 -1590
rect 3025 -1911 3347 -1910
rect 2735 -2038 2862 -2022
rect 2735 -2162 2839 -2038
rect 2735 -2178 2862 -2162
rect 2306 -2290 2628 -2289
rect 2306 -2610 2307 -2290
rect 2627 -2610 2628 -2290
rect 2306 -2611 2628 -2610
rect 2016 -2738 2143 -2722
rect 2016 -2862 2120 -2738
rect 2016 -2878 2143 -2862
rect 1587 -2990 1909 -2989
rect 1587 -3310 1588 -2990
rect 1908 -3310 1909 -2990
rect 1587 -3311 1909 -3310
rect 1297 -3438 1424 -3422
rect 1297 -3500 1401 -3438
rect 1696 -3500 1800 -3311
rect 2016 -3422 2063 -2878
rect 2127 -3422 2143 -2878
rect 2415 -2989 2519 -2611
rect 2735 -2722 2782 -2178
rect 2846 -2722 2862 -2178
rect 3134 -2289 3238 -1911
rect 3454 -2022 3501 -1478
rect 3565 -2022 3581 -1478
rect 3454 -2038 3581 -2022
rect 3454 -2162 3558 -2038
rect 3454 -2178 3581 -2162
rect 3025 -2290 3347 -2289
rect 3025 -2610 3026 -2290
rect 3346 -2610 3347 -2290
rect 3025 -2611 3347 -2610
rect 2735 -2738 2862 -2722
rect 2735 -2862 2839 -2738
rect 2735 -2878 2862 -2862
rect 2306 -2990 2628 -2989
rect 2306 -3310 2307 -2990
rect 2627 -3310 2628 -2990
rect 2306 -3311 2628 -3310
rect 2016 -3438 2143 -3422
rect 2016 -3500 2120 -3438
rect 2415 -3500 2519 -3311
rect 2735 -3422 2782 -2878
rect 2846 -3422 2862 -2878
rect 3134 -2989 3238 -2611
rect 3454 -2722 3501 -2178
rect 3565 -2722 3581 -2178
rect 3454 -2738 3581 -2722
rect 3454 -2862 3558 -2738
rect 3454 -2878 3581 -2862
rect 3025 -2990 3347 -2989
rect 3025 -3310 3026 -2990
rect 3346 -3310 3347 -2990
rect 3025 -3311 3347 -3310
rect 2735 -3438 2862 -3422
rect 2735 -3500 2839 -3438
rect 3134 -3500 3238 -3311
rect 3454 -3422 3501 -2878
rect 3565 -3422 3581 -2878
rect 3454 -3438 3581 -3422
rect 3454 -3500 3558 -3438
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 2886 2850 3486 3450
string parameters w 2.00 l 2.00 val 5.36 carea 1.00 cperi 0.17 nx 10 ny 10 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
