magic
tech sky130A
magscale 1 2
timestamp 1621213367
<< xpolycontact >>
rect -6829 3152 -6259 3584
rect -6829 -3584 -6259 -3152
rect -6011 3152 -5441 3584
rect -6011 -3584 -5441 -3152
rect -5193 3152 -4623 3584
rect -5193 -3584 -4623 -3152
rect -4375 3152 -3805 3584
rect -4375 -3584 -3805 -3152
rect -3557 3152 -2987 3584
rect -3557 -3584 -2987 -3152
rect -2739 3152 -2169 3584
rect -2739 -3584 -2169 -3152
rect -1921 3152 -1351 3584
rect -1921 -3584 -1351 -3152
rect -1103 3152 -533 3584
rect -1103 -3584 -533 -3152
rect -285 3152 285 3584
rect -285 -3584 285 -3152
rect 533 3152 1103 3584
rect 533 -3584 1103 -3152
rect 1351 3152 1921 3584
rect 1351 -3584 1921 -3152
rect 2169 3152 2739 3584
rect 2169 -3584 2739 -3152
rect 2987 3152 3557 3584
rect 2987 -3584 3557 -3152
rect 3805 3152 4375 3584
rect 3805 -3584 4375 -3152
rect 4623 3152 5193 3584
rect 4623 -3584 5193 -3152
rect 5441 3152 6011 3584
rect 5441 -3584 6011 -3152
rect 6259 3152 6829 3584
rect 6259 -3584 6829 -3152
<< xpolyres >>
rect -6829 -3152 -6259 3152
rect -6011 -3152 -5441 3152
rect -5193 -3152 -4623 3152
rect -4375 -3152 -3805 3152
rect -3557 -3152 -2987 3152
rect -2739 -3152 -2169 3152
rect -1921 -3152 -1351 3152
rect -1103 -3152 -533 3152
rect -285 -3152 285 3152
rect 533 -3152 1103 3152
rect 1351 -3152 1921 3152
rect 2169 -3152 2739 3152
rect 2987 -3152 3557 3152
rect 3805 -3152 4375 3152
rect 4623 -3152 5193 3152
rect 5441 -3152 6011 3152
rect 6259 -3152 6829 3152
<< res2p85 >>
rect -6831 -3154 -6257 3154
rect -6013 -3154 -5439 3154
rect -5195 -3154 -4621 3154
rect -4377 -3154 -3803 3154
rect -3559 -3154 -2985 3154
rect -2741 -3154 -2167 3154
rect -1923 -3154 -1349 3154
rect -1105 -3154 -531 3154
rect -287 -3154 287 3154
rect 531 -3154 1105 3154
rect 1349 -3154 1923 3154
rect 2167 -3154 2741 3154
rect 2985 -3154 3559 3154
rect 3803 -3154 4377 3154
rect 4621 -3154 5195 3154
rect 5439 -3154 6013 3154
rect 6257 -3154 6831 3154
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_2p85
string parameters w 2.850 l 31.52 m 1 nx 17 wmin 2.850 lmin 0.50 rho 2000 val 22.132k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 2.850 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 0 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
