magic
tech sky130A
timestamp 1621229569
<< nmoslvt >>
rect -100 -1350 100 1350
<< ndiff >>
rect -129 1344 -100 1350
rect -129 -1344 -123 1344
rect -106 -1344 -100 1344
rect -129 -1350 -100 -1344
rect 100 1344 129 1350
rect 100 -1344 106 1344
rect 123 -1344 129 1344
rect 100 -1350 129 -1344
<< ndiffc >>
rect -123 -1344 -106 1344
rect 106 -1344 123 1344
<< poly >>
rect -100 1386 100 1394
rect -100 1369 -92 1386
rect 92 1369 100 1386
rect -100 1350 100 1369
rect -100 -1369 100 -1350
rect -100 -1386 -92 -1369
rect 92 -1386 100 -1369
rect -100 -1394 100 -1386
<< polycont >>
rect -92 1369 92 1386
rect -92 -1386 92 -1369
<< locali >>
rect -100 1369 -92 1386
rect 92 1369 100 1386
rect -123 1344 -106 1352
rect -123 -1352 -106 -1344
rect 106 1344 123 1352
rect 106 -1352 123 -1344
rect -100 -1386 -92 -1369
rect 92 -1386 100 -1369
<< viali >>
rect -92 1369 92 1386
rect -123 -1344 -106 1344
rect 106 -1344 123 1344
rect -92 -1386 92 -1369
<< metal1 >>
rect -98 1386 98 1389
rect -98 1369 -92 1386
rect 92 1369 98 1386
rect -98 1366 98 1369
rect -126 1344 -103 1350
rect -126 -1344 -123 1344
rect -106 -1344 -103 1344
rect -126 -1350 -103 -1344
rect 103 1344 126 1350
rect 103 -1344 106 1344
rect 123 -1344 126 1344
rect 103 -1350 126 -1344
rect -98 -1369 98 -1366
rect -98 -1386 -92 -1369
rect 92 -1386 98 -1369
rect -98 -1389 98 -1386
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string parameters w 27 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
