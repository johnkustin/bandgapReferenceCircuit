magic
tech sky130A
magscale 1 2
timestamp 1621231188
<< psubdiff >>
rect -17894 9382 -11418 9394
rect -17894 9050 -17882 9382
rect -11430 9050 -11418 9382
rect -17894 9038 -11418 9050
<< psubdiffcont >>
rect -17882 9050 -11430 9382
<< locali >>
rect -17898 9388 -11414 9398
rect -17898 9044 -17888 9388
rect -11424 9044 -11414 9388
rect -17898 9034 -11414 9044
<< viali >>
rect -17888 9382 -11424 9388
rect -17888 9050 -17882 9382
rect -17882 9050 -11430 9382
rect -11430 9050 -11424 9382
rect -17888 9044 -11424 9050
<< metal1 >>
rect -8104 15426 -7556 16438
rect 9804 13500 10508 15196
rect -2890 12808 10508 13500
rect 9278 12640 10226 12646
rect 9278 12122 9286 12640
rect 10220 12122 10226 12640
rect -8390 11860 -6390 11902
rect -8390 11410 -8384 11860
rect -6396 11410 -6390 11860
rect -9908 11104 -9776 11110
rect -9908 10690 -9902 11104
rect -9782 10690 -9776 11104
rect -8390 10996 -6390 11410
rect 5310 11860 7310 11902
rect 5310 11410 5316 11860
rect 7304 11410 7310 11860
rect 5310 10996 7310 11410
rect -10364 10398 -10232 10684
rect -10364 10106 -10358 10398
rect -10238 10106 -10232 10398
rect -17900 9388 -11412 9400
rect -17900 9044 -17888 9388
rect -11424 9044 -11412 9388
rect -17900 8832 -11412 9044
rect -19254 8502 -17208 8710
rect -17894 8038 -11418 8394
rect -18930 5002 -18724 5008
rect -18930 4944 -18924 5002
rect -18730 4944 -18724 5002
rect -18930 1358 -18724 4944
rect -17894 4282 -17686 8038
rect -11626 4282 -11418 8038
rect -10364 6866 -10232 10106
rect -9908 7006 -9776 10690
rect -5690 9502 -3690 10408
rect 2610 9502 4610 10408
rect -9908 6926 -9902 7006
rect -9782 6926 -9776 7006
rect -9908 6920 -9776 6926
rect -10364 6786 -10358 6866
rect -10248 6786 -10232 6866
rect -10364 6780 -10232 6786
rect -9496 4630 -9016 4636
rect -9496 4376 -9490 4630
rect -9022 4376 -9016 4630
rect -9496 1536 -9016 4376
rect 9278 2220 10226 12122
rect 11440 10396 12144 15196
rect 11440 10108 11448 10396
rect 12138 10108 12144 10396
rect 11440 10102 12144 10108
rect -9496 1388 -9490 1536
rect -9022 1388 -9016 1536
rect -9496 1382 -9016 1388
rect -18930 1244 -18924 1358
rect -18730 1244 -18724 1358
rect -18930 1238 -18724 1244
<< via1 >>
rect 9286 12122 10220 12640
rect -8384 11410 -6396 11860
rect -9902 10690 -9782 11104
rect 5316 11410 7304 11860
rect -10358 10106 -10238 10398
rect -18924 4944 -18730 5002
rect -9902 6926 -9782 7006
rect -10358 6786 -10248 6866
rect -9490 4376 -9022 4630
rect 10628 11410 11320 11860
rect 11448 10108 12138 10396
rect -9490 1388 -9022 1536
rect -18924 1244 -18730 1358
<< metal2 >>
rect 5714 12646 6416 14640
rect 5714 12640 10226 12646
rect 5714 12122 9286 12640
rect 10220 12122 10226 12640
rect 5714 12116 10226 12122
rect -9906 11860 11340 11868
rect -9906 11410 -8384 11860
rect -6396 11410 5316 11860
rect 7304 11410 10628 11860
rect 11320 11410 11340 11860
rect -9906 11110 11340 11410
rect -9908 11104 11340 11110
rect -9908 10690 -9902 11104
rect -9782 10690 11340 11104
rect -9908 10686 11340 10690
rect -9908 10684 -9776 10686
rect -10364 10398 12144 10402
rect -10364 10106 -10358 10398
rect -10238 10396 12144 10398
rect -10238 10108 11448 10396
rect 12138 10108 12144 10396
rect -10238 10106 12144 10108
rect -10364 9802 12144 10106
rect -14276 6926 -9902 7006
rect -9782 6926 -9776 7006
rect -14848 6786 -10358 6866
rect -10248 6786 -10242 6866
rect -19536 5002 -18724 5008
rect -19536 4944 -18924 5002
rect -18730 4944 -18724 5002
rect -19536 4938 -18724 4944
rect -21317 4664 -12946 4798
rect -11488 4630 -9016 4636
rect -11488 4376 -9490 4630
rect -9022 4376 -9016 4630
rect -11488 4370 -9016 4376
rect -19268 1438 -19266 1562
rect -10006 1438 -10002 1562
rect -9496 1536 -8010 1542
rect -9496 1388 -9490 1536
rect -9022 1388 -8010 1536
rect -9496 1382 -8010 1388
rect -18930 1362 -18724 1364
rect -18930 1358 -17838 1362
rect -18930 1244 -18924 1358
rect -18730 1244 -17838 1358
rect -18930 1238 -17838 1244
rect -9504 1324 8454 1334
rect -9504 1006 -9494 1324
rect 8444 1006 8454 1324
rect -9504 998 8454 1006
<< via2 >>
rect -19258 1442 -10012 1556
rect -9494 1006 8444 1324
<< metal3 >>
rect -19266 1556 8465 1562
rect -19266 1442 -19258 1556
rect -10012 1442 8465 1556
rect -20266 1324 8465 1442
rect -20266 1006 -9494 1324
rect 8444 1006 8465 1324
rect -20266 1000 8465 1006
use sky130_fd_pr__nfet_01v8_lvt_5FLLME  sky130_fd_pr__nfet_01v8_lvt_5FLLME_0
timestamp 1621229569
transform 0 1 -14507 -1 0 8606
box -258 -2757 258 2757
use currentmirror  currentmirror_0
timestamp 1621228141
transform 1 0 -8490 0 -1 9302
box -1748 -4198 17156 8302
use bandgapcorev3  bandgapcorev3_0
timestamp 1621229569
transform 0 1 30186 -1 0 28802
box 5270 -39968 26884 -11302
use ampcurrentsource  ampcurrentsource_0
timestamp 1621192096
transform 1 0 -21372 0 1 5166
box -498 -438 2400 694
use amplifier  amplifier_0
timestamp 1621192096
transform 1 0 -16310 0 -1 6762
box -3090 -244 6438 5762
<< labels >>
flabel metal1 -19254 8502 -18792 8700 1 FreeSans 1600 0 0 0 porst
flabel metal1 -2858 12824 1810 13500 1 FreeSans 1600 0 0 0 Vbg
port 1 n
flabel metal3 -20266 1000 -19556 1422 1 FreeSans 1600 0 0 0 VDD!
<< end >>
