magic
tech sky130A
magscale 1 2
timestamp 1621270775
<< error_s >>
rect 106 -1406 112 -1400
rect 2088 -1406 2094 -1400
rect 100 -1412 106 -1406
rect 2094 -1412 2100 -1406
rect 100 -1694 106 -1688
rect 2094 -1694 2100 -1688
rect 106 -1700 112 -1694
rect 2088 -1700 2094 -1694
<< nwell >>
rect -1110 7700 -358 7702
rect -1110 -200 -212 7700
rect 98 -200 120 7700
rect 4800 -200 5600 7700
rect 10300 -200 11100 7700
rect 15800 -200 15810 7700
rect 16180 7588 16226 7690
rect 16266 -198 17156 7702
<< nsubdiff >>
rect -1010 7200 -410 7400
rect -1010 200 -810 7200
rect -610 200 -410 7200
rect -1010 0 -410 200
rect 4900 7200 5500 7400
rect 4900 200 5100 7200
rect 5300 200 5500 7200
rect 4900 0 5500 200
rect 10400 7200 11000 7400
rect 10400 200 10600 7200
rect 10800 200 11000 7200
rect 10400 0 11000 200
rect 16356 7202 16956 7402
rect 16356 202 16556 7202
rect 16756 202 16956 7202
rect 16356 2 16956 202
<< nsubdiffcont >>
rect -810 200 -610 7200
rect 5100 200 5300 7200
rect 10600 200 10800 7200
rect 16556 202 16756 7202
<< locali >>
rect -1010 8200 -410 8300
rect -1010 8100 -910 8200
rect -510 8100 -410 8200
rect -1010 7200 -410 8100
rect -1010 200 -810 7200
rect -610 200 -410 7200
rect -1010 0 -410 200
rect 4900 8200 5500 8300
rect 4900 8100 5000 8200
rect 5400 8100 5500 8200
rect 4900 7200 5500 8100
rect 4900 200 5100 7200
rect 5300 200 5500 7200
rect 4900 0 5500 200
rect 10400 8200 11000 8300
rect 10400 8100 10500 8200
rect 10900 8100 11000 8200
rect 10400 7200 11000 8100
rect 10400 200 10600 7200
rect 10800 200 11000 7200
rect 10400 0 11000 200
rect 16356 8202 16956 8302
rect 16356 8102 16456 8202
rect 16856 8102 16956 8202
rect 16356 7202 16956 8102
rect 16356 202 16556 7202
rect 16756 202 16956 7202
rect 16356 2 16956 202
<< viali >>
rect -910 8100 -510 8200
rect 5000 8100 5400 8200
rect 10500 8100 10900 8200
rect 16456 8102 16856 8202
<< metal1 >>
rect -1010 8200 142 8300
rect -1010 8100 -910 8200
rect -510 8100 142 8200
rect -1010 8000 142 8100
rect 4900 8200 5500 8300
rect 4900 8100 5000 8200
rect 5400 8100 5500 8200
rect -316 7648 142 8000
rect 560 8060 680 8080
rect 560 7980 580 8060
rect 660 7980 680 8060
rect 560 7960 680 7980
rect 1480 8060 1600 8080
rect 1480 7980 1500 8060
rect 1580 7980 1600 8060
rect 1480 7960 1600 7980
rect 2400 8060 2520 8080
rect 2400 7980 2420 8060
rect 2500 7980 2520 8060
rect 2400 7960 2520 7980
rect 3320 8060 3440 8080
rect 3320 7980 3340 8060
rect 3420 7980 3440 8060
rect 3320 7960 3440 7980
rect 4240 8060 4360 8080
rect 4240 7980 4260 8060
rect 4340 7980 4360 8060
rect 4900 8000 5500 8100
rect 10400 8200 11000 8300
rect 10400 8100 10500 8200
rect 10900 8100 11000 8200
rect 6060 8060 6180 8080
rect 4240 7960 4360 7980
rect 6060 7980 6080 8060
rect 6160 7980 6180 8060
rect 6060 7960 6180 7980
rect 6980 8060 7100 8080
rect 6980 7980 7000 8060
rect 7080 7980 7100 8060
rect 6980 7960 7100 7980
rect 7900 8060 8020 8080
rect 7900 7980 7920 8060
rect 8000 7980 8020 8060
rect 7900 7960 8020 7980
rect 8820 8060 8940 8080
rect 8820 7980 8840 8060
rect 8920 7980 8940 8060
rect 8820 7960 8940 7980
rect 9740 8060 9860 8080
rect 9740 7980 9760 8060
rect 9840 7980 9860 8060
rect 10400 8000 11000 8100
rect 15768 8202 16956 8302
rect 15768 8102 16456 8202
rect 16856 8102 16956 8202
rect 11560 8060 11680 8080
rect 9740 7960 9860 7980
rect 11560 7980 11580 8060
rect 11660 7980 11680 8060
rect 11560 7960 11680 7980
rect 12480 8060 12600 8080
rect 12480 7980 12500 8060
rect 12580 7980 12600 8060
rect 12480 7960 12600 7980
rect 13400 8060 13520 8080
rect 13400 7980 13420 8060
rect 13500 7980 13520 8060
rect 13400 7960 13520 7980
rect 14320 8060 14440 8080
rect 14320 7980 14340 8060
rect 14420 7980 14440 8060
rect 14320 7960 14440 7980
rect 15240 8060 15360 8080
rect 15240 7980 15260 8060
rect 15340 7980 15360 8060
rect 15240 7960 15360 7980
rect 15768 8002 16956 8102
rect -316 7642 -168 7648
rect 24 7642 142 7648
rect 300 7900 480 7920
rect 300 7780 320 7900
rect 460 7780 480 7900
rect -316 7600 -270 7642
rect 300 7640 480 7780
rect -316 7596 -276 7600
rect -316 -132 -270 7596
rect 142 -100 188 7606
rect 600 7580 640 7960
rect 760 7900 940 7920
rect 760 7780 780 7900
rect 920 7780 940 7900
rect 760 7640 940 7780
rect 1220 7900 1400 7920
rect 1220 7780 1240 7900
rect 1380 7780 1400 7900
rect 1220 7640 1400 7780
rect 1520 7580 1560 7960
rect 1680 7900 1860 7920
rect 1680 7780 1700 7900
rect 1840 7780 1860 7900
rect 1680 7640 1860 7780
rect 2140 7900 2320 7920
rect 2140 7780 2160 7900
rect 2300 7780 2320 7900
rect 2140 7640 2320 7780
rect 2440 7580 2480 7960
rect 2600 7900 2780 7920
rect 2600 7780 2620 7900
rect 2760 7780 2780 7900
rect 2600 7640 2780 7780
rect 3060 7900 3240 7920
rect 3060 7780 3080 7900
rect 3220 7780 3240 7900
rect 3060 7640 3240 7780
rect 3340 7580 3380 7960
rect 3520 7900 3700 7920
rect 3520 7780 3540 7900
rect 3680 7780 3700 7900
rect 3520 7640 3700 7780
rect 3980 7900 4160 7920
rect 3980 7780 4000 7900
rect 4140 7780 4160 7900
rect 3980 7640 4160 7780
rect 4260 7580 4300 7960
rect 4440 7900 4620 7920
rect 4440 7780 4460 7900
rect 4600 7780 4620 7900
rect 4440 7640 4620 7780
rect 5800 7900 5980 7920
rect 5800 7780 5820 7900
rect 5960 7780 5980 7900
rect 5800 7640 5980 7780
rect 6100 7580 6140 7960
rect 6260 7900 6440 7920
rect 6260 7780 6280 7900
rect 6420 7780 6440 7900
rect 6260 7640 6440 7780
rect 6720 7900 6900 7920
rect 6720 7780 6740 7900
rect 6880 7780 6900 7900
rect 6720 7640 6900 7780
rect 7020 7580 7060 7960
rect 7180 7900 7360 7920
rect 7180 7780 7200 7900
rect 7340 7780 7360 7900
rect 7180 7640 7360 7780
rect 7640 7900 7820 7920
rect 7640 7780 7660 7900
rect 7800 7780 7820 7900
rect 7640 7640 7820 7780
rect 7940 7580 7980 7960
rect 8100 7900 8280 7920
rect 8100 7780 8120 7900
rect 8260 7780 8280 7900
rect 8100 7640 8280 7780
rect 8560 7900 8740 7920
rect 8560 7780 8580 7900
rect 8720 7780 8740 7900
rect 8560 7640 8740 7780
rect 8840 7580 8880 7960
rect 9020 7900 9200 7920
rect 9020 7780 9040 7900
rect 9180 7780 9200 7900
rect 9020 7640 9200 7780
rect 9480 7900 9660 7920
rect 9480 7780 9500 7900
rect 9640 7780 9660 7900
rect 9480 7640 9660 7780
rect 9760 7580 9800 7960
rect 9940 7900 10120 7920
rect 9940 7780 9960 7900
rect 10100 7780 10120 7900
rect 9940 7640 10120 7780
rect 11300 7900 11480 7920
rect 11300 7780 11320 7900
rect 11460 7780 11480 7900
rect 11300 7640 11480 7780
rect 11600 7580 11640 7960
rect 11760 7900 11940 7920
rect 11760 7780 11780 7900
rect 11920 7780 11940 7900
rect 11760 7640 11940 7780
rect 12220 7900 12400 7920
rect 12220 7780 12240 7900
rect 12380 7780 12400 7900
rect 12220 7640 12400 7780
rect 12520 7580 12560 7960
rect 12680 7900 12860 7920
rect 12680 7780 12700 7900
rect 12840 7780 12860 7900
rect 12680 7640 12860 7780
rect 13140 7900 13320 7920
rect 13140 7780 13160 7900
rect 13300 7780 13320 7900
rect 13140 7640 13320 7780
rect 13440 7580 13480 7960
rect 13600 7900 13780 7920
rect 13600 7780 13620 7900
rect 13760 7780 13780 7900
rect 13600 7640 13780 7780
rect 14060 7900 14240 7920
rect 14060 7780 14080 7900
rect 14220 7780 14240 7900
rect 14060 7640 14240 7780
rect 14340 7580 14380 7960
rect 14520 7900 14700 7920
rect 14520 7780 14540 7900
rect 14680 7780 14700 7900
rect 14520 7640 14700 7780
rect 14980 7900 15160 7920
rect 14980 7780 15000 7900
rect 15140 7780 15160 7900
rect 14980 7640 15160 7780
rect 15260 7580 15300 7960
rect 15440 7900 15620 7920
rect 15440 7780 15460 7900
rect 15600 7780 15620 7900
rect 15440 7640 15620 7780
rect 15768 7642 16226 8002
rect 140 -132 188 -100
rect 140 -200 180 -132
rect 1060 -200 1100 -120
rect 1980 -200 2020 -100
rect 2880 -200 2940 -120
rect 3800 -200 3860 -100
rect 4720 -200 4780 -100
rect 5640 -198 5680 -120
rect 6560 -198 6600 -120
rect 7480 -198 7520 -100
rect 8400 -198 8440 -100
rect 9300 -198 9360 -100
rect 10220 -198 10280 -100
rect 100 -1406 2100 -200
rect 2800 -806 4800 -200
rect 2800 -1094 2806 -806
rect 4794 -1094 4800 -806
rect 2800 -1100 4800 -1094
rect 100 -1694 106 -1406
rect 2094 -1694 2100 -1406
rect 100 -1800 2100 -1694
rect 5600 -4198 10300 -198
rect 11140 -200 11180 -100
rect 12060 -200 12100 -100
rect 12980 -200 13020 -100
rect 13880 -200 13940 -100
rect 15722 -120 15768 7606
rect 16180 7588 16226 7642
rect 14800 -200 14860 -120
rect 15720 -132 15768 -120
rect 16183 -129 16223 7588
rect 15720 -200 15760 -132
rect 11100 -806 13100 -200
rect 11100 -1094 11106 -806
rect 13094 -1094 13100 -806
rect 11100 -1100 13100 -1094
rect 13800 -1406 15800 -200
rect 13800 -1694 13806 -1406
rect 15794 -1694 15800 -1406
rect 13800 -1800 15800 -1694
<< via1 >>
rect -910 8100 -510 8200
rect 5000 8100 5400 8200
rect 580 7980 660 8060
rect 1500 7980 1580 8060
rect 2420 7980 2500 8060
rect 3340 7980 3420 8060
rect 4260 7980 4340 8060
rect 10500 8100 10900 8200
rect 6080 7980 6160 8060
rect 7000 7980 7080 8060
rect 7920 7980 8000 8060
rect 8840 7980 8920 8060
rect 9760 7980 9840 8060
rect 16456 8102 16856 8202
rect 11580 7980 11660 8060
rect 12500 7980 12580 8060
rect 13420 7980 13500 8060
rect 14340 7980 14420 8060
rect 15260 7980 15340 8060
rect 320 7780 460 7900
rect 780 7780 920 7900
rect 1240 7780 1380 7900
rect 1700 7780 1840 7900
rect 2160 7780 2300 7900
rect 2620 7780 2760 7900
rect 3080 7780 3220 7900
rect 3540 7780 3680 7900
rect 4000 7780 4140 7900
rect 4460 7780 4600 7900
rect 5820 7780 5960 7900
rect 6280 7780 6420 7900
rect 6740 7780 6880 7900
rect 7200 7780 7340 7900
rect 7660 7780 7800 7900
rect 8120 7780 8260 7900
rect 8580 7780 8720 7900
rect 9040 7780 9180 7900
rect 9500 7780 9640 7900
rect 9960 7780 10100 7900
rect 11320 7780 11460 7900
rect 11780 7780 11920 7900
rect 12240 7780 12380 7900
rect 12700 7780 12840 7900
rect 13160 7780 13300 7900
rect 13620 7780 13760 7900
rect 14080 7780 14220 7900
rect 14540 7780 14680 7900
rect 15000 7780 15140 7900
rect 15460 7780 15600 7900
rect 2806 -1094 4794 -806
rect 106 -1694 2094 -1406
rect 11106 -1094 13094 -806
rect 13806 -1694 15794 -1406
<< metal2 >>
rect -1010 8200 -410 8300
rect -1010 8100 -910 8200
rect -510 8100 -410 8200
rect -1010 8000 -410 8100
rect 4900 8200 5500 8300
rect 4900 8100 5000 8200
rect 5400 8100 5500 8200
rect 560 8060 680 8080
rect 560 7980 580 8060
rect 660 7980 680 8060
rect 560 7960 680 7980
rect 1480 8060 1600 8080
rect 1480 7980 1500 8060
rect 1580 7980 1600 8060
rect 1480 7960 1600 7980
rect 2400 8060 2520 8080
rect 2400 7980 2420 8060
rect 2500 7980 2520 8060
rect 2400 7960 2520 7980
rect 3320 8060 3440 8080
rect 3320 7980 3340 8060
rect 3420 7980 3440 8060
rect 3320 7960 3440 7980
rect 4240 8060 4360 8080
rect 4240 7980 4260 8060
rect 4340 7980 4360 8060
rect 4900 8000 5500 8100
rect 10400 8200 11000 8300
rect 10400 8100 10500 8200
rect 10900 8100 11000 8200
rect 6060 8060 6180 8080
rect 4240 7960 4360 7980
rect 6060 7980 6080 8060
rect 6160 7980 6180 8060
rect 6060 7960 6180 7980
rect 6980 8060 7100 8080
rect 6980 7980 7000 8060
rect 7080 7980 7100 8060
rect 6980 7960 7100 7980
rect 7900 8060 8020 8080
rect 7900 7980 7920 8060
rect 8000 7980 8020 8060
rect 7900 7960 8020 7980
rect 8820 8060 8940 8080
rect 8820 7980 8840 8060
rect 8920 7980 8940 8060
rect 8820 7960 8940 7980
rect 9740 8060 9860 8080
rect 9740 7980 9760 8060
rect 9840 7980 9860 8060
rect 10400 8000 11000 8100
rect 16356 8202 16956 8302
rect 16356 8102 16456 8202
rect 16856 8102 16956 8202
rect 11560 8060 11680 8080
rect 9740 7960 9860 7980
rect 11560 7980 11580 8060
rect 11660 7980 11680 8060
rect 11560 7960 11680 7980
rect 12480 8060 12600 8080
rect 12480 7980 12500 8060
rect 12580 7980 12600 8060
rect 12480 7960 12600 7980
rect 13400 8060 13520 8080
rect 13400 7980 13420 8060
rect 13500 7980 13520 8060
rect 13400 7960 13520 7980
rect 14320 8060 14440 8080
rect 14320 7980 14340 8060
rect 14420 7980 14440 8060
rect 14320 7960 14440 7980
rect 15240 8060 15360 8080
rect 15240 7980 15260 8060
rect 15340 7980 15360 8060
rect 16356 8002 16956 8102
rect 15240 7960 15360 7980
rect 300 7900 15620 7920
rect 300 7780 320 7900
rect 460 7780 780 7900
rect 920 7780 1240 7900
rect 1380 7780 1700 7900
rect 1840 7780 2160 7900
rect 2300 7780 2620 7900
rect 2760 7780 3080 7900
rect 3220 7780 3540 7900
rect 3680 7780 4000 7900
rect 4140 7780 4460 7900
rect 4600 7780 5820 7900
rect 5960 7780 6280 7900
rect 6420 7780 6740 7900
rect 6880 7780 7200 7900
rect 7340 7780 7660 7900
rect 7800 7780 8120 7900
rect 8260 7780 8580 7900
rect 8720 7780 9040 7900
rect 9180 7780 9500 7900
rect 9640 7780 9960 7900
rect 10100 7780 11320 7900
rect 11460 7780 11780 7900
rect 11920 7780 12240 7900
rect 12380 7780 12700 7900
rect 12840 7780 13160 7900
rect 13300 7780 13620 7900
rect 13760 7780 14080 7900
rect 14220 7780 14540 7900
rect 14680 7780 15000 7900
rect 15140 7780 15460 7900
rect 15600 7780 15620 7900
rect 300 7760 15620 7780
rect -1748 -806 13100 -800
rect -1748 -1094 2806 -806
rect 4794 -1094 11106 -806
rect 13094 -1094 13100 -806
rect -1748 -1100 13100 -1094
rect 2500 -1406 15800 -1400
rect 2500 -1694 13806 -1406
rect 15794 -1694 15800 -1406
rect 2500 -1700 15800 -1694
<< via2 >>
rect -910 8100 -510 8200
rect 5000 8100 5400 8200
rect 580 7980 660 8060
rect 1500 7980 1580 8060
rect 2420 7980 2500 8060
rect 3340 7980 3420 8060
rect 4260 7980 4340 8060
rect 10500 8100 10900 8200
rect 6080 7980 6160 8060
rect 7000 7980 7080 8060
rect 7920 7980 8000 8060
rect 8840 7980 8920 8060
rect 9760 7980 9840 8060
rect 16456 8102 16856 8202
rect 11580 7980 11660 8060
rect 12500 7980 12580 8060
rect 13420 7980 13500 8060
rect 14340 7980 14420 8060
rect 15260 7980 15340 8060
<< metal3 >>
rect -1010 8202 16956 8302
rect -1010 8200 16456 8202
rect -1010 8100 -910 8200
rect -510 8100 5000 8200
rect 5400 8100 10500 8200
rect 10900 8102 16456 8200
rect 16856 8102 16956 8202
rect 10900 8100 16956 8102
rect -1010 8060 16956 8100
rect -1010 7980 580 8060
rect 660 7980 1500 8060
rect 1580 7980 2420 8060
rect 2500 7980 3340 8060
rect 3420 7980 4260 8060
rect 4340 7980 6080 8060
rect 6160 7980 7000 8060
rect 7080 7980 7920 8060
rect 8000 7980 8840 8060
rect 8920 7980 9760 8060
rect 9840 7980 11580 8060
rect 11660 7980 12500 8060
rect 12580 7980 13420 8060
rect 13500 7980 14340 8060
rect 14420 7980 15260 8060
rect 15340 7980 16956 8060
rect -1010 7962 16956 7980
rect -1010 7960 16358 7962
use sky130_fd_pr__pfet_01v8_lvt_8QZ6MX  sky130_fd_pr__pfet_01v8_lvt_8QZ6MX_1
timestamp 1621270775
transform 1 0 7955 0 1 3768
box -2355 -3968 2355 3934
use sky130_fd_pr__pfet_01v8_lvt_E8HSF7  sky130_fd_pr__pfet_01v8_lvt_E8HSF7_0
timestamp 1621270775
transform 1 0 2226 0 1 3768
box -2584 -3968 2584 3934
use sky130_fd_pr__pfet_01v8_lvt_E8HSF7  sky130_fd_pr__pfet_01v8_lvt_E8HSF7_1
timestamp 1621270775
transform 1 0 13684 0 1 3768
box -2584 -3968 2584 3934
<< labels >>
rlabel via1 372 7840 418 7884 1 Vgate
port 1 n
rlabel metal3 1094 8122 1228 8240 1 VDD!
port 0 n
flabel metal1 7900 -400 8200 -300 1 FreeSans 1600 0 0 0 Vbg
port 2 n
flabel metal2 7900 -1000 8100 -900 1 FreeSans 1600 0 0 0 Vb
port 4 n
flabel metal2 7900 -1600 8100 -1500 1 FreeSans 1600 0 0 0 Va
port 3 n
<< end >>
