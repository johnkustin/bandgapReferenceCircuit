magic
tech sky130A
magscale 1 2
timestamp 1621288169
<< pwell >>
rect 16568 -11403 26872 -11302
rect 16568 -12489 16669 -11403
rect 17755 -12489 17957 -11403
rect 19043 -12489 19245 -11403
rect 20331 -12489 20533 -11403
rect 21619 -12489 21821 -11403
rect 22907 -12489 23109 -11403
rect 24195 -12489 24397 -11403
rect 25483 -12489 25685 -11403
rect 26771 -12489 26872 -11403
rect 16568 -12691 26872 -12489
rect 16568 -13777 16669 -12691
rect 17755 -13777 17957 -12691
rect 19043 -13777 19245 -12691
rect 20331 -13777 20533 -12691
rect 21619 -13777 21821 -12691
rect 22907 -13777 23109 -12691
rect 24195 -13777 24397 -12691
rect 25483 -13777 25685 -12691
rect 26771 -13777 26872 -12691
rect 16568 -13979 26872 -13777
rect 16568 -15065 16669 -13979
rect 17755 -15065 17957 -13979
rect 19043 -15065 19245 -13979
rect 20331 -15065 20533 -13979
rect 21619 -15065 21821 -13979
rect 22907 -15065 23109 -13979
rect 24195 -15065 24397 -13979
rect 25483 -15065 25685 -13979
rect 26771 -15065 26872 -13979
rect 16568 -15267 26872 -15065
rect 16568 -16353 16669 -15267
rect 17755 -16353 17957 -15267
rect 19043 -16353 19245 -15267
rect 20331 -16353 20533 -15267
rect 21619 -16353 21821 -15267
rect 22907 -16353 23109 -15267
rect 24195 -16353 24397 -15267
rect 25483 -16353 25685 -15267
rect 26771 -16353 26872 -15267
rect 16568 -16555 26872 -16353
rect 16568 -17641 16669 -16555
rect 17755 -17641 17957 -16555
rect 19043 -17641 19245 -16555
rect 20331 -17641 20533 -16555
rect 21619 -17641 21821 -16555
rect 22907 -17641 23109 -16555
rect 24195 -17641 24397 -16555
rect 25483 -17641 25685 -16555
rect 26771 -17641 26872 -16555
rect 16568 -17742 26872 -17641
<< nbase >>
rect 16695 -12463 17729 -11429
rect 17983 -12463 19017 -11429
rect 19271 -12463 20305 -11429
rect 20559 -12463 21593 -11429
rect 21847 -12463 22881 -11429
rect 23135 -12463 24169 -11429
rect 24423 -12463 25457 -11429
rect 25711 -12463 26745 -11429
rect 16695 -13751 17729 -12717
rect 17983 -13751 19017 -12717
rect 19271 -13751 20305 -12717
rect 20559 -13751 21593 -12717
rect 21847 -13751 22881 -12717
rect 23135 -13751 24169 -12717
rect 24423 -13751 25457 -12717
rect 25711 -13751 26745 -12717
rect 16695 -15039 17729 -14005
rect 17983 -15039 19017 -14005
rect 19271 -15039 20305 -14005
rect 20559 -15039 21593 -14005
rect 21847 -15039 22881 -14005
rect 23135 -15039 24169 -14005
rect 24423 -15039 25457 -14005
rect 25711 -15039 26745 -14005
rect 16695 -16327 17729 -15293
rect 17983 -16327 19017 -15293
rect 19271 -16327 20305 -15293
rect 20559 -16327 21593 -15293
rect 21847 -16327 22881 -15293
rect 23135 -16327 24169 -15293
rect 24423 -16327 25457 -15293
rect 25711 -16327 26745 -15293
rect 16695 -17615 17729 -16581
rect 17983 -17615 19017 -16581
rect 19271 -17615 20305 -16581
rect 20559 -17615 21593 -16581
rect 21847 -17615 22881 -16581
rect 23135 -17615 24169 -16581
rect 24423 -17615 25457 -16581
rect 25711 -17615 26745 -16581
<< pdiff >>
rect 16872 -11660 17552 -11606
rect 16872 -11694 16926 -11660
rect 16960 -11694 17016 -11660
rect 17050 -11694 17106 -11660
rect 17140 -11694 17196 -11660
rect 17230 -11694 17286 -11660
rect 17320 -11694 17376 -11660
rect 17410 -11694 17466 -11660
rect 17500 -11694 17552 -11660
rect 16872 -11750 17552 -11694
rect 16872 -11784 16926 -11750
rect 16960 -11784 17016 -11750
rect 17050 -11784 17106 -11750
rect 17140 -11784 17196 -11750
rect 17230 -11784 17286 -11750
rect 17320 -11784 17376 -11750
rect 17410 -11784 17466 -11750
rect 17500 -11784 17552 -11750
rect 16872 -11840 17552 -11784
rect 16872 -11874 16926 -11840
rect 16960 -11874 17016 -11840
rect 17050 -11874 17106 -11840
rect 17140 -11874 17196 -11840
rect 17230 -11874 17286 -11840
rect 17320 -11874 17376 -11840
rect 17410 -11874 17466 -11840
rect 17500 -11874 17552 -11840
rect 16872 -11930 17552 -11874
rect 16872 -11964 16926 -11930
rect 16960 -11964 17016 -11930
rect 17050 -11964 17106 -11930
rect 17140 -11964 17196 -11930
rect 17230 -11964 17286 -11930
rect 17320 -11964 17376 -11930
rect 17410 -11964 17466 -11930
rect 17500 -11964 17552 -11930
rect 16872 -12020 17552 -11964
rect 16872 -12054 16926 -12020
rect 16960 -12054 17016 -12020
rect 17050 -12054 17106 -12020
rect 17140 -12054 17196 -12020
rect 17230 -12054 17286 -12020
rect 17320 -12054 17376 -12020
rect 17410 -12054 17466 -12020
rect 17500 -12054 17552 -12020
rect 16872 -12110 17552 -12054
rect 16872 -12144 16926 -12110
rect 16960 -12144 17016 -12110
rect 17050 -12144 17106 -12110
rect 17140 -12144 17196 -12110
rect 17230 -12144 17286 -12110
rect 17320 -12144 17376 -12110
rect 17410 -12144 17466 -12110
rect 17500 -12144 17552 -12110
rect 16872 -12200 17552 -12144
rect 16872 -12234 16926 -12200
rect 16960 -12234 17016 -12200
rect 17050 -12234 17106 -12200
rect 17140 -12234 17196 -12200
rect 17230 -12234 17286 -12200
rect 17320 -12234 17376 -12200
rect 17410 -12234 17466 -12200
rect 17500 -12234 17552 -12200
rect 16872 -12286 17552 -12234
rect 18160 -11660 18840 -11606
rect 18160 -11694 18214 -11660
rect 18248 -11694 18304 -11660
rect 18338 -11694 18394 -11660
rect 18428 -11694 18484 -11660
rect 18518 -11694 18574 -11660
rect 18608 -11694 18664 -11660
rect 18698 -11694 18754 -11660
rect 18788 -11694 18840 -11660
rect 18160 -11750 18840 -11694
rect 18160 -11784 18214 -11750
rect 18248 -11784 18304 -11750
rect 18338 -11784 18394 -11750
rect 18428 -11784 18484 -11750
rect 18518 -11784 18574 -11750
rect 18608 -11784 18664 -11750
rect 18698 -11784 18754 -11750
rect 18788 -11784 18840 -11750
rect 18160 -11840 18840 -11784
rect 18160 -11874 18214 -11840
rect 18248 -11874 18304 -11840
rect 18338 -11874 18394 -11840
rect 18428 -11874 18484 -11840
rect 18518 -11874 18574 -11840
rect 18608 -11874 18664 -11840
rect 18698 -11874 18754 -11840
rect 18788 -11874 18840 -11840
rect 18160 -11930 18840 -11874
rect 18160 -11964 18214 -11930
rect 18248 -11964 18304 -11930
rect 18338 -11964 18394 -11930
rect 18428 -11964 18484 -11930
rect 18518 -11964 18574 -11930
rect 18608 -11964 18664 -11930
rect 18698 -11964 18754 -11930
rect 18788 -11964 18840 -11930
rect 18160 -12020 18840 -11964
rect 18160 -12054 18214 -12020
rect 18248 -12054 18304 -12020
rect 18338 -12054 18394 -12020
rect 18428 -12054 18484 -12020
rect 18518 -12054 18574 -12020
rect 18608 -12054 18664 -12020
rect 18698 -12054 18754 -12020
rect 18788 -12054 18840 -12020
rect 18160 -12110 18840 -12054
rect 18160 -12144 18214 -12110
rect 18248 -12144 18304 -12110
rect 18338 -12144 18394 -12110
rect 18428 -12144 18484 -12110
rect 18518 -12144 18574 -12110
rect 18608 -12144 18664 -12110
rect 18698 -12144 18754 -12110
rect 18788 -12144 18840 -12110
rect 18160 -12200 18840 -12144
rect 18160 -12234 18214 -12200
rect 18248 -12234 18304 -12200
rect 18338 -12234 18394 -12200
rect 18428 -12234 18484 -12200
rect 18518 -12234 18574 -12200
rect 18608 -12234 18664 -12200
rect 18698 -12234 18754 -12200
rect 18788 -12234 18840 -12200
rect 18160 -12286 18840 -12234
rect 19448 -11660 20128 -11606
rect 19448 -11694 19502 -11660
rect 19536 -11694 19592 -11660
rect 19626 -11694 19682 -11660
rect 19716 -11694 19772 -11660
rect 19806 -11694 19862 -11660
rect 19896 -11694 19952 -11660
rect 19986 -11694 20042 -11660
rect 20076 -11694 20128 -11660
rect 19448 -11750 20128 -11694
rect 19448 -11784 19502 -11750
rect 19536 -11784 19592 -11750
rect 19626 -11784 19682 -11750
rect 19716 -11784 19772 -11750
rect 19806 -11784 19862 -11750
rect 19896 -11784 19952 -11750
rect 19986 -11784 20042 -11750
rect 20076 -11784 20128 -11750
rect 19448 -11840 20128 -11784
rect 19448 -11874 19502 -11840
rect 19536 -11874 19592 -11840
rect 19626 -11874 19682 -11840
rect 19716 -11874 19772 -11840
rect 19806 -11874 19862 -11840
rect 19896 -11874 19952 -11840
rect 19986 -11874 20042 -11840
rect 20076 -11874 20128 -11840
rect 19448 -11930 20128 -11874
rect 19448 -11964 19502 -11930
rect 19536 -11964 19592 -11930
rect 19626 -11964 19682 -11930
rect 19716 -11964 19772 -11930
rect 19806 -11964 19862 -11930
rect 19896 -11964 19952 -11930
rect 19986 -11964 20042 -11930
rect 20076 -11964 20128 -11930
rect 19448 -12020 20128 -11964
rect 19448 -12054 19502 -12020
rect 19536 -12054 19592 -12020
rect 19626 -12054 19682 -12020
rect 19716 -12054 19772 -12020
rect 19806 -12054 19862 -12020
rect 19896 -12054 19952 -12020
rect 19986 -12054 20042 -12020
rect 20076 -12054 20128 -12020
rect 19448 -12110 20128 -12054
rect 19448 -12144 19502 -12110
rect 19536 -12144 19592 -12110
rect 19626 -12144 19682 -12110
rect 19716 -12144 19772 -12110
rect 19806 -12144 19862 -12110
rect 19896 -12144 19952 -12110
rect 19986 -12144 20042 -12110
rect 20076 -12144 20128 -12110
rect 19448 -12200 20128 -12144
rect 19448 -12234 19502 -12200
rect 19536 -12234 19592 -12200
rect 19626 -12234 19682 -12200
rect 19716 -12234 19772 -12200
rect 19806 -12234 19862 -12200
rect 19896 -12234 19952 -12200
rect 19986 -12234 20042 -12200
rect 20076 -12234 20128 -12200
rect 19448 -12286 20128 -12234
rect 20736 -11660 21416 -11606
rect 20736 -11694 20790 -11660
rect 20824 -11694 20880 -11660
rect 20914 -11694 20970 -11660
rect 21004 -11694 21060 -11660
rect 21094 -11694 21150 -11660
rect 21184 -11694 21240 -11660
rect 21274 -11694 21330 -11660
rect 21364 -11694 21416 -11660
rect 20736 -11750 21416 -11694
rect 20736 -11784 20790 -11750
rect 20824 -11784 20880 -11750
rect 20914 -11784 20970 -11750
rect 21004 -11784 21060 -11750
rect 21094 -11784 21150 -11750
rect 21184 -11784 21240 -11750
rect 21274 -11784 21330 -11750
rect 21364 -11784 21416 -11750
rect 20736 -11840 21416 -11784
rect 20736 -11874 20790 -11840
rect 20824 -11874 20880 -11840
rect 20914 -11874 20970 -11840
rect 21004 -11874 21060 -11840
rect 21094 -11874 21150 -11840
rect 21184 -11874 21240 -11840
rect 21274 -11874 21330 -11840
rect 21364 -11874 21416 -11840
rect 20736 -11930 21416 -11874
rect 20736 -11964 20790 -11930
rect 20824 -11964 20880 -11930
rect 20914 -11964 20970 -11930
rect 21004 -11964 21060 -11930
rect 21094 -11964 21150 -11930
rect 21184 -11964 21240 -11930
rect 21274 -11964 21330 -11930
rect 21364 -11964 21416 -11930
rect 20736 -12020 21416 -11964
rect 20736 -12054 20790 -12020
rect 20824 -12054 20880 -12020
rect 20914 -12054 20970 -12020
rect 21004 -12054 21060 -12020
rect 21094 -12054 21150 -12020
rect 21184 -12054 21240 -12020
rect 21274 -12054 21330 -12020
rect 21364 -12054 21416 -12020
rect 20736 -12110 21416 -12054
rect 20736 -12144 20790 -12110
rect 20824 -12144 20880 -12110
rect 20914 -12144 20970 -12110
rect 21004 -12144 21060 -12110
rect 21094 -12144 21150 -12110
rect 21184 -12144 21240 -12110
rect 21274 -12144 21330 -12110
rect 21364 -12144 21416 -12110
rect 20736 -12200 21416 -12144
rect 20736 -12234 20790 -12200
rect 20824 -12234 20880 -12200
rect 20914 -12234 20970 -12200
rect 21004 -12234 21060 -12200
rect 21094 -12234 21150 -12200
rect 21184 -12234 21240 -12200
rect 21274 -12234 21330 -12200
rect 21364 -12234 21416 -12200
rect 20736 -12286 21416 -12234
rect 22024 -11660 22704 -11606
rect 22024 -11694 22078 -11660
rect 22112 -11694 22168 -11660
rect 22202 -11694 22258 -11660
rect 22292 -11694 22348 -11660
rect 22382 -11694 22438 -11660
rect 22472 -11694 22528 -11660
rect 22562 -11694 22618 -11660
rect 22652 -11694 22704 -11660
rect 22024 -11750 22704 -11694
rect 22024 -11784 22078 -11750
rect 22112 -11784 22168 -11750
rect 22202 -11784 22258 -11750
rect 22292 -11784 22348 -11750
rect 22382 -11784 22438 -11750
rect 22472 -11784 22528 -11750
rect 22562 -11784 22618 -11750
rect 22652 -11784 22704 -11750
rect 22024 -11840 22704 -11784
rect 22024 -11874 22078 -11840
rect 22112 -11874 22168 -11840
rect 22202 -11874 22258 -11840
rect 22292 -11874 22348 -11840
rect 22382 -11874 22438 -11840
rect 22472 -11874 22528 -11840
rect 22562 -11874 22618 -11840
rect 22652 -11874 22704 -11840
rect 22024 -11930 22704 -11874
rect 22024 -11964 22078 -11930
rect 22112 -11964 22168 -11930
rect 22202 -11964 22258 -11930
rect 22292 -11964 22348 -11930
rect 22382 -11964 22438 -11930
rect 22472 -11964 22528 -11930
rect 22562 -11964 22618 -11930
rect 22652 -11964 22704 -11930
rect 22024 -12020 22704 -11964
rect 22024 -12054 22078 -12020
rect 22112 -12054 22168 -12020
rect 22202 -12054 22258 -12020
rect 22292 -12054 22348 -12020
rect 22382 -12054 22438 -12020
rect 22472 -12054 22528 -12020
rect 22562 -12054 22618 -12020
rect 22652 -12054 22704 -12020
rect 22024 -12110 22704 -12054
rect 22024 -12144 22078 -12110
rect 22112 -12144 22168 -12110
rect 22202 -12144 22258 -12110
rect 22292 -12144 22348 -12110
rect 22382 -12144 22438 -12110
rect 22472 -12144 22528 -12110
rect 22562 -12144 22618 -12110
rect 22652 -12144 22704 -12110
rect 22024 -12200 22704 -12144
rect 22024 -12234 22078 -12200
rect 22112 -12234 22168 -12200
rect 22202 -12234 22258 -12200
rect 22292 -12234 22348 -12200
rect 22382 -12234 22438 -12200
rect 22472 -12234 22528 -12200
rect 22562 -12234 22618 -12200
rect 22652 -12234 22704 -12200
rect 22024 -12286 22704 -12234
rect 23312 -11660 23992 -11606
rect 23312 -11694 23366 -11660
rect 23400 -11694 23456 -11660
rect 23490 -11694 23546 -11660
rect 23580 -11694 23636 -11660
rect 23670 -11694 23726 -11660
rect 23760 -11694 23816 -11660
rect 23850 -11694 23906 -11660
rect 23940 -11694 23992 -11660
rect 23312 -11750 23992 -11694
rect 23312 -11784 23366 -11750
rect 23400 -11784 23456 -11750
rect 23490 -11784 23546 -11750
rect 23580 -11784 23636 -11750
rect 23670 -11784 23726 -11750
rect 23760 -11784 23816 -11750
rect 23850 -11784 23906 -11750
rect 23940 -11784 23992 -11750
rect 23312 -11840 23992 -11784
rect 23312 -11874 23366 -11840
rect 23400 -11874 23456 -11840
rect 23490 -11874 23546 -11840
rect 23580 -11874 23636 -11840
rect 23670 -11874 23726 -11840
rect 23760 -11874 23816 -11840
rect 23850 -11874 23906 -11840
rect 23940 -11874 23992 -11840
rect 23312 -11930 23992 -11874
rect 23312 -11964 23366 -11930
rect 23400 -11964 23456 -11930
rect 23490 -11964 23546 -11930
rect 23580 -11964 23636 -11930
rect 23670 -11964 23726 -11930
rect 23760 -11964 23816 -11930
rect 23850 -11964 23906 -11930
rect 23940 -11964 23992 -11930
rect 23312 -12020 23992 -11964
rect 23312 -12054 23366 -12020
rect 23400 -12054 23456 -12020
rect 23490 -12054 23546 -12020
rect 23580 -12054 23636 -12020
rect 23670 -12054 23726 -12020
rect 23760 -12054 23816 -12020
rect 23850 -12054 23906 -12020
rect 23940 -12054 23992 -12020
rect 23312 -12110 23992 -12054
rect 23312 -12144 23366 -12110
rect 23400 -12144 23456 -12110
rect 23490 -12144 23546 -12110
rect 23580 -12144 23636 -12110
rect 23670 -12144 23726 -12110
rect 23760 -12144 23816 -12110
rect 23850 -12144 23906 -12110
rect 23940 -12144 23992 -12110
rect 23312 -12200 23992 -12144
rect 23312 -12234 23366 -12200
rect 23400 -12234 23456 -12200
rect 23490 -12234 23546 -12200
rect 23580 -12234 23636 -12200
rect 23670 -12234 23726 -12200
rect 23760 -12234 23816 -12200
rect 23850 -12234 23906 -12200
rect 23940 -12234 23992 -12200
rect 23312 -12286 23992 -12234
rect 24600 -11660 25280 -11606
rect 24600 -11694 24654 -11660
rect 24688 -11694 24744 -11660
rect 24778 -11694 24834 -11660
rect 24868 -11694 24924 -11660
rect 24958 -11694 25014 -11660
rect 25048 -11694 25104 -11660
rect 25138 -11694 25194 -11660
rect 25228 -11694 25280 -11660
rect 24600 -11750 25280 -11694
rect 24600 -11784 24654 -11750
rect 24688 -11784 24744 -11750
rect 24778 -11784 24834 -11750
rect 24868 -11784 24924 -11750
rect 24958 -11784 25014 -11750
rect 25048 -11784 25104 -11750
rect 25138 -11784 25194 -11750
rect 25228 -11784 25280 -11750
rect 24600 -11840 25280 -11784
rect 24600 -11874 24654 -11840
rect 24688 -11874 24744 -11840
rect 24778 -11874 24834 -11840
rect 24868 -11874 24924 -11840
rect 24958 -11874 25014 -11840
rect 25048 -11874 25104 -11840
rect 25138 -11874 25194 -11840
rect 25228 -11874 25280 -11840
rect 24600 -11930 25280 -11874
rect 24600 -11964 24654 -11930
rect 24688 -11964 24744 -11930
rect 24778 -11964 24834 -11930
rect 24868 -11964 24924 -11930
rect 24958 -11964 25014 -11930
rect 25048 -11964 25104 -11930
rect 25138 -11964 25194 -11930
rect 25228 -11964 25280 -11930
rect 24600 -12020 25280 -11964
rect 24600 -12054 24654 -12020
rect 24688 -12054 24744 -12020
rect 24778 -12054 24834 -12020
rect 24868 -12054 24924 -12020
rect 24958 -12054 25014 -12020
rect 25048 -12054 25104 -12020
rect 25138 -12054 25194 -12020
rect 25228 -12054 25280 -12020
rect 24600 -12110 25280 -12054
rect 24600 -12144 24654 -12110
rect 24688 -12144 24744 -12110
rect 24778 -12144 24834 -12110
rect 24868 -12144 24924 -12110
rect 24958 -12144 25014 -12110
rect 25048 -12144 25104 -12110
rect 25138 -12144 25194 -12110
rect 25228 -12144 25280 -12110
rect 24600 -12200 25280 -12144
rect 24600 -12234 24654 -12200
rect 24688 -12234 24744 -12200
rect 24778 -12234 24834 -12200
rect 24868 -12234 24924 -12200
rect 24958 -12234 25014 -12200
rect 25048 -12234 25104 -12200
rect 25138 -12234 25194 -12200
rect 25228 -12234 25280 -12200
rect 24600 -12286 25280 -12234
rect 25888 -11660 26568 -11606
rect 25888 -11694 25942 -11660
rect 25976 -11694 26032 -11660
rect 26066 -11694 26122 -11660
rect 26156 -11694 26212 -11660
rect 26246 -11694 26302 -11660
rect 26336 -11694 26392 -11660
rect 26426 -11694 26482 -11660
rect 26516 -11694 26568 -11660
rect 25888 -11750 26568 -11694
rect 25888 -11784 25942 -11750
rect 25976 -11784 26032 -11750
rect 26066 -11784 26122 -11750
rect 26156 -11784 26212 -11750
rect 26246 -11784 26302 -11750
rect 26336 -11784 26392 -11750
rect 26426 -11784 26482 -11750
rect 26516 -11784 26568 -11750
rect 25888 -11840 26568 -11784
rect 25888 -11874 25942 -11840
rect 25976 -11874 26032 -11840
rect 26066 -11874 26122 -11840
rect 26156 -11874 26212 -11840
rect 26246 -11874 26302 -11840
rect 26336 -11874 26392 -11840
rect 26426 -11874 26482 -11840
rect 26516 -11874 26568 -11840
rect 25888 -11930 26568 -11874
rect 25888 -11964 25942 -11930
rect 25976 -11964 26032 -11930
rect 26066 -11964 26122 -11930
rect 26156 -11964 26212 -11930
rect 26246 -11964 26302 -11930
rect 26336 -11964 26392 -11930
rect 26426 -11964 26482 -11930
rect 26516 -11964 26568 -11930
rect 25888 -12020 26568 -11964
rect 25888 -12054 25942 -12020
rect 25976 -12054 26032 -12020
rect 26066 -12054 26122 -12020
rect 26156 -12054 26212 -12020
rect 26246 -12054 26302 -12020
rect 26336 -12054 26392 -12020
rect 26426 -12054 26482 -12020
rect 26516 -12054 26568 -12020
rect 25888 -12110 26568 -12054
rect 25888 -12144 25942 -12110
rect 25976 -12144 26032 -12110
rect 26066 -12144 26122 -12110
rect 26156 -12144 26212 -12110
rect 26246 -12144 26302 -12110
rect 26336 -12144 26392 -12110
rect 26426 -12144 26482 -12110
rect 26516 -12144 26568 -12110
rect 25888 -12200 26568 -12144
rect 25888 -12234 25942 -12200
rect 25976 -12234 26032 -12200
rect 26066 -12234 26122 -12200
rect 26156 -12234 26212 -12200
rect 26246 -12234 26302 -12200
rect 26336 -12234 26392 -12200
rect 26426 -12234 26482 -12200
rect 26516 -12234 26568 -12200
rect 25888 -12286 26568 -12234
rect 16872 -12948 17552 -12894
rect 16872 -12982 16926 -12948
rect 16960 -12982 17016 -12948
rect 17050 -12982 17106 -12948
rect 17140 -12982 17196 -12948
rect 17230 -12982 17286 -12948
rect 17320 -12982 17376 -12948
rect 17410 -12982 17466 -12948
rect 17500 -12982 17552 -12948
rect 16872 -13038 17552 -12982
rect 16872 -13072 16926 -13038
rect 16960 -13072 17016 -13038
rect 17050 -13072 17106 -13038
rect 17140 -13072 17196 -13038
rect 17230 -13072 17286 -13038
rect 17320 -13072 17376 -13038
rect 17410 -13072 17466 -13038
rect 17500 -13072 17552 -13038
rect 16872 -13128 17552 -13072
rect 16872 -13162 16926 -13128
rect 16960 -13162 17016 -13128
rect 17050 -13162 17106 -13128
rect 17140 -13162 17196 -13128
rect 17230 -13162 17286 -13128
rect 17320 -13162 17376 -13128
rect 17410 -13162 17466 -13128
rect 17500 -13162 17552 -13128
rect 16872 -13218 17552 -13162
rect 16872 -13252 16926 -13218
rect 16960 -13252 17016 -13218
rect 17050 -13252 17106 -13218
rect 17140 -13252 17196 -13218
rect 17230 -13252 17286 -13218
rect 17320 -13252 17376 -13218
rect 17410 -13252 17466 -13218
rect 17500 -13252 17552 -13218
rect 16872 -13308 17552 -13252
rect 16872 -13342 16926 -13308
rect 16960 -13342 17016 -13308
rect 17050 -13342 17106 -13308
rect 17140 -13342 17196 -13308
rect 17230 -13342 17286 -13308
rect 17320 -13342 17376 -13308
rect 17410 -13342 17466 -13308
rect 17500 -13342 17552 -13308
rect 16872 -13398 17552 -13342
rect 16872 -13432 16926 -13398
rect 16960 -13432 17016 -13398
rect 17050 -13432 17106 -13398
rect 17140 -13432 17196 -13398
rect 17230 -13432 17286 -13398
rect 17320 -13432 17376 -13398
rect 17410 -13432 17466 -13398
rect 17500 -13432 17552 -13398
rect 16872 -13488 17552 -13432
rect 16872 -13522 16926 -13488
rect 16960 -13522 17016 -13488
rect 17050 -13522 17106 -13488
rect 17140 -13522 17196 -13488
rect 17230 -13522 17286 -13488
rect 17320 -13522 17376 -13488
rect 17410 -13522 17466 -13488
rect 17500 -13522 17552 -13488
rect 16872 -13574 17552 -13522
rect 18160 -12948 18840 -12894
rect 18160 -12982 18214 -12948
rect 18248 -12982 18304 -12948
rect 18338 -12982 18394 -12948
rect 18428 -12982 18484 -12948
rect 18518 -12982 18574 -12948
rect 18608 -12982 18664 -12948
rect 18698 -12982 18754 -12948
rect 18788 -12982 18840 -12948
rect 18160 -13038 18840 -12982
rect 18160 -13072 18214 -13038
rect 18248 -13072 18304 -13038
rect 18338 -13072 18394 -13038
rect 18428 -13072 18484 -13038
rect 18518 -13072 18574 -13038
rect 18608 -13072 18664 -13038
rect 18698 -13072 18754 -13038
rect 18788 -13072 18840 -13038
rect 18160 -13128 18840 -13072
rect 18160 -13162 18214 -13128
rect 18248 -13162 18304 -13128
rect 18338 -13162 18394 -13128
rect 18428 -13162 18484 -13128
rect 18518 -13162 18574 -13128
rect 18608 -13162 18664 -13128
rect 18698 -13162 18754 -13128
rect 18788 -13162 18840 -13128
rect 18160 -13218 18840 -13162
rect 18160 -13252 18214 -13218
rect 18248 -13252 18304 -13218
rect 18338 -13252 18394 -13218
rect 18428 -13252 18484 -13218
rect 18518 -13252 18574 -13218
rect 18608 -13252 18664 -13218
rect 18698 -13252 18754 -13218
rect 18788 -13252 18840 -13218
rect 18160 -13308 18840 -13252
rect 18160 -13342 18214 -13308
rect 18248 -13342 18304 -13308
rect 18338 -13342 18394 -13308
rect 18428 -13342 18484 -13308
rect 18518 -13342 18574 -13308
rect 18608 -13342 18664 -13308
rect 18698 -13342 18754 -13308
rect 18788 -13342 18840 -13308
rect 18160 -13398 18840 -13342
rect 18160 -13432 18214 -13398
rect 18248 -13432 18304 -13398
rect 18338 -13432 18394 -13398
rect 18428 -13432 18484 -13398
rect 18518 -13432 18574 -13398
rect 18608 -13432 18664 -13398
rect 18698 -13432 18754 -13398
rect 18788 -13432 18840 -13398
rect 18160 -13488 18840 -13432
rect 18160 -13522 18214 -13488
rect 18248 -13522 18304 -13488
rect 18338 -13522 18394 -13488
rect 18428 -13522 18484 -13488
rect 18518 -13522 18574 -13488
rect 18608 -13522 18664 -13488
rect 18698 -13522 18754 -13488
rect 18788 -13522 18840 -13488
rect 18160 -13574 18840 -13522
rect 19448 -12948 20128 -12894
rect 19448 -12982 19502 -12948
rect 19536 -12982 19592 -12948
rect 19626 -12982 19682 -12948
rect 19716 -12982 19772 -12948
rect 19806 -12982 19862 -12948
rect 19896 -12982 19952 -12948
rect 19986 -12982 20042 -12948
rect 20076 -12982 20128 -12948
rect 19448 -13038 20128 -12982
rect 19448 -13072 19502 -13038
rect 19536 -13072 19592 -13038
rect 19626 -13072 19682 -13038
rect 19716 -13072 19772 -13038
rect 19806 -13072 19862 -13038
rect 19896 -13072 19952 -13038
rect 19986 -13072 20042 -13038
rect 20076 -13072 20128 -13038
rect 19448 -13128 20128 -13072
rect 19448 -13162 19502 -13128
rect 19536 -13162 19592 -13128
rect 19626 -13162 19682 -13128
rect 19716 -13162 19772 -13128
rect 19806 -13162 19862 -13128
rect 19896 -13162 19952 -13128
rect 19986 -13162 20042 -13128
rect 20076 -13162 20128 -13128
rect 19448 -13218 20128 -13162
rect 19448 -13252 19502 -13218
rect 19536 -13252 19592 -13218
rect 19626 -13252 19682 -13218
rect 19716 -13252 19772 -13218
rect 19806 -13252 19862 -13218
rect 19896 -13252 19952 -13218
rect 19986 -13252 20042 -13218
rect 20076 -13252 20128 -13218
rect 19448 -13308 20128 -13252
rect 19448 -13342 19502 -13308
rect 19536 -13342 19592 -13308
rect 19626 -13342 19682 -13308
rect 19716 -13342 19772 -13308
rect 19806 -13342 19862 -13308
rect 19896 -13342 19952 -13308
rect 19986 -13342 20042 -13308
rect 20076 -13342 20128 -13308
rect 19448 -13398 20128 -13342
rect 19448 -13432 19502 -13398
rect 19536 -13432 19592 -13398
rect 19626 -13432 19682 -13398
rect 19716 -13432 19772 -13398
rect 19806 -13432 19862 -13398
rect 19896 -13432 19952 -13398
rect 19986 -13432 20042 -13398
rect 20076 -13432 20128 -13398
rect 19448 -13488 20128 -13432
rect 19448 -13522 19502 -13488
rect 19536 -13522 19592 -13488
rect 19626 -13522 19682 -13488
rect 19716 -13522 19772 -13488
rect 19806 -13522 19862 -13488
rect 19896 -13522 19952 -13488
rect 19986 -13522 20042 -13488
rect 20076 -13522 20128 -13488
rect 19448 -13574 20128 -13522
rect 20736 -12948 21416 -12894
rect 20736 -12982 20790 -12948
rect 20824 -12982 20880 -12948
rect 20914 -12982 20970 -12948
rect 21004 -12982 21060 -12948
rect 21094 -12982 21150 -12948
rect 21184 -12982 21240 -12948
rect 21274 -12982 21330 -12948
rect 21364 -12982 21416 -12948
rect 20736 -13038 21416 -12982
rect 20736 -13072 20790 -13038
rect 20824 -13072 20880 -13038
rect 20914 -13072 20970 -13038
rect 21004 -13072 21060 -13038
rect 21094 -13072 21150 -13038
rect 21184 -13072 21240 -13038
rect 21274 -13072 21330 -13038
rect 21364 -13072 21416 -13038
rect 20736 -13128 21416 -13072
rect 20736 -13162 20790 -13128
rect 20824 -13162 20880 -13128
rect 20914 -13162 20970 -13128
rect 21004 -13162 21060 -13128
rect 21094 -13162 21150 -13128
rect 21184 -13162 21240 -13128
rect 21274 -13162 21330 -13128
rect 21364 -13162 21416 -13128
rect 20736 -13218 21416 -13162
rect 20736 -13252 20790 -13218
rect 20824 -13252 20880 -13218
rect 20914 -13252 20970 -13218
rect 21004 -13252 21060 -13218
rect 21094 -13252 21150 -13218
rect 21184 -13252 21240 -13218
rect 21274 -13252 21330 -13218
rect 21364 -13252 21416 -13218
rect 20736 -13308 21416 -13252
rect 20736 -13342 20790 -13308
rect 20824 -13342 20880 -13308
rect 20914 -13342 20970 -13308
rect 21004 -13342 21060 -13308
rect 21094 -13342 21150 -13308
rect 21184 -13342 21240 -13308
rect 21274 -13342 21330 -13308
rect 21364 -13342 21416 -13308
rect 20736 -13398 21416 -13342
rect 20736 -13432 20790 -13398
rect 20824 -13432 20880 -13398
rect 20914 -13432 20970 -13398
rect 21004 -13432 21060 -13398
rect 21094 -13432 21150 -13398
rect 21184 -13432 21240 -13398
rect 21274 -13432 21330 -13398
rect 21364 -13432 21416 -13398
rect 20736 -13488 21416 -13432
rect 20736 -13522 20790 -13488
rect 20824 -13522 20880 -13488
rect 20914 -13522 20970 -13488
rect 21004 -13522 21060 -13488
rect 21094 -13522 21150 -13488
rect 21184 -13522 21240 -13488
rect 21274 -13522 21330 -13488
rect 21364 -13522 21416 -13488
rect 20736 -13574 21416 -13522
rect 22024 -12948 22704 -12894
rect 22024 -12982 22078 -12948
rect 22112 -12982 22168 -12948
rect 22202 -12982 22258 -12948
rect 22292 -12982 22348 -12948
rect 22382 -12982 22438 -12948
rect 22472 -12982 22528 -12948
rect 22562 -12982 22618 -12948
rect 22652 -12982 22704 -12948
rect 22024 -13038 22704 -12982
rect 22024 -13072 22078 -13038
rect 22112 -13072 22168 -13038
rect 22202 -13072 22258 -13038
rect 22292 -13072 22348 -13038
rect 22382 -13072 22438 -13038
rect 22472 -13072 22528 -13038
rect 22562 -13072 22618 -13038
rect 22652 -13072 22704 -13038
rect 22024 -13128 22704 -13072
rect 22024 -13162 22078 -13128
rect 22112 -13162 22168 -13128
rect 22202 -13162 22258 -13128
rect 22292 -13162 22348 -13128
rect 22382 -13162 22438 -13128
rect 22472 -13162 22528 -13128
rect 22562 -13162 22618 -13128
rect 22652 -13162 22704 -13128
rect 22024 -13218 22704 -13162
rect 22024 -13252 22078 -13218
rect 22112 -13252 22168 -13218
rect 22202 -13252 22258 -13218
rect 22292 -13252 22348 -13218
rect 22382 -13252 22438 -13218
rect 22472 -13252 22528 -13218
rect 22562 -13252 22618 -13218
rect 22652 -13252 22704 -13218
rect 22024 -13308 22704 -13252
rect 22024 -13342 22078 -13308
rect 22112 -13342 22168 -13308
rect 22202 -13342 22258 -13308
rect 22292 -13342 22348 -13308
rect 22382 -13342 22438 -13308
rect 22472 -13342 22528 -13308
rect 22562 -13342 22618 -13308
rect 22652 -13342 22704 -13308
rect 22024 -13398 22704 -13342
rect 22024 -13432 22078 -13398
rect 22112 -13432 22168 -13398
rect 22202 -13432 22258 -13398
rect 22292 -13432 22348 -13398
rect 22382 -13432 22438 -13398
rect 22472 -13432 22528 -13398
rect 22562 -13432 22618 -13398
rect 22652 -13432 22704 -13398
rect 22024 -13488 22704 -13432
rect 22024 -13522 22078 -13488
rect 22112 -13522 22168 -13488
rect 22202 -13522 22258 -13488
rect 22292 -13522 22348 -13488
rect 22382 -13522 22438 -13488
rect 22472 -13522 22528 -13488
rect 22562 -13522 22618 -13488
rect 22652 -13522 22704 -13488
rect 22024 -13574 22704 -13522
rect 23312 -12948 23992 -12894
rect 23312 -12982 23366 -12948
rect 23400 -12982 23456 -12948
rect 23490 -12982 23546 -12948
rect 23580 -12982 23636 -12948
rect 23670 -12982 23726 -12948
rect 23760 -12982 23816 -12948
rect 23850 -12982 23906 -12948
rect 23940 -12982 23992 -12948
rect 23312 -13038 23992 -12982
rect 23312 -13072 23366 -13038
rect 23400 -13072 23456 -13038
rect 23490 -13072 23546 -13038
rect 23580 -13072 23636 -13038
rect 23670 -13072 23726 -13038
rect 23760 -13072 23816 -13038
rect 23850 -13072 23906 -13038
rect 23940 -13072 23992 -13038
rect 23312 -13128 23992 -13072
rect 23312 -13162 23366 -13128
rect 23400 -13162 23456 -13128
rect 23490 -13162 23546 -13128
rect 23580 -13162 23636 -13128
rect 23670 -13162 23726 -13128
rect 23760 -13162 23816 -13128
rect 23850 -13162 23906 -13128
rect 23940 -13162 23992 -13128
rect 23312 -13218 23992 -13162
rect 23312 -13252 23366 -13218
rect 23400 -13252 23456 -13218
rect 23490 -13252 23546 -13218
rect 23580 -13252 23636 -13218
rect 23670 -13252 23726 -13218
rect 23760 -13252 23816 -13218
rect 23850 -13252 23906 -13218
rect 23940 -13252 23992 -13218
rect 23312 -13308 23992 -13252
rect 23312 -13342 23366 -13308
rect 23400 -13342 23456 -13308
rect 23490 -13342 23546 -13308
rect 23580 -13342 23636 -13308
rect 23670 -13342 23726 -13308
rect 23760 -13342 23816 -13308
rect 23850 -13342 23906 -13308
rect 23940 -13342 23992 -13308
rect 23312 -13398 23992 -13342
rect 23312 -13432 23366 -13398
rect 23400 -13432 23456 -13398
rect 23490 -13432 23546 -13398
rect 23580 -13432 23636 -13398
rect 23670 -13432 23726 -13398
rect 23760 -13432 23816 -13398
rect 23850 -13432 23906 -13398
rect 23940 -13432 23992 -13398
rect 23312 -13488 23992 -13432
rect 23312 -13522 23366 -13488
rect 23400 -13522 23456 -13488
rect 23490 -13522 23546 -13488
rect 23580 -13522 23636 -13488
rect 23670 -13522 23726 -13488
rect 23760 -13522 23816 -13488
rect 23850 -13522 23906 -13488
rect 23940 -13522 23992 -13488
rect 23312 -13574 23992 -13522
rect 24600 -12948 25280 -12894
rect 24600 -12982 24654 -12948
rect 24688 -12982 24744 -12948
rect 24778 -12982 24834 -12948
rect 24868 -12982 24924 -12948
rect 24958 -12982 25014 -12948
rect 25048 -12982 25104 -12948
rect 25138 -12982 25194 -12948
rect 25228 -12982 25280 -12948
rect 24600 -13038 25280 -12982
rect 24600 -13072 24654 -13038
rect 24688 -13072 24744 -13038
rect 24778 -13072 24834 -13038
rect 24868 -13072 24924 -13038
rect 24958 -13072 25014 -13038
rect 25048 -13072 25104 -13038
rect 25138 -13072 25194 -13038
rect 25228 -13072 25280 -13038
rect 24600 -13128 25280 -13072
rect 24600 -13162 24654 -13128
rect 24688 -13162 24744 -13128
rect 24778 -13162 24834 -13128
rect 24868 -13162 24924 -13128
rect 24958 -13162 25014 -13128
rect 25048 -13162 25104 -13128
rect 25138 -13162 25194 -13128
rect 25228 -13162 25280 -13128
rect 24600 -13218 25280 -13162
rect 24600 -13252 24654 -13218
rect 24688 -13252 24744 -13218
rect 24778 -13252 24834 -13218
rect 24868 -13252 24924 -13218
rect 24958 -13252 25014 -13218
rect 25048 -13252 25104 -13218
rect 25138 -13252 25194 -13218
rect 25228 -13252 25280 -13218
rect 24600 -13308 25280 -13252
rect 24600 -13342 24654 -13308
rect 24688 -13342 24744 -13308
rect 24778 -13342 24834 -13308
rect 24868 -13342 24924 -13308
rect 24958 -13342 25014 -13308
rect 25048 -13342 25104 -13308
rect 25138 -13342 25194 -13308
rect 25228 -13342 25280 -13308
rect 24600 -13398 25280 -13342
rect 24600 -13432 24654 -13398
rect 24688 -13432 24744 -13398
rect 24778 -13432 24834 -13398
rect 24868 -13432 24924 -13398
rect 24958 -13432 25014 -13398
rect 25048 -13432 25104 -13398
rect 25138 -13432 25194 -13398
rect 25228 -13432 25280 -13398
rect 24600 -13488 25280 -13432
rect 24600 -13522 24654 -13488
rect 24688 -13522 24744 -13488
rect 24778 -13522 24834 -13488
rect 24868 -13522 24924 -13488
rect 24958 -13522 25014 -13488
rect 25048 -13522 25104 -13488
rect 25138 -13522 25194 -13488
rect 25228 -13522 25280 -13488
rect 24600 -13574 25280 -13522
rect 25888 -12948 26568 -12894
rect 25888 -12982 25942 -12948
rect 25976 -12982 26032 -12948
rect 26066 -12982 26122 -12948
rect 26156 -12982 26212 -12948
rect 26246 -12982 26302 -12948
rect 26336 -12982 26392 -12948
rect 26426 -12982 26482 -12948
rect 26516 -12982 26568 -12948
rect 25888 -13038 26568 -12982
rect 25888 -13072 25942 -13038
rect 25976 -13072 26032 -13038
rect 26066 -13072 26122 -13038
rect 26156 -13072 26212 -13038
rect 26246 -13072 26302 -13038
rect 26336 -13072 26392 -13038
rect 26426 -13072 26482 -13038
rect 26516 -13072 26568 -13038
rect 25888 -13128 26568 -13072
rect 25888 -13162 25942 -13128
rect 25976 -13162 26032 -13128
rect 26066 -13162 26122 -13128
rect 26156 -13162 26212 -13128
rect 26246 -13162 26302 -13128
rect 26336 -13162 26392 -13128
rect 26426 -13162 26482 -13128
rect 26516 -13162 26568 -13128
rect 25888 -13218 26568 -13162
rect 25888 -13252 25942 -13218
rect 25976 -13252 26032 -13218
rect 26066 -13252 26122 -13218
rect 26156 -13252 26212 -13218
rect 26246 -13252 26302 -13218
rect 26336 -13252 26392 -13218
rect 26426 -13252 26482 -13218
rect 26516 -13252 26568 -13218
rect 25888 -13308 26568 -13252
rect 25888 -13342 25942 -13308
rect 25976 -13342 26032 -13308
rect 26066 -13342 26122 -13308
rect 26156 -13342 26212 -13308
rect 26246 -13342 26302 -13308
rect 26336 -13342 26392 -13308
rect 26426 -13342 26482 -13308
rect 26516 -13342 26568 -13308
rect 25888 -13398 26568 -13342
rect 25888 -13432 25942 -13398
rect 25976 -13432 26032 -13398
rect 26066 -13432 26122 -13398
rect 26156 -13432 26212 -13398
rect 26246 -13432 26302 -13398
rect 26336 -13432 26392 -13398
rect 26426 -13432 26482 -13398
rect 26516 -13432 26568 -13398
rect 25888 -13488 26568 -13432
rect 25888 -13522 25942 -13488
rect 25976 -13522 26032 -13488
rect 26066 -13522 26122 -13488
rect 26156 -13522 26212 -13488
rect 26246 -13522 26302 -13488
rect 26336 -13522 26392 -13488
rect 26426 -13522 26482 -13488
rect 26516 -13522 26568 -13488
rect 25888 -13574 26568 -13522
rect 16872 -14236 17552 -14182
rect 16872 -14270 16926 -14236
rect 16960 -14270 17016 -14236
rect 17050 -14270 17106 -14236
rect 17140 -14270 17196 -14236
rect 17230 -14270 17286 -14236
rect 17320 -14270 17376 -14236
rect 17410 -14270 17466 -14236
rect 17500 -14270 17552 -14236
rect 16872 -14326 17552 -14270
rect 16872 -14360 16926 -14326
rect 16960 -14360 17016 -14326
rect 17050 -14360 17106 -14326
rect 17140 -14360 17196 -14326
rect 17230 -14360 17286 -14326
rect 17320 -14360 17376 -14326
rect 17410 -14360 17466 -14326
rect 17500 -14360 17552 -14326
rect 16872 -14416 17552 -14360
rect 16872 -14450 16926 -14416
rect 16960 -14450 17016 -14416
rect 17050 -14450 17106 -14416
rect 17140 -14450 17196 -14416
rect 17230 -14450 17286 -14416
rect 17320 -14450 17376 -14416
rect 17410 -14450 17466 -14416
rect 17500 -14450 17552 -14416
rect 16872 -14506 17552 -14450
rect 16872 -14540 16926 -14506
rect 16960 -14540 17016 -14506
rect 17050 -14540 17106 -14506
rect 17140 -14540 17196 -14506
rect 17230 -14540 17286 -14506
rect 17320 -14540 17376 -14506
rect 17410 -14540 17466 -14506
rect 17500 -14540 17552 -14506
rect 16872 -14596 17552 -14540
rect 16872 -14630 16926 -14596
rect 16960 -14630 17016 -14596
rect 17050 -14630 17106 -14596
rect 17140 -14630 17196 -14596
rect 17230 -14630 17286 -14596
rect 17320 -14630 17376 -14596
rect 17410 -14630 17466 -14596
rect 17500 -14630 17552 -14596
rect 16872 -14686 17552 -14630
rect 16872 -14720 16926 -14686
rect 16960 -14720 17016 -14686
rect 17050 -14720 17106 -14686
rect 17140 -14720 17196 -14686
rect 17230 -14720 17286 -14686
rect 17320 -14720 17376 -14686
rect 17410 -14720 17466 -14686
rect 17500 -14720 17552 -14686
rect 16872 -14776 17552 -14720
rect 16872 -14810 16926 -14776
rect 16960 -14810 17016 -14776
rect 17050 -14810 17106 -14776
rect 17140 -14810 17196 -14776
rect 17230 -14810 17286 -14776
rect 17320 -14810 17376 -14776
rect 17410 -14810 17466 -14776
rect 17500 -14810 17552 -14776
rect 16872 -14862 17552 -14810
rect 18160 -14236 18840 -14182
rect 18160 -14270 18214 -14236
rect 18248 -14270 18304 -14236
rect 18338 -14270 18394 -14236
rect 18428 -14270 18484 -14236
rect 18518 -14270 18574 -14236
rect 18608 -14270 18664 -14236
rect 18698 -14270 18754 -14236
rect 18788 -14270 18840 -14236
rect 18160 -14326 18840 -14270
rect 18160 -14360 18214 -14326
rect 18248 -14360 18304 -14326
rect 18338 -14360 18394 -14326
rect 18428 -14360 18484 -14326
rect 18518 -14360 18574 -14326
rect 18608 -14360 18664 -14326
rect 18698 -14360 18754 -14326
rect 18788 -14360 18840 -14326
rect 18160 -14416 18840 -14360
rect 18160 -14450 18214 -14416
rect 18248 -14450 18304 -14416
rect 18338 -14450 18394 -14416
rect 18428 -14450 18484 -14416
rect 18518 -14450 18574 -14416
rect 18608 -14450 18664 -14416
rect 18698 -14450 18754 -14416
rect 18788 -14450 18840 -14416
rect 18160 -14506 18840 -14450
rect 18160 -14540 18214 -14506
rect 18248 -14540 18304 -14506
rect 18338 -14540 18394 -14506
rect 18428 -14540 18484 -14506
rect 18518 -14540 18574 -14506
rect 18608 -14540 18664 -14506
rect 18698 -14540 18754 -14506
rect 18788 -14540 18840 -14506
rect 18160 -14596 18840 -14540
rect 18160 -14630 18214 -14596
rect 18248 -14630 18304 -14596
rect 18338 -14630 18394 -14596
rect 18428 -14630 18484 -14596
rect 18518 -14630 18574 -14596
rect 18608 -14630 18664 -14596
rect 18698 -14630 18754 -14596
rect 18788 -14630 18840 -14596
rect 18160 -14686 18840 -14630
rect 18160 -14720 18214 -14686
rect 18248 -14720 18304 -14686
rect 18338 -14720 18394 -14686
rect 18428 -14720 18484 -14686
rect 18518 -14720 18574 -14686
rect 18608 -14720 18664 -14686
rect 18698 -14720 18754 -14686
rect 18788 -14720 18840 -14686
rect 18160 -14776 18840 -14720
rect 18160 -14810 18214 -14776
rect 18248 -14810 18304 -14776
rect 18338 -14810 18394 -14776
rect 18428 -14810 18484 -14776
rect 18518 -14810 18574 -14776
rect 18608 -14810 18664 -14776
rect 18698 -14810 18754 -14776
rect 18788 -14810 18840 -14776
rect 18160 -14862 18840 -14810
rect 19448 -14236 20128 -14182
rect 19448 -14270 19502 -14236
rect 19536 -14270 19592 -14236
rect 19626 -14270 19682 -14236
rect 19716 -14270 19772 -14236
rect 19806 -14270 19862 -14236
rect 19896 -14270 19952 -14236
rect 19986 -14270 20042 -14236
rect 20076 -14270 20128 -14236
rect 19448 -14326 20128 -14270
rect 19448 -14360 19502 -14326
rect 19536 -14360 19592 -14326
rect 19626 -14360 19682 -14326
rect 19716 -14360 19772 -14326
rect 19806 -14360 19862 -14326
rect 19896 -14360 19952 -14326
rect 19986 -14360 20042 -14326
rect 20076 -14360 20128 -14326
rect 19448 -14416 20128 -14360
rect 19448 -14450 19502 -14416
rect 19536 -14450 19592 -14416
rect 19626 -14450 19682 -14416
rect 19716 -14450 19772 -14416
rect 19806 -14450 19862 -14416
rect 19896 -14450 19952 -14416
rect 19986 -14450 20042 -14416
rect 20076 -14450 20128 -14416
rect 19448 -14506 20128 -14450
rect 19448 -14540 19502 -14506
rect 19536 -14540 19592 -14506
rect 19626 -14540 19682 -14506
rect 19716 -14540 19772 -14506
rect 19806 -14540 19862 -14506
rect 19896 -14540 19952 -14506
rect 19986 -14540 20042 -14506
rect 20076 -14540 20128 -14506
rect 19448 -14596 20128 -14540
rect 19448 -14630 19502 -14596
rect 19536 -14630 19592 -14596
rect 19626 -14630 19682 -14596
rect 19716 -14630 19772 -14596
rect 19806 -14630 19862 -14596
rect 19896 -14630 19952 -14596
rect 19986 -14630 20042 -14596
rect 20076 -14630 20128 -14596
rect 19448 -14686 20128 -14630
rect 19448 -14720 19502 -14686
rect 19536 -14720 19592 -14686
rect 19626 -14720 19682 -14686
rect 19716 -14720 19772 -14686
rect 19806 -14720 19862 -14686
rect 19896 -14720 19952 -14686
rect 19986 -14720 20042 -14686
rect 20076 -14720 20128 -14686
rect 19448 -14776 20128 -14720
rect 19448 -14810 19502 -14776
rect 19536 -14810 19592 -14776
rect 19626 -14810 19682 -14776
rect 19716 -14810 19772 -14776
rect 19806 -14810 19862 -14776
rect 19896 -14810 19952 -14776
rect 19986 -14810 20042 -14776
rect 20076 -14810 20128 -14776
rect 19448 -14862 20128 -14810
rect 20736 -14236 21416 -14182
rect 20736 -14270 20790 -14236
rect 20824 -14270 20880 -14236
rect 20914 -14270 20970 -14236
rect 21004 -14270 21060 -14236
rect 21094 -14270 21150 -14236
rect 21184 -14270 21240 -14236
rect 21274 -14270 21330 -14236
rect 21364 -14270 21416 -14236
rect 20736 -14326 21416 -14270
rect 20736 -14360 20790 -14326
rect 20824 -14360 20880 -14326
rect 20914 -14360 20970 -14326
rect 21004 -14360 21060 -14326
rect 21094 -14360 21150 -14326
rect 21184 -14360 21240 -14326
rect 21274 -14360 21330 -14326
rect 21364 -14360 21416 -14326
rect 20736 -14416 21416 -14360
rect 20736 -14450 20790 -14416
rect 20824 -14450 20880 -14416
rect 20914 -14450 20970 -14416
rect 21004 -14450 21060 -14416
rect 21094 -14450 21150 -14416
rect 21184 -14450 21240 -14416
rect 21274 -14450 21330 -14416
rect 21364 -14450 21416 -14416
rect 20736 -14506 21416 -14450
rect 20736 -14540 20790 -14506
rect 20824 -14540 20880 -14506
rect 20914 -14540 20970 -14506
rect 21004 -14540 21060 -14506
rect 21094 -14540 21150 -14506
rect 21184 -14540 21240 -14506
rect 21274 -14540 21330 -14506
rect 21364 -14540 21416 -14506
rect 20736 -14596 21416 -14540
rect 20736 -14630 20790 -14596
rect 20824 -14630 20880 -14596
rect 20914 -14630 20970 -14596
rect 21004 -14630 21060 -14596
rect 21094 -14630 21150 -14596
rect 21184 -14630 21240 -14596
rect 21274 -14630 21330 -14596
rect 21364 -14630 21416 -14596
rect 20736 -14686 21416 -14630
rect 20736 -14720 20790 -14686
rect 20824 -14720 20880 -14686
rect 20914 -14720 20970 -14686
rect 21004 -14720 21060 -14686
rect 21094 -14720 21150 -14686
rect 21184 -14720 21240 -14686
rect 21274 -14720 21330 -14686
rect 21364 -14720 21416 -14686
rect 20736 -14776 21416 -14720
rect 20736 -14810 20790 -14776
rect 20824 -14810 20880 -14776
rect 20914 -14810 20970 -14776
rect 21004 -14810 21060 -14776
rect 21094 -14810 21150 -14776
rect 21184 -14810 21240 -14776
rect 21274 -14810 21330 -14776
rect 21364 -14810 21416 -14776
rect 20736 -14862 21416 -14810
rect 22024 -14236 22704 -14182
rect 22024 -14270 22078 -14236
rect 22112 -14270 22168 -14236
rect 22202 -14270 22258 -14236
rect 22292 -14270 22348 -14236
rect 22382 -14270 22438 -14236
rect 22472 -14270 22528 -14236
rect 22562 -14270 22618 -14236
rect 22652 -14270 22704 -14236
rect 22024 -14326 22704 -14270
rect 22024 -14360 22078 -14326
rect 22112 -14360 22168 -14326
rect 22202 -14360 22258 -14326
rect 22292 -14360 22348 -14326
rect 22382 -14360 22438 -14326
rect 22472 -14360 22528 -14326
rect 22562 -14360 22618 -14326
rect 22652 -14360 22704 -14326
rect 22024 -14416 22704 -14360
rect 22024 -14450 22078 -14416
rect 22112 -14450 22168 -14416
rect 22202 -14450 22258 -14416
rect 22292 -14450 22348 -14416
rect 22382 -14450 22438 -14416
rect 22472 -14450 22528 -14416
rect 22562 -14450 22618 -14416
rect 22652 -14450 22704 -14416
rect 22024 -14506 22704 -14450
rect 22024 -14540 22078 -14506
rect 22112 -14540 22168 -14506
rect 22202 -14540 22258 -14506
rect 22292 -14540 22348 -14506
rect 22382 -14540 22438 -14506
rect 22472 -14540 22528 -14506
rect 22562 -14540 22618 -14506
rect 22652 -14540 22704 -14506
rect 22024 -14596 22704 -14540
rect 22024 -14630 22078 -14596
rect 22112 -14630 22168 -14596
rect 22202 -14630 22258 -14596
rect 22292 -14630 22348 -14596
rect 22382 -14630 22438 -14596
rect 22472 -14630 22528 -14596
rect 22562 -14630 22618 -14596
rect 22652 -14630 22704 -14596
rect 22024 -14686 22704 -14630
rect 22024 -14720 22078 -14686
rect 22112 -14720 22168 -14686
rect 22202 -14720 22258 -14686
rect 22292 -14720 22348 -14686
rect 22382 -14720 22438 -14686
rect 22472 -14720 22528 -14686
rect 22562 -14720 22618 -14686
rect 22652 -14720 22704 -14686
rect 22024 -14776 22704 -14720
rect 22024 -14810 22078 -14776
rect 22112 -14810 22168 -14776
rect 22202 -14810 22258 -14776
rect 22292 -14810 22348 -14776
rect 22382 -14810 22438 -14776
rect 22472 -14810 22528 -14776
rect 22562 -14810 22618 -14776
rect 22652 -14810 22704 -14776
rect 22024 -14862 22704 -14810
rect 23312 -14236 23992 -14182
rect 23312 -14270 23366 -14236
rect 23400 -14270 23456 -14236
rect 23490 -14270 23546 -14236
rect 23580 -14270 23636 -14236
rect 23670 -14270 23726 -14236
rect 23760 -14270 23816 -14236
rect 23850 -14270 23906 -14236
rect 23940 -14270 23992 -14236
rect 23312 -14326 23992 -14270
rect 23312 -14360 23366 -14326
rect 23400 -14360 23456 -14326
rect 23490 -14360 23546 -14326
rect 23580 -14360 23636 -14326
rect 23670 -14360 23726 -14326
rect 23760 -14360 23816 -14326
rect 23850 -14360 23906 -14326
rect 23940 -14360 23992 -14326
rect 23312 -14416 23992 -14360
rect 23312 -14450 23366 -14416
rect 23400 -14450 23456 -14416
rect 23490 -14450 23546 -14416
rect 23580 -14450 23636 -14416
rect 23670 -14450 23726 -14416
rect 23760 -14450 23816 -14416
rect 23850 -14450 23906 -14416
rect 23940 -14450 23992 -14416
rect 23312 -14506 23992 -14450
rect 23312 -14540 23366 -14506
rect 23400 -14540 23456 -14506
rect 23490 -14540 23546 -14506
rect 23580 -14540 23636 -14506
rect 23670 -14540 23726 -14506
rect 23760 -14540 23816 -14506
rect 23850 -14540 23906 -14506
rect 23940 -14540 23992 -14506
rect 23312 -14596 23992 -14540
rect 23312 -14630 23366 -14596
rect 23400 -14630 23456 -14596
rect 23490 -14630 23546 -14596
rect 23580 -14630 23636 -14596
rect 23670 -14630 23726 -14596
rect 23760 -14630 23816 -14596
rect 23850 -14630 23906 -14596
rect 23940 -14630 23992 -14596
rect 23312 -14686 23992 -14630
rect 23312 -14720 23366 -14686
rect 23400 -14720 23456 -14686
rect 23490 -14720 23546 -14686
rect 23580 -14720 23636 -14686
rect 23670 -14720 23726 -14686
rect 23760 -14720 23816 -14686
rect 23850 -14720 23906 -14686
rect 23940 -14720 23992 -14686
rect 23312 -14776 23992 -14720
rect 23312 -14810 23366 -14776
rect 23400 -14810 23456 -14776
rect 23490 -14810 23546 -14776
rect 23580 -14810 23636 -14776
rect 23670 -14810 23726 -14776
rect 23760 -14810 23816 -14776
rect 23850 -14810 23906 -14776
rect 23940 -14810 23992 -14776
rect 23312 -14862 23992 -14810
rect 24600 -14236 25280 -14182
rect 24600 -14270 24654 -14236
rect 24688 -14270 24744 -14236
rect 24778 -14270 24834 -14236
rect 24868 -14270 24924 -14236
rect 24958 -14270 25014 -14236
rect 25048 -14270 25104 -14236
rect 25138 -14270 25194 -14236
rect 25228 -14270 25280 -14236
rect 24600 -14326 25280 -14270
rect 24600 -14360 24654 -14326
rect 24688 -14360 24744 -14326
rect 24778 -14360 24834 -14326
rect 24868 -14360 24924 -14326
rect 24958 -14360 25014 -14326
rect 25048 -14360 25104 -14326
rect 25138 -14360 25194 -14326
rect 25228 -14360 25280 -14326
rect 24600 -14416 25280 -14360
rect 24600 -14450 24654 -14416
rect 24688 -14450 24744 -14416
rect 24778 -14450 24834 -14416
rect 24868 -14450 24924 -14416
rect 24958 -14450 25014 -14416
rect 25048 -14450 25104 -14416
rect 25138 -14450 25194 -14416
rect 25228 -14450 25280 -14416
rect 24600 -14506 25280 -14450
rect 24600 -14540 24654 -14506
rect 24688 -14540 24744 -14506
rect 24778 -14540 24834 -14506
rect 24868 -14540 24924 -14506
rect 24958 -14540 25014 -14506
rect 25048 -14540 25104 -14506
rect 25138 -14540 25194 -14506
rect 25228 -14540 25280 -14506
rect 24600 -14596 25280 -14540
rect 24600 -14630 24654 -14596
rect 24688 -14630 24744 -14596
rect 24778 -14630 24834 -14596
rect 24868 -14630 24924 -14596
rect 24958 -14630 25014 -14596
rect 25048 -14630 25104 -14596
rect 25138 -14630 25194 -14596
rect 25228 -14630 25280 -14596
rect 24600 -14686 25280 -14630
rect 24600 -14720 24654 -14686
rect 24688 -14720 24744 -14686
rect 24778 -14720 24834 -14686
rect 24868 -14720 24924 -14686
rect 24958 -14720 25014 -14686
rect 25048 -14720 25104 -14686
rect 25138 -14720 25194 -14686
rect 25228 -14720 25280 -14686
rect 24600 -14776 25280 -14720
rect 24600 -14810 24654 -14776
rect 24688 -14810 24744 -14776
rect 24778 -14810 24834 -14776
rect 24868 -14810 24924 -14776
rect 24958 -14810 25014 -14776
rect 25048 -14810 25104 -14776
rect 25138 -14810 25194 -14776
rect 25228 -14810 25280 -14776
rect 24600 -14862 25280 -14810
rect 25888 -14236 26568 -14182
rect 25888 -14270 25942 -14236
rect 25976 -14270 26032 -14236
rect 26066 -14270 26122 -14236
rect 26156 -14270 26212 -14236
rect 26246 -14270 26302 -14236
rect 26336 -14270 26392 -14236
rect 26426 -14270 26482 -14236
rect 26516 -14270 26568 -14236
rect 25888 -14326 26568 -14270
rect 25888 -14360 25942 -14326
rect 25976 -14360 26032 -14326
rect 26066 -14360 26122 -14326
rect 26156 -14360 26212 -14326
rect 26246 -14360 26302 -14326
rect 26336 -14360 26392 -14326
rect 26426 -14360 26482 -14326
rect 26516 -14360 26568 -14326
rect 25888 -14416 26568 -14360
rect 25888 -14450 25942 -14416
rect 25976 -14450 26032 -14416
rect 26066 -14450 26122 -14416
rect 26156 -14450 26212 -14416
rect 26246 -14450 26302 -14416
rect 26336 -14450 26392 -14416
rect 26426 -14450 26482 -14416
rect 26516 -14450 26568 -14416
rect 25888 -14506 26568 -14450
rect 25888 -14540 25942 -14506
rect 25976 -14540 26032 -14506
rect 26066 -14540 26122 -14506
rect 26156 -14540 26212 -14506
rect 26246 -14540 26302 -14506
rect 26336 -14540 26392 -14506
rect 26426 -14540 26482 -14506
rect 26516 -14540 26568 -14506
rect 25888 -14596 26568 -14540
rect 25888 -14630 25942 -14596
rect 25976 -14630 26032 -14596
rect 26066 -14630 26122 -14596
rect 26156 -14630 26212 -14596
rect 26246 -14630 26302 -14596
rect 26336 -14630 26392 -14596
rect 26426 -14630 26482 -14596
rect 26516 -14630 26568 -14596
rect 25888 -14686 26568 -14630
rect 25888 -14720 25942 -14686
rect 25976 -14720 26032 -14686
rect 26066 -14720 26122 -14686
rect 26156 -14720 26212 -14686
rect 26246 -14720 26302 -14686
rect 26336 -14720 26392 -14686
rect 26426 -14720 26482 -14686
rect 26516 -14720 26568 -14686
rect 25888 -14776 26568 -14720
rect 25888 -14810 25942 -14776
rect 25976 -14810 26032 -14776
rect 26066 -14810 26122 -14776
rect 26156 -14810 26212 -14776
rect 26246 -14810 26302 -14776
rect 26336 -14810 26392 -14776
rect 26426 -14810 26482 -14776
rect 26516 -14810 26568 -14776
rect 25888 -14862 26568 -14810
rect 16872 -15524 17552 -15470
rect 16872 -15558 16926 -15524
rect 16960 -15558 17016 -15524
rect 17050 -15558 17106 -15524
rect 17140 -15558 17196 -15524
rect 17230 -15558 17286 -15524
rect 17320 -15558 17376 -15524
rect 17410 -15558 17466 -15524
rect 17500 -15558 17552 -15524
rect 16872 -15614 17552 -15558
rect 16872 -15648 16926 -15614
rect 16960 -15648 17016 -15614
rect 17050 -15648 17106 -15614
rect 17140 -15648 17196 -15614
rect 17230 -15648 17286 -15614
rect 17320 -15648 17376 -15614
rect 17410 -15648 17466 -15614
rect 17500 -15648 17552 -15614
rect 16872 -15704 17552 -15648
rect 16872 -15738 16926 -15704
rect 16960 -15738 17016 -15704
rect 17050 -15738 17106 -15704
rect 17140 -15738 17196 -15704
rect 17230 -15738 17286 -15704
rect 17320 -15738 17376 -15704
rect 17410 -15738 17466 -15704
rect 17500 -15738 17552 -15704
rect 16872 -15794 17552 -15738
rect 16872 -15828 16926 -15794
rect 16960 -15828 17016 -15794
rect 17050 -15828 17106 -15794
rect 17140 -15828 17196 -15794
rect 17230 -15828 17286 -15794
rect 17320 -15828 17376 -15794
rect 17410 -15828 17466 -15794
rect 17500 -15828 17552 -15794
rect 16872 -15884 17552 -15828
rect 16872 -15918 16926 -15884
rect 16960 -15918 17016 -15884
rect 17050 -15918 17106 -15884
rect 17140 -15918 17196 -15884
rect 17230 -15918 17286 -15884
rect 17320 -15918 17376 -15884
rect 17410 -15918 17466 -15884
rect 17500 -15918 17552 -15884
rect 16872 -15974 17552 -15918
rect 16872 -16008 16926 -15974
rect 16960 -16008 17016 -15974
rect 17050 -16008 17106 -15974
rect 17140 -16008 17196 -15974
rect 17230 -16008 17286 -15974
rect 17320 -16008 17376 -15974
rect 17410 -16008 17466 -15974
rect 17500 -16008 17552 -15974
rect 16872 -16064 17552 -16008
rect 16872 -16098 16926 -16064
rect 16960 -16098 17016 -16064
rect 17050 -16098 17106 -16064
rect 17140 -16098 17196 -16064
rect 17230 -16098 17286 -16064
rect 17320 -16098 17376 -16064
rect 17410 -16098 17466 -16064
rect 17500 -16098 17552 -16064
rect 16872 -16150 17552 -16098
rect 18160 -15524 18840 -15470
rect 18160 -15558 18214 -15524
rect 18248 -15558 18304 -15524
rect 18338 -15558 18394 -15524
rect 18428 -15558 18484 -15524
rect 18518 -15558 18574 -15524
rect 18608 -15558 18664 -15524
rect 18698 -15558 18754 -15524
rect 18788 -15558 18840 -15524
rect 18160 -15614 18840 -15558
rect 18160 -15648 18214 -15614
rect 18248 -15648 18304 -15614
rect 18338 -15648 18394 -15614
rect 18428 -15648 18484 -15614
rect 18518 -15648 18574 -15614
rect 18608 -15648 18664 -15614
rect 18698 -15648 18754 -15614
rect 18788 -15648 18840 -15614
rect 18160 -15704 18840 -15648
rect 18160 -15738 18214 -15704
rect 18248 -15738 18304 -15704
rect 18338 -15738 18394 -15704
rect 18428 -15738 18484 -15704
rect 18518 -15738 18574 -15704
rect 18608 -15738 18664 -15704
rect 18698 -15738 18754 -15704
rect 18788 -15738 18840 -15704
rect 18160 -15794 18840 -15738
rect 18160 -15828 18214 -15794
rect 18248 -15828 18304 -15794
rect 18338 -15828 18394 -15794
rect 18428 -15828 18484 -15794
rect 18518 -15828 18574 -15794
rect 18608 -15828 18664 -15794
rect 18698 -15828 18754 -15794
rect 18788 -15828 18840 -15794
rect 18160 -15884 18840 -15828
rect 18160 -15918 18214 -15884
rect 18248 -15918 18304 -15884
rect 18338 -15918 18394 -15884
rect 18428 -15918 18484 -15884
rect 18518 -15918 18574 -15884
rect 18608 -15918 18664 -15884
rect 18698 -15918 18754 -15884
rect 18788 -15918 18840 -15884
rect 18160 -15974 18840 -15918
rect 18160 -16008 18214 -15974
rect 18248 -16008 18304 -15974
rect 18338 -16008 18394 -15974
rect 18428 -16008 18484 -15974
rect 18518 -16008 18574 -15974
rect 18608 -16008 18664 -15974
rect 18698 -16008 18754 -15974
rect 18788 -16008 18840 -15974
rect 18160 -16064 18840 -16008
rect 18160 -16098 18214 -16064
rect 18248 -16098 18304 -16064
rect 18338 -16098 18394 -16064
rect 18428 -16098 18484 -16064
rect 18518 -16098 18574 -16064
rect 18608 -16098 18664 -16064
rect 18698 -16098 18754 -16064
rect 18788 -16098 18840 -16064
rect 18160 -16150 18840 -16098
rect 19448 -15524 20128 -15470
rect 19448 -15558 19502 -15524
rect 19536 -15558 19592 -15524
rect 19626 -15558 19682 -15524
rect 19716 -15558 19772 -15524
rect 19806 -15558 19862 -15524
rect 19896 -15558 19952 -15524
rect 19986 -15558 20042 -15524
rect 20076 -15558 20128 -15524
rect 19448 -15614 20128 -15558
rect 19448 -15648 19502 -15614
rect 19536 -15648 19592 -15614
rect 19626 -15648 19682 -15614
rect 19716 -15648 19772 -15614
rect 19806 -15648 19862 -15614
rect 19896 -15648 19952 -15614
rect 19986 -15648 20042 -15614
rect 20076 -15648 20128 -15614
rect 19448 -15704 20128 -15648
rect 19448 -15738 19502 -15704
rect 19536 -15738 19592 -15704
rect 19626 -15738 19682 -15704
rect 19716 -15738 19772 -15704
rect 19806 -15738 19862 -15704
rect 19896 -15738 19952 -15704
rect 19986 -15738 20042 -15704
rect 20076 -15738 20128 -15704
rect 19448 -15794 20128 -15738
rect 19448 -15828 19502 -15794
rect 19536 -15828 19592 -15794
rect 19626 -15828 19682 -15794
rect 19716 -15828 19772 -15794
rect 19806 -15828 19862 -15794
rect 19896 -15828 19952 -15794
rect 19986 -15828 20042 -15794
rect 20076 -15828 20128 -15794
rect 19448 -15884 20128 -15828
rect 19448 -15918 19502 -15884
rect 19536 -15918 19592 -15884
rect 19626 -15918 19682 -15884
rect 19716 -15918 19772 -15884
rect 19806 -15918 19862 -15884
rect 19896 -15918 19952 -15884
rect 19986 -15918 20042 -15884
rect 20076 -15918 20128 -15884
rect 19448 -15974 20128 -15918
rect 19448 -16008 19502 -15974
rect 19536 -16008 19592 -15974
rect 19626 -16008 19682 -15974
rect 19716 -16008 19772 -15974
rect 19806 -16008 19862 -15974
rect 19896 -16008 19952 -15974
rect 19986 -16008 20042 -15974
rect 20076 -16008 20128 -15974
rect 19448 -16064 20128 -16008
rect 19448 -16098 19502 -16064
rect 19536 -16098 19592 -16064
rect 19626 -16098 19682 -16064
rect 19716 -16098 19772 -16064
rect 19806 -16098 19862 -16064
rect 19896 -16098 19952 -16064
rect 19986 -16098 20042 -16064
rect 20076 -16098 20128 -16064
rect 19448 -16150 20128 -16098
rect 20736 -15524 21416 -15470
rect 20736 -15558 20790 -15524
rect 20824 -15558 20880 -15524
rect 20914 -15558 20970 -15524
rect 21004 -15558 21060 -15524
rect 21094 -15558 21150 -15524
rect 21184 -15558 21240 -15524
rect 21274 -15558 21330 -15524
rect 21364 -15558 21416 -15524
rect 20736 -15614 21416 -15558
rect 20736 -15648 20790 -15614
rect 20824 -15648 20880 -15614
rect 20914 -15648 20970 -15614
rect 21004 -15648 21060 -15614
rect 21094 -15648 21150 -15614
rect 21184 -15648 21240 -15614
rect 21274 -15648 21330 -15614
rect 21364 -15648 21416 -15614
rect 20736 -15704 21416 -15648
rect 20736 -15738 20790 -15704
rect 20824 -15738 20880 -15704
rect 20914 -15738 20970 -15704
rect 21004 -15738 21060 -15704
rect 21094 -15738 21150 -15704
rect 21184 -15738 21240 -15704
rect 21274 -15738 21330 -15704
rect 21364 -15738 21416 -15704
rect 20736 -15794 21416 -15738
rect 20736 -15828 20790 -15794
rect 20824 -15828 20880 -15794
rect 20914 -15828 20970 -15794
rect 21004 -15828 21060 -15794
rect 21094 -15828 21150 -15794
rect 21184 -15828 21240 -15794
rect 21274 -15828 21330 -15794
rect 21364 -15828 21416 -15794
rect 20736 -15884 21416 -15828
rect 20736 -15918 20790 -15884
rect 20824 -15918 20880 -15884
rect 20914 -15918 20970 -15884
rect 21004 -15918 21060 -15884
rect 21094 -15918 21150 -15884
rect 21184 -15918 21240 -15884
rect 21274 -15918 21330 -15884
rect 21364 -15918 21416 -15884
rect 20736 -15974 21416 -15918
rect 20736 -16008 20790 -15974
rect 20824 -16008 20880 -15974
rect 20914 -16008 20970 -15974
rect 21004 -16008 21060 -15974
rect 21094 -16008 21150 -15974
rect 21184 -16008 21240 -15974
rect 21274 -16008 21330 -15974
rect 21364 -16008 21416 -15974
rect 20736 -16064 21416 -16008
rect 20736 -16098 20790 -16064
rect 20824 -16098 20880 -16064
rect 20914 -16098 20970 -16064
rect 21004 -16098 21060 -16064
rect 21094 -16098 21150 -16064
rect 21184 -16098 21240 -16064
rect 21274 -16098 21330 -16064
rect 21364 -16098 21416 -16064
rect 20736 -16150 21416 -16098
rect 22024 -15524 22704 -15470
rect 22024 -15558 22078 -15524
rect 22112 -15558 22168 -15524
rect 22202 -15558 22258 -15524
rect 22292 -15558 22348 -15524
rect 22382 -15558 22438 -15524
rect 22472 -15558 22528 -15524
rect 22562 -15558 22618 -15524
rect 22652 -15558 22704 -15524
rect 22024 -15614 22704 -15558
rect 22024 -15648 22078 -15614
rect 22112 -15648 22168 -15614
rect 22202 -15648 22258 -15614
rect 22292 -15648 22348 -15614
rect 22382 -15648 22438 -15614
rect 22472 -15648 22528 -15614
rect 22562 -15648 22618 -15614
rect 22652 -15648 22704 -15614
rect 22024 -15704 22704 -15648
rect 22024 -15738 22078 -15704
rect 22112 -15738 22168 -15704
rect 22202 -15738 22258 -15704
rect 22292 -15738 22348 -15704
rect 22382 -15738 22438 -15704
rect 22472 -15738 22528 -15704
rect 22562 -15738 22618 -15704
rect 22652 -15738 22704 -15704
rect 22024 -15794 22704 -15738
rect 22024 -15828 22078 -15794
rect 22112 -15828 22168 -15794
rect 22202 -15828 22258 -15794
rect 22292 -15828 22348 -15794
rect 22382 -15828 22438 -15794
rect 22472 -15828 22528 -15794
rect 22562 -15828 22618 -15794
rect 22652 -15828 22704 -15794
rect 22024 -15884 22704 -15828
rect 22024 -15918 22078 -15884
rect 22112 -15918 22168 -15884
rect 22202 -15918 22258 -15884
rect 22292 -15918 22348 -15884
rect 22382 -15918 22438 -15884
rect 22472 -15918 22528 -15884
rect 22562 -15918 22618 -15884
rect 22652 -15918 22704 -15884
rect 22024 -15974 22704 -15918
rect 22024 -16008 22078 -15974
rect 22112 -16008 22168 -15974
rect 22202 -16008 22258 -15974
rect 22292 -16008 22348 -15974
rect 22382 -16008 22438 -15974
rect 22472 -16008 22528 -15974
rect 22562 -16008 22618 -15974
rect 22652 -16008 22704 -15974
rect 22024 -16064 22704 -16008
rect 22024 -16098 22078 -16064
rect 22112 -16098 22168 -16064
rect 22202 -16098 22258 -16064
rect 22292 -16098 22348 -16064
rect 22382 -16098 22438 -16064
rect 22472 -16098 22528 -16064
rect 22562 -16098 22618 -16064
rect 22652 -16098 22704 -16064
rect 22024 -16150 22704 -16098
rect 23312 -15524 23992 -15470
rect 23312 -15558 23366 -15524
rect 23400 -15558 23456 -15524
rect 23490 -15558 23546 -15524
rect 23580 -15558 23636 -15524
rect 23670 -15558 23726 -15524
rect 23760 -15558 23816 -15524
rect 23850 -15558 23906 -15524
rect 23940 -15558 23992 -15524
rect 23312 -15614 23992 -15558
rect 23312 -15648 23366 -15614
rect 23400 -15648 23456 -15614
rect 23490 -15648 23546 -15614
rect 23580 -15648 23636 -15614
rect 23670 -15648 23726 -15614
rect 23760 -15648 23816 -15614
rect 23850 -15648 23906 -15614
rect 23940 -15648 23992 -15614
rect 23312 -15704 23992 -15648
rect 23312 -15738 23366 -15704
rect 23400 -15738 23456 -15704
rect 23490 -15738 23546 -15704
rect 23580 -15738 23636 -15704
rect 23670 -15738 23726 -15704
rect 23760 -15738 23816 -15704
rect 23850 -15738 23906 -15704
rect 23940 -15738 23992 -15704
rect 23312 -15794 23992 -15738
rect 23312 -15828 23366 -15794
rect 23400 -15828 23456 -15794
rect 23490 -15828 23546 -15794
rect 23580 -15828 23636 -15794
rect 23670 -15828 23726 -15794
rect 23760 -15828 23816 -15794
rect 23850 -15828 23906 -15794
rect 23940 -15828 23992 -15794
rect 23312 -15884 23992 -15828
rect 23312 -15918 23366 -15884
rect 23400 -15918 23456 -15884
rect 23490 -15918 23546 -15884
rect 23580 -15918 23636 -15884
rect 23670 -15918 23726 -15884
rect 23760 -15918 23816 -15884
rect 23850 -15918 23906 -15884
rect 23940 -15918 23992 -15884
rect 23312 -15974 23992 -15918
rect 23312 -16008 23366 -15974
rect 23400 -16008 23456 -15974
rect 23490 -16008 23546 -15974
rect 23580 -16008 23636 -15974
rect 23670 -16008 23726 -15974
rect 23760 -16008 23816 -15974
rect 23850 -16008 23906 -15974
rect 23940 -16008 23992 -15974
rect 23312 -16064 23992 -16008
rect 23312 -16098 23366 -16064
rect 23400 -16098 23456 -16064
rect 23490 -16098 23546 -16064
rect 23580 -16098 23636 -16064
rect 23670 -16098 23726 -16064
rect 23760 -16098 23816 -16064
rect 23850 -16098 23906 -16064
rect 23940 -16098 23992 -16064
rect 23312 -16150 23992 -16098
rect 24600 -15524 25280 -15470
rect 24600 -15558 24654 -15524
rect 24688 -15558 24744 -15524
rect 24778 -15558 24834 -15524
rect 24868 -15558 24924 -15524
rect 24958 -15558 25014 -15524
rect 25048 -15558 25104 -15524
rect 25138 -15558 25194 -15524
rect 25228 -15558 25280 -15524
rect 24600 -15614 25280 -15558
rect 24600 -15648 24654 -15614
rect 24688 -15648 24744 -15614
rect 24778 -15648 24834 -15614
rect 24868 -15648 24924 -15614
rect 24958 -15648 25014 -15614
rect 25048 -15648 25104 -15614
rect 25138 -15648 25194 -15614
rect 25228 -15648 25280 -15614
rect 24600 -15704 25280 -15648
rect 24600 -15738 24654 -15704
rect 24688 -15738 24744 -15704
rect 24778 -15738 24834 -15704
rect 24868 -15738 24924 -15704
rect 24958 -15738 25014 -15704
rect 25048 -15738 25104 -15704
rect 25138 -15738 25194 -15704
rect 25228 -15738 25280 -15704
rect 24600 -15794 25280 -15738
rect 24600 -15828 24654 -15794
rect 24688 -15828 24744 -15794
rect 24778 -15828 24834 -15794
rect 24868 -15828 24924 -15794
rect 24958 -15828 25014 -15794
rect 25048 -15828 25104 -15794
rect 25138 -15828 25194 -15794
rect 25228 -15828 25280 -15794
rect 24600 -15884 25280 -15828
rect 24600 -15918 24654 -15884
rect 24688 -15918 24744 -15884
rect 24778 -15918 24834 -15884
rect 24868 -15918 24924 -15884
rect 24958 -15918 25014 -15884
rect 25048 -15918 25104 -15884
rect 25138 -15918 25194 -15884
rect 25228 -15918 25280 -15884
rect 24600 -15974 25280 -15918
rect 24600 -16008 24654 -15974
rect 24688 -16008 24744 -15974
rect 24778 -16008 24834 -15974
rect 24868 -16008 24924 -15974
rect 24958 -16008 25014 -15974
rect 25048 -16008 25104 -15974
rect 25138 -16008 25194 -15974
rect 25228 -16008 25280 -15974
rect 24600 -16064 25280 -16008
rect 24600 -16098 24654 -16064
rect 24688 -16098 24744 -16064
rect 24778 -16098 24834 -16064
rect 24868 -16098 24924 -16064
rect 24958 -16098 25014 -16064
rect 25048 -16098 25104 -16064
rect 25138 -16098 25194 -16064
rect 25228 -16098 25280 -16064
rect 24600 -16150 25280 -16098
rect 25888 -15524 26568 -15470
rect 25888 -15558 25942 -15524
rect 25976 -15558 26032 -15524
rect 26066 -15558 26122 -15524
rect 26156 -15558 26212 -15524
rect 26246 -15558 26302 -15524
rect 26336 -15558 26392 -15524
rect 26426 -15558 26482 -15524
rect 26516 -15558 26568 -15524
rect 25888 -15614 26568 -15558
rect 25888 -15648 25942 -15614
rect 25976 -15648 26032 -15614
rect 26066 -15648 26122 -15614
rect 26156 -15648 26212 -15614
rect 26246 -15648 26302 -15614
rect 26336 -15648 26392 -15614
rect 26426 -15648 26482 -15614
rect 26516 -15648 26568 -15614
rect 25888 -15704 26568 -15648
rect 25888 -15738 25942 -15704
rect 25976 -15738 26032 -15704
rect 26066 -15738 26122 -15704
rect 26156 -15738 26212 -15704
rect 26246 -15738 26302 -15704
rect 26336 -15738 26392 -15704
rect 26426 -15738 26482 -15704
rect 26516 -15738 26568 -15704
rect 25888 -15794 26568 -15738
rect 25888 -15828 25942 -15794
rect 25976 -15828 26032 -15794
rect 26066 -15828 26122 -15794
rect 26156 -15828 26212 -15794
rect 26246 -15828 26302 -15794
rect 26336 -15828 26392 -15794
rect 26426 -15828 26482 -15794
rect 26516 -15828 26568 -15794
rect 25888 -15884 26568 -15828
rect 25888 -15918 25942 -15884
rect 25976 -15918 26032 -15884
rect 26066 -15918 26122 -15884
rect 26156 -15918 26212 -15884
rect 26246 -15918 26302 -15884
rect 26336 -15918 26392 -15884
rect 26426 -15918 26482 -15884
rect 26516 -15918 26568 -15884
rect 25888 -15974 26568 -15918
rect 25888 -16008 25942 -15974
rect 25976 -16008 26032 -15974
rect 26066 -16008 26122 -15974
rect 26156 -16008 26212 -15974
rect 26246 -16008 26302 -15974
rect 26336 -16008 26392 -15974
rect 26426 -16008 26482 -15974
rect 26516 -16008 26568 -15974
rect 25888 -16064 26568 -16008
rect 25888 -16098 25942 -16064
rect 25976 -16098 26032 -16064
rect 26066 -16098 26122 -16064
rect 26156 -16098 26212 -16064
rect 26246 -16098 26302 -16064
rect 26336 -16098 26392 -16064
rect 26426 -16098 26482 -16064
rect 26516 -16098 26568 -16064
rect 25888 -16150 26568 -16098
rect 16872 -16812 17552 -16758
rect 16872 -16846 16926 -16812
rect 16960 -16846 17016 -16812
rect 17050 -16846 17106 -16812
rect 17140 -16846 17196 -16812
rect 17230 -16846 17286 -16812
rect 17320 -16846 17376 -16812
rect 17410 -16846 17466 -16812
rect 17500 -16846 17552 -16812
rect 16872 -16902 17552 -16846
rect 16872 -16936 16926 -16902
rect 16960 -16936 17016 -16902
rect 17050 -16936 17106 -16902
rect 17140 -16936 17196 -16902
rect 17230 -16936 17286 -16902
rect 17320 -16936 17376 -16902
rect 17410 -16936 17466 -16902
rect 17500 -16936 17552 -16902
rect 16872 -16992 17552 -16936
rect 16872 -17026 16926 -16992
rect 16960 -17026 17016 -16992
rect 17050 -17026 17106 -16992
rect 17140 -17026 17196 -16992
rect 17230 -17026 17286 -16992
rect 17320 -17026 17376 -16992
rect 17410 -17026 17466 -16992
rect 17500 -17026 17552 -16992
rect 16872 -17082 17552 -17026
rect 16872 -17116 16926 -17082
rect 16960 -17116 17016 -17082
rect 17050 -17116 17106 -17082
rect 17140 -17116 17196 -17082
rect 17230 -17116 17286 -17082
rect 17320 -17116 17376 -17082
rect 17410 -17116 17466 -17082
rect 17500 -17116 17552 -17082
rect 16872 -17172 17552 -17116
rect 16872 -17206 16926 -17172
rect 16960 -17206 17016 -17172
rect 17050 -17206 17106 -17172
rect 17140 -17206 17196 -17172
rect 17230 -17206 17286 -17172
rect 17320 -17206 17376 -17172
rect 17410 -17206 17466 -17172
rect 17500 -17206 17552 -17172
rect 16872 -17262 17552 -17206
rect 16872 -17296 16926 -17262
rect 16960 -17296 17016 -17262
rect 17050 -17296 17106 -17262
rect 17140 -17296 17196 -17262
rect 17230 -17296 17286 -17262
rect 17320 -17296 17376 -17262
rect 17410 -17296 17466 -17262
rect 17500 -17296 17552 -17262
rect 16872 -17352 17552 -17296
rect 16872 -17386 16926 -17352
rect 16960 -17386 17016 -17352
rect 17050 -17386 17106 -17352
rect 17140 -17386 17196 -17352
rect 17230 -17386 17286 -17352
rect 17320 -17386 17376 -17352
rect 17410 -17386 17466 -17352
rect 17500 -17386 17552 -17352
rect 16872 -17438 17552 -17386
rect 18160 -16812 18840 -16758
rect 18160 -16846 18214 -16812
rect 18248 -16846 18304 -16812
rect 18338 -16846 18394 -16812
rect 18428 -16846 18484 -16812
rect 18518 -16846 18574 -16812
rect 18608 -16846 18664 -16812
rect 18698 -16846 18754 -16812
rect 18788 -16846 18840 -16812
rect 18160 -16902 18840 -16846
rect 18160 -16936 18214 -16902
rect 18248 -16936 18304 -16902
rect 18338 -16936 18394 -16902
rect 18428 -16936 18484 -16902
rect 18518 -16936 18574 -16902
rect 18608 -16936 18664 -16902
rect 18698 -16936 18754 -16902
rect 18788 -16936 18840 -16902
rect 18160 -16992 18840 -16936
rect 18160 -17026 18214 -16992
rect 18248 -17026 18304 -16992
rect 18338 -17026 18394 -16992
rect 18428 -17026 18484 -16992
rect 18518 -17026 18574 -16992
rect 18608 -17026 18664 -16992
rect 18698 -17026 18754 -16992
rect 18788 -17026 18840 -16992
rect 18160 -17082 18840 -17026
rect 18160 -17116 18214 -17082
rect 18248 -17116 18304 -17082
rect 18338 -17116 18394 -17082
rect 18428 -17116 18484 -17082
rect 18518 -17116 18574 -17082
rect 18608 -17116 18664 -17082
rect 18698 -17116 18754 -17082
rect 18788 -17116 18840 -17082
rect 18160 -17172 18840 -17116
rect 18160 -17206 18214 -17172
rect 18248 -17206 18304 -17172
rect 18338 -17206 18394 -17172
rect 18428 -17206 18484 -17172
rect 18518 -17206 18574 -17172
rect 18608 -17206 18664 -17172
rect 18698 -17206 18754 -17172
rect 18788 -17206 18840 -17172
rect 18160 -17262 18840 -17206
rect 18160 -17296 18214 -17262
rect 18248 -17296 18304 -17262
rect 18338 -17296 18394 -17262
rect 18428 -17296 18484 -17262
rect 18518 -17296 18574 -17262
rect 18608 -17296 18664 -17262
rect 18698 -17296 18754 -17262
rect 18788 -17296 18840 -17262
rect 18160 -17352 18840 -17296
rect 18160 -17386 18214 -17352
rect 18248 -17386 18304 -17352
rect 18338 -17386 18394 -17352
rect 18428 -17386 18484 -17352
rect 18518 -17386 18574 -17352
rect 18608 -17386 18664 -17352
rect 18698 -17386 18754 -17352
rect 18788 -17386 18840 -17352
rect 18160 -17438 18840 -17386
rect 19448 -16812 20128 -16758
rect 19448 -16846 19502 -16812
rect 19536 -16846 19592 -16812
rect 19626 -16846 19682 -16812
rect 19716 -16846 19772 -16812
rect 19806 -16846 19862 -16812
rect 19896 -16846 19952 -16812
rect 19986 -16846 20042 -16812
rect 20076 -16846 20128 -16812
rect 19448 -16902 20128 -16846
rect 19448 -16936 19502 -16902
rect 19536 -16936 19592 -16902
rect 19626 -16936 19682 -16902
rect 19716 -16936 19772 -16902
rect 19806 -16936 19862 -16902
rect 19896 -16936 19952 -16902
rect 19986 -16936 20042 -16902
rect 20076 -16936 20128 -16902
rect 19448 -16992 20128 -16936
rect 19448 -17026 19502 -16992
rect 19536 -17026 19592 -16992
rect 19626 -17026 19682 -16992
rect 19716 -17026 19772 -16992
rect 19806 -17026 19862 -16992
rect 19896 -17026 19952 -16992
rect 19986 -17026 20042 -16992
rect 20076 -17026 20128 -16992
rect 19448 -17082 20128 -17026
rect 19448 -17116 19502 -17082
rect 19536 -17116 19592 -17082
rect 19626 -17116 19682 -17082
rect 19716 -17116 19772 -17082
rect 19806 -17116 19862 -17082
rect 19896 -17116 19952 -17082
rect 19986 -17116 20042 -17082
rect 20076 -17116 20128 -17082
rect 19448 -17172 20128 -17116
rect 19448 -17206 19502 -17172
rect 19536 -17206 19592 -17172
rect 19626 -17206 19682 -17172
rect 19716 -17206 19772 -17172
rect 19806 -17206 19862 -17172
rect 19896 -17206 19952 -17172
rect 19986 -17206 20042 -17172
rect 20076 -17206 20128 -17172
rect 19448 -17262 20128 -17206
rect 19448 -17296 19502 -17262
rect 19536 -17296 19592 -17262
rect 19626 -17296 19682 -17262
rect 19716 -17296 19772 -17262
rect 19806 -17296 19862 -17262
rect 19896 -17296 19952 -17262
rect 19986 -17296 20042 -17262
rect 20076 -17296 20128 -17262
rect 19448 -17352 20128 -17296
rect 19448 -17386 19502 -17352
rect 19536 -17386 19592 -17352
rect 19626 -17386 19682 -17352
rect 19716 -17386 19772 -17352
rect 19806 -17386 19862 -17352
rect 19896 -17386 19952 -17352
rect 19986 -17386 20042 -17352
rect 20076 -17386 20128 -17352
rect 19448 -17438 20128 -17386
rect 20736 -16812 21416 -16758
rect 20736 -16846 20790 -16812
rect 20824 -16846 20880 -16812
rect 20914 -16846 20970 -16812
rect 21004 -16846 21060 -16812
rect 21094 -16846 21150 -16812
rect 21184 -16846 21240 -16812
rect 21274 -16846 21330 -16812
rect 21364 -16846 21416 -16812
rect 20736 -16902 21416 -16846
rect 20736 -16936 20790 -16902
rect 20824 -16936 20880 -16902
rect 20914 -16936 20970 -16902
rect 21004 -16936 21060 -16902
rect 21094 -16936 21150 -16902
rect 21184 -16936 21240 -16902
rect 21274 -16936 21330 -16902
rect 21364 -16936 21416 -16902
rect 20736 -16992 21416 -16936
rect 20736 -17026 20790 -16992
rect 20824 -17026 20880 -16992
rect 20914 -17026 20970 -16992
rect 21004 -17026 21060 -16992
rect 21094 -17026 21150 -16992
rect 21184 -17026 21240 -16992
rect 21274 -17026 21330 -16992
rect 21364 -17026 21416 -16992
rect 20736 -17082 21416 -17026
rect 20736 -17116 20790 -17082
rect 20824 -17116 20880 -17082
rect 20914 -17116 20970 -17082
rect 21004 -17116 21060 -17082
rect 21094 -17116 21150 -17082
rect 21184 -17116 21240 -17082
rect 21274 -17116 21330 -17082
rect 21364 -17116 21416 -17082
rect 20736 -17172 21416 -17116
rect 20736 -17206 20790 -17172
rect 20824 -17206 20880 -17172
rect 20914 -17206 20970 -17172
rect 21004 -17206 21060 -17172
rect 21094 -17206 21150 -17172
rect 21184 -17206 21240 -17172
rect 21274 -17206 21330 -17172
rect 21364 -17206 21416 -17172
rect 20736 -17262 21416 -17206
rect 20736 -17296 20790 -17262
rect 20824 -17296 20880 -17262
rect 20914 -17296 20970 -17262
rect 21004 -17296 21060 -17262
rect 21094 -17296 21150 -17262
rect 21184 -17296 21240 -17262
rect 21274 -17296 21330 -17262
rect 21364 -17296 21416 -17262
rect 20736 -17352 21416 -17296
rect 20736 -17386 20790 -17352
rect 20824 -17386 20880 -17352
rect 20914 -17386 20970 -17352
rect 21004 -17386 21060 -17352
rect 21094 -17386 21150 -17352
rect 21184 -17386 21240 -17352
rect 21274 -17386 21330 -17352
rect 21364 -17386 21416 -17352
rect 20736 -17438 21416 -17386
rect 22024 -16812 22704 -16758
rect 22024 -16846 22078 -16812
rect 22112 -16846 22168 -16812
rect 22202 -16846 22258 -16812
rect 22292 -16846 22348 -16812
rect 22382 -16846 22438 -16812
rect 22472 -16846 22528 -16812
rect 22562 -16846 22618 -16812
rect 22652 -16846 22704 -16812
rect 22024 -16902 22704 -16846
rect 22024 -16936 22078 -16902
rect 22112 -16936 22168 -16902
rect 22202 -16936 22258 -16902
rect 22292 -16936 22348 -16902
rect 22382 -16936 22438 -16902
rect 22472 -16936 22528 -16902
rect 22562 -16936 22618 -16902
rect 22652 -16936 22704 -16902
rect 22024 -16992 22704 -16936
rect 22024 -17026 22078 -16992
rect 22112 -17026 22168 -16992
rect 22202 -17026 22258 -16992
rect 22292 -17026 22348 -16992
rect 22382 -17026 22438 -16992
rect 22472 -17026 22528 -16992
rect 22562 -17026 22618 -16992
rect 22652 -17026 22704 -16992
rect 22024 -17082 22704 -17026
rect 22024 -17116 22078 -17082
rect 22112 -17116 22168 -17082
rect 22202 -17116 22258 -17082
rect 22292 -17116 22348 -17082
rect 22382 -17116 22438 -17082
rect 22472 -17116 22528 -17082
rect 22562 -17116 22618 -17082
rect 22652 -17116 22704 -17082
rect 22024 -17172 22704 -17116
rect 22024 -17206 22078 -17172
rect 22112 -17206 22168 -17172
rect 22202 -17206 22258 -17172
rect 22292 -17206 22348 -17172
rect 22382 -17206 22438 -17172
rect 22472 -17206 22528 -17172
rect 22562 -17206 22618 -17172
rect 22652 -17206 22704 -17172
rect 22024 -17262 22704 -17206
rect 22024 -17296 22078 -17262
rect 22112 -17296 22168 -17262
rect 22202 -17296 22258 -17262
rect 22292 -17296 22348 -17262
rect 22382 -17296 22438 -17262
rect 22472 -17296 22528 -17262
rect 22562 -17296 22618 -17262
rect 22652 -17296 22704 -17262
rect 22024 -17352 22704 -17296
rect 22024 -17386 22078 -17352
rect 22112 -17386 22168 -17352
rect 22202 -17386 22258 -17352
rect 22292 -17386 22348 -17352
rect 22382 -17386 22438 -17352
rect 22472 -17386 22528 -17352
rect 22562 -17386 22618 -17352
rect 22652 -17386 22704 -17352
rect 22024 -17438 22704 -17386
rect 23312 -16812 23992 -16758
rect 23312 -16846 23366 -16812
rect 23400 -16846 23456 -16812
rect 23490 -16846 23546 -16812
rect 23580 -16846 23636 -16812
rect 23670 -16846 23726 -16812
rect 23760 -16846 23816 -16812
rect 23850 -16846 23906 -16812
rect 23940 -16846 23992 -16812
rect 23312 -16902 23992 -16846
rect 23312 -16936 23366 -16902
rect 23400 -16936 23456 -16902
rect 23490 -16936 23546 -16902
rect 23580 -16936 23636 -16902
rect 23670 -16936 23726 -16902
rect 23760 -16936 23816 -16902
rect 23850 -16936 23906 -16902
rect 23940 -16936 23992 -16902
rect 23312 -16992 23992 -16936
rect 23312 -17026 23366 -16992
rect 23400 -17026 23456 -16992
rect 23490 -17026 23546 -16992
rect 23580 -17026 23636 -16992
rect 23670 -17026 23726 -16992
rect 23760 -17026 23816 -16992
rect 23850 -17026 23906 -16992
rect 23940 -17026 23992 -16992
rect 23312 -17082 23992 -17026
rect 23312 -17116 23366 -17082
rect 23400 -17116 23456 -17082
rect 23490 -17116 23546 -17082
rect 23580 -17116 23636 -17082
rect 23670 -17116 23726 -17082
rect 23760 -17116 23816 -17082
rect 23850 -17116 23906 -17082
rect 23940 -17116 23992 -17082
rect 23312 -17172 23992 -17116
rect 23312 -17206 23366 -17172
rect 23400 -17206 23456 -17172
rect 23490 -17206 23546 -17172
rect 23580 -17206 23636 -17172
rect 23670 -17206 23726 -17172
rect 23760 -17206 23816 -17172
rect 23850 -17206 23906 -17172
rect 23940 -17206 23992 -17172
rect 23312 -17262 23992 -17206
rect 23312 -17296 23366 -17262
rect 23400 -17296 23456 -17262
rect 23490 -17296 23546 -17262
rect 23580 -17296 23636 -17262
rect 23670 -17296 23726 -17262
rect 23760 -17296 23816 -17262
rect 23850 -17296 23906 -17262
rect 23940 -17296 23992 -17262
rect 23312 -17352 23992 -17296
rect 23312 -17386 23366 -17352
rect 23400 -17386 23456 -17352
rect 23490 -17386 23546 -17352
rect 23580 -17386 23636 -17352
rect 23670 -17386 23726 -17352
rect 23760 -17386 23816 -17352
rect 23850 -17386 23906 -17352
rect 23940 -17386 23992 -17352
rect 23312 -17438 23992 -17386
rect 24600 -16812 25280 -16758
rect 24600 -16846 24654 -16812
rect 24688 -16846 24744 -16812
rect 24778 -16846 24834 -16812
rect 24868 -16846 24924 -16812
rect 24958 -16846 25014 -16812
rect 25048 -16846 25104 -16812
rect 25138 -16846 25194 -16812
rect 25228 -16846 25280 -16812
rect 24600 -16902 25280 -16846
rect 24600 -16936 24654 -16902
rect 24688 -16936 24744 -16902
rect 24778 -16936 24834 -16902
rect 24868 -16936 24924 -16902
rect 24958 -16936 25014 -16902
rect 25048 -16936 25104 -16902
rect 25138 -16936 25194 -16902
rect 25228 -16936 25280 -16902
rect 24600 -16992 25280 -16936
rect 24600 -17026 24654 -16992
rect 24688 -17026 24744 -16992
rect 24778 -17026 24834 -16992
rect 24868 -17026 24924 -16992
rect 24958 -17026 25014 -16992
rect 25048 -17026 25104 -16992
rect 25138 -17026 25194 -16992
rect 25228 -17026 25280 -16992
rect 24600 -17082 25280 -17026
rect 24600 -17116 24654 -17082
rect 24688 -17116 24744 -17082
rect 24778 -17116 24834 -17082
rect 24868 -17116 24924 -17082
rect 24958 -17116 25014 -17082
rect 25048 -17116 25104 -17082
rect 25138 -17116 25194 -17082
rect 25228 -17116 25280 -17082
rect 24600 -17172 25280 -17116
rect 24600 -17206 24654 -17172
rect 24688 -17206 24744 -17172
rect 24778 -17206 24834 -17172
rect 24868 -17206 24924 -17172
rect 24958 -17206 25014 -17172
rect 25048 -17206 25104 -17172
rect 25138 -17206 25194 -17172
rect 25228 -17206 25280 -17172
rect 24600 -17262 25280 -17206
rect 24600 -17296 24654 -17262
rect 24688 -17296 24744 -17262
rect 24778 -17296 24834 -17262
rect 24868 -17296 24924 -17262
rect 24958 -17296 25014 -17262
rect 25048 -17296 25104 -17262
rect 25138 -17296 25194 -17262
rect 25228 -17296 25280 -17262
rect 24600 -17352 25280 -17296
rect 24600 -17386 24654 -17352
rect 24688 -17386 24744 -17352
rect 24778 -17386 24834 -17352
rect 24868 -17386 24924 -17352
rect 24958 -17386 25014 -17352
rect 25048 -17386 25104 -17352
rect 25138 -17386 25194 -17352
rect 25228 -17386 25280 -17352
rect 24600 -17438 25280 -17386
rect 25888 -16811 26568 -16757
rect 25888 -16846 25942 -16811
rect 25976 -16846 26032 -16811
rect 26066 -16846 26122 -16811
rect 26156 -16846 26212 -16811
rect 26246 -16846 26302 -16811
rect 26336 -16846 26392 -16811
rect 26426 -16846 26482 -16811
rect 26516 -16846 26568 -16811
rect 25888 -16901 26568 -16846
rect 25888 -16936 25942 -16901
rect 25976 -16936 26032 -16901
rect 26066 -16936 26122 -16901
rect 26156 -16936 26212 -16901
rect 26246 -16936 26302 -16901
rect 26336 -16936 26392 -16901
rect 26426 -16936 26482 -16901
rect 26516 -16936 26568 -16901
rect 25888 -16991 26568 -16936
rect 25888 -17026 25942 -16991
rect 25976 -17026 26032 -16991
rect 26066 -17026 26122 -16991
rect 26156 -17026 26212 -16991
rect 26246 -17026 26302 -16991
rect 26336 -17026 26392 -16991
rect 26426 -17026 26482 -16991
rect 26516 -17026 26568 -16991
rect 25888 -17081 26568 -17026
rect 25888 -17116 25942 -17081
rect 25976 -17116 26032 -17081
rect 26066 -17116 26122 -17081
rect 26156 -17116 26212 -17081
rect 26246 -17116 26302 -17081
rect 26336 -17116 26392 -17081
rect 26426 -17116 26482 -17081
rect 26516 -17116 26568 -17081
rect 25888 -17171 26568 -17116
rect 25888 -17206 25942 -17171
rect 25976 -17206 26032 -17171
rect 26066 -17206 26122 -17171
rect 26156 -17206 26212 -17171
rect 26246 -17206 26302 -17171
rect 26336 -17206 26392 -17171
rect 26426 -17206 26482 -17171
rect 26516 -17206 26568 -17171
rect 25888 -17261 26568 -17206
rect 25888 -17296 25942 -17261
rect 25976 -17296 26032 -17261
rect 26066 -17296 26122 -17261
rect 26156 -17296 26212 -17261
rect 26246 -17296 26302 -17261
rect 26336 -17296 26392 -17261
rect 26426 -17296 26482 -17261
rect 26516 -17296 26568 -17261
rect 25888 -17351 26568 -17296
rect 25888 -17386 25942 -17351
rect 25976 -17386 26032 -17351
rect 26066 -17386 26122 -17351
rect 26156 -17386 26212 -17351
rect 26246 -17386 26302 -17351
rect 26336 -17386 26392 -17351
rect 26426 -17386 26482 -17351
rect 26516 -17386 26568 -17351
rect 25888 -17438 26568 -17386
<< pdiffc >>
rect 16926 -11694 16960 -11660
rect 17016 -11694 17050 -11660
rect 17106 -11694 17140 -11660
rect 17196 -11694 17230 -11660
rect 17286 -11694 17320 -11660
rect 17376 -11694 17410 -11660
rect 17466 -11694 17500 -11660
rect 16926 -11784 16960 -11750
rect 17016 -11784 17050 -11750
rect 17106 -11784 17140 -11750
rect 17196 -11784 17230 -11750
rect 17286 -11784 17320 -11750
rect 17376 -11784 17410 -11750
rect 17466 -11784 17500 -11750
rect 16926 -11874 16960 -11840
rect 17016 -11874 17050 -11840
rect 17106 -11874 17140 -11840
rect 17196 -11874 17230 -11840
rect 17286 -11874 17320 -11840
rect 17376 -11874 17410 -11840
rect 17466 -11874 17500 -11840
rect 16926 -11964 16960 -11930
rect 17016 -11964 17050 -11930
rect 17106 -11964 17140 -11930
rect 17196 -11964 17230 -11930
rect 17286 -11964 17320 -11930
rect 17376 -11964 17410 -11930
rect 17466 -11964 17500 -11930
rect 16926 -12054 16960 -12020
rect 17016 -12054 17050 -12020
rect 17106 -12054 17140 -12020
rect 17196 -12054 17230 -12020
rect 17286 -12054 17320 -12020
rect 17376 -12054 17410 -12020
rect 17466 -12054 17500 -12020
rect 16926 -12144 16960 -12110
rect 17016 -12144 17050 -12110
rect 17106 -12144 17140 -12110
rect 17196 -12144 17230 -12110
rect 17286 -12144 17320 -12110
rect 17376 -12144 17410 -12110
rect 17466 -12144 17500 -12110
rect 16926 -12234 16960 -12200
rect 17016 -12234 17050 -12200
rect 17106 -12234 17140 -12200
rect 17196 -12234 17230 -12200
rect 17286 -12234 17320 -12200
rect 17376 -12234 17410 -12200
rect 17466 -12234 17500 -12200
rect 18214 -11694 18248 -11660
rect 18304 -11694 18338 -11660
rect 18394 -11694 18428 -11660
rect 18484 -11694 18518 -11660
rect 18574 -11694 18608 -11660
rect 18664 -11694 18698 -11660
rect 18754 -11694 18788 -11660
rect 18214 -11784 18248 -11750
rect 18304 -11784 18338 -11750
rect 18394 -11784 18428 -11750
rect 18484 -11784 18518 -11750
rect 18574 -11784 18608 -11750
rect 18664 -11784 18698 -11750
rect 18754 -11784 18788 -11750
rect 18214 -11874 18248 -11840
rect 18304 -11874 18338 -11840
rect 18394 -11874 18428 -11840
rect 18484 -11874 18518 -11840
rect 18574 -11874 18608 -11840
rect 18664 -11874 18698 -11840
rect 18754 -11874 18788 -11840
rect 18214 -11964 18248 -11930
rect 18304 -11964 18338 -11930
rect 18394 -11964 18428 -11930
rect 18484 -11964 18518 -11930
rect 18574 -11964 18608 -11930
rect 18664 -11964 18698 -11930
rect 18754 -11964 18788 -11930
rect 18214 -12054 18248 -12020
rect 18304 -12054 18338 -12020
rect 18394 -12054 18428 -12020
rect 18484 -12054 18518 -12020
rect 18574 -12054 18608 -12020
rect 18664 -12054 18698 -12020
rect 18754 -12054 18788 -12020
rect 18214 -12144 18248 -12110
rect 18304 -12144 18338 -12110
rect 18394 -12144 18428 -12110
rect 18484 -12144 18518 -12110
rect 18574 -12144 18608 -12110
rect 18664 -12144 18698 -12110
rect 18754 -12144 18788 -12110
rect 18214 -12234 18248 -12200
rect 18304 -12234 18338 -12200
rect 18394 -12234 18428 -12200
rect 18484 -12234 18518 -12200
rect 18574 -12234 18608 -12200
rect 18664 -12234 18698 -12200
rect 18754 -12234 18788 -12200
rect 19502 -11694 19536 -11660
rect 19592 -11694 19626 -11660
rect 19682 -11694 19716 -11660
rect 19772 -11694 19806 -11660
rect 19862 -11694 19896 -11660
rect 19952 -11694 19986 -11660
rect 20042 -11694 20076 -11660
rect 19502 -11784 19536 -11750
rect 19592 -11784 19626 -11750
rect 19682 -11784 19716 -11750
rect 19772 -11784 19806 -11750
rect 19862 -11784 19896 -11750
rect 19952 -11784 19986 -11750
rect 20042 -11784 20076 -11750
rect 19502 -11874 19536 -11840
rect 19592 -11874 19626 -11840
rect 19682 -11874 19716 -11840
rect 19772 -11874 19806 -11840
rect 19862 -11874 19896 -11840
rect 19952 -11874 19986 -11840
rect 20042 -11874 20076 -11840
rect 19502 -11964 19536 -11930
rect 19592 -11964 19626 -11930
rect 19682 -11964 19716 -11930
rect 19772 -11964 19806 -11930
rect 19862 -11964 19896 -11930
rect 19952 -11964 19986 -11930
rect 20042 -11964 20076 -11930
rect 19502 -12054 19536 -12020
rect 19592 -12054 19626 -12020
rect 19682 -12054 19716 -12020
rect 19772 -12054 19806 -12020
rect 19862 -12054 19896 -12020
rect 19952 -12054 19986 -12020
rect 20042 -12054 20076 -12020
rect 19502 -12144 19536 -12110
rect 19592 -12144 19626 -12110
rect 19682 -12144 19716 -12110
rect 19772 -12144 19806 -12110
rect 19862 -12144 19896 -12110
rect 19952 -12144 19986 -12110
rect 20042 -12144 20076 -12110
rect 19502 -12234 19536 -12200
rect 19592 -12234 19626 -12200
rect 19682 -12234 19716 -12200
rect 19772 -12234 19806 -12200
rect 19862 -12234 19896 -12200
rect 19952 -12234 19986 -12200
rect 20042 -12234 20076 -12200
rect 20790 -11694 20824 -11660
rect 20880 -11694 20914 -11660
rect 20970 -11694 21004 -11660
rect 21060 -11694 21094 -11660
rect 21150 -11694 21184 -11660
rect 21240 -11694 21274 -11660
rect 21330 -11694 21364 -11660
rect 20790 -11784 20824 -11750
rect 20880 -11784 20914 -11750
rect 20970 -11784 21004 -11750
rect 21060 -11784 21094 -11750
rect 21150 -11784 21184 -11750
rect 21240 -11784 21274 -11750
rect 21330 -11784 21364 -11750
rect 20790 -11874 20824 -11840
rect 20880 -11874 20914 -11840
rect 20970 -11874 21004 -11840
rect 21060 -11874 21094 -11840
rect 21150 -11874 21184 -11840
rect 21240 -11874 21274 -11840
rect 21330 -11874 21364 -11840
rect 20790 -11964 20824 -11930
rect 20880 -11964 20914 -11930
rect 20970 -11964 21004 -11930
rect 21060 -11964 21094 -11930
rect 21150 -11964 21184 -11930
rect 21240 -11964 21274 -11930
rect 21330 -11964 21364 -11930
rect 20790 -12054 20824 -12020
rect 20880 -12054 20914 -12020
rect 20970 -12054 21004 -12020
rect 21060 -12054 21094 -12020
rect 21150 -12054 21184 -12020
rect 21240 -12054 21274 -12020
rect 21330 -12054 21364 -12020
rect 20790 -12144 20824 -12110
rect 20880 -12144 20914 -12110
rect 20970 -12144 21004 -12110
rect 21060 -12144 21094 -12110
rect 21150 -12144 21184 -12110
rect 21240 -12144 21274 -12110
rect 21330 -12144 21364 -12110
rect 20790 -12234 20824 -12200
rect 20880 -12234 20914 -12200
rect 20970 -12234 21004 -12200
rect 21060 -12234 21094 -12200
rect 21150 -12234 21184 -12200
rect 21240 -12234 21274 -12200
rect 21330 -12234 21364 -12200
rect 22078 -11694 22112 -11660
rect 22168 -11694 22202 -11660
rect 22258 -11694 22292 -11660
rect 22348 -11694 22382 -11660
rect 22438 -11694 22472 -11660
rect 22528 -11694 22562 -11660
rect 22618 -11694 22652 -11660
rect 22078 -11784 22112 -11750
rect 22168 -11784 22202 -11750
rect 22258 -11784 22292 -11750
rect 22348 -11784 22382 -11750
rect 22438 -11784 22472 -11750
rect 22528 -11784 22562 -11750
rect 22618 -11784 22652 -11750
rect 22078 -11874 22112 -11840
rect 22168 -11874 22202 -11840
rect 22258 -11874 22292 -11840
rect 22348 -11874 22382 -11840
rect 22438 -11874 22472 -11840
rect 22528 -11874 22562 -11840
rect 22618 -11874 22652 -11840
rect 22078 -11964 22112 -11930
rect 22168 -11964 22202 -11930
rect 22258 -11964 22292 -11930
rect 22348 -11964 22382 -11930
rect 22438 -11964 22472 -11930
rect 22528 -11964 22562 -11930
rect 22618 -11964 22652 -11930
rect 22078 -12054 22112 -12020
rect 22168 -12054 22202 -12020
rect 22258 -12054 22292 -12020
rect 22348 -12054 22382 -12020
rect 22438 -12054 22472 -12020
rect 22528 -12054 22562 -12020
rect 22618 -12054 22652 -12020
rect 22078 -12144 22112 -12110
rect 22168 -12144 22202 -12110
rect 22258 -12144 22292 -12110
rect 22348 -12144 22382 -12110
rect 22438 -12144 22472 -12110
rect 22528 -12144 22562 -12110
rect 22618 -12144 22652 -12110
rect 22078 -12234 22112 -12200
rect 22168 -12234 22202 -12200
rect 22258 -12234 22292 -12200
rect 22348 -12234 22382 -12200
rect 22438 -12234 22472 -12200
rect 22528 -12234 22562 -12200
rect 22618 -12234 22652 -12200
rect 23366 -11694 23400 -11660
rect 23456 -11694 23490 -11660
rect 23546 -11694 23580 -11660
rect 23636 -11694 23670 -11660
rect 23726 -11694 23760 -11660
rect 23816 -11694 23850 -11660
rect 23906 -11694 23940 -11660
rect 23366 -11784 23400 -11750
rect 23456 -11784 23490 -11750
rect 23546 -11784 23580 -11750
rect 23636 -11784 23670 -11750
rect 23726 -11784 23760 -11750
rect 23816 -11784 23850 -11750
rect 23906 -11784 23940 -11750
rect 23366 -11874 23400 -11840
rect 23456 -11874 23490 -11840
rect 23546 -11874 23580 -11840
rect 23636 -11874 23670 -11840
rect 23726 -11874 23760 -11840
rect 23816 -11874 23850 -11840
rect 23906 -11874 23940 -11840
rect 23366 -11964 23400 -11930
rect 23456 -11964 23490 -11930
rect 23546 -11964 23580 -11930
rect 23636 -11964 23670 -11930
rect 23726 -11964 23760 -11930
rect 23816 -11964 23850 -11930
rect 23906 -11964 23940 -11930
rect 23366 -12054 23400 -12020
rect 23456 -12054 23490 -12020
rect 23546 -12054 23580 -12020
rect 23636 -12054 23670 -12020
rect 23726 -12054 23760 -12020
rect 23816 -12054 23850 -12020
rect 23906 -12054 23940 -12020
rect 23366 -12144 23400 -12110
rect 23456 -12144 23490 -12110
rect 23546 -12144 23580 -12110
rect 23636 -12144 23670 -12110
rect 23726 -12144 23760 -12110
rect 23816 -12144 23850 -12110
rect 23906 -12144 23940 -12110
rect 23366 -12234 23400 -12200
rect 23456 -12234 23490 -12200
rect 23546 -12234 23580 -12200
rect 23636 -12234 23670 -12200
rect 23726 -12234 23760 -12200
rect 23816 -12234 23850 -12200
rect 23906 -12234 23940 -12200
rect 24654 -11694 24688 -11660
rect 24744 -11694 24778 -11660
rect 24834 -11694 24868 -11660
rect 24924 -11694 24958 -11660
rect 25014 -11694 25048 -11660
rect 25104 -11694 25138 -11660
rect 25194 -11694 25228 -11660
rect 24654 -11784 24688 -11750
rect 24744 -11784 24778 -11750
rect 24834 -11784 24868 -11750
rect 24924 -11784 24958 -11750
rect 25014 -11784 25048 -11750
rect 25104 -11784 25138 -11750
rect 25194 -11784 25228 -11750
rect 24654 -11874 24688 -11840
rect 24744 -11874 24778 -11840
rect 24834 -11874 24868 -11840
rect 24924 -11874 24958 -11840
rect 25014 -11874 25048 -11840
rect 25104 -11874 25138 -11840
rect 25194 -11874 25228 -11840
rect 24654 -11964 24688 -11930
rect 24744 -11964 24778 -11930
rect 24834 -11964 24868 -11930
rect 24924 -11964 24958 -11930
rect 25014 -11964 25048 -11930
rect 25104 -11964 25138 -11930
rect 25194 -11964 25228 -11930
rect 24654 -12054 24688 -12020
rect 24744 -12054 24778 -12020
rect 24834 -12054 24868 -12020
rect 24924 -12054 24958 -12020
rect 25014 -12054 25048 -12020
rect 25104 -12054 25138 -12020
rect 25194 -12054 25228 -12020
rect 24654 -12144 24688 -12110
rect 24744 -12144 24778 -12110
rect 24834 -12144 24868 -12110
rect 24924 -12144 24958 -12110
rect 25014 -12144 25048 -12110
rect 25104 -12144 25138 -12110
rect 25194 -12144 25228 -12110
rect 24654 -12234 24688 -12200
rect 24744 -12234 24778 -12200
rect 24834 -12234 24868 -12200
rect 24924 -12234 24958 -12200
rect 25014 -12234 25048 -12200
rect 25104 -12234 25138 -12200
rect 25194 -12234 25228 -12200
rect 25942 -11694 25976 -11660
rect 26032 -11694 26066 -11660
rect 26122 -11694 26156 -11660
rect 26212 -11694 26246 -11660
rect 26302 -11694 26336 -11660
rect 26392 -11694 26426 -11660
rect 26482 -11694 26516 -11660
rect 25942 -11784 25976 -11750
rect 26032 -11784 26066 -11750
rect 26122 -11784 26156 -11750
rect 26212 -11784 26246 -11750
rect 26302 -11784 26336 -11750
rect 26392 -11784 26426 -11750
rect 26482 -11784 26516 -11750
rect 25942 -11874 25976 -11840
rect 26032 -11874 26066 -11840
rect 26122 -11874 26156 -11840
rect 26212 -11874 26246 -11840
rect 26302 -11874 26336 -11840
rect 26392 -11874 26426 -11840
rect 26482 -11874 26516 -11840
rect 25942 -11964 25976 -11930
rect 26032 -11964 26066 -11930
rect 26122 -11964 26156 -11930
rect 26212 -11964 26246 -11930
rect 26302 -11964 26336 -11930
rect 26392 -11964 26426 -11930
rect 26482 -11964 26516 -11930
rect 25942 -12054 25976 -12020
rect 26032 -12054 26066 -12020
rect 26122 -12054 26156 -12020
rect 26212 -12054 26246 -12020
rect 26302 -12054 26336 -12020
rect 26392 -12054 26426 -12020
rect 26482 -12054 26516 -12020
rect 25942 -12144 25976 -12110
rect 26032 -12144 26066 -12110
rect 26122 -12144 26156 -12110
rect 26212 -12144 26246 -12110
rect 26302 -12144 26336 -12110
rect 26392 -12144 26426 -12110
rect 26482 -12144 26516 -12110
rect 25942 -12234 25976 -12200
rect 26032 -12234 26066 -12200
rect 26122 -12234 26156 -12200
rect 26212 -12234 26246 -12200
rect 26302 -12234 26336 -12200
rect 26392 -12234 26426 -12200
rect 26482 -12234 26516 -12200
rect 16926 -12982 16960 -12948
rect 17016 -12982 17050 -12948
rect 17106 -12982 17140 -12948
rect 17196 -12982 17230 -12948
rect 17286 -12982 17320 -12948
rect 17376 -12982 17410 -12948
rect 17466 -12982 17500 -12948
rect 16926 -13072 16960 -13038
rect 17016 -13072 17050 -13038
rect 17106 -13072 17140 -13038
rect 17196 -13072 17230 -13038
rect 17286 -13072 17320 -13038
rect 17376 -13072 17410 -13038
rect 17466 -13072 17500 -13038
rect 16926 -13162 16960 -13128
rect 17016 -13162 17050 -13128
rect 17106 -13162 17140 -13128
rect 17196 -13162 17230 -13128
rect 17286 -13162 17320 -13128
rect 17376 -13162 17410 -13128
rect 17466 -13162 17500 -13128
rect 16926 -13252 16960 -13218
rect 17016 -13252 17050 -13218
rect 17106 -13252 17140 -13218
rect 17196 -13252 17230 -13218
rect 17286 -13252 17320 -13218
rect 17376 -13252 17410 -13218
rect 17466 -13252 17500 -13218
rect 16926 -13342 16960 -13308
rect 17016 -13342 17050 -13308
rect 17106 -13342 17140 -13308
rect 17196 -13342 17230 -13308
rect 17286 -13342 17320 -13308
rect 17376 -13342 17410 -13308
rect 17466 -13342 17500 -13308
rect 16926 -13432 16960 -13398
rect 17016 -13432 17050 -13398
rect 17106 -13432 17140 -13398
rect 17196 -13432 17230 -13398
rect 17286 -13432 17320 -13398
rect 17376 -13432 17410 -13398
rect 17466 -13432 17500 -13398
rect 16926 -13522 16960 -13488
rect 17016 -13522 17050 -13488
rect 17106 -13522 17140 -13488
rect 17196 -13522 17230 -13488
rect 17286 -13522 17320 -13488
rect 17376 -13522 17410 -13488
rect 17466 -13522 17500 -13488
rect 18214 -12982 18248 -12948
rect 18304 -12982 18338 -12948
rect 18394 -12982 18428 -12948
rect 18484 -12982 18518 -12948
rect 18574 -12982 18608 -12948
rect 18664 -12982 18698 -12948
rect 18754 -12982 18788 -12948
rect 18214 -13072 18248 -13038
rect 18304 -13072 18338 -13038
rect 18394 -13072 18428 -13038
rect 18484 -13072 18518 -13038
rect 18574 -13072 18608 -13038
rect 18664 -13072 18698 -13038
rect 18754 -13072 18788 -13038
rect 18214 -13162 18248 -13128
rect 18304 -13162 18338 -13128
rect 18394 -13162 18428 -13128
rect 18484 -13162 18518 -13128
rect 18574 -13162 18608 -13128
rect 18664 -13162 18698 -13128
rect 18754 -13162 18788 -13128
rect 18214 -13252 18248 -13218
rect 18304 -13252 18338 -13218
rect 18394 -13252 18428 -13218
rect 18484 -13252 18518 -13218
rect 18574 -13252 18608 -13218
rect 18664 -13252 18698 -13218
rect 18754 -13252 18788 -13218
rect 18214 -13342 18248 -13308
rect 18304 -13342 18338 -13308
rect 18394 -13342 18428 -13308
rect 18484 -13342 18518 -13308
rect 18574 -13342 18608 -13308
rect 18664 -13342 18698 -13308
rect 18754 -13342 18788 -13308
rect 18214 -13432 18248 -13398
rect 18304 -13432 18338 -13398
rect 18394 -13432 18428 -13398
rect 18484 -13432 18518 -13398
rect 18574 -13432 18608 -13398
rect 18664 -13432 18698 -13398
rect 18754 -13432 18788 -13398
rect 18214 -13522 18248 -13488
rect 18304 -13522 18338 -13488
rect 18394 -13522 18428 -13488
rect 18484 -13522 18518 -13488
rect 18574 -13522 18608 -13488
rect 18664 -13522 18698 -13488
rect 18754 -13522 18788 -13488
rect 19502 -12982 19536 -12948
rect 19592 -12982 19626 -12948
rect 19682 -12982 19716 -12948
rect 19772 -12982 19806 -12948
rect 19862 -12982 19896 -12948
rect 19952 -12982 19986 -12948
rect 20042 -12982 20076 -12948
rect 19502 -13072 19536 -13038
rect 19592 -13072 19626 -13038
rect 19682 -13072 19716 -13038
rect 19772 -13072 19806 -13038
rect 19862 -13072 19896 -13038
rect 19952 -13072 19986 -13038
rect 20042 -13072 20076 -13038
rect 19502 -13162 19536 -13128
rect 19592 -13162 19626 -13128
rect 19682 -13162 19716 -13128
rect 19772 -13162 19806 -13128
rect 19862 -13162 19896 -13128
rect 19952 -13162 19986 -13128
rect 20042 -13162 20076 -13128
rect 19502 -13252 19536 -13218
rect 19592 -13252 19626 -13218
rect 19682 -13252 19716 -13218
rect 19772 -13252 19806 -13218
rect 19862 -13252 19896 -13218
rect 19952 -13252 19986 -13218
rect 20042 -13252 20076 -13218
rect 19502 -13342 19536 -13308
rect 19592 -13342 19626 -13308
rect 19682 -13342 19716 -13308
rect 19772 -13342 19806 -13308
rect 19862 -13342 19896 -13308
rect 19952 -13342 19986 -13308
rect 20042 -13342 20076 -13308
rect 19502 -13432 19536 -13398
rect 19592 -13432 19626 -13398
rect 19682 -13432 19716 -13398
rect 19772 -13432 19806 -13398
rect 19862 -13432 19896 -13398
rect 19952 -13432 19986 -13398
rect 20042 -13432 20076 -13398
rect 19502 -13522 19536 -13488
rect 19592 -13522 19626 -13488
rect 19682 -13522 19716 -13488
rect 19772 -13522 19806 -13488
rect 19862 -13522 19896 -13488
rect 19952 -13522 19986 -13488
rect 20042 -13522 20076 -13488
rect 20790 -12982 20824 -12948
rect 20880 -12982 20914 -12948
rect 20970 -12982 21004 -12948
rect 21060 -12982 21094 -12948
rect 21150 -12982 21184 -12948
rect 21240 -12982 21274 -12948
rect 21330 -12982 21364 -12948
rect 20790 -13072 20824 -13038
rect 20880 -13072 20914 -13038
rect 20970 -13072 21004 -13038
rect 21060 -13072 21094 -13038
rect 21150 -13072 21184 -13038
rect 21240 -13072 21274 -13038
rect 21330 -13072 21364 -13038
rect 20790 -13162 20824 -13128
rect 20880 -13162 20914 -13128
rect 20970 -13162 21004 -13128
rect 21060 -13162 21094 -13128
rect 21150 -13162 21184 -13128
rect 21240 -13162 21274 -13128
rect 21330 -13162 21364 -13128
rect 20790 -13252 20824 -13218
rect 20880 -13252 20914 -13218
rect 20970 -13252 21004 -13218
rect 21060 -13252 21094 -13218
rect 21150 -13252 21184 -13218
rect 21240 -13252 21274 -13218
rect 21330 -13252 21364 -13218
rect 20790 -13342 20824 -13308
rect 20880 -13342 20914 -13308
rect 20970 -13342 21004 -13308
rect 21060 -13342 21094 -13308
rect 21150 -13342 21184 -13308
rect 21240 -13342 21274 -13308
rect 21330 -13342 21364 -13308
rect 20790 -13432 20824 -13398
rect 20880 -13432 20914 -13398
rect 20970 -13432 21004 -13398
rect 21060 -13432 21094 -13398
rect 21150 -13432 21184 -13398
rect 21240 -13432 21274 -13398
rect 21330 -13432 21364 -13398
rect 20790 -13522 20824 -13488
rect 20880 -13522 20914 -13488
rect 20970 -13522 21004 -13488
rect 21060 -13522 21094 -13488
rect 21150 -13522 21184 -13488
rect 21240 -13522 21274 -13488
rect 21330 -13522 21364 -13488
rect 22078 -12982 22112 -12948
rect 22168 -12982 22202 -12948
rect 22258 -12982 22292 -12948
rect 22348 -12982 22382 -12948
rect 22438 -12982 22472 -12948
rect 22528 -12982 22562 -12948
rect 22618 -12982 22652 -12948
rect 22078 -13072 22112 -13038
rect 22168 -13072 22202 -13038
rect 22258 -13072 22292 -13038
rect 22348 -13072 22382 -13038
rect 22438 -13072 22472 -13038
rect 22528 -13072 22562 -13038
rect 22618 -13072 22652 -13038
rect 22078 -13162 22112 -13128
rect 22168 -13162 22202 -13128
rect 22258 -13162 22292 -13128
rect 22348 -13162 22382 -13128
rect 22438 -13162 22472 -13128
rect 22528 -13162 22562 -13128
rect 22618 -13162 22652 -13128
rect 22078 -13252 22112 -13218
rect 22168 -13252 22202 -13218
rect 22258 -13252 22292 -13218
rect 22348 -13252 22382 -13218
rect 22438 -13252 22472 -13218
rect 22528 -13252 22562 -13218
rect 22618 -13252 22652 -13218
rect 22078 -13342 22112 -13308
rect 22168 -13342 22202 -13308
rect 22258 -13342 22292 -13308
rect 22348 -13342 22382 -13308
rect 22438 -13342 22472 -13308
rect 22528 -13342 22562 -13308
rect 22618 -13342 22652 -13308
rect 22078 -13432 22112 -13398
rect 22168 -13432 22202 -13398
rect 22258 -13432 22292 -13398
rect 22348 -13432 22382 -13398
rect 22438 -13432 22472 -13398
rect 22528 -13432 22562 -13398
rect 22618 -13432 22652 -13398
rect 22078 -13522 22112 -13488
rect 22168 -13522 22202 -13488
rect 22258 -13522 22292 -13488
rect 22348 -13522 22382 -13488
rect 22438 -13522 22472 -13488
rect 22528 -13522 22562 -13488
rect 22618 -13522 22652 -13488
rect 23366 -12982 23400 -12948
rect 23456 -12982 23490 -12948
rect 23546 -12982 23580 -12948
rect 23636 -12982 23670 -12948
rect 23726 -12982 23760 -12948
rect 23816 -12982 23850 -12948
rect 23906 -12982 23940 -12948
rect 23366 -13072 23400 -13038
rect 23456 -13072 23490 -13038
rect 23546 -13072 23580 -13038
rect 23636 -13072 23670 -13038
rect 23726 -13072 23760 -13038
rect 23816 -13072 23850 -13038
rect 23906 -13072 23940 -13038
rect 23366 -13162 23400 -13128
rect 23456 -13162 23490 -13128
rect 23546 -13162 23580 -13128
rect 23636 -13162 23670 -13128
rect 23726 -13162 23760 -13128
rect 23816 -13162 23850 -13128
rect 23906 -13162 23940 -13128
rect 23366 -13252 23400 -13218
rect 23456 -13252 23490 -13218
rect 23546 -13252 23580 -13218
rect 23636 -13252 23670 -13218
rect 23726 -13252 23760 -13218
rect 23816 -13252 23850 -13218
rect 23906 -13252 23940 -13218
rect 23366 -13342 23400 -13308
rect 23456 -13342 23490 -13308
rect 23546 -13342 23580 -13308
rect 23636 -13342 23670 -13308
rect 23726 -13342 23760 -13308
rect 23816 -13342 23850 -13308
rect 23906 -13342 23940 -13308
rect 23366 -13432 23400 -13398
rect 23456 -13432 23490 -13398
rect 23546 -13432 23580 -13398
rect 23636 -13432 23670 -13398
rect 23726 -13432 23760 -13398
rect 23816 -13432 23850 -13398
rect 23906 -13432 23940 -13398
rect 23366 -13522 23400 -13488
rect 23456 -13522 23490 -13488
rect 23546 -13522 23580 -13488
rect 23636 -13522 23670 -13488
rect 23726 -13522 23760 -13488
rect 23816 -13522 23850 -13488
rect 23906 -13522 23940 -13488
rect 24654 -12982 24688 -12948
rect 24744 -12982 24778 -12948
rect 24834 -12982 24868 -12948
rect 24924 -12982 24958 -12948
rect 25014 -12982 25048 -12948
rect 25104 -12982 25138 -12948
rect 25194 -12982 25228 -12948
rect 24654 -13072 24688 -13038
rect 24744 -13072 24778 -13038
rect 24834 -13072 24868 -13038
rect 24924 -13072 24958 -13038
rect 25014 -13072 25048 -13038
rect 25104 -13072 25138 -13038
rect 25194 -13072 25228 -13038
rect 24654 -13162 24688 -13128
rect 24744 -13162 24778 -13128
rect 24834 -13162 24868 -13128
rect 24924 -13162 24958 -13128
rect 25014 -13162 25048 -13128
rect 25104 -13162 25138 -13128
rect 25194 -13162 25228 -13128
rect 24654 -13252 24688 -13218
rect 24744 -13252 24778 -13218
rect 24834 -13252 24868 -13218
rect 24924 -13252 24958 -13218
rect 25014 -13252 25048 -13218
rect 25104 -13252 25138 -13218
rect 25194 -13252 25228 -13218
rect 24654 -13342 24688 -13308
rect 24744 -13342 24778 -13308
rect 24834 -13342 24868 -13308
rect 24924 -13342 24958 -13308
rect 25014 -13342 25048 -13308
rect 25104 -13342 25138 -13308
rect 25194 -13342 25228 -13308
rect 24654 -13432 24688 -13398
rect 24744 -13432 24778 -13398
rect 24834 -13432 24868 -13398
rect 24924 -13432 24958 -13398
rect 25014 -13432 25048 -13398
rect 25104 -13432 25138 -13398
rect 25194 -13432 25228 -13398
rect 24654 -13522 24688 -13488
rect 24744 -13522 24778 -13488
rect 24834 -13522 24868 -13488
rect 24924 -13522 24958 -13488
rect 25014 -13522 25048 -13488
rect 25104 -13522 25138 -13488
rect 25194 -13522 25228 -13488
rect 25942 -12982 25976 -12948
rect 26032 -12982 26066 -12948
rect 26122 -12982 26156 -12948
rect 26212 -12982 26246 -12948
rect 26302 -12982 26336 -12948
rect 26392 -12982 26426 -12948
rect 26482 -12982 26516 -12948
rect 25942 -13072 25976 -13038
rect 26032 -13072 26066 -13038
rect 26122 -13072 26156 -13038
rect 26212 -13072 26246 -13038
rect 26302 -13072 26336 -13038
rect 26392 -13072 26426 -13038
rect 26482 -13072 26516 -13038
rect 25942 -13162 25976 -13128
rect 26032 -13162 26066 -13128
rect 26122 -13162 26156 -13128
rect 26212 -13162 26246 -13128
rect 26302 -13162 26336 -13128
rect 26392 -13162 26426 -13128
rect 26482 -13162 26516 -13128
rect 25942 -13252 25976 -13218
rect 26032 -13252 26066 -13218
rect 26122 -13252 26156 -13218
rect 26212 -13252 26246 -13218
rect 26302 -13252 26336 -13218
rect 26392 -13252 26426 -13218
rect 26482 -13252 26516 -13218
rect 25942 -13342 25976 -13308
rect 26032 -13342 26066 -13308
rect 26122 -13342 26156 -13308
rect 26212 -13342 26246 -13308
rect 26302 -13342 26336 -13308
rect 26392 -13342 26426 -13308
rect 26482 -13342 26516 -13308
rect 25942 -13432 25976 -13398
rect 26032 -13432 26066 -13398
rect 26122 -13432 26156 -13398
rect 26212 -13432 26246 -13398
rect 26302 -13432 26336 -13398
rect 26392 -13432 26426 -13398
rect 26482 -13432 26516 -13398
rect 25942 -13522 25976 -13488
rect 26032 -13522 26066 -13488
rect 26122 -13522 26156 -13488
rect 26212 -13522 26246 -13488
rect 26302 -13522 26336 -13488
rect 26392 -13522 26426 -13488
rect 26482 -13522 26516 -13488
rect 16926 -14270 16960 -14236
rect 17016 -14270 17050 -14236
rect 17106 -14270 17140 -14236
rect 17196 -14270 17230 -14236
rect 17286 -14270 17320 -14236
rect 17376 -14270 17410 -14236
rect 17466 -14270 17500 -14236
rect 16926 -14360 16960 -14326
rect 17016 -14360 17050 -14326
rect 17106 -14360 17140 -14326
rect 17196 -14360 17230 -14326
rect 17286 -14360 17320 -14326
rect 17376 -14360 17410 -14326
rect 17466 -14360 17500 -14326
rect 16926 -14450 16960 -14416
rect 17016 -14450 17050 -14416
rect 17106 -14450 17140 -14416
rect 17196 -14450 17230 -14416
rect 17286 -14450 17320 -14416
rect 17376 -14450 17410 -14416
rect 17466 -14450 17500 -14416
rect 16926 -14540 16960 -14506
rect 17016 -14540 17050 -14506
rect 17106 -14540 17140 -14506
rect 17196 -14540 17230 -14506
rect 17286 -14540 17320 -14506
rect 17376 -14540 17410 -14506
rect 17466 -14540 17500 -14506
rect 16926 -14630 16960 -14596
rect 17016 -14630 17050 -14596
rect 17106 -14630 17140 -14596
rect 17196 -14630 17230 -14596
rect 17286 -14630 17320 -14596
rect 17376 -14630 17410 -14596
rect 17466 -14630 17500 -14596
rect 16926 -14720 16960 -14686
rect 17016 -14720 17050 -14686
rect 17106 -14720 17140 -14686
rect 17196 -14720 17230 -14686
rect 17286 -14720 17320 -14686
rect 17376 -14720 17410 -14686
rect 17466 -14720 17500 -14686
rect 16926 -14810 16960 -14776
rect 17016 -14810 17050 -14776
rect 17106 -14810 17140 -14776
rect 17196 -14810 17230 -14776
rect 17286 -14810 17320 -14776
rect 17376 -14810 17410 -14776
rect 17466 -14810 17500 -14776
rect 18214 -14270 18248 -14236
rect 18304 -14270 18338 -14236
rect 18394 -14270 18428 -14236
rect 18484 -14270 18518 -14236
rect 18574 -14270 18608 -14236
rect 18664 -14270 18698 -14236
rect 18754 -14270 18788 -14236
rect 18214 -14360 18248 -14326
rect 18304 -14360 18338 -14326
rect 18394 -14360 18428 -14326
rect 18484 -14360 18518 -14326
rect 18574 -14360 18608 -14326
rect 18664 -14360 18698 -14326
rect 18754 -14360 18788 -14326
rect 18214 -14450 18248 -14416
rect 18304 -14450 18338 -14416
rect 18394 -14450 18428 -14416
rect 18484 -14450 18518 -14416
rect 18574 -14450 18608 -14416
rect 18664 -14450 18698 -14416
rect 18754 -14450 18788 -14416
rect 18214 -14540 18248 -14506
rect 18304 -14540 18338 -14506
rect 18394 -14540 18428 -14506
rect 18484 -14540 18518 -14506
rect 18574 -14540 18608 -14506
rect 18664 -14540 18698 -14506
rect 18754 -14540 18788 -14506
rect 18214 -14630 18248 -14596
rect 18304 -14630 18338 -14596
rect 18394 -14630 18428 -14596
rect 18484 -14630 18518 -14596
rect 18574 -14630 18608 -14596
rect 18664 -14630 18698 -14596
rect 18754 -14630 18788 -14596
rect 18214 -14720 18248 -14686
rect 18304 -14720 18338 -14686
rect 18394 -14720 18428 -14686
rect 18484 -14720 18518 -14686
rect 18574 -14720 18608 -14686
rect 18664 -14720 18698 -14686
rect 18754 -14720 18788 -14686
rect 18214 -14810 18248 -14776
rect 18304 -14810 18338 -14776
rect 18394 -14810 18428 -14776
rect 18484 -14810 18518 -14776
rect 18574 -14810 18608 -14776
rect 18664 -14810 18698 -14776
rect 18754 -14810 18788 -14776
rect 19502 -14270 19536 -14236
rect 19592 -14270 19626 -14236
rect 19682 -14270 19716 -14236
rect 19772 -14270 19806 -14236
rect 19862 -14270 19896 -14236
rect 19952 -14270 19986 -14236
rect 20042 -14270 20076 -14236
rect 19502 -14360 19536 -14326
rect 19592 -14360 19626 -14326
rect 19682 -14360 19716 -14326
rect 19772 -14360 19806 -14326
rect 19862 -14360 19896 -14326
rect 19952 -14360 19986 -14326
rect 20042 -14360 20076 -14326
rect 19502 -14450 19536 -14416
rect 19592 -14450 19626 -14416
rect 19682 -14450 19716 -14416
rect 19772 -14450 19806 -14416
rect 19862 -14450 19896 -14416
rect 19952 -14450 19986 -14416
rect 20042 -14450 20076 -14416
rect 19502 -14540 19536 -14506
rect 19592 -14540 19626 -14506
rect 19682 -14540 19716 -14506
rect 19772 -14540 19806 -14506
rect 19862 -14540 19896 -14506
rect 19952 -14540 19986 -14506
rect 20042 -14540 20076 -14506
rect 19502 -14630 19536 -14596
rect 19592 -14630 19626 -14596
rect 19682 -14630 19716 -14596
rect 19772 -14630 19806 -14596
rect 19862 -14630 19896 -14596
rect 19952 -14630 19986 -14596
rect 20042 -14630 20076 -14596
rect 19502 -14720 19536 -14686
rect 19592 -14720 19626 -14686
rect 19682 -14720 19716 -14686
rect 19772 -14720 19806 -14686
rect 19862 -14720 19896 -14686
rect 19952 -14720 19986 -14686
rect 20042 -14720 20076 -14686
rect 19502 -14810 19536 -14776
rect 19592 -14810 19626 -14776
rect 19682 -14810 19716 -14776
rect 19772 -14810 19806 -14776
rect 19862 -14810 19896 -14776
rect 19952 -14810 19986 -14776
rect 20042 -14810 20076 -14776
rect 20790 -14270 20824 -14236
rect 20880 -14270 20914 -14236
rect 20970 -14270 21004 -14236
rect 21060 -14270 21094 -14236
rect 21150 -14270 21184 -14236
rect 21240 -14270 21274 -14236
rect 21330 -14270 21364 -14236
rect 20790 -14360 20824 -14326
rect 20880 -14360 20914 -14326
rect 20970 -14360 21004 -14326
rect 21060 -14360 21094 -14326
rect 21150 -14360 21184 -14326
rect 21240 -14360 21274 -14326
rect 21330 -14360 21364 -14326
rect 20790 -14450 20824 -14416
rect 20880 -14450 20914 -14416
rect 20970 -14450 21004 -14416
rect 21060 -14450 21094 -14416
rect 21150 -14450 21184 -14416
rect 21240 -14450 21274 -14416
rect 21330 -14450 21364 -14416
rect 20790 -14540 20824 -14506
rect 20880 -14540 20914 -14506
rect 20970 -14540 21004 -14506
rect 21060 -14540 21094 -14506
rect 21150 -14540 21184 -14506
rect 21240 -14540 21274 -14506
rect 21330 -14540 21364 -14506
rect 20790 -14630 20824 -14596
rect 20880 -14630 20914 -14596
rect 20970 -14630 21004 -14596
rect 21060 -14630 21094 -14596
rect 21150 -14630 21184 -14596
rect 21240 -14630 21274 -14596
rect 21330 -14630 21364 -14596
rect 20790 -14720 20824 -14686
rect 20880 -14720 20914 -14686
rect 20970 -14720 21004 -14686
rect 21060 -14720 21094 -14686
rect 21150 -14720 21184 -14686
rect 21240 -14720 21274 -14686
rect 21330 -14720 21364 -14686
rect 20790 -14810 20824 -14776
rect 20880 -14810 20914 -14776
rect 20970 -14810 21004 -14776
rect 21060 -14810 21094 -14776
rect 21150 -14810 21184 -14776
rect 21240 -14810 21274 -14776
rect 21330 -14810 21364 -14776
rect 22078 -14270 22112 -14236
rect 22168 -14270 22202 -14236
rect 22258 -14270 22292 -14236
rect 22348 -14270 22382 -14236
rect 22438 -14270 22472 -14236
rect 22528 -14270 22562 -14236
rect 22618 -14270 22652 -14236
rect 22078 -14360 22112 -14326
rect 22168 -14360 22202 -14326
rect 22258 -14360 22292 -14326
rect 22348 -14360 22382 -14326
rect 22438 -14360 22472 -14326
rect 22528 -14360 22562 -14326
rect 22618 -14360 22652 -14326
rect 22078 -14450 22112 -14416
rect 22168 -14450 22202 -14416
rect 22258 -14450 22292 -14416
rect 22348 -14450 22382 -14416
rect 22438 -14450 22472 -14416
rect 22528 -14450 22562 -14416
rect 22618 -14450 22652 -14416
rect 22078 -14540 22112 -14506
rect 22168 -14540 22202 -14506
rect 22258 -14540 22292 -14506
rect 22348 -14540 22382 -14506
rect 22438 -14540 22472 -14506
rect 22528 -14540 22562 -14506
rect 22618 -14540 22652 -14506
rect 22078 -14630 22112 -14596
rect 22168 -14630 22202 -14596
rect 22258 -14630 22292 -14596
rect 22348 -14630 22382 -14596
rect 22438 -14630 22472 -14596
rect 22528 -14630 22562 -14596
rect 22618 -14630 22652 -14596
rect 22078 -14720 22112 -14686
rect 22168 -14720 22202 -14686
rect 22258 -14720 22292 -14686
rect 22348 -14720 22382 -14686
rect 22438 -14720 22472 -14686
rect 22528 -14720 22562 -14686
rect 22618 -14720 22652 -14686
rect 22078 -14810 22112 -14776
rect 22168 -14810 22202 -14776
rect 22258 -14810 22292 -14776
rect 22348 -14810 22382 -14776
rect 22438 -14810 22472 -14776
rect 22528 -14810 22562 -14776
rect 22618 -14810 22652 -14776
rect 23366 -14270 23400 -14236
rect 23456 -14270 23490 -14236
rect 23546 -14270 23580 -14236
rect 23636 -14270 23670 -14236
rect 23726 -14270 23760 -14236
rect 23816 -14270 23850 -14236
rect 23906 -14270 23940 -14236
rect 23366 -14360 23400 -14326
rect 23456 -14360 23490 -14326
rect 23546 -14360 23580 -14326
rect 23636 -14360 23670 -14326
rect 23726 -14360 23760 -14326
rect 23816 -14360 23850 -14326
rect 23906 -14360 23940 -14326
rect 23366 -14450 23400 -14416
rect 23456 -14450 23490 -14416
rect 23546 -14450 23580 -14416
rect 23636 -14450 23670 -14416
rect 23726 -14450 23760 -14416
rect 23816 -14450 23850 -14416
rect 23906 -14450 23940 -14416
rect 23366 -14540 23400 -14506
rect 23456 -14540 23490 -14506
rect 23546 -14540 23580 -14506
rect 23636 -14540 23670 -14506
rect 23726 -14540 23760 -14506
rect 23816 -14540 23850 -14506
rect 23906 -14540 23940 -14506
rect 23366 -14630 23400 -14596
rect 23456 -14630 23490 -14596
rect 23546 -14630 23580 -14596
rect 23636 -14630 23670 -14596
rect 23726 -14630 23760 -14596
rect 23816 -14630 23850 -14596
rect 23906 -14630 23940 -14596
rect 23366 -14720 23400 -14686
rect 23456 -14720 23490 -14686
rect 23546 -14720 23580 -14686
rect 23636 -14720 23670 -14686
rect 23726 -14720 23760 -14686
rect 23816 -14720 23850 -14686
rect 23906 -14720 23940 -14686
rect 23366 -14810 23400 -14776
rect 23456 -14810 23490 -14776
rect 23546 -14810 23580 -14776
rect 23636 -14810 23670 -14776
rect 23726 -14810 23760 -14776
rect 23816 -14810 23850 -14776
rect 23906 -14810 23940 -14776
rect 24654 -14270 24688 -14236
rect 24744 -14270 24778 -14236
rect 24834 -14270 24868 -14236
rect 24924 -14270 24958 -14236
rect 25014 -14270 25048 -14236
rect 25104 -14270 25138 -14236
rect 25194 -14270 25228 -14236
rect 24654 -14360 24688 -14326
rect 24744 -14360 24778 -14326
rect 24834 -14360 24868 -14326
rect 24924 -14360 24958 -14326
rect 25014 -14360 25048 -14326
rect 25104 -14360 25138 -14326
rect 25194 -14360 25228 -14326
rect 24654 -14450 24688 -14416
rect 24744 -14450 24778 -14416
rect 24834 -14450 24868 -14416
rect 24924 -14450 24958 -14416
rect 25014 -14450 25048 -14416
rect 25104 -14450 25138 -14416
rect 25194 -14450 25228 -14416
rect 24654 -14540 24688 -14506
rect 24744 -14540 24778 -14506
rect 24834 -14540 24868 -14506
rect 24924 -14540 24958 -14506
rect 25014 -14540 25048 -14506
rect 25104 -14540 25138 -14506
rect 25194 -14540 25228 -14506
rect 24654 -14630 24688 -14596
rect 24744 -14630 24778 -14596
rect 24834 -14630 24868 -14596
rect 24924 -14630 24958 -14596
rect 25014 -14630 25048 -14596
rect 25104 -14630 25138 -14596
rect 25194 -14630 25228 -14596
rect 24654 -14720 24688 -14686
rect 24744 -14720 24778 -14686
rect 24834 -14720 24868 -14686
rect 24924 -14720 24958 -14686
rect 25014 -14720 25048 -14686
rect 25104 -14720 25138 -14686
rect 25194 -14720 25228 -14686
rect 24654 -14810 24688 -14776
rect 24744 -14810 24778 -14776
rect 24834 -14810 24868 -14776
rect 24924 -14810 24958 -14776
rect 25014 -14810 25048 -14776
rect 25104 -14810 25138 -14776
rect 25194 -14810 25228 -14776
rect 25942 -14270 25976 -14236
rect 26032 -14270 26066 -14236
rect 26122 -14270 26156 -14236
rect 26212 -14270 26246 -14236
rect 26302 -14270 26336 -14236
rect 26392 -14270 26426 -14236
rect 26482 -14270 26516 -14236
rect 25942 -14360 25976 -14326
rect 26032 -14360 26066 -14326
rect 26122 -14360 26156 -14326
rect 26212 -14360 26246 -14326
rect 26302 -14360 26336 -14326
rect 26392 -14360 26426 -14326
rect 26482 -14360 26516 -14326
rect 25942 -14450 25976 -14416
rect 26032 -14450 26066 -14416
rect 26122 -14450 26156 -14416
rect 26212 -14450 26246 -14416
rect 26302 -14450 26336 -14416
rect 26392 -14450 26426 -14416
rect 26482 -14450 26516 -14416
rect 25942 -14540 25976 -14506
rect 26032 -14540 26066 -14506
rect 26122 -14540 26156 -14506
rect 26212 -14540 26246 -14506
rect 26302 -14540 26336 -14506
rect 26392 -14540 26426 -14506
rect 26482 -14540 26516 -14506
rect 25942 -14630 25976 -14596
rect 26032 -14630 26066 -14596
rect 26122 -14630 26156 -14596
rect 26212 -14630 26246 -14596
rect 26302 -14630 26336 -14596
rect 26392 -14630 26426 -14596
rect 26482 -14630 26516 -14596
rect 25942 -14720 25976 -14686
rect 26032 -14720 26066 -14686
rect 26122 -14720 26156 -14686
rect 26212 -14720 26246 -14686
rect 26302 -14720 26336 -14686
rect 26392 -14720 26426 -14686
rect 26482 -14720 26516 -14686
rect 25942 -14810 25976 -14776
rect 26032 -14810 26066 -14776
rect 26122 -14810 26156 -14776
rect 26212 -14810 26246 -14776
rect 26302 -14810 26336 -14776
rect 26392 -14810 26426 -14776
rect 26482 -14810 26516 -14776
rect 16926 -15558 16960 -15524
rect 17016 -15558 17050 -15524
rect 17106 -15558 17140 -15524
rect 17196 -15558 17230 -15524
rect 17286 -15558 17320 -15524
rect 17376 -15558 17410 -15524
rect 17466 -15558 17500 -15524
rect 16926 -15648 16960 -15614
rect 17016 -15648 17050 -15614
rect 17106 -15648 17140 -15614
rect 17196 -15648 17230 -15614
rect 17286 -15648 17320 -15614
rect 17376 -15648 17410 -15614
rect 17466 -15648 17500 -15614
rect 16926 -15738 16960 -15704
rect 17016 -15738 17050 -15704
rect 17106 -15738 17140 -15704
rect 17196 -15738 17230 -15704
rect 17286 -15738 17320 -15704
rect 17376 -15738 17410 -15704
rect 17466 -15738 17500 -15704
rect 16926 -15828 16960 -15794
rect 17016 -15828 17050 -15794
rect 17106 -15828 17140 -15794
rect 17196 -15828 17230 -15794
rect 17286 -15828 17320 -15794
rect 17376 -15828 17410 -15794
rect 17466 -15828 17500 -15794
rect 16926 -15918 16960 -15884
rect 17016 -15918 17050 -15884
rect 17106 -15918 17140 -15884
rect 17196 -15918 17230 -15884
rect 17286 -15918 17320 -15884
rect 17376 -15918 17410 -15884
rect 17466 -15918 17500 -15884
rect 16926 -16008 16960 -15974
rect 17016 -16008 17050 -15974
rect 17106 -16008 17140 -15974
rect 17196 -16008 17230 -15974
rect 17286 -16008 17320 -15974
rect 17376 -16008 17410 -15974
rect 17466 -16008 17500 -15974
rect 16926 -16098 16960 -16064
rect 17016 -16098 17050 -16064
rect 17106 -16098 17140 -16064
rect 17196 -16098 17230 -16064
rect 17286 -16098 17320 -16064
rect 17376 -16098 17410 -16064
rect 17466 -16098 17500 -16064
rect 18214 -15558 18248 -15524
rect 18304 -15558 18338 -15524
rect 18394 -15558 18428 -15524
rect 18484 -15558 18518 -15524
rect 18574 -15558 18608 -15524
rect 18664 -15558 18698 -15524
rect 18754 -15558 18788 -15524
rect 18214 -15648 18248 -15614
rect 18304 -15648 18338 -15614
rect 18394 -15648 18428 -15614
rect 18484 -15648 18518 -15614
rect 18574 -15648 18608 -15614
rect 18664 -15648 18698 -15614
rect 18754 -15648 18788 -15614
rect 18214 -15738 18248 -15704
rect 18304 -15738 18338 -15704
rect 18394 -15738 18428 -15704
rect 18484 -15738 18518 -15704
rect 18574 -15738 18608 -15704
rect 18664 -15738 18698 -15704
rect 18754 -15738 18788 -15704
rect 18214 -15828 18248 -15794
rect 18304 -15828 18338 -15794
rect 18394 -15828 18428 -15794
rect 18484 -15828 18518 -15794
rect 18574 -15828 18608 -15794
rect 18664 -15828 18698 -15794
rect 18754 -15828 18788 -15794
rect 18214 -15918 18248 -15884
rect 18304 -15918 18338 -15884
rect 18394 -15918 18428 -15884
rect 18484 -15918 18518 -15884
rect 18574 -15918 18608 -15884
rect 18664 -15918 18698 -15884
rect 18754 -15918 18788 -15884
rect 18214 -16008 18248 -15974
rect 18304 -16008 18338 -15974
rect 18394 -16008 18428 -15974
rect 18484 -16008 18518 -15974
rect 18574 -16008 18608 -15974
rect 18664 -16008 18698 -15974
rect 18754 -16008 18788 -15974
rect 18214 -16098 18248 -16064
rect 18304 -16098 18338 -16064
rect 18394 -16098 18428 -16064
rect 18484 -16098 18518 -16064
rect 18574 -16098 18608 -16064
rect 18664 -16098 18698 -16064
rect 18754 -16098 18788 -16064
rect 19502 -15558 19536 -15524
rect 19592 -15558 19626 -15524
rect 19682 -15558 19716 -15524
rect 19772 -15558 19806 -15524
rect 19862 -15558 19896 -15524
rect 19952 -15558 19986 -15524
rect 20042 -15558 20076 -15524
rect 19502 -15648 19536 -15614
rect 19592 -15648 19626 -15614
rect 19682 -15648 19716 -15614
rect 19772 -15648 19806 -15614
rect 19862 -15648 19896 -15614
rect 19952 -15648 19986 -15614
rect 20042 -15648 20076 -15614
rect 19502 -15738 19536 -15704
rect 19592 -15738 19626 -15704
rect 19682 -15738 19716 -15704
rect 19772 -15738 19806 -15704
rect 19862 -15738 19896 -15704
rect 19952 -15738 19986 -15704
rect 20042 -15738 20076 -15704
rect 19502 -15828 19536 -15794
rect 19592 -15828 19626 -15794
rect 19682 -15828 19716 -15794
rect 19772 -15828 19806 -15794
rect 19862 -15828 19896 -15794
rect 19952 -15828 19986 -15794
rect 20042 -15828 20076 -15794
rect 19502 -15918 19536 -15884
rect 19592 -15918 19626 -15884
rect 19682 -15918 19716 -15884
rect 19772 -15918 19806 -15884
rect 19862 -15918 19896 -15884
rect 19952 -15918 19986 -15884
rect 20042 -15918 20076 -15884
rect 19502 -16008 19536 -15974
rect 19592 -16008 19626 -15974
rect 19682 -16008 19716 -15974
rect 19772 -16008 19806 -15974
rect 19862 -16008 19896 -15974
rect 19952 -16008 19986 -15974
rect 20042 -16008 20076 -15974
rect 19502 -16098 19536 -16064
rect 19592 -16098 19626 -16064
rect 19682 -16098 19716 -16064
rect 19772 -16098 19806 -16064
rect 19862 -16098 19896 -16064
rect 19952 -16098 19986 -16064
rect 20042 -16098 20076 -16064
rect 20790 -15558 20824 -15524
rect 20880 -15558 20914 -15524
rect 20970 -15558 21004 -15524
rect 21060 -15558 21094 -15524
rect 21150 -15558 21184 -15524
rect 21240 -15558 21274 -15524
rect 21330 -15558 21364 -15524
rect 20790 -15648 20824 -15614
rect 20880 -15648 20914 -15614
rect 20970 -15648 21004 -15614
rect 21060 -15648 21094 -15614
rect 21150 -15648 21184 -15614
rect 21240 -15648 21274 -15614
rect 21330 -15648 21364 -15614
rect 20790 -15738 20824 -15704
rect 20880 -15738 20914 -15704
rect 20970 -15738 21004 -15704
rect 21060 -15738 21094 -15704
rect 21150 -15738 21184 -15704
rect 21240 -15738 21274 -15704
rect 21330 -15738 21364 -15704
rect 20790 -15828 20824 -15794
rect 20880 -15828 20914 -15794
rect 20970 -15828 21004 -15794
rect 21060 -15828 21094 -15794
rect 21150 -15828 21184 -15794
rect 21240 -15828 21274 -15794
rect 21330 -15828 21364 -15794
rect 20790 -15918 20824 -15884
rect 20880 -15918 20914 -15884
rect 20970 -15918 21004 -15884
rect 21060 -15918 21094 -15884
rect 21150 -15918 21184 -15884
rect 21240 -15918 21274 -15884
rect 21330 -15918 21364 -15884
rect 20790 -16008 20824 -15974
rect 20880 -16008 20914 -15974
rect 20970 -16008 21004 -15974
rect 21060 -16008 21094 -15974
rect 21150 -16008 21184 -15974
rect 21240 -16008 21274 -15974
rect 21330 -16008 21364 -15974
rect 20790 -16098 20824 -16064
rect 20880 -16098 20914 -16064
rect 20970 -16098 21004 -16064
rect 21060 -16098 21094 -16064
rect 21150 -16098 21184 -16064
rect 21240 -16098 21274 -16064
rect 21330 -16098 21364 -16064
rect 22078 -15558 22112 -15524
rect 22168 -15558 22202 -15524
rect 22258 -15558 22292 -15524
rect 22348 -15558 22382 -15524
rect 22438 -15558 22472 -15524
rect 22528 -15558 22562 -15524
rect 22618 -15558 22652 -15524
rect 22078 -15648 22112 -15614
rect 22168 -15648 22202 -15614
rect 22258 -15648 22292 -15614
rect 22348 -15648 22382 -15614
rect 22438 -15648 22472 -15614
rect 22528 -15648 22562 -15614
rect 22618 -15648 22652 -15614
rect 22078 -15738 22112 -15704
rect 22168 -15738 22202 -15704
rect 22258 -15738 22292 -15704
rect 22348 -15738 22382 -15704
rect 22438 -15738 22472 -15704
rect 22528 -15738 22562 -15704
rect 22618 -15738 22652 -15704
rect 22078 -15828 22112 -15794
rect 22168 -15828 22202 -15794
rect 22258 -15828 22292 -15794
rect 22348 -15828 22382 -15794
rect 22438 -15828 22472 -15794
rect 22528 -15828 22562 -15794
rect 22618 -15828 22652 -15794
rect 22078 -15918 22112 -15884
rect 22168 -15918 22202 -15884
rect 22258 -15918 22292 -15884
rect 22348 -15918 22382 -15884
rect 22438 -15918 22472 -15884
rect 22528 -15918 22562 -15884
rect 22618 -15918 22652 -15884
rect 22078 -16008 22112 -15974
rect 22168 -16008 22202 -15974
rect 22258 -16008 22292 -15974
rect 22348 -16008 22382 -15974
rect 22438 -16008 22472 -15974
rect 22528 -16008 22562 -15974
rect 22618 -16008 22652 -15974
rect 22078 -16098 22112 -16064
rect 22168 -16098 22202 -16064
rect 22258 -16098 22292 -16064
rect 22348 -16098 22382 -16064
rect 22438 -16098 22472 -16064
rect 22528 -16098 22562 -16064
rect 22618 -16098 22652 -16064
rect 23366 -15558 23400 -15524
rect 23456 -15558 23490 -15524
rect 23546 -15558 23580 -15524
rect 23636 -15558 23670 -15524
rect 23726 -15558 23760 -15524
rect 23816 -15558 23850 -15524
rect 23906 -15558 23940 -15524
rect 23366 -15648 23400 -15614
rect 23456 -15648 23490 -15614
rect 23546 -15648 23580 -15614
rect 23636 -15648 23670 -15614
rect 23726 -15648 23760 -15614
rect 23816 -15648 23850 -15614
rect 23906 -15648 23940 -15614
rect 23366 -15738 23400 -15704
rect 23456 -15738 23490 -15704
rect 23546 -15738 23580 -15704
rect 23636 -15738 23670 -15704
rect 23726 -15738 23760 -15704
rect 23816 -15738 23850 -15704
rect 23906 -15738 23940 -15704
rect 23366 -15828 23400 -15794
rect 23456 -15828 23490 -15794
rect 23546 -15828 23580 -15794
rect 23636 -15828 23670 -15794
rect 23726 -15828 23760 -15794
rect 23816 -15828 23850 -15794
rect 23906 -15828 23940 -15794
rect 23366 -15918 23400 -15884
rect 23456 -15918 23490 -15884
rect 23546 -15918 23580 -15884
rect 23636 -15918 23670 -15884
rect 23726 -15918 23760 -15884
rect 23816 -15918 23850 -15884
rect 23906 -15918 23940 -15884
rect 23366 -16008 23400 -15974
rect 23456 -16008 23490 -15974
rect 23546 -16008 23580 -15974
rect 23636 -16008 23670 -15974
rect 23726 -16008 23760 -15974
rect 23816 -16008 23850 -15974
rect 23906 -16008 23940 -15974
rect 23366 -16098 23400 -16064
rect 23456 -16098 23490 -16064
rect 23546 -16098 23580 -16064
rect 23636 -16098 23670 -16064
rect 23726 -16098 23760 -16064
rect 23816 -16098 23850 -16064
rect 23906 -16098 23940 -16064
rect 24654 -15558 24688 -15524
rect 24744 -15558 24778 -15524
rect 24834 -15558 24868 -15524
rect 24924 -15558 24958 -15524
rect 25014 -15558 25048 -15524
rect 25104 -15558 25138 -15524
rect 25194 -15558 25228 -15524
rect 24654 -15648 24688 -15614
rect 24744 -15648 24778 -15614
rect 24834 -15648 24868 -15614
rect 24924 -15648 24958 -15614
rect 25014 -15648 25048 -15614
rect 25104 -15648 25138 -15614
rect 25194 -15648 25228 -15614
rect 24654 -15738 24688 -15704
rect 24744 -15738 24778 -15704
rect 24834 -15738 24868 -15704
rect 24924 -15738 24958 -15704
rect 25014 -15738 25048 -15704
rect 25104 -15738 25138 -15704
rect 25194 -15738 25228 -15704
rect 24654 -15828 24688 -15794
rect 24744 -15828 24778 -15794
rect 24834 -15828 24868 -15794
rect 24924 -15828 24958 -15794
rect 25014 -15828 25048 -15794
rect 25104 -15828 25138 -15794
rect 25194 -15828 25228 -15794
rect 24654 -15918 24688 -15884
rect 24744 -15918 24778 -15884
rect 24834 -15918 24868 -15884
rect 24924 -15918 24958 -15884
rect 25014 -15918 25048 -15884
rect 25104 -15918 25138 -15884
rect 25194 -15918 25228 -15884
rect 24654 -16008 24688 -15974
rect 24744 -16008 24778 -15974
rect 24834 -16008 24868 -15974
rect 24924 -16008 24958 -15974
rect 25014 -16008 25048 -15974
rect 25104 -16008 25138 -15974
rect 25194 -16008 25228 -15974
rect 24654 -16098 24688 -16064
rect 24744 -16098 24778 -16064
rect 24834 -16098 24868 -16064
rect 24924 -16098 24958 -16064
rect 25014 -16098 25048 -16064
rect 25104 -16098 25138 -16064
rect 25194 -16098 25228 -16064
rect 25942 -15558 25976 -15524
rect 26032 -15558 26066 -15524
rect 26122 -15558 26156 -15524
rect 26212 -15558 26246 -15524
rect 26302 -15558 26336 -15524
rect 26392 -15558 26426 -15524
rect 26482 -15558 26516 -15524
rect 25942 -15648 25976 -15614
rect 26032 -15648 26066 -15614
rect 26122 -15648 26156 -15614
rect 26212 -15648 26246 -15614
rect 26302 -15648 26336 -15614
rect 26392 -15648 26426 -15614
rect 26482 -15648 26516 -15614
rect 25942 -15738 25976 -15704
rect 26032 -15738 26066 -15704
rect 26122 -15738 26156 -15704
rect 26212 -15738 26246 -15704
rect 26302 -15738 26336 -15704
rect 26392 -15738 26426 -15704
rect 26482 -15738 26516 -15704
rect 25942 -15828 25976 -15794
rect 26032 -15828 26066 -15794
rect 26122 -15828 26156 -15794
rect 26212 -15828 26246 -15794
rect 26302 -15828 26336 -15794
rect 26392 -15828 26426 -15794
rect 26482 -15828 26516 -15794
rect 25942 -15918 25976 -15884
rect 26032 -15918 26066 -15884
rect 26122 -15918 26156 -15884
rect 26212 -15918 26246 -15884
rect 26302 -15918 26336 -15884
rect 26392 -15918 26426 -15884
rect 26482 -15918 26516 -15884
rect 25942 -16008 25976 -15974
rect 26032 -16008 26066 -15974
rect 26122 -16008 26156 -15974
rect 26212 -16008 26246 -15974
rect 26302 -16008 26336 -15974
rect 26392 -16008 26426 -15974
rect 26482 -16008 26516 -15974
rect 25942 -16098 25976 -16064
rect 26032 -16098 26066 -16064
rect 26122 -16098 26156 -16064
rect 26212 -16098 26246 -16064
rect 26302 -16098 26336 -16064
rect 26392 -16098 26426 -16064
rect 26482 -16098 26516 -16064
rect 16926 -16846 16960 -16812
rect 17016 -16846 17050 -16812
rect 17106 -16846 17140 -16812
rect 17196 -16846 17230 -16812
rect 17286 -16846 17320 -16812
rect 17376 -16846 17410 -16812
rect 17466 -16846 17500 -16812
rect 16926 -16936 16960 -16902
rect 17016 -16936 17050 -16902
rect 17106 -16936 17140 -16902
rect 17196 -16936 17230 -16902
rect 17286 -16936 17320 -16902
rect 17376 -16936 17410 -16902
rect 17466 -16936 17500 -16902
rect 16926 -17026 16960 -16992
rect 17016 -17026 17050 -16992
rect 17106 -17026 17140 -16992
rect 17196 -17026 17230 -16992
rect 17286 -17026 17320 -16992
rect 17376 -17026 17410 -16992
rect 17466 -17026 17500 -16992
rect 16926 -17116 16960 -17082
rect 17016 -17116 17050 -17082
rect 17106 -17116 17140 -17082
rect 17196 -17116 17230 -17082
rect 17286 -17116 17320 -17082
rect 17376 -17116 17410 -17082
rect 17466 -17116 17500 -17082
rect 16926 -17206 16960 -17172
rect 17016 -17206 17050 -17172
rect 17106 -17206 17140 -17172
rect 17196 -17206 17230 -17172
rect 17286 -17206 17320 -17172
rect 17376 -17206 17410 -17172
rect 17466 -17206 17500 -17172
rect 16926 -17296 16960 -17262
rect 17016 -17296 17050 -17262
rect 17106 -17296 17140 -17262
rect 17196 -17296 17230 -17262
rect 17286 -17296 17320 -17262
rect 17376 -17296 17410 -17262
rect 17466 -17296 17500 -17262
rect 16926 -17386 16960 -17352
rect 17016 -17386 17050 -17352
rect 17106 -17386 17140 -17352
rect 17196 -17386 17230 -17352
rect 17286 -17386 17320 -17352
rect 17376 -17386 17410 -17352
rect 17466 -17386 17500 -17352
rect 18214 -16846 18248 -16812
rect 18304 -16846 18338 -16812
rect 18394 -16846 18428 -16812
rect 18484 -16846 18518 -16812
rect 18574 -16846 18608 -16812
rect 18664 -16846 18698 -16812
rect 18754 -16846 18788 -16812
rect 18214 -16936 18248 -16902
rect 18304 -16936 18338 -16902
rect 18394 -16936 18428 -16902
rect 18484 -16936 18518 -16902
rect 18574 -16936 18608 -16902
rect 18664 -16936 18698 -16902
rect 18754 -16936 18788 -16902
rect 18214 -17026 18248 -16992
rect 18304 -17026 18338 -16992
rect 18394 -17026 18428 -16992
rect 18484 -17026 18518 -16992
rect 18574 -17026 18608 -16992
rect 18664 -17026 18698 -16992
rect 18754 -17026 18788 -16992
rect 18214 -17116 18248 -17082
rect 18304 -17116 18338 -17082
rect 18394 -17116 18428 -17082
rect 18484 -17116 18518 -17082
rect 18574 -17116 18608 -17082
rect 18664 -17116 18698 -17082
rect 18754 -17116 18788 -17082
rect 18214 -17206 18248 -17172
rect 18304 -17206 18338 -17172
rect 18394 -17206 18428 -17172
rect 18484 -17206 18518 -17172
rect 18574 -17206 18608 -17172
rect 18664 -17206 18698 -17172
rect 18754 -17206 18788 -17172
rect 18214 -17296 18248 -17262
rect 18304 -17296 18338 -17262
rect 18394 -17296 18428 -17262
rect 18484 -17296 18518 -17262
rect 18574 -17296 18608 -17262
rect 18664 -17296 18698 -17262
rect 18754 -17296 18788 -17262
rect 18214 -17386 18248 -17352
rect 18304 -17386 18338 -17352
rect 18394 -17386 18428 -17352
rect 18484 -17386 18518 -17352
rect 18574 -17386 18608 -17352
rect 18664 -17386 18698 -17352
rect 18754 -17386 18788 -17352
rect 19502 -16846 19536 -16812
rect 19592 -16846 19626 -16812
rect 19682 -16846 19716 -16812
rect 19772 -16846 19806 -16812
rect 19862 -16846 19896 -16812
rect 19952 -16846 19986 -16812
rect 20042 -16846 20076 -16812
rect 19502 -16936 19536 -16902
rect 19592 -16936 19626 -16902
rect 19682 -16936 19716 -16902
rect 19772 -16936 19806 -16902
rect 19862 -16936 19896 -16902
rect 19952 -16936 19986 -16902
rect 20042 -16936 20076 -16902
rect 19502 -17026 19536 -16992
rect 19592 -17026 19626 -16992
rect 19682 -17026 19716 -16992
rect 19772 -17026 19806 -16992
rect 19862 -17026 19896 -16992
rect 19952 -17026 19986 -16992
rect 20042 -17026 20076 -16992
rect 19502 -17116 19536 -17082
rect 19592 -17116 19626 -17082
rect 19682 -17116 19716 -17082
rect 19772 -17116 19806 -17082
rect 19862 -17116 19896 -17082
rect 19952 -17116 19986 -17082
rect 20042 -17116 20076 -17082
rect 19502 -17206 19536 -17172
rect 19592 -17206 19626 -17172
rect 19682 -17206 19716 -17172
rect 19772 -17206 19806 -17172
rect 19862 -17206 19896 -17172
rect 19952 -17206 19986 -17172
rect 20042 -17206 20076 -17172
rect 19502 -17296 19536 -17262
rect 19592 -17296 19626 -17262
rect 19682 -17296 19716 -17262
rect 19772 -17296 19806 -17262
rect 19862 -17296 19896 -17262
rect 19952 -17296 19986 -17262
rect 20042 -17296 20076 -17262
rect 19502 -17386 19536 -17352
rect 19592 -17386 19626 -17352
rect 19682 -17386 19716 -17352
rect 19772 -17386 19806 -17352
rect 19862 -17386 19896 -17352
rect 19952 -17386 19986 -17352
rect 20042 -17386 20076 -17352
rect 20790 -16846 20824 -16812
rect 20880 -16846 20914 -16812
rect 20970 -16846 21004 -16812
rect 21060 -16846 21094 -16812
rect 21150 -16846 21184 -16812
rect 21240 -16846 21274 -16812
rect 21330 -16846 21364 -16812
rect 20790 -16936 20824 -16902
rect 20880 -16936 20914 -16902
rect 20970 -16936 21004 -16902
rect 21060 -16936 21094 -16902
rect 21150 -16936 21184 -16902
rect 21240 -16936 21274 -16902
rect 21330 -16936 21364 -16902
rect 20790 -17026 20824 -16992
rect 20880 -17026 20914 -16992
rect 20970 -17026 21004 -16992
rect 21060 -17026 21094 -16992
rect 21150 -17026 21184 -16992
rect 21240 -17026 21274 -16992
rect 21330 -17026 21364 -16992
rect 20790 -17116 20824 -17082
rect 20880 -17116 20914 -17082
rect 20970 -17116 21004 -17082
rect 21060 -17116 21094 -17082
rect 21150 -17116 21184 -17082
rect 21240 -17116 21274 -17082
rect 21330 -17116 21364 -17082
rect 20790 -17206 20824 -17172
rect 20880 -17206 20914 -17172
rect 20970 -17206 21004 -17172
rect 21060 -17206 21094 -17172
rect 21150 -17206 21184 -17172
rect 21240 -17206 21274 -17172
rect 21330 -17206 21364 -17172
rect 20790 -17296 20824 -17262
rect 20880 -17296 20914 -17262
rect 20970 -17296 21004 -17262
rect 21060 -17296 21094 -17262
rect 21150 -17296 21184 -17262
rect 21240 -17296 21274 -17262
rect 21330 -17296 21364 -17262
rect 20790 -17386 20824 -17352
rect 20880 -17386 20914 -17352
rect 20970 -17386 21004 -17352
rect 21060 -17386 21094 -17352
rect 21150 -17386 21184 -17352
rect 21240 -17386 21274 -17352
rect 21330 -17386 21364 -17352
rect 22078 -16846 22112 -16812
rect 22168 -16846 22202 -16812
rect 22258 -16846 22292 -16812
rect 22348 -16846 22382 -16812
rect 22438 -16846 22472 -16812
rect 22528 -16846 22562 -16812
rect 22618 -16846 22652 -16812
rect 22078 -16936 22112 -16902
rect 22168 -16936 22202 -16902
rect 22258 -16936 22292 -16902
rect 22348 -16936 22382 -16902
rect 22438 -16936 22472 -16902
rect 22528 -16936 22562 -16902
rect 22618 -16936 22652 -16902
rect 22078 -17026 22112 -16992
rect 22168 -17026 22202 -16992
rect 22258 -17026 22292 -16992
rect 22348 -17026 22382 -16992
rect 22438 -17026 22472 -16992
rect 22528 -17026 22562 -16992
rect 22618 -17026 22652 -16992
rect 22078 -17116 22112 -17082
rect 22168 -17116 22202 -17082
rect 22258 -17116 22292 -17082
rect 22348 -17116 22382 -17082
rect 22438 -17116 22472 -17082
rect 22528 -17116 22562 -17082
rect 22618 -17116 22652 -17082
rect 22078 -17206 22112 -17172
rect 22168 -17206 22202 -17172
rect 22258 -17206 22292 -17172
rect 22348 -17206 22382 -17172
rect 22438 -17206 22472 -17172
rect 22528 -17206 22562 -17172
rect 22618 -17206 22652 -17172
rect 22078 -17296 22112 -17262
rect 22168 -17296 22202 -17262
rect 22258 -17296 22292 -17262
rect 22348 -17296 22382 -17262
rect 22438 -17296 22472 -17262
rect 22528 -17296 22562 -17262
rect 22618 -17296 22652 -17262
rect 22078 -17386 22112 -17352
rect 22168 -17386 22202 -17352
rect 22258 -17386 22292 -17352
rect 22348 -17386 22382 -17352
rect 22438 -17386 22472 -17352
rect 22528 -17386 22562 -17352
rect 22618 -17386 22652 -17352
rect 23366 -16846 23400 -16812
rect 23456 -16846 23490 -16812
rect 23546 -16846 23580 -16812
rect 23636 -16846 23670 -16812
rect 23726 -16846 23760 -16812
rect 23816 -16846 23850 -16812
rect 23906 -16846 23940 -16812
rect 23366 -16936 23400 -16902
rect 23456 -16936 23490 -16902
rect 23546 -16936 23580 -16902
rect 23636 -16936 23670 -16902
rect 23726 -16936 23760 -16902
rect 23816 -16936 23850 -16902
rect 23906 -16936 23940 -16902
rect 23366 -17026 23400 -16992
rect 23456 -17026 23490 -16992
rect 23546 -17026 23580 -16992
rect 23636 -17026 23670 -16992
rect 23726 -17026 23760 -16992
rect 23816 -17026 23850 -16992
rect 23906 -17026 23940 -16992
rect 23366 -17116 23400 -17082
rect 23456 -17116 23490 -17082
rect 23546 -17116 23580 -17082
rect 23636 -17116 23670 -17082
rect 23726 -17116 23760 -17082
rect 23816 -17116 23850 -17082
rect 23906 -17116 23940 -17082
rect 23366 -17206 23400 -17172
rect 23456 -17206 23490 -17172
rect 23546 -17206 23580 -17172
rect 23636 -17206 23670 -17172
rect 23726 -17206 23760 -17172
rect 23816 -17206 23850 -17172
rect 23906 -17206 23940 -17172
rect 23366 -17296 23400 -17262
rect 23456 -17296 23490 -17262
rect 23546 -17296 23580 -17262
rect 23636 -17296 23670 -17262
rect 23726 -17296 23760 -17262
rect 23816 -17296 23850 -17262
rect 23906 -17296 23940 -17262
rect 23366 -17386 23400 -17352
rect 23456 -17386 23490 -17352
rect 23546 -17386 23580 -17352
rect 23636 -17386 23670 -17352
rect 23726 -17386 23760 -17352
rect 23816 -17386 23850 -17352
rect 23906 -17386 23940 -17352
rect 24654 -16846 24688 -16812
rect 24744 -16846 24778 -16812
rect 24834 -16846 24868 -16812
rect 24924 -16846 24958 -16812
rect 25014 -16846 25048 -16812
rect 25104 -16846 25138 -16812
rect 25194 -16846 25228 -16812
rect 24654 -16936 24688 -16902
rect 24744 -16936 24778 -16902
rect 24834 -16936 24868 -16902
rect 24924 -16936 24958 -16902
rect 25014 -16936 25048 -16902
rect 25104 -16936 25138 -16902
rect 25194 -16936 25228 -16902
rect 24654 -17026 24688 -16992
rect 24744 -17026 24778 -16992
rect 24834 -17026 24868 -16992
rect 24924 -17026 24958 -16992
rect 25014 -17026 25048 -16992
rect 25104 -17026 25138 -16992
rect 25194 -17026 25228 -16992
rect 24654 -17116 24688 -17082
rect 24744 -17116 24778 -17082
rect 24834 -17116 24868 -17082
rect 24924 -17116 24958 -17082
rect 25014 -17116 25048 -17082
rect 25104 -17116 25138 -17082
rect 25194 -17116 25228 -17082
rect 24654 -17206 24688 -17172
rect 24744 -17206 24778 -17172
rect 24834 -17206 24868 -17172
rect 24924 -17206 24958 -17172
rect 25014 -17206 25048 -17172
rect 25104 -17206 25138 -17172
rect 25194 -17206 25228 -17172
rect 24654 -17296 24688 -17262
rect 24744 -17296 24778 -17262
rect 24834 -17296 24868 -17262
rect 24924 -17296 24958 -17262
rect 25014 -17296 25048 -17262
rect 25104 -17296 25138 -17262
rect 25194 -17296 25228 -17262
rect 24654 -17386 24688 -17352
rect 24744 -17386 24778 -17352
rect 24834 -17386 24868 -17352
rect 24924 -17386 24958 -17352
rect 25014 -17386 25048 -17352
rect 25104 -17386 25138 -17352
rect 25194 -17386 25228 -17352
rect 25942 -16846 25976 -16811
rect 26032 -16846 26066 -16811
rect 26122 -16846 26156 -16811
rect 26212 -16846 26246 -16811
rect 26302 -16846 26336 -16811
rect 26392 -16846 26426 -16811
rect 26482 -16846 26516 -16811
rect 25942 -16936 25976 -16901
rect 26032 -16936 26066 -16901
rect 26122 -16936 26156 -16901
rect 26212 -16936 26246 -16901
rect 26302 -16936 26336 -16901
rect 26392 -16936 26426 -16901
rect 26482 -16936 26516 -16901
rect 25942 -17026 25976 -16991
rect 26032 -17026 26066 -16991
rect 26122 -17026 26156 -16991
rect 26212 -17026 26246 -16991
rect 26302 -17026 26336 -16991
rect 26392 -17026 26426 -16991
rect 26482 -17026 26516 -16991
rect 25942 -17116 25976 -17081
rect 26032 -17116 26066 -17081
rect 26122 -17116 26156 -17081
rect 26212 -17116 26246 -17081
rect 26302 -17116 26336 -17081
rect 26392 -17116 26426 -17081
rect 26482 -17116 26516 -17081
rect 25942 -17206 25976 -17171
rect 26032 -17206 26066 -17171
rect 26122 -17206 26156 -17171
rect 26212 -17206 26246 -17171
rect 26302 -17206 26336 -17171
rect 26392 -17206 26426 -17171
rect 26482 -17206 26516 -17171
rect 25942 -17296 25976 -17261
rect 26032 -17296 26066 -17261
rect 26122 -17296 26156 -17261
rect 26212 -17296 26246 -17261
rect 26302 -17296 26336 -17261
rect 26392 -17296 26426 -17261
rect 26482 -17296 26516 -17261
rect 25942 -17386 25976 -17351
rect 26032 -17386 26066 -17351
rect 26122 -17386 26156 -17351
rect 26212 -17386 26246 -17351
rect 26302 -17386 26336 -17351
rect 26392 -17386 26426 -17351
rect 26482 -17386 26516 -17351
<< psubdiff >>
rect 16568 -11336 26872 -11302
rect 16568 -11370 16684 -11336
rect 16718 -11370 16774 -11336
rect 16808 -11370 16864 -11336
rect 16898 -11370 16954 -11336
rect 16988 -11370 17044 -11336
rect 17078 -11370 17134 -11336
rect 17168 -11370 17224 -11336
rect 17258 -11370 17314 -11336
rect 17348 -11370 17404 -11336
rect 17438 -11370 17494 -11336
rect 17528 -11370 17584 -11336
rect 17618 -11370 17674 -11336
rect 17708 -11370 17764 -11336
rect 17798 -11370 17972 -11336
rect 18006 -11370 18062 -11336
rect 18096 -11370 18152 -11336
rect 18186 -11370 18242 -11336
rect 18276 -11370 18332 -11336
rect 18366 -11370 18422 -11336
rect 18456 -11370 18512 -11336
rect 18546 -11370 18602 -11336
rect 18636 -11370 18692 -11336
rect 18726 -11370 18782 -11336
rect 18816 -11370 18872 -11336
rect 18906 -11370 18962 -11336
rect 18996 -11370 19052 -11336
rect 19086 -11370 19260 -11336
rect 19294 -11370 19350 -11336
rect 19384 -11370 19440 -11336
rect 19474 -11370 19530 -11336
rect 19564 -11370 19620 -11336
rect 19654 -11370 19710 -11336
rect 19744 -11370 19800 -11336
rect 19834 -11370 19890 -11336
rect 19924 -11370 19980 -11336
rect 20014 -11370 20070 -11336
rect 20104 -11370 20160 -11336
rect 20194 -11370 20250 -11336
rect 20284 -11370 20340 -11336
rect 20374 -11370 20548 -11336
rect 20582 -11370 20638 -11336
rect 20672 -11370 20728 -11336
rect 20762 -11370 20818 -11336
rect 20852 -11370 20908 -11336
rect 20942 -11370 20998 -11336
rect 21032 -11370 21088 -11336
rect 21122 -11370 21178 -11336
rect 21212 -11370 21268 -11336
rect 21302 -11370 21358 -11336
rect 21392 -11370 21448 -11336
rect 21482 -11370 21538 -11336
rect 21572 -11370 21628 -11336
rect 21662 -11370 21836 -11336
rect 21870 -11370 21926 -11336
rect 21960 -11370 22016 -11336
rect 22050 -11370 22106 -11336
rect 22140 -11370 22196 -11336
rect 22230 -11370 22286 -11336
rect 22320 -11370 22376 -11336
rect 22410 -11370 22466 -11336
rect 22500 -11370 22556 -11336
rect 22590 -11370 22646 -11336
rect 22680 -11370 22736 -11336
rect 22770 -11370 22826 -11336
rect 22860 -11370 22916 -11336
rect 22950 -11370 23124 -11336
rect 23158 -11370 23214 -11336
rect 23248 -11370 23304 -11336
rect 23338 -11370 23394 -11336
rect 23428 -11370 23484 -11336
rect 23518 -11370 23574 -11336
rect 23608 -11370 23664 -11336
rect 23698 -11370 23754 -11336
rect 23788 -11370 23844 -11336
rect 23878 -11370 23934 -11336
rect 23968 -11370 24024 -11336
rect 24058 -11370 24114 -11336
rect 24148 -11370 24204 -11336
rect 24238 -11370 24412 -11336
rect 24446 -11370 24502 -11336
rect 24536 -11370 24592 -11336
rect 24626 -11370 24682 -11336
rect 24716 -11370 24772 -11336
rect 24806 -11370 24862 -11336
rect 24896 -11370 24952 -11336
rect 24986 -11370 25042 -11336
rect 25076 -11370 25132 -11336
rect 25166 -11370 25222 -11336
rect 25256 -11370 25312 -11336
rect 25346 -11370 25402 -11336
rect 25436 -11370 25492 -11336
rect 25526 -11370 25700 -11336
rect 25734 -11370 25790 -11336
rect 25824 -11370 25880 -11336
rect 25914 -11370 25970 -11336
rect 26004 -11370 26060 -11336
rect 26094 -11370 26150 -11336
rect 26184 -11370 26240 -11336
rect 26274 -11370 26330 -11336
rect 26364 -11370 26420 -11336
rect 26454 -11370 26510 -11336
rect 26544 -11370 26600 -11336
rect 26634 -11370 26690 -11336
rect 26724 -11370 26780 -11336
rect 26814 -11370 26872 -11336
rect 16568 -11403 26872 -11370
rect 16568 -11432 16669 -11403
rect 16568 -11466 16600 -11432
rect 16634 -11466 16669 -11432
rect 17755 -11432 17957 -11403
rect 16568 -11522 16669 -11466
rect 16568 -11556 16600 -11522
rect 16634 -11556 16669 -11522
rect 16568 -11612 16669 -11556
rect 16568 -11646 16600 -11612
rect 16634 -11646 16669 -11612
rect 16568 -11702 16669 -11646
rect 16568 -11736 16600 -11702
rect 16634 -11736 16669 -11702
rect 16568 -11792 16669 -11736
rect 16568 -11826 16600 -11792
rect 16634 -11826 16669 -11792
rect 16568 -11882 16669 -11826
rect 16568 -11916 16600 -11882
rect 16634 -11916 16669 -11882
rect 16568 -11972 16669 -11916
rect 16568 -12006 16600 -11972
rect 16634 -12006 16669 -11972
rect 16568 -12062 16669 -12006
rect 16568 -12096 16600 -12062
rect 16634 -12096 16669 -12062
rect 16568 -12152 16669 -12096
rect 16568 -12186 16600 -12152
rect 16634 -12186 16669 -12152
rect 16568 -12242 16669 -12186
rect 16568 -12276 16600 -12242
rect 16634 -12276 16669 -12242
rect 16568 -12332 16669 -12276
rect 16568 -12366 16600 -12332
rect 16634 -12366 16669 -12332
rect 16568 -12422 16669 -12366
rect 16568 -12456 16600 -12422
rect 16634 -12456 16669 -12422
rect 17755 -11466 17787 -11432
rect 17821 -11466 17888 -11432
rect 17922 -11466 17957 -11432
rect 19043 -11432 19245 -11403
rect 17755 -11522 17957 -11466
rect 17755 -11556 17787 -11522
rect 17821 -11556 17888 -11522
rect 17922 -11556 17957 -11522
rect 17755 -11612 17957 -11556
rect 17755 -11646 17787 -11612
rect 17821 -11646 17888 -11612
rect 17922 -11646 17957 -11612
rect 17755 -11702 17957 -11646
rect 17755 -11736 17787 -11702
rect 17821 -11736 17888 -11702
rect 17922 -11736 17957 -11702
rect 17755 -11792 17957 -11736
rect 17755 -11826 17787 -11792
rect 17821 -11826 17888 -11792
rect 17922 -11826 17957 -11792
rect 17755 -11882 17957 -11826
rect 17755 -11916 17787 -11882
rect 17821 -11916 17888 -11882
rect 17922 -11916 17957 -11882
rect 17755 -11972 17957 -11916
rect 17755 -12006 17787 -11972
rect 17821 -12006 17888 -11972
rect 17922 -12006 17957 -11972
rect 17755 -12062 17957 -12006
rect 17755 -12096 17787 -12062
rect 17821 -12096 17888 -12062
rect 17922 -12096 17957 -12062
rect 17755 -12152 17957 -12096
rect 17755 -12186 17787 -12152
rect 17821 -12186 17888 -12152
rect 17922 -12186 17957 -12152
rect 17755 -12242 17957 -12186
rect 17755 -12276 17787 -12242
rect 17821 -12276 17888 -12242
rect 17922 -12276 17957 -12242
rect 17755 -12332 17957 -12276
rect 17755 -12366 17787 -12332
rect 17821 -12366 17888 -12332
rect 17922 -12366 17957 -12332
rect 17755 -12422 17957 -12366
rect 16568 -12489 16669 -12456
rect 17755 -12456 17787 -12422
rect 17821 -12456 17888 -12422
rect 17922 -12456 17957 -12422
rect 19043 -11466 19075 -11432
rect 19109 -11466 19176 -11432
rect 19210 -11466 19245 -11432
rect 20331 -11432 20533 -11403
rect 19043 -11522 19245 -11466
rect 19043 -11556 19075 -11522
rect 19109 -11556 19176 -11522
rect 19210 -11556 19245 -11522
rect 19043 -11612 19245 -11556
rect 19043 -11646 19075 -11612
rect 19109 -11646 19176 -11612
rect 19210 -11646 19245 -11612
rect 19043 -11702 19245 -11646
rect 19043 -11736 19075 -11702
rect 19109 -11736 19176 -11702
rect 19210 -11736 19245 -11702
rect 19043 -11792 19245 -11736
rect 19043 -11826 19075 -11792
rect 19109 -11826 19176 -11792
rect 19210 -11826 19245 -11792
rect 19043 -11882 19245 -11826
rect 19043 -11916 19075 -11882
rect 19109 -11916 19176 -11882
rect 19210 -11916 19245 -11882
rect 19043 -11972 19245 -11916
rect 19043 -12006 19075 -11972
rect 19109 -12006 19176 -11972
rect 19210 -12006 19245 -11972
rect 19043 -12062 19245 -12006
rect 19043 -12096 19075 -12062
rect 19109 -12096 19176 -12062
rect 19210 -12096 19245 -12062
rect 19043 -12152 19245 -12096
rect 19043 -12186 19075 -12152
rect 19109 -12186 19176 -12152
rect 19210 -12186 19245 -12152
rect 19043 -12242 19245 -12186
rect 19043 -12276 19075 -12242
rect 19109 -12276 19176 -12242
rect 19210 -12276 19245 -12242
rect 19043 -12332 19245 -12276
rect 19043 -12366 19075 -12332
rect 19109 -12366 19176 -12332
rect 19210 -12366 19245 -12332
rect 19043 -12422 19245 -12366
rect 17755 -12489 17957 -12456
rect 19043 -12456 19075 -12422
rect 19109 -12456 19176 -12422
rect 19210 -12456 19245 -12422
rect 20331 -11466 20363 -11432
rect 20397 -11466 20464 -11432
rect 20498 -11466 20533 -11432
rect 21619 -11432 21821 -11403
rect 20331 -11522 20533 -11466
rect 20331 -11556 20363 -11522
rect 20397 -11556 20464 -11522
rect 20498 -11556 20533 -11522
rect 20331 -11612 20533 -11556
rect 20331 -11646 20363 -11612
rect 20397 -11646 20464 -11612
rect 20498 -11646 20533 -11612
rect 20331 -11702 20533 -11646
rect 20331 -11736 20363 -11702
rect 20397 -11736 20464 -11702
rect 20498 -11736 20533 -11702
rect 20331 -11792 20533 -11736
rect 20331 -11826 20363 -11792
rect 20397 -11826 20464 -11792
rect 20498 -11826 20533 -11792
rect 20331 -11882 20533 -11826
rect 20331 -11916 20363 -11882
rect 20397 -11916 20464 -11882
rect 20498 -11916 20533 -11882
rect 20331 -11972 20533 -11916
rect 20331 -12006 20363 -11972
rect 20397 -12006 20464 -11972
rect 20498 -12006 20533 -11972
rect 20331 -12062 20533 -12006
rect 20331 -12096 20363 -12062
rect 20397 -12096 20464 -12062
rect 20498 -12096 20533 -12062
rect 20331 -12152 20533 -12096
rect 20331 -12186 20363 -12152
rect 20397 -12186 20464 -12152
rect 20498 -12186 20533 -12152
rect 20331 -12242 20533 -12186
rect 20331 -12276 20363 -12242
rect 20397 -12276 20464 -12242
rect 20498 -12276 20533 -12242
rect 20331 -12332 20533 -12276
rect 20331 -12366 20363 -12332
rect 20397 -12366 20464 -12332
rect 20498 -12366 20533 -12332
rect 20331 -12422 20533 -12366
rect 19043 -12489 19245 -12456
rect 20331 -12456 20363 -12422
rect 20397 -12456 20464 -12422
rect 20498 -12456 20533 -12422
rect 21619 -11466 21651 -11432
rect 21685 -11466 21752 -11432
rect 21786 -11466 21821 -11432
rect 22907 -11432 23109 -11403
rect 21619 -11522 21821 -11466
rect 21619 -11556 21651 -11522
rect 21685 -11556 21752 -11522
rect 21786 -11556 21821 -11522
rect 21619 -11612 21821 -11556
rect 21619 -11646 21651 -11612
rect 21685 -11646 21752 -11612
rect 21786 -11646 21821 -11612
rect 21619 -11702 21821 -11646
rect 21619 -11736 21651 -11702
rect 21685 -11736 21752 -11702
rect 21786 -11736 21821 -11702
rect 21619 -11792 21821 -11736
rect 21619 -11826 21651 -11792
rect 21685 -11826 21752 -11792
rect 21786 -11826 21821 -11792
rect 21619 -11882 21821 -11826
rect 21619 -11916 21651 -11882
rect 21685 -11916 21752 -11882
rect 21786 -11916 21821 -11882
rect 21619 -11972 21821 -11916
rect 21619 -12006 21651 -11972
rect 21685 -12006 21752 -11972
rect 21786 -12006 21821 -11972
rect 21619 -12062 21821 -12006
rect 21619 -12096 21651 -12062
rect 21685 -12096 21752 -12062
rect 21786 -12096 21821 -12062
rect 21619 -12152 21821 -12096
rect 21619 -12186 21651 -12152
rect 21685 -12186 21752 -12152
rect 21786 -12186 21821 -12152
rect 21619 -12242 21821 -12186
rect 21619 -12276 21651 -12242
rect 21685 -12276 21752 -12242
rect 21786 -12276 21821 -12242
rect 21619 -12332 21821 -12276
rect 21619 -12366 21651 -12332
rect 21685 -12366 21752 -12332
rect 21786 -12366 21821 -12332
rect 21619 -12422 21821 -12366
rect 20331 -12489 20533 -12456
rect 21619 -12456 21651 -12422
rect 21685 -12456 21752 -12422
rect 21786 -12456 21821 -12422
rect 22907 -11466 22939 -11432
rect 22973 -11466 23040 -11432
rect 23074 -11466 23109 -11432
rect 24195 -11432 24397 -11403
rect 22907 -11522 23109 -11466
rect 22907 -11556 22939 -11522
rect 22973 -11556 23040 -11522
rect 23074 -11556 23109 -11522
rect 22907 -11612 23109 -11556
rect 22907 -11646 22939 -11612
rect 22973 -11646 23040 -11612
rect 23074 -11646 23109 -11612
rect 22907 -11702 23109 -11646
rect 22907 -11736 22939 -11702
rect 22973 -11736 23040 -11702
rect 23074 -11736 23109 -11702
rect 22907 -11792 23109 -11736
rect 22907 -11826 22939 -11792
rect 22973 -11826 23040 -11792
rect 23074 -11826 23109 -11792
rect 22907 -11882 23109 -11826
rect 22907 -11916 22939 -11882
rect 22973 -11916 23040 -11882
rect 23074 -11916 23109 -11882
rect 22907 -11972 23109 -11916
rect 22907 -12006 22939 -11972
rect 22973 -12006 23040 -11972
rect 23074 -12006 23109 -11972
rect 22907 -12062 23109 -12006
rect 22907 -12096 22939 -12062
rect 22973 -12096 23040 -12062
rect 23074 -12096 23109 -12062
rect 22907 -12152 23109 -12096
rect 22907 -12186 22939 -12152
rect 22973 -12186 23040 -12152
rect 23074 -12186 23109 -12152
rect 22907 -12242 23109 -12186
rect 22907 -12276 22939 -12242
rect 22973 -12276 23040 -12242
rect 23074 -12276 23109 -12242
rect 22907 -12332 23109 -12276
rect 22907 -12366 22939 -12332
rect 22973 -12366 23040 -12332
rect 23074 -12366 23109 -12332
rect 22907 -12422 23109 -12366
rect 21619 -12489 21821 -12456
rect 22907 -12456 22939 -12422
rect 22973 -12456 23040 -12422
rect 23074 -12456 23109 -12422
rect 24195 -11466 24227 -11432
rect 24261 -11466 24328 -11432
rect 24362 -11466 24397 -11432
rect 25483 -11432 25685 -11403
rect 24195 -11522 24397 -11466
rect 24195 -11556 24227 -11522
rect 24261 -11556 24328 -11522
rect 24362 -11556 24397 -11522
rect 24195 -11612 24397 -11556
rect 24195 -11646 24227 -11612
rect 24261 -11646 24328 -11612
rect 24362 -11646 24397 -11612
rect 24195 -11702 24397 -11646
rect 24195 -11736 24227 -11702
rect 24261 -11736 24328 -11702
rect 24362 -11736 24397 -11702
rect 24195 -11792 24397 -11736
rect 24195 -11826 24227 -11792
rect 24261 -11826 24328 -11792
rect 24362 -11826 24397 -11792
rect 24195 -11882 24397 -11826
rect 24195 -11916 24227 -11882
rect 24261 -11916 24328 -11882
rect 24362 -11916 24397 -11882
rect 24195 -11972 24397 -11916
rect 24195 -12006 24227 -11972
rect 24261 -12006 24328 -11972
rect 24362 -12006 24397 -11972
rect 24195 -12062 24397 -12006
rect 24195 -12096 24227 -12062
rect 24261 -12096 24328 -12062
rect 24362 -12096 24397 -12062
rect 24195 -12152 24397 -12096
rect 24195 -12186 24227 -12152
rect 24261 -12186 24328 -12152
rect 24362 -12186 24397 -12152
rect 24195 -12242 24397 -12186
rect 24195 -12276 24227 -12242
rect 24261 -12276 24328 -12242
rect 24362 -12276 24397 -12242
rect 24195 -12332 24397 -12276
rect 24195 -12366 24227 -12332
rect 24261 -12366 24328 -12332
rect 24362 -12366 24397 -12332
rect 24195 -12422 24397 -12366
rect 22907 -12489 23109 -12456
rect 24195 -12456 24227 -12422
rect 24261 -12456 24328 -12422
rect 24362 -12456 24397 -12422
rect 25483 -11466 25515 -11432
rect 25549 -11466 25616 -11432
rect 25650 -11466 25685 -11432
rect 26771 -11432 26872 -11403
rect 25483 -11522 25685 -11466
rect 25483 -11556 25515 -11522
rect 25549 -11556 25616 -11522
rect 25650 -11556 25685 -11522
rect 25483 -11612 25685 -11556
rect 25483 -11646 25515 -11612
rect 25549 -11646 25616 -11612
rect 25650 -11646 25685 -11612
rect 25483 -11702 25685 -11646
rect 25483 -11736 25515 -11702
rect 25549 -11736 25616 -11702
rect 25650 -11736 25685 -11702
rect 25483 -11792 25685 -11736
rect 25483 -11826 25515 -11792
rect 25549 -11826 25616 -11792
rect 25650 -11826 25685 -11792
rect 25483 -11882 25685 -11826
rect 25483 -11916 25515 -11882
rect 25549 -11916 25616 -11882
rect 25650 -11916 25685 -11882
rect 25483 -11972 25685 -11916
rect 25483 -12006 25515 -11972
rect 25549 -12006 25616 -11972
rect 25650 -12006 25685 -11972
rect 25483 -12062 25685 -12006
rect 25483 -12096 25515 -12062
rect 25549 -12096 25616 -12062
rect 25650 -12096 25685 -12062
rect 25483 -12152 25685 -12096
rect 25483 -12186 25515 -12152
rect 25549 -12186 25616 -12152
rect 25650 -12186 25685 -12152
rect 25483 -12242 25685 -12186
rect 25483 -12276 25515 -12242
rect 25549 -12276 25616 -12242
rect 25650 -12276 25685 -12242
rect 25483 -12332 25685 -12276
rect 25483 -12366 25515 -12332
rect 25549 -12366 25616 -12332
rect 25650 -12366 25685 -12332
rect 25483 -12422 25685 -12366
rect 24195 -12489 24397 -12456
rect 25483 -12456 25515 -12422
rect 25549 -12456 25616 -12422
rect 25650 -12456 25685 -12422
rect 26771 -11466 26803 -11432
rect 26837 -11466 26872 -11432
rect 26771 -11522 26872 -11466
rect 26771 -11556 26803 -11522
rect 26837 -11556 26872 -11522
rect 26771 -11612 26872 -11556
rect 26771 -11646 26803 -11612
rect 26837 -11646 26872 -11612
rect 26771 -11702 26872 -11646
rect 26771 -11736 26803 -11702
rect 26837 -11736 26872 -11702
rect 26771 -11792 26872 -11736
rect 26771 -11826 26803 -11792
rect 26837 -11826 26872 -11792
rect 26771 -11882 26872 -11826
rect 26771 -11916 26803 -11882
rect 26837 -11916 26872 -11882
rect 26771 -11972 26872 -11916
rect 26771 -12006 26803 -11972
rect 26837 -12006 26872 -11972
rect 26771 -12062 26872 -12006
rect 26771 -12096 26803 -12062
rect 26837 -12096 26872 -12062
rect 26771 -12152 26872 -12096
rect 26771 -12186 26803 -12152
rect 26837 -12186 26872 -12152
rect 26771 -12242 26872 -12186
rect 26771 -12276 26803 -12242
rect 26837 -12276 26872 -12242
rect 26771 -12332 26872 -12276
rect 26771 -12366 26803 -12332
rect 26837 -12366 26872 -12332
rect 26771 -12422 26872 -12366
rect 25483 -12489 25685 -12456
rect 26771 -12456 26803 -12422
rect 26837 -12456 26872 -12422
rect 26771 -12489 26872 -12456
rect 16568 -12523 26872 -12489
rect 16568 -12557 16684 -12523
rect 16718 -12557 16774 -12523
rect 16808 -12557 16864 -12523
rect 16898 -12557 16954 -12523
rect 16988 -12557 17044 -12523
rect 17078 -12557 17134 -12523
rect 17168 -12557 17224 -12523
rect 17258 -12557 17314 -12523
rect 17348 -12557 17404 -12523
rect 17438 -12557 17494 -12523
rect 17528 -12557 17584 -12523
rect 17618 -12557 17674 -12523
rect 17708 -12557 17764 -12523
rect 17798 -12557 17972 -12523
rect 18006 -12557 18062 -12523
rect 18096 -12557 18152 -12523
rect 18186 -12557 18242 -12523
rect 18276 -12557 18332 -12523
rect 18366 -12557 18422 -12523
rect 18456 -12557 18512 -12523
rect 18546 -12557 18602 -12523
rect 18636 -12557 18692 -12523
rect 18726 -12557 18782 -12523
rect 18816 -12557 18872 -12523
rect 18906 -12557 18962 -12523
rect 18996 -12557 19052 -12523
rect 19086 -12557 19260 -12523
rect 19294 -12557 19350 -12523
rect 19384 -12557 19440 -12523
rect 19474 -12557 19530 -12523
rect 19564 -12557 19620 -12523
rect 19654 -12557 19710 -12523
rect 19744 -12557 19800 -12523
rect 19834 -12557 19890 -12523
rect 19924 -12557 19980 -12523
rect 20014 -12557 20070 -12523
rect 20104 -12557 20160 -12523
rect 20194 -12557 20250 -12523
rect 20284 -12557 20340 -12523
rect 20374 -12557 20548 -12523
rect 20582 -12557 20638 -12523
rect 20672 -12557 20728 -12523
rect 20762 -12557 20818 -12523
rect 20852 -12557 20908 -12523
rect 20942 -12557 20998 -12523
rect 21032 -12557 21088 -12523
rect 21122 -12557 21178 -12523
rect 21212 -12557 21268 -12523
rect 21302 -12557 21358 -12523
rect 21392 -12557 21448 -12523
rect 21482 -12557 21538 -12523
rect 21572 -12557 21628 -12523
rect 21662 -12557 21836 -12523
rect 21870 -12557 21926 -12523
rect 21960 -12557 22016 -12523
rect 22050 -12557 22106 -12523
rect 22140 -12557 22196 -12523
rect 22230 -12557 22286 -12523
rect 22320 -12557 22376 -12523
rect 22410 -12557 22466 -12523
rect 22500 -12557 22556 -12523
rect 22590 -12557 22646 -12523
rect 22680 -12557 22736 -12523
rect 22770 -12557 22826 -12523
rect 22860 -12557 22916 -12523
rect 22950 -12557 23124 -12523
rect 23158 -12557 23214 -12523
rect 23248 -12557 23304 -12523
rect 23338 -12557 23394 -12523
rect 23428 -12557 23484 -12523
rect 23518 -12557 23574 -12523
rect 23608 -12557 23664 -12523
rect 23698 -12557 23754 -12523
rect 23788 -12557 23844 -12523
rect 23878 -12557 23934 -12523
rect 23968 -12557 24024 -12523
rect 24058 -12557 24114 -12523
rect 24148 -12557 24204 -12523
rect 24238 -12557 24412 -12523
rect 24446 -12557 24502 -12523
rect 24536 -12557 24592 -12523
rect 24626 -12557 24682 -12523
rect 24716 -12557 24772 -12523
rect 24806 -12557 24862 -12523
rect 24896 -12557 24952 -12523
rect 24986 -12557 25042 -12523
rect 25076 -12557 25132 -12523
rect 25166 -12557 25222 -12523
rect 25256 -12557 25312 -12523
rect 25346 -12557 25402 -12523
rect 25436 -12557 25492 -12523
rect 25526 -12557 25700 -12523
rect 25734 -12557 25790 -12523
rect 25824 -12557 25880 -12523
rect 25914 -12557 25970 -12523
rect 26004 -12557 26060 -12523
rect 26094 -12557 26150 -12523
rect 26184 -12557 26240 -12523
rect 26274 -12557 26330 -12523
rect 26364 -12557 26420 -12523
rect 26454 -12557 26510 -12523
rect 26544 -12557 26600 -12523
rect 26634 -12557 26690 -12523
rect 26724 -12557 26780 -12523
rect 26814 -12557 26872 -12523
rect 16568 -12624 26872 -12557
rect 16568 -12658 16684 -12624
rect 16718 -12658 16774 -12624
rect 16808 -12658 16864 -12624
rect 16898 -12658 16954 -12624
rect 16988 -12658 17044 -12624
rect 17078 -12658 17134 -12624
rect 17168 -12658 17224 -12624
rect 17258 -12658 17314 -12624
rect 17348 -12658 17404 -12624
rect 17438 -12658 17494 -12624
rect 17528 -12658 17584 -12624
rect 17618 -12658 17674 -12624
rect 17708 -12658 17764 -12624
rect 17798 -12658 17972 -12624
rect 18006 -12658 18062 -12624
rect 18096 -12658 18152 -12624
rect 18186 -12658 18242 -12624
rect 18276 -12658 18332 -12624
rect 18366 -12658 18422 -12624
rect 18456 -12658 18512 -12624
rect 18546 -12658 18602 -12624
rect 18636 -12658 18692 -12624
rect 18726 -12658 18782 -12624
rect 18816 -12658 18872 -12624
rect 18906 -12658 18962 -12624
rect 18996 -12658 19052 -12624
rect 19086 -12658 19260 -12624
rect 19294 -12658 19350 -12624
rect 19384 -12658 19440 -12624
rect 19474 -12658 19530 -12624
rect 19564 -12658 19620 -12624
rect 19654 -12658 19710 -12624
rect 19744 -12658 19800 -12624
rect 19834 -12658 19890 -12624
rect 19924 -12658 19980 -12624
rect 20014 -12658 20070 -12624
rect 20104 -12658 20160 -12624
rect 20194 -12658 20250 -12624
rect 20284 -12658 20340 -12624
rect 20374 -12658 20548 -12624
rect 20582 -12658 20638 -12624
rect 20672 -12658 20728 -12624
rect 20762 -12658 20818 -12624
rect 20852 -12658 20908 -12624
rect 20942 -12658 20998 -12624
rect 21032 -12658 21088 -12624
rect 21122 -12658 21178 -12624
rect 21212 -12658 21268 -12624
rect 21302 -12658 21358 -12624
rect 21392 -12658 21448 -12624
rect 21482 -12658 21538 -12624
rect 21572 -12658 21628 -12624
rect 21662 -12658 21836 -12624
rect 21870 -12658 21926 -12624
rect 21960 -12658 22016 -12624
rect 22050 -12658 22106 -12624
rect 22140 -12658 22196 -12624
rect 22230 -12658 22286 -12624
rect 22320 -12658 22376 -12624
rect 22410 -12658 22466 -12624
rect 22500 -12658 22556 -12624
rect 22590 -12658 22646 -12624
rect 22680 -12658 22736 -12624
rect 22770 -12658 22826 -12624
rect 22860 -12658 22916 -12624
rect 22950 -12658 23124 -12624
rect 23158 -12658 23214 -12624
rect 23248 -12658 23304 -12624
rect 23338 -12658 23394 -12624
rect 23428 -12658 23484 -12624
rect 23518 -12658 23574 -12624
rect 23608 -12658 23664 -12624
rect 23698 -12658 23754 -12624
rect 23788 -12658 23844 -12624
rect 23878 -12658 23934 -12624
rect 23968 -12658 24024 -12624
rect 24058 -12658 24114 -12624
rect 24148 -12658 24204 -12624
rect 24238 -12658 24412 -12624
rect 24446 -12658 24502 -12624
rect 24536 -12658 24592 -12624
rect 24626 -12658 24682 -12624
rect 24716 -12658 24772 -12624
rect 24806 -12658 24862 -12624
rect 24896 -12658 24952 -12624
rect 24986 -12658 25042 -12624
rect 25076 -12658 25132 -12624
rect 25166 -12658 25222 -12624
rect 25256 -12658 25312 -12624
rect 25346 -12658 25402 -12624
rect 25436 -12658 25492 -12624
rect 25526 -12658 25700 -12624
rect 25734 -12658 25790 -12624
rect 25824 -12658 25880 -12624
rect 25914 -12658 25970 -12624
rect 26004 -12658 26060 -12624
rect 26094 -12658 26150 -12624
rect 26184 -12658 26240 -12624
rect 26274 -12658 26330 -12624
rect 26364 -12658 26420 -12624
rect 26454 -12658 26510 -12624
rect 26544 -12658 26600 -12624
rect 26634 -12658 26690 -12624
rect 26724 -12658 26780 -12624
rect 26814 -12658 26872 -12624
rect 16568 -12691 26872 -12658
rect 16568 -12720 16669 -12691
rect 16568 -12754 16600 -12720
rect 16634 -12754 16669 -12720
rect 17755 -12720 17957 -12691
rect 16568 -12810 16669 -12754
rect 16568 -12844 16600 -12810
rect 16634 -12844 16669 -12810
rect 16568 -12900 16669 -12844
rect 16568 -12934 16600 -12900
rect 16634 -12934 16669 -12900
rect 16568 -12990 16669 -12934
rect 16568 -13024 16600 -12990
rect 16634 -13024 16669 -12990
rect 16568 -13080 16669 -13024
rect 16568 -13114 16600 -13080
rect 16634 -13114 16669 -13080
rect 16568 -13170 16669 -13114
rect 16568 -13204 16600 -13170
rect 16634 -13204 16669 -13170
rect 16568 -13260 16669 -13204
rect 16568 -13294 16600 -13260
rect 16634 -13294 16669 -13260
rect 16568 -13350 16669 -13294
rect 16568 -13384 16600 -13350
rect 16634 -13384 16669 -13350
rect 16568 -13440 16669 -13384
rect 16568 -13474 16600 -13440
rect 16634 -13474 16669 -13440
rect 16568 -13530 16669 -13474
rect 16568 -13564 16600 -13530
rect 16634 -13564 16669 -13530
rect 16568 -13620 16669 -13564
rect 16568 -13654 16600 -13620
rect 16634 -13654 16669 -13620
rect 16568 -13710 16669 -13654
rect 16568 -13744 16600 -13710
rect 16634 -13744 16669 -13710
rect 17755 -12754 17787 -12720
rect 17821 -12754 17888 -12720
rect 17922 -12754 17957 -12720
rect 19043 -12720 19245 -12691
rect 17755 -12810 17957 -12754
rect 17755 -12844 17787 -12810
rect 17821 -12844 17888 -12810
rect 17922 -12844 17957 -12810
rect 17755 -12900 17957 -12844
rect 17755 -12934 17787 -12900
rect 17821 -12934 17888 -12900
rect 17922 -12934 17957 -12900
rect 17755 -12990 17957 -12934
rect 17755 -13024 17787 -12990
rect 17821 -13024 17888 -12990
rect 17922 -13024 17957 -12990
rect 17755 -13080 17957 -13024
rect 17755 -13114 17787 -13080
rect 17821 -13114 17888 -13080
rect 17922 -13114 17957 -13080
rect 17755 -13170 17957 -13114
rect 17755 -13204 17787 -13170
rect 17821 -13204 17888 -13170
rect 17922 -13204 17957 -13170
rect 17755 -13260 17957 -13204
rect 17755 -13294 17787 -13260
rect 17821 -13294 17888 -13260
rect 17922 -13294 17957 -13260
rect 17755 -13350 17957 -13294
rect 17755 -13384 17787 -13350
rect 17821 -13384 17888 -13350
rect 17922 -13384 17957 -13350
rect 17755 -13440 17957 -13384
rect 17755 -13474 17787 -13440
rect 17821 -13474 17888 -13440
rect 17922 -13474 17957 -13440
rect 17755 -13530 17957 -13474
rect 17755 -13564 17787 -13530
rect 17821 -13564 17888 -13530
rect 17922 -13564 17957 -13530
rect 17755 -13620 17957 -13564
rect 17755 -13654 17787 -13620
rect 17821 -13654 17888 -13620
rect 17922 -13654 17957 -13620
rect 17755 -13710 17957 -13654
rect 16568 -13777 16669 -13744
rect 17755 -13744 17787 -13710
rect 17821 -13744 17888 -13710
rect 17922 -13744 17957 -13710
rect 19043 -12754 19075 -12720
rect 19109 -12754 19176 -12720
rect 19210 -12754 19245 -12720
rect 20331 -12720 20533 -12691
rect 19043 -12810 19245 -12754
rect 19043 -12844 19075 -12810
rect 19109 -12844 19176 -12810
rect 19210 -12844 19245 -12810
rect 19043 -12900 19245 -12844
rect 19043 -12934 19075 -12900
rect 19109 -12934 19176 -12900
rect 19210 -12934 19245 -12900
rect 19043 -12990 19245 -12934
rect 19043 -13024 19075 -12990
rect 19109 -13024 19176 -12990
rect 19210 -13024 19245 -12990
rect 19043 -13080 19245 -13024
rect 19043 -13114 19075 -13080
rect 19109 -13114 19176 -13080
rect 19210 -13114 19245 -13080
rect 19043 -13170 19245 -13114
rect 19043 -13204 19075 -13170
rect 19109 -13204 19176 -13170
rect 19210 -13204 19245 -13170
rect 19043 -13260 19245 -13204
rect 19043 -13294 19075 -13260
rect 19109 -13294 19176 -13260
rect 19210 -13294 19245 -13260
rect 19043 -13350 19245 -13294
rect 19043 -13384 19075 -13350
rect 19109 -13384 19176 -13350
rect 19210 -13384 19245 -13350
rect 19043 -13440 19245 -13384
rect 19043 -13474 19075 -13440
rect 19109 -13474 19176 -13440
rect 19210 -13474 19245 -13440
rect 19043 -13530 19245 -13474
rect 19043 -13564 19075 -13530
rect 19109 -13564 19176 -13530
rect 19210 -13564 19245 -13530
rect 19043 -13620 19245 -13564
rect 19043 -13654 19075 -13620
rect 19109 -13654 19176 -13620
rect 19210 -13654 19245 -13620
rect 19043 -13710 19245 -13654
rect 17755 -13777 17957 -13744
rect 19043 -13744 19075 -13710
rect 19109 -13744 19176 -13710
rect 19210 -13744 19245 -13710
rect 20331 -12754 20363 -12720
rect 20397 -12754 20464 -12720
rect 20498 -12754 20533 -12720
rect 21619 -12720 21821 -12691
rect 20331 -12810 20533 -12754
rect 20331 -12844 20363 -12810
rect 20397 -12844 20464 -12810
rect 20498 -12844 20533 -12810
rect 20331 -12900 20533 -12844
rect 20331 -12934 20363 -12900
rect 20397 -12934 20464 -12900
rect 20498 -12934 20533 -12900
rect 20331 -12990 20533 -12934
rect 20331 -13024 20363 -12990
rect 20397 -13024 20464 -12990
rect 20498 -13024 20533 -12990
rect 20331 -13080 20533 -13024
rect 20331 -13114 20363 -13080
rect 20397 -13114 20464 -13080
rect 20498 -13114 20533 -13080
rect 20331 -13170 20533 -13114
rect 20331 -13204 20363 -13170
rect 20397 -13204 20464 -13170
rect 20498 -13204 20533 -13170
rect 20331 -13260 20533 -13204
rect 20331 -13294 20363 -13260
rect 20397 -13294 20464 -13260
rect 20498 -13294 20533 -13260
rect 20331 -13350 20533 -13294
rect 20331 -13384 20363 -13350
rect 20397 -13384 20464 -13350
rect 20498 -13384 20533 -13350
rect 20331 -13440 20533 -13384
rect 20331 -13474 20363 -13440
rect 20397 -13474 20464 -13440
rect 20498 -13474 20533 -13440
rect 20331 -13530 20533 -13474
rect 20331 -13564 20363 -13530
rect 20397 -13564 20464 -13530
rect 20498 -13564 20533 -13530
rect 20331 -13620 20533 -13564
rect 20331 -13654 20363 -13620
rect 20397 -13654 20464 -13620
rect 20498 -13654 20533 -13620
rect 20331 -13710 20533 -13654
rect 19043 -13777 19245 -13744
rect 20331 -13744 20363 -13710
rect 20397 -13744 20464 -13710
rect 20498 -13744 20533 -13710
rect 21619 -12754 21651 -12720
rect 21685 -12754 21752 -12720
rect 21786 -12754 21821 -12720
rect 22907 -12720 23109 -12691
rect 21619 -12810 21821 -12754
rect 21619 -12844 21651 -12810
rect 21685 -12844 21752 -12810
rect 21786 -12844 21821 -12810
rect 21619 -12900 21821 -12844
rect 21619 -12934 21651 -12900
rect 21685 -12934 21752 -12900
rect 21786 -12934 21821 -12900
rect 21619 -12990 21821 -12934
rect 21619 -13024 21651 -12990
rect 21685 -13024 21752 -12990
rect 21786 -13024 21821 -12990
rect 21619 -13080 21821 -13024
rect 21619 -13114 21651 -13080
rect 21685 -13114 21752 -13080
rect 21786 -13114 21821 -13080
rect 21619 -13170 21821 -13114
rect 21619 -13204 21651 -13170
rect 21685 -13204 21752 -13170
rect 21786 -13204 21821 -13170
rect 21619 -13260 21821 -13204
rect 21619 -13294 21651 -13260
rect 21685 -13294 21752 -13260
rect 21786 -13294 21821 -13260
rect 21619 -13350 21821 -13294
rect 21619 -13384 21651 -13350
rect 21685 -13384 21752 -13350
rect 21786 -13384 21821 -13350
rect 21619 -13440 21821 -13384
rect 21619 -13474 21651 -13440
rect 21685 -13474 21752 -13440
rect 21786 -13474 21821 -13440
rect 21619 -13530 21821 -13474
rect 21619 -13564 21651 -13530
rect 21685 -13564 21752 -13530
rect 21786 -13564 21821 -13530
rect 21619 -13620 21821 -13564
rect 21619 -13654 21651 -13620
rect 21685 -13654 21752 -13620
rect 21786 -13654 21821 -13620
rect 21619 -13710 21821 -13654
rect 20331 -13777 20533 -13744
rect 21619 -13744 21651 -13710
rect 21685 -13744 21752 -13710
rect 21786 -13744 21821 -13710
rect 22907 -12754 22939 -12720
rect 22973 -12754 23040 -12720
rect 23074 -12754 23109 -12720
rect 24195 -12720 24397 -12691
rect 22907 -12810 23109 -12754
rect 22907 -12844 22939 -12810
rect 22973 -12844 23040 -12810
rect 23074 -12844 23109 -12810
rect 22907 -12900 23109 -12844
rect 22907 -12934 22939 -12900
rect 22973 -12934 23040 -12900
rect 23074 -12934 23109 -12900
rect 22907 -12990 23109 -12934
rect 22907 -13024 22939 -12990
rect 22973 -13024 23040 -12990
rect 23074 -13024 23109 -12990
rect 22907 -13080 23109 -13024
rect 22907 -13114 22939 -13080
rect 22973 -13114 23040 -13080
rect 23074 -13114 23109 -13080
rect 22907 -13170 23109 -13114
rect 22907 -13204 22939 -13170
rect 22973 -13204 23040 -13170
rect 23074 -13204 23109 -13170
rect 22907 -13260 23109 -13204
rect 22907 -13294 22939 -13260
rect 22973 -13294 23040 -13260
rect 23074 -13294 23109 -13260
rect 22907 -13350 23109 -13294
rect 22907 -13384 22939 -13350
rect 22973 -13384 23040 -13350
rect 23074 -13384 23109 -13350
rect 22907 -13440 23109 -13384
rect 22907 -13474 22939 -13440
rect 22973 -13474 23040 -13440
rect 23074 -13474 23109 -13440
rect 22907 -13530 23109 -13474
rect 22907 -13564 22939 -13530
rect 22973 -13564 23040 -13530
rect 23074 -13564 23109 -13530
rect 22907 -13620 23109 -13564
rect 22907 -13654 22939 -13620
rect 22973 -13654 23040 -13620
rect 23074 -13654 23109 -13620
rect 22907 -13710 23109 -13654
rect 21619 -13777 21821 -13744
rect 22907 -13744 22939 -13710
rect 22973 -13744 23040 -13710
rect 23074 -13744 23109 -13710
rect 24195 -12754 24227 -12720
rect 24261 -12754 24328 -12720
rect 24362 -12754 24397 -12720
rect 25483 -12720 25685 -12691
rect 24195 -12810 24397 -12754
rect 24195 -12844 24227 -12810
rect 24261 -12844 24328 -12810
rect 24362 -12844 24397 -12810
rect 24195 -12900 24397 -12844
rect 24195 -12934 24227 -12900
rect 24261 -12934 24328 -12900
rect 24362 -12934 24397 -12900
rect 24195 -12990 24397 -12934
rect 24195 -13024 24227 -12990
rect 24261 -13024 24328 -12990
rect 24362 -13024 24397 -12990
rect 24195 -13080 24397 -13024
rect 24195 -13114 24227 -13080
rect 24261 -13114 24328 -13080
rect 24362 -13114 24397 -13080
rect 24195 -13170 24397 -13114
rect 24195 -13204 24227 -13170
rect 24261 -13204 24328 -13170
rect 24362 -13204 24397 -13170
rect 24195 -13260 24397 -13204
rect 24195 -13294 24227 -13260
rect 24261 -13294 24328 -13260
rect 24362 -13294 24397 -13260
rect 24195 -13350 24397 -13294
rect 24195 -13384 24227 -13350
rect 24261 -13384 24328 -13350
rect 24362 -13384 24397 -13350
rect 24195 -13440 24397 -13384
rect 24195 -13474 24227 -13440
rect 24261 -13474 24328 -13440
rect 24362 -13474 24397 -13440
rect 24195 -13530 24397 -13474
rect 24195 -13564 24227 -13530
rect 24261 -13564 24328 -13530
rect 24362 -13564 24397 -13530
rect 24195 -13620 24397 -13564
rect 24195 -13654 24227 -13620
rect 24261 -13654 24328 -13620
rect 24362 -13654 24397 -13620
rect 24195 -13710 24397 -13654
rect 22907 -13777 23109 -13744
rect 24195 -13744 24227 -13710
rect 24261 -13744 24328 -13710
rect 24362 -13744 24397 -13710
rect 25483 -12754 25515 -12720
rect 25549 -12754 25616 -12720
rect 25650 -12754 25685 -12720
rect 26771 -12720 26872 -12691
rect 25483 -12810 25685 -12754
rect 25483 -12844 25515 -12810
rect 25549 -12844 25616 -12810
rect 25650 -12844 25685 -12810
rect 25483 -12900 25685 -12844
rect 25483 -12934 25515 -12900
rect 25549 -12934 25616 -12900
rect 25650 -12934 25685 -12900
rect 25483 -12990 25685 -12934
rect 25483 -13024 25515 -12990
rect 25549 -13024 25616 -12990
rect 25650 -13024 25685 -12990
rect 25483 -13080 25685 -13024
rect 25483 -13114 25515 -13080
rect 25549 -13114 25616 -13080
rect 25650 -13114 25685 -13080
rect 25483 -13170 25685 -13114
rect 25483 -13204 25515 -13170
rect 25549 -13204 25616 -13170
rect 25650 -13204 25685 -13170
rect 25483 -13260 25685 -13204
rect 25483 -13294 25515 -13260
rect 25549 -13294 25616 -13260
rect 25650 -13294 25685 -13260
rect 25483 -13350 25685 -13294
rect 25483 -13384 25515 -13350
rect 25549 -13384 25616 -13350
rect 25650 -13384 25685 -13350
rect 25483 -13440 25685 -13384
rect 25483 -13474 25515 -13440
rect 25549 -13474 25616 -13440
rect 25650 -13474 25685 -13440
rect 25483 -13530 25685 -13474
rect 25483 -13564 25515 -13530
rect 25549 -13564 25616 -13530
rect 25650 -13564 25685 -13530
rect 25483 -13620 25685 -13564
rect 25483 -13654 25515 -13620
rect 25549 -13654 25616 -13620
rect 25650 -13654 25685 -13620
rect 25483 -13710 25685 -13654
rect 24195 -13777 24397 -13744
rect 25483 -13744 25515 -13710
rect 25549 -13744 25616 -13710
rect 25650 -13744 25685 -13710
rect 26771 -12754 26803 -12720
rect 26837 -12754 26872 -12720
rect 26771 -12810 26872 -12754
rect 26771 -12844 26803 -12810
rect 26837 -12844 26872 -12810
rect 26771 -12900 26872 -12844
rect 26771 -12934 26803 -12900
rect 26837 -12934 26872 -12900
rect 26771 -12990 26872 -12934
rect 26771 -13024 26803 -12990
rect 26837 -13024 26872 -12990
rect 26771 -13080 26872 -13024
rect 26771 -13114 26803 -13080
rect 26837 -13114 26872 -13080
rect 26771 -13170 26872 -13114
rect 26771 -13204 26803 -13170
rect 26837 -13204 26872 -13170
rect 26771 -13260 26872 -13204
rect 26771 -13294 26803 -13260
rect 26837 -13294 26872 -13260
rect 26771 -13350 26872 -13294
rect 26771 -13384 26803 -13350
rect 26837 -13384 26872 -13350
rect 26771 -13440 26872 -13384
rect 26771 -13474 26803 -13440
rect 26837 -13474 26872 -13440
rect 26771 -13530 26872 -13474
rect 26771 -13564 26803 -13530
rect 26837 -13564 26872 -13530
rect 26771 -13620 26872 -13564
rect 26771 -13654 26803 -13620
rect 26837 -13654 26872 -13620
rect 26771 -13710 26872 -13654
rect 25483 -13777 25685 -13744
rect 26771 -13744 26803 -13710
rect 26837 -13744 26872 -13710
rect 26771 -13777 26872 -13744
rect 16568 -13811 26872 -13777
rect 16568 -13845 16684 -13811
rect 16718 -13845 16774 -13811
rect 16808 -13845 16864 -13811
rect 16898 -13845 16954 -13811
rect 16988 -13845 17044 -13811
rect 17078 -13845 17134 -13811
rect 17168 -13845 17224 -13811
rect 17258 -13845 17314 -13811
rect 17348 -13845 17404 -13811
rect 17438 -13845 17494 -13811
rect 17528 -13845 17584 -13811
rect 17618 -13845 17674 -13811
rect 17708 -13845 17764 -13811
rect 17798 -13845 17972 -13811
rect 18006 -13845 18062 -13811
rect 18096 -13845 18152 -13811
rect 18186 -13845 18242 -13811
rect 18276 -13845 18332 -13811
rect 18366 -13845 18422 -13811
rect 18456 -13845 18512 -13811
rect 18546 -13845 18602 -13811
rect 18636 -13845 18692 -13811
rect 18726 -13845 18782 -13811
rect 18816 -13845 18872 -13811
rect 18906 -13845 18962 -13811
rect 18996 -13845 19052 -13811
rect 19086 -13845 19260 -13811
rect 19294 -13845 19350 -13811
rect 19384 -13845 19440 -13811
rect 19474 -13845 19530 -13811
rect 19564 -13845 19620 -13811
rect 19654 -13845 19710 -13811
rect 19744 -13845 19800 -13811
rect 19834 -13845 19890 -13811
rect 19924 -13845 19980 -13811
rect 20014 -13845 20070 -13811
rect 20104 -13845 20160 -13811
rect 20194 -13845 20250 -13811
rect 20284 -13845 20340 -13811
rect 20374 -13845 20548 -13811
rect 20582 -13845 20638 -13811
rect 20672 -13845 20728 -13811
rect 20762 -13845 20818 -13811
rect 20852 -13845 20908 -13811
rect 20942 -13845 20998 -13811
rect 21032 -13845 21088 -13811
rect 21122 -13845 21178 -13811
rect 21212 -13845 21268 -13811
rect 21302 -13845 21358 -13811
rect 21392 -13845 21448 -13811
rect 21482 -13845 21538 -13811
rect 21572 -13845 21628 -13811
rect 21662 -13845 21836 -13811
rect 21870 -13845 21926 -13811
rect 21960 -13845 22016 -13811
rect 22050 -13845 22106 -13811
rect 22140 -13845 22196 -13811
rect 22230 -13845 22286 -13811
rect 22320 -13845 22376 -13811
rect 22410 -13845 22466 -13811
rect 22500 -13845 22556 -13811
rect 22590 -13845 22646 -13811
rect 22680 -13845 22736 -13811
rect 22770 -13845 22826 -13811
rect 22860 -13845 22916 -13811
rect 22950 -13845 23124 -13811
rect 23158 -13845 23214 -13811
rect 23248 -13845 23304 -13811
rect 23338 -13845 23394 -13811
rect 23428 -13845 23484 -13811
rect 23518 -13845 23574 -13811
rect 23608 -13845 23664 -13811
rect 23698 -13845 23754 -13811
rect 23788 -13845 23844 -13811
rect 23878 -13845 23934 -13811
rect 23968 -13845 24024 -13811
rect 24058 -13845 24114 -13811
rect 24148 -13845 24204 -13811
rect 24238 -13845 24412 -13811
rect 24446 -13845 24502 -13811
rect 24536 -13845 24592 -13811
rect 24626 -13845 24682 -13811
rect 24716 -13845 24772 -13811
rect 24806 -13845 24862 -13811
rect 24896 -13845 24952 -13811
rect 24986 -13845 25042 -13811
rect 25076 -13845 25132 -13811
rect 25166 -13845 25222 -13811
rect 25256 -13845 25312 -13811
rect 25346 -13845 25402 -13811
rect 25436 -13845 25492 -13811
rect 25526 -13845 25700 -13811
rect 25734 -13845 25790 -13811
rect 25824 -13845 25880 -13811
rect 25914 -13845 25970 -13811
rect 26004 -13845 26060 -13811
rect 26094 -13845 26150 -13811
rect 26184 -13845 26240 -13811
rect 26274 -13845 26330 -13811
rect 26364 -13845 26420 -13811
rect 26454 -13845 26510 -13811
rect 26544 -13845 26600 -13811
rect 26634 -13845 26690 -13811
rect 26724 -13845 26780 -13811
rect 26814 -13845 26872 -13811
rect 16568 -13912 26872 -13845
rect 16568 -13946 16684 -13912
rect 16718 -13946 16774 -13912
rect 16808 -13946 16864 -13912
rect 16898 -13946 16954 -13912
rect 16988 -13946 17044 -13912
rect 17078 -13946 17134 -13912
rect 17168 -13946 17224 -13912
rect 17258 -13946 17314 -13912
rect 17348 -13946 17404 -13912
rect 17438 -13946 17494 -13912
rect 17528 -13946 17584 -13912
rect 17618 -13946 17674 -13912
rect 17708 -13946 17764 -13912
rect 17798 -13946 17972 -13912
rect 18006 -13946 18062 -13912
rect 18096 -13946 18152 -13912
rect 18186 -13946 18242 -13912
rect 18276 -13946 18332 -13912
rect 18366 -13946 18422 -13912
rect 18456 -13946 18512 -13912
rect 18546 -13946 18602 -13912
rect 18636 -13946 18692 -13912
rect 18726 -13946 18782 -13912
rect 18816 -13946 18872 -13912
rect 18906 -13946 18962 -13912
rect 18996 -13946 19052 -13912
rect 19086 -13946 19260 -13912
rect 19294 -13946 19350 -13912
rect 19384 -13946 19440 -13912
rect 19474 -13946 19530 -13912
rect 19564 -13946 19620 -13912
rect 19654 -13946 19710 -13912
rect 19744 -13946 19800 -13912
rect 19834 -13946 19890 -13912
rect 19924 -13946 19980 -13912
rect 20014 -13946 20070 -13912
rect 20104 -13946 20160 -13912
rect 20194 -13946 20250 -13912
rect 20284 -13946 20340 -13912
rect 20374 -13946 20548 -13912
rect 20582 -13946 20638 -13912
rect 20672 -13946 20728 -13912
rect 20762 -13946 20818 -13912
rect 20852 -13946 20908 -13912
rect 20942 -13946 20998 -13912
rect 21032 -13946 21088 -13912
rect 21122 -13946 21178 -13912
rect 21212 -13946 21268 -13912
rect 21302 -13946 21358 -13912
rect 21392 -13946 21448 -13912
rect 21482 -13946 21538 -13912
rect 21572 -13946 21628 -13912
rect 21662 -13946 21836 -13912
rect 21870 -13946 21926 -13912
rect 21960 -13946 22016 -13912
rect 22050 -13946 22106 -13912
rect 22140 -13946 22196 -13912
rect 22230 -13946 22286 -13912
rect 22320 -13946 22376 -13912
rect 22410 -13946 22466 -13912
rect 22500 -13946 22556 -13912
rect 22590 -13946 22646 -13912
rect 22680 -13946 22736 -13912
rect 22770 -13946 22826 -13912
rect 22860 -13946 22916 -13912
rect 22950 -13946 23124 -13912
rect 23158 -13946 23214 -13912
rect 23248 -13946 23304 -13912
rect 23338 -13946 23394 -13912
rect 23428 -13946 23484 -13912
rect 23518 -13946 23574 -13912
rect 23608 -13946 23664 -13912
rect 23698 -13946 23754 -13912
rect 23788 -13946 23844 -13912
rect 23878 -13946 23934 -13912
rect 23968 -13946 24024 -13912
rect 24058 -13946 24114 -13912
rect 24148 -13946 24204 -13912
rect 24238 -13946 24412 -13912
rect 24446 -13946 24502 -13912
rect 24536 -13946 24592 -13912
rect 24626 -13946 24682 -13912
rect 24716 -13946 24772 -13912
rect 24806 -13946 24862 -13912
rect 24896 -13946 24952 -13912
rect 24986 -13946 25042 -13912
rect 25076 -13946 25132 -13912
rect 25166 -13946 25222 -13912
rect 25256 -13946 25312 -13912
rect 25346 -13946 25402 -13912
rect 25436 -13946 25492 -13912
rect 25526 -13946 25700 -13912
rect 25734 -13946 25790 -13912
rect 25824 -13946 25880 -13912
rect 25914 -13946 25970 -13912
rect 26004 -13946 26060 -13912
rect 26094 -13946 26150 -13912
rect 26184 -13946 26240 -13912
rect 26274 -13946 26330 -13912
rect 26364 -13946 26420 -13912
rect 26454 -13946 26510 -13912
rect 26544 -13946 26600 -13912
rect 26634 -13946 26690 -13912
rect 26724 -13946 26780 -13912
rect 26814 -13946 26872 -13912
rect 16568 -13979 26872 -13946
rect 16568 -14008 16669 -13979
rect 16568 -14042 16600 -14008
rect 16634 -14042 16669 -14008
rect 17755 -14008 17957 -13979
rect 16568 -14098 16669 -14042
rect 16568 -14132 16600 -14098
rect 16634 -14132 16669 -14098
rect 16568 -14188 16669 -14132
rect 16568 -14222 16600 -14188
rect 16634 -14222 16669 -14188
rect 16568 -14278 16669 -14222
rect 16568 -14312 16600 -14278
rect 16634 -14312 16669 -14278
rect 16568 -14368 16669 -14312
rect 16568 -14402 16600 -14368
rect 16634 -14402 16669 -14368
rect 16568 -14458 16669 -14402
rect 16568 -14492 16600 -14458
rect 16634 -14492 16669 -14458
rect 16568 -14548 16669 -14492
rect 16568 -14582 16600 -14548
rect 16634 -14582 16669 -14548
rect 16568 -14638 16669 -14582
rect 16568 -14672 16600 -14638
rect 16634 -14672 16669 -14638
rect 16568 -14728 16669 -14672
rect 16568 -14762 16600 -14728
rect 16634 -14762 16669 -14728
rect 16568 -14818 16669 -14762
rect 16568 -14852 16600 -14818
rect 16634 -14852 16669 -14818
rect 16568 -14908 16669 -14852
rect 16568 -14942 16600 -14908
rect 16634 -14942 16669 -14908
rect 16568 -14998 16669 -14942
rect 16568 -15032 16600 -14998
rect 16634 -15032 16669 -14998
rect 17755 -14042 17787 -14008
rect 17821 -14042 17888 -14008
rect 17922 -14042 17957 -14008
rect 19043 -14008 19245 -13979
rect 17755 -14098 17957 -14042
rect 17755 -14132 17787 -14098
rect 17821 -14132 17888 -14098
rect 17922 -14132 17957 -14098
rect 17755 -14188 17957 -14132
rect 17755 -14222 17787 -14188
rect 17821 -14222 17888 -14188
rect 17922 -14222 17957 -14188
rect 17755 -14278 17957 -14222
rect 17755 -14312 17787 -14278
rect 17821 -14312 17888 -14278
rect 17922 -14312 17957 -14278
rect 17755 -14368 17957 -14312
rect 17755 -14402 17787 -14368
rect 17821 -14402 17888 -14368
rect 17922 -14402 17957 -14368
rect 17755 -14458 17957 -14402
rect 17755 -14492 17787 -14458
rect 17821 -14492 17888 -14458
rect 17922 -14492 17957 -14458
rect 17755 -14548 17957 -14492
rect 17755 -14582 17787 -14548
rect 17821 -14582 17888 -14548
rect 17922 -14582 17957 -14548
rect 17755 -14638 17957 -14582
rect 17755 -14672 17787 -14638
rect 17821 -14672 17888 -14638
rect 17922 -14672 17957 -14638
rect 17755 -14728 17957 -14672
rect 17755 -14762 17787 -14728
rect 17821 -14762 17888 -14728
rect 17922 -14762 17957 -14728
rect 17755 -14818 17957 -14762
rect 17755 -14852 17787 -14818
rect 17821 -14852 17888 -14818
rect 17922 -14852 17957 -14818
rect 17755 -14908 17957 -14852
rect 17755 -14942 17787 -14908
rect 17821 -14942 17888 -14908
rect 17922 -14942 17957 -14908
rect 17755 -14998 17957 -14942
rect 16568 -15065 16669 -15032
rect 17755 -15032 17787 -14998
rect 17821 -15032 17888 -14998
rect 17922 -15032 17957 -14998
rect 19043 -14042 19075 -14008
rect 19109 -14042 19176 -14008
rect 19210 -14042 19245 -14008
rect 20331 -14008 20533 -13979
rect 19043 -14098 19245 -14042
rect 19043 -14132 19075 -14098
rect 19109 -14132 19176 -14098
rect 19210 -14132 19245 -14098
rect 19043 -14188 19245 -14132
rect 19043 -14222 19075 -14188
rect 19109 -14222 19176 -14188
rect 19210 -14222 19245 -14188
rect 19043 -14278 19245 -14222
rect 19043 -14312 19075 -14278
rect 19109 -14312 19176 -14278
rect 19210 -14312 19245 -14278
rect 19043 -14368 19245 -14312
rect 19043 -14402 19075 -14368
rect 19109 -14402 19176 -14368
rect 19210 -14402 19245 -14368
rect 19043 -14458 19245 -14402
rect 19043 -14492 19075 -14458
rect 19109 -14492 19176 -14458
rect 19210 -14492 19245 -14458
rect 19043 -14548 19245 -14492
rect 19043 -14582 19075 -14548
rect 19109 -14582 19176 -14548
rect 19210 -14582 19245 -14548
rect 19043 -14638 19245 -14582
rect 19043 -14672 19075 -14638
rect 19109 -14672 19176 -14638
rect 19210 -14672 19245 -14638
rect 19043 -14728 19245 -14672
rect 19043 -14762 19075 -14728
rect 19109 -14762 19176 -14728
rect 19210 -14762 19245 -14728
rect 19043 -14818 19245 -14762
rect 19043 -14852 19075 -14818
rect 19109 -14852 19176 -14818
rect 19210 -14852 19245 -14818
rect 19043 -14908 19245 -14852
rect 19043 -14942 19075 -14908
rect 19109 -14942 19176 -14908
rect 19210 -14942 19245 -14908
rect 19043 -14998 19245 -14942
rect 17755 -15065 17957 -15032
rect 19043 -15032 19075 -14998
rect 19109 -15032 19176 -14998
rect 19210 -15032 19245 -14998
rect 20331 -14042 20363 -14008
rect 20397 -14042 20464 -14008
rect 20498 -14042 20533 -14008
rect 21619 -14008 21821 -13979
rect 20331 -14098 20533 -14042
rect 20331 -14132 20363 -14098
rect 20397 -14132 20464 -14098
rect 20498 -14132 20533 -14098
rect 20331 -14188 20533 -14132
rect 20331 -14222 20363 -14188
rect 20397 -14222 20464 -14188
rect 20498 -14222 20533 -14188
rect 20331 -14278 20533 -14222
rect 20331 -14312 20363 -14278
rect 20397 -14312 20464 -14278
rect 20498 -14312 20533 -14278
rect 20331 -14368 20533 -14312
rect 20331 -14402 20363 -14368
rect 20397 -14402 20464 -14368
rect 20498 -14402 20533 -14368
rect 20331 -14458 20533 -14402
rect 20331 -14492 20363 -14458
rect 20397 -14492 20464 -14458
rect 20498 -14492 20533 -14458
rect 20331 -14548 20533 -14492
rect 20331 -14582 20363 -14548
rect 20397 -14582 20464 -14548
rect 20498 -14582 20533 -14548
rect 20331 -14638 20533 -14582
rect 20331 -14672 20363 -14638
rect 20397 -14672 20464 -14638
rect 20498 -14672 20533 -14638
rect 20331 -14728 20533 -14672
rect 20331 -14762 20363 -14728
rect 20397 -14762 20464 -14728
rect 20498 -14762 20533 -14728
rect 20331 -14818 20533 -14762
rect 20331 -14852 20363 -14818
rect 20397 -14852 20464 -14818
rect 20498 -14852 20533 -14818
rect 20331 -14908 20533 -14852
rect 20331 -14942 20363 -14908
rect 20397 -14942 20464 -14908
rect 20498 -14942 20533 -14908
rect 20331 -14998 20533 -14942
rect 19043 -15065 19245 -15032
rect 20331 -15032 20363 -14998
rect 20397 -15032 20464 -14998
rect 20498 -15032 20533 -14998
rect 21619 -14042 21651 -14008
rect 21685 -14042 21752 -14008
rect 21786 -14042 21821 -14008
rect 22907 -14008 23109 -13979
rect 21619 -14098 21821 -14042
rect 21619 -14132 21651 -14098
rect 21685 -14132 21752 -14098
rect 21786 -14132 21821 -14098
rect 21619 -14188 21821 -14132
rect 21619 -14222 21651 -14188
rect 21685 -14222 21752 -14188
rect 21786 -14222 21821 -14188
rect 21619 -14278 21821 -14222
rect 21619 -14312 21651 -14278
rect 21685 -14312 21752 -14278
rect 21786 -14312 21821 -14278
rect 21619 -14368 21821 -14312
rect 21619 -14402 21651 -14368
rect 21685 -14402 21752 -14368
rect 21786 -14402 21821 -14368
rect 21619 -14458 21821 -14402
rect 21619 -14492 21651 -14458
rect 21685 -14492 21752 -14458
rect 21786 -14492 21821 -14458
rect 21619 -14548 21821 -14492
rect 21619 -14582 21651 -14548
rect 21685 -14582 21752 -14548
rect 21786 -14582 21821 -14548
rect 21619 -14638 21821 -14582
rect 21619 -14672 21651 -14638
rect 21685 -14672 21752 -14638
rect 21786 -14672 21821 -14638
rect 21619 -14728 21821 -14672
rect 21619 -14762 21651 -14728
rect 21685 -14762 21752 -14728
rect 21786 -14762 21821 -14728
rect 21619 -14818 21821 -14762
rect 21619 -14852 21651 -14818
rect 21685 -14852 21752 -14818
rect 21786 -14852 21821 -14818
rect 21619 -14908 21821 -14852
rect 21619 -14942 21651 -14908
rect 21685 -14942 21752 -14908
rect 21786 -14942 21821 -14908
rect 21619 -14998 21821 -14942
rect 20331 -15065 20533 -15032
rect 21619 -15032 21651 -14998
rect 21685 -15032 21752 -14998
rect 21786 -15032 21821 -14998
rect 22907 -14042 22939 -14008
rect 22973 -14042 23040 -14008
rect 23074 -14042 23109 -14008
rect 24195 -14008 24397 -13979
rect 22907 -14098 23109 -14042
rect 22907 -14132 22939 -14098
rect 22973 -14132 23040 -14098
rect 23074 -14132 23109 -14098
rect 22907 -14188 23109 -14132
rect 22907 -14222 22939 -14188
rect 22973 -14222 23040 -14188
rect 23074 -14222 23109 -14188
rect 22907 -14278 23109 -14222
rect 22907 -14312 22939 -14278
rect 22973 -14312 23040 -14278
rect 23074 -14312 23109 -14278
rect 22907 -14368 23109 -14312
rect 22907 -14402 22939 -14368
rect 22973 -14402 23040 -14368
rect 23074 -14402 23109 -14368
rect 22907 -14458 23109 -14402
rect 22907 -14492 22939 -14458
rect 22973 -14492 23040 -14458
rect 23074 -14492 23109 -14458
rect 22907 -14548 23109 -14492
rect 22907 -14582 22939 -14548
rect 22973 -14582 23040 -14548
rect 23074 -14582 23109 -14548
rect 22907 -14638 23109 -14582
rect 22907 -14672 22939 -14638
rect 22973 -14672 23040 -14638
rect 23074 -14672 23109 -14638
rect 22907 -14728 23109 -14672
rect 22907 -14762 22939 -14728
rect 22973 -14762 23040 -14728
rect 23074 -14762 23109 -14728
rect 22907 -14818 23109 -14762
rect 22907 -14852 22939 -14818
rect 22973 -14852 23040 -14818
rect 23074 -14852 23109 -14818
rect 22907 -14908 23109 -14852
rect 22907 -14942 22939 -14908
rect 22973 -14942 23040 -14908
rect 23074 -14942 23109 -14908
rect 22907 -14998 23109 -14942
rect 21619 -15065 21821 -15032
rect 22907 -15032 22939 -14998
rect 22973 -15032 23040 -14998
rect 23074 -15032 23109 -14998
rect 24195 -14042 24227 -14008
rect 24261 -14042 24328 -14008
rect 24362 -14042 24397 -14008
rect 25483 -14008 25685 -13979
rect 24195 -14098 24397 -14042
rect 24195 -14132 24227 -14098
rect 24261 -14132 24328 -14098
rect 24362 -14132 24397 -14098
rect 24195 -14188 24397 -14132
rect 24195 -14222 24227 -14188
rect 24261 -14222 24328 -14188
rect 24362 -14222 24397 -14188
rect 24195 -14278 24397 -14222
rect 24195 -14312 24227 -14278
rect 24261 -14312 24328 -14278
rect 24362 -14312 24397 -14278
rect 24195 -14368 24397 -14312
rect 24195 -14402 24227 -14368
rect 24261 -14402 24328 -14368
rect 24362 -14402 24397 -14368
rect 24195 -14458 24397 -14402
rect 24195 -14492 24227 -14458
rect 24261 -14492 24328 -14458
rect 24362 -14492 24397 -14458
rect 24195 -14548 24397 -14492
rect 24195 -14582 24227 -14548
rect 24261 -14582 24328 -14548
rect 24362 -14582 24397 -14548
rect 24195 -14638 24397 -14582
rect 24195 -14672 24227 -14638
rect 24261 -14672 24328 -14638
rect 24362 -14672 24397 -14638
rect 24195 -14728 24397 -14672
rect 24195 -14762 24227 -14728
rect 24261 -14762 24328 -14728
rect 24362 -14762 24397 -14728
rect 24195 -14818 24397 -14762
rect 24195 -14852 24227 -14818
rect 24261 -14852 24328 -14818
rect 24362 -14852 24397 -14818
rect 24195 -14908 24397 -14852
rect 24195 -14942 24227 -14908
rect 24261 -14942 24328 -14908
rect 24362 -14942 24397 -14908
rect 24195 -14998 24397 -14942
rect 22907 -15065 23109 -15032
rect 24195 -15032 24227 -14998
rect 24261 -15032 24328 -14998
rect 24362 -15032 24397 -14998
rect 25483 -14042 25515 -14008
rect 25549 -14042 25616 -14008
rect 25650 -14042 25685 -14008
rect 26771 -14008 26872 -13979
rect 25483 -14098 25685 -14042
rect 25483 -14132 25515 -14098
rect 25549 -14132 25616 -14098
rect 25650 -14132 25685 -14098
rect 25483 -14188 25685 -14132
rect 25483 -14222 25515 -14188
rect 25549 -14222 25616 -14188
rect 25650 -14222 25685 -14188
rect 25483 -14278 25685 -14222
rect 25483 -14312 25515 -14278
rect 25549 -14312 25616 -14278
rect 25650 -14312 25685 -14278
rect 25483 -14368 25685 -14312
rect 25483 -14402 25515 -14368
rect 25549 -14402 25616 -14368
rect 25650 -14402 25685 -14368
rect 25483 -14458 25685 -14402
rect 25483 -14492 25515 -14458
rect 25549 -14492 25616 -14458
rect 25650 -14492 25685 -14458
rect 25483 -14548 25685 -14492
rect 25483 -14582 25515 -14548
rect 25549 -14582 25616 -14548
rect 25650 -14582 25685 -14548
rect 25483 -14638 25685 -14582
rect 25483 -14672 25515 -14638
rect 25549 -14672 25616 -14638
rect 25650 -14672 25685 -14638
rect 25483 -14728 25685 -14672
rect 25483 -14762 25515 -14728
rect 25549 -14762 25616 -14728
rect 25650 -14762 25685 -14728
rect 25483 -14818 25685 -14762
rect 25483 -14852 25515 -14818
rect 25549 -14852 25616 -14818
rect 25650 -14852 25685 -14818
rect 25483 -14908 25685 -14852
rect 25483 -14942 25515 -14908
rect 25549 -14942 25616 -14908
rect 25650 -14942 25685 -14908
rect 25483 -14998 25685 -14942
rect 24195 -15065 24397 -15032
rect 25483 -15032 25515 -14998
rect 25549 -15032 25616 -14998
rect 25650 -15032 25685 -14998
rect 26771 -14042 26803 -14008
rect 26837 -14042 26872 -14008
rect 26771 -14098 26872 -14042
rect 26771 -14132 26803 -14098
rect 26837 -14132 26872 -14098
rect 26771 -14188 26872 -14132
rect 26771 -14222 26803 -14188
rect 26837 -14222 26872 -14188
rect 26771 -14278 26872 -14222
rect 26771 -14312 26803 -14278
rect 26837 -14312 26872 -14278
rect 26771 -14368 26872 -14312
rect 26771 -14402 26803 -14368
rect 26837 -14402 26872 -14368
rect 26771 -14458 26872 -14402
rect 26771 -14492 26803 -14458
rect 26837 -14492 26872 -14458
rect 26771 -14548 26872 -14492
rect 26771 -14582 26803 -14548
rect 26837 -14582 26872 -14548
rect 26771 -14638 26872 -14582
rect 26771 -14672 26803 -14638
rect 26837 -14672 26872 -14638
rect 26771 -14728 26872 -14672
rect 26771 -14762 26803 -14728
rect 26837 -14762 26872 -14728
rect 26771 -14818 26872 -14762
rect 26771 -14852 26803 -14818
rect 26837 -14852 26872 -14818
rect 26771 -14908 26872 -14852
rect 26771 -14942 26803 -14908
rect 26837 -14942 26872 -14908
rect 26771 -14998 26872 -14942
rect 25483 -15065 25685 -15032
rect 26771 -15032 26803 -14998
rect 26837 -15032 26872 -14998
rect 26771 -15065 26872 -15032
rect 16568 -15099 26872 -15065
rect 16568 -15133 16684 -15099
rect 16718 -15133 16774 -15099
rect 16808 -15133 16864 -15099
rect 16898 -15133 16954 -15099
rect 16988 -15133 17044 -15099
rect 17078 -15133 17134 -15099
rect 17168 -15133 17224 -15099
rect 17258 -15133 17314 -15099
rect 17348 -15133 17404 -15099
rect 17438 -15133 17494 -15099
rect 17528 -15133 17584 -15099
rect 17618 -15133 17674 -15099
rect 17708 -15133 17764 -15099
rect 17798 -15133 17972 -15099
rect 18006 -15133 18062 -15099
rect 18096 -15133 18152 -15099
rect 18186 -15133 18242 -15099
rect 18276 -15133 18332 -15099
rect 18366 -15133 18422 -15099
rect 18456 -15133 18512 -15099
rect 18546 -15133 18602 -15099
rect 18636 -15133 18692 -15099
rect 18726 -15133 18782 -15099
rect 18816 -15133 18872 -15099
rect 18906 -15133 18962 -15099
rect 18996 -15133 19052 -15099
rect 19086 -15133 19260 -15099
rect 19294 -15133 19350 -15099
rect 19384 -15133 19440 -15099
rect 19474 -15133 19530 -15099
rect 19564 -15133 19620 -15099
rect 19654 -15133 19710 -15099
rect 19744 -15133 19800 -15099
rect 19834 -15133 19890 -15099
rect 19924 -15133 19980 -15099
rect 20014 -15133 20070 -15099
rect 20104 -15133 20160 -15099
rect 20194 -15133 20250 -15099
rect 20284 -15133 20340 -15099
rect 20374 -15133 20548 -15099
rect 20582 -15133 20638 -15099
rect 20672 -15133 20728 -15099
rect 20762 -15133 20818 -15099
rect 20852 -15133 20908 -15099
rect 20942 -15133 20998 -15099
rect 21032 -15133 21088 -15099
rect 21122 -15133 21178 -15099
rect 21212 -15133 21268 -15099
rect 21302 -15133 21358 -15099
rect 21392 -15133 21448 -15099
rect 21482 -15133 21538 -15099
rect 21572 -15133 21628 -15099
rect 21662 -15133 21836 -15099
rect 21870 -15133 21926 -15099
rect 21960 -15133 22016 -15099
rect 22050 -15133 22106 -15099
rect 22140 -15133 22196 -15099
rect 22230 -15133 22286 -15099
rect 22320 -15133 22376 -15099
rect 22410 -15133 22466 -15099
rect 22500 -15133 22556 -15099
rect 22590 -15133 22646 -15099
rect 22680 -15133 22736 -15099
rect 22770 -15133 22826 -15099
rect 22860 -15133 22916 -15099
rect 22950 -15133 23124 -15099
rect 23158 -15133 23214 -15099
rect 23248 -15133 23304 -15099
rect 23338 -15133 23394 -15099
rect 23428 -15133 23484 -15099
rect 23518 -15133 23574 -15099
rect 23608 -15133 23664 -15099
rect 23698 -15133 23754 -15099
rect 23788 -15133 23844 -15099
rect 23878 -15133 23934 -15099
rect 23968 -15133 24024 -15099
rect 24058 -15133 24114 -15099
rect 24148 -15133 24204 -15099
rect 24238 -15133 24412 -15099
rect 24446 -15133 24502 -15099
rect 24536 -15133 24592 -15099
rect 24626 -15133 24682 -15099
rect 24716 -15133 24772 -15099
rect 24806 -15133 24862 -15099
rect 24896 -15133 24952 -15099
rect 24986 -15133 25042 -15099
rect 25076 -15133 25132 -15099
rect 25166 -15133 25222 -15099
rect 25256 -15133 25312 -15099
rect 25346 -15133 25402 -15099
rect 25436 -15133 25492 -15099
rect 25526 -15133 25700 -15099
rect 25734 -15133 25790 -15099
rect 25824 -15133 25880 -15099
rect 25914 -15133 25970 -15099
rect 26004 -15133 26060 -15099
rect 26094 -15133 26150 -15099
rect 26184 -15133 26240 -15099
rect 26274 -15133 26330 -15099
rect 26364 -15133 26420 -15099
rect 26454 -15133 26510 -15099
rect 26544 -15133 26600 -15099
rect 26634 -15133 26690 -15099
rect 26724 -15133 26780 -15099
rect 26814 -15133 26872 -15099
rect 16568 -15200 26872 -15133
rect 16568 -15234 16684 -15200
rect 16718 -15234 16774 -15200
rect 16808 -15234 16864 -15200
rect 16898 -15234 16954 -15200
rect 16988 -15234 17044 -15200
rect 17078 -15234 17134 -15200
rect 17168 -15234 17224 -15200
rect 17258 -15234 17314 -15200
rect 17348 -15234 17404 -15200
rect 17438 -15234 17494 -15200
rect 17528 -15234 17584 -15200
rect 17618 -15234 17674 -15200
rect 17708 -15234 17764 -15200
rect 17798 -15234 17972 -15200
rect 18006 -15234 18062 -15200
rect 18096 -15234 18152 -15200
rect 18186 -15234 18242 -15200
rect 18276 -15234 18332 -15200
rect 18366 -15234 18422 -15200
rect 18456 -15234 18512 -15200
rect 18546 -15234 18602 -15200
rect 18636 -15234 18692 -15200
rect 18726 -15234 18782 -15200
rect 18816 -15234 18872 -15200
rect 18906 -15234 18962 -15200
rect 18996 -15234 19052 -15200
rect 19086 -15234 19260 -15200
rect 19294 -15234 19350 -15200
rect 19384 -15234 19440 -15200
rect 19474 -15234 19530 -15200
rect 19564 -15234 19620 -15200
rect 19654 -15234 19710 -15200
rect 19744 -15234 19800 -15200
rect 19834 -15234 19890 -15200
rect 19924 -15234 19980 -15200
rect 20014 -15234 20070 -15200
rect 20104 -15234 20160 -15200
rect 20194 -15234 20250 -15200
rect 20284 -15234 20340 -15200
rect 20374 -15234 20548 -15200
rect 20582 -15234 20638 -15200
rect 20672 -15234 20728 -15200
rect 20762 -15234 20818 -15200
rect 20852 -15234 20908 -15200
rect 20942 -15234 20998 -15200
rect 21032 -15234 21088 -15200
rect 21122 -15234 21178 -15200
rect 21212 -15234 21268 -15200
rect 21302 -15234 21358 -15200
rect 21392 -15234 21448 -15200
rect 21482 -15234 21538 -15200
rect 21572 -15234 21628 -15200
rect 21662 -15234 21836 -15200
rect 21870 -15234 21926 -15200
rect 21960 -15234 22016 -15200
rect 22050 -15234 22106 -15200
rect 22140 -15234 22196 -15200
rect 22230 -15234 22286 -15200
rect 22320 -15234 22376 -15200
rect 22410 -15234 22466 -15200
rect 22500 -15234 22556 -15200
rect 22590 -15234 22646 -15200
rect 22680 -15234 22736 -15200
rect 22770 -15234 22826 -15200
rect 22860 -15234 22916 -15200
rect 22950 -15234 23124 -15200
rect 23158 -15234 23214 -15200
rect 23248 -15234 23304 -15200
rect 23338 -15234 23394 -15200
rect 23428 -15234 23484 -15200
rect 23518 -15234 23574 -15200
rect 23608 -15234 23664 -15200
rect 23698 -15234 23754 -15200
rect 23788 -15234 23844 -15200
rect 23878 -15234 23934 -15200
rect 23968 -15234 24024 -15200
rect 24058 -15234 24114 -15200
rect 24148 -15234 24204 -15200
rect 24238 -15234 24412 -15200
rect 24446 -15234 24502 -15200
rect 24536 -15234 24592 -15200
rect 24626 -15234 24682 -15200
rect 24716 -15234 24772 -15200
rect 24806 -15234 24862 -15200
rect 24896 -15234 24952 -15200
rect 24986 -15234 25042 -15200
rect 25076 -15234 25132 -15200
rect 25166 -15234 25222 -15200
rect 25256 -15234 25312 -15200
rect 25346 -15234 25402 -15200
rect 25436 -15234 25492 -15200
rect 25526 -15234 25700 -15200
rect 25734 -15234 25790 -15200
rect 25824 -15234 25880 -15200
rect 25914 -15234 25970 -15200
rect 26004 -15234 26060 -15200
rect 26094 -15234 26150 -15200
rect 26184 -15234 26240 -15200
rect 26274 -15234 26330 -15200
rect 26364 -15234 26420 -15200
rect 26454 -15234 26510 -15200
rect 26544 -15234 26600 -15200
rect 26634 -15234 26690 -15200
rect 26724 -15234 26780 -15200
rect 26814 -15234 26872 -15200
rect 16568 -15267 26872 -15234
rect 16568 -15296 16669 -15267
rect 16568 -15330 16600 -15296
rect 16634 -15330 16669 -15296
rect 17755 -15296 17957 -15267
rect 16568 -15386 16669 -15330
rect 16568 -15420 16600 -15386
rect 16634 -15420 16669 -15386
rect 16568 -15476 16669 -15420
rect 16568 -15510 16600 -15476
rect 16634 -15510 16669 -15476
rect 16568 -15566 16669 -15510
rect 16568 -15600 16600 -15566
rect 16634 -15600 16669 -15566
rect 16568 -15656 16669 -15600
rect 16568 -15690 16600 -15656
rect 16634 -15690 16669 -15656
rect 16568 -15746 16669 -15690
rect 16568 -15780 16600 -15746
rect 16634 -15780 16669 -15746
rect 16568 -15836 16669 -15780
rect 16568 -15870 16600 -15836
rect 16634 -15870 16669 -15836
rect 16568 -15926 16669 -15870
rect 16568 -15960 16600 -15926
rect 16634 -15960 16669 -15926
rect 16568 -16016 16669 -15960
rect 16568 -16050 16600 -16016
rect 16634 -16050 16669 -16016
rect 16568 -16106 16669 -16050
rect 16568 -16140 16600 -16106
rect 16634 -16140 16669 -16106
rect 16568 -16196 16669 -16140
rect 16568 -16230 16600 -16196
rect 16634 -16230 16669 -16196
rect 16568 -16286 16669 -16230
rect 16568 -16320 16600 -16286
rect 16634 -16320 16669 -16286
rect 17755 -15330 17787 -15296
rect 17821 -15330 17888 -15296
rect 17922 -15330 17957 -15296
rect 19043 -15296 19245 -15267
rect 17755 -15386 17957 -15330
rect 17755 -15420 17787 -15386
rect 17821 -15420 17888 -15386
rect 17922 -15420 17957 -15386
rect 17755 -15476 17957 -15420
rect 17755 -15510 17787 -15476
rect 17821 -15510 17888 -15476
rect 17922 -15510 17957 -15476
rect 17755 -15566 17957 -15510
rect 17755 -15600 17787 -15566
rect 17821 -15600 17888 -15566
rect 17922 -15600 17957 -15566
rect 17755 -15656 17957 -15600
rect 17755 -15690 17787 -15656
rect 17821 -15690 17888 -15656
rect 17922 -15690 17957 -15656
rect 17755 -15746 17957 -15690
rect 17755 -15780 17787 -15746
rect 17821 -15780 17888 -15746
rect 17922 -15780 17957 -15746
rect 17755 -15836 17957 -15780
rect 17755 -15870 17787 -15836
rect 17821 -15870 17888 -15836
rect 17922 -15870 17957 -15836
rect 17755 -15926 17957 -15870
rect 17755 -15960 17787 -15926
rect 17821 -15960 17888 -15926
rect 17922 -15960 17957 -15926
rect 17755 -16016 17957 -15960
rect 17755 -16050 17787 -16016
rect 17821 -16050 17888 -16016
rect 17922 -16050 17957 -16016
rect 17755 -16106 17957 -16050
rect 17755 -16140 17787 -16106
rect 17821 -16140 17888 -16106
rect 17922 -16140 17957 -16106
rect 17755 -16196 17957 -16140
rect 17755 -16230 17787 -16196
rect 17821 -16230 17888 -16196
rect 17922 -16230 17957 -16196
rect 17755 -16286 17957 -16230
rect 16568 -16353 16669 -16320
rect 17755 -16320 17787 -16286
rect 17821 -16320 17888 -16286
rect 17922 -16320 17957 -16286
rect 19043 -15330 19075 -15296
rect 19109 -15330 19176 -15296
rect 19210 -15330 19245 -15296
rect 20331 -15296 20533 -15267
rect 19043 -15386 19245 -15330
rect 19043 -15420 19075 -15386
rect 19109 -15420 19176 -15386
rect 19210 -15420 19245 -15386
rect 19043 -15476 19245 -15420
rect 19043 -15510 19075 -15476
rect 19109 -15510 19176 -15476
rect 19210 -15510 19245 -15476
rect 19043 -15566 19245 -15510
rect 19043 -15600 19075 -15566
rect 19109 -15600 19176 -15566
rect 19210 -15600 19245 -15566
rect 19043 -15656 19245 -15600
rect 19043 -15690 19075 -15656
rect 19109 -15690 19176 -15656
rect 19210 -15690 19245 -15656
rect 19043 -15746 19245 -15690
rect 19043 -15780 19075 -15746
rect 19109 -15780 19176 -15746
rect 19210 -15780 19245 -15746
rect 19043 -15836 19245 -15780
rect 19043 -15870 19075 -15836
rect 19109 -15870 19176 -15836
rect 19210 -15870 19245 -15836
rect 19043 -15926 19245 -15870
rect 19043 -15960 19075 -15926
rect 19109 -15960 19176 -15926
rect 19210 -15960 19245 -15926
rect 19043 -16016 19245 -15960
rect 19043 -16050 19075 -16016
rect 19109 -16050 19176 -16016
rect 19210 -16050 19245 -16016
rect 19043 -16106 19245 -16050
rect 19043 -16140 19075 -16106
rect 19109 -16140 19176 -16106
rect 19210 -16140 19245 -16106
rect 19043 -16196 19245 -16140
rect 19043 -16230 19075 -16196
rect 19109 -16230 19176 -16196
rect 19210 -16230 19245 -16196
rect 19043 -16286 19245 -16230
rect 17755 -16353 17957 -16320
rect 19043 -16320 19075 -16286
rect 19109 -16320 19176 -16286
rect 19210 -16320 19245 -16286
rect 20331 -15330 20363 -15296
rect 20397 -15330 20464 -15296
rect 20498 -15330 20533 -15296
rect 21619 -15296 21821 -15267
rect 20331 -15386 20533 -15330
rect 20331 -15420 20363 -15386
rect 20397 -15420 20464 -15386
rect 20498 -15420 20533 -15386
rect 20331 -15476 20533 -15420
rect 20331 -15510 20363 -15476
rect 20397 -15510 20464 -15476
rect 20498 -15510 20533 -15476
rect 20331 -15566 20533 -15510
rect 20331 -15600 20363 -15566
rect 20397 -15600 20464 -15566
rect 20498 -15600 20533 -15566
rect 20331 -15656 20533 -15600
rect 20331 -15690 20363 -15656
rect 20397 -15690 20464 -15656
rect 20498 -15690 20533 -15656
rect 20331 -15746 20533 -15690
rect 20331 -15780 20363 -15746
rect 20397 -15780 20464 -15746
rect 20498 -15780 20533 -15746
rect 20331 -15836 20533 -15780
rect 20331 -15870 20363 -15836
rect 20397 -15870 20464 -15836
rect 20498 -15870 20533 -15836
rect 20331 -15926 20533 -15870
rect 20331 -15960 20363 -15926
rect 20397 -15960 20464 -15926
rect 20498 -15960 20533 -15926
rect 20331 -16016 20533 -15960
rect 20331 -16050 20363 -16016
rect 20397 -16050 20464 -16016
rect 20498 -16050 20533 -16016
rect 20331 -16106 20533 -16050
rect 20331 -16140 20363 -16106
rect 20397 -16140 20464 -16106
rect 20498 -16140 20533 -16106
rect 20331 -16196 20533 -16140
rect 20331 -16230 20363 -16196
rect 20397 -16230 20464 -16196
rect 20498 -16230 20533 -16196
rect 20331 -16286 20533 -16230
rect 19043 -16353 19245 -16320
rect 20331 -16320 20363 -16286
rect 20397 -16320 20464 -16286
rect 20498 -16320 20533 -16286
rect 21619 -15330 21651 -15296
rect 21685 -15330 21752 -15296
rect 21786 -15330 21821 -15296
rect 22907 -15296 23109 -15267
rect 21619 -15386 21821 -15330
rect 21619 -15420 21651 -15386
rect 21685 -15420 21752 -15386
rect 21786 -15420 21821 -15386
rect 21619 -15476 21821 -15420
rect 21619 -15510 21651 -15476
rect 21685 -15510 21752 -15476
rect 21786 -15510 21821 -15476
rect 21619 -15566 21821 -15510
rect 21619 -15600 21651 -15566
rect 21685 -15600 21752 -15566
rect 21786 -15600 21821 -15566
rect 21619 -15656 21821 -15600
rect 21619 -15690 21651 -15656
rect 21685 -15690 21752 -15656
rect 21786 -15690 21821 -15656
rect 21619 -15746 21821 -15690
rect 21619 -15780 21651 -15746
rect 21685 -15780 21752 -15746
rect 21786 -15780 21821 -15746
rect 21619 -15836 21821 -15780
rect 21619 -15870 21651 -15836
rect 21685 -15870 21752 -15836
rect 21786 -15870 21821 -15836
rect 21619 -15926 21821 -15870
rect 21619 -15960 21651 -15926
rect 21685 -15960 21752 -15926
rect 21786 -15960 21821 -15926
rect 21619 -16016 21821 -15960
rect 21619 -16050 21651 -16016
rect 21685 -16050 21752 -16016
rect 21786 -16050 21821 -16016
rect 21619 -16106 21821 -16050
rect 21619 -16140 21651 -16106
rect 21685 -16140 21752 -16106
rect 21786 -16140 21821 -16106
rect 21619 -16196 21821 -16140
rect 21619 -16230 21651 -16196
rect 21685 -16230 21752 -16196
rect 21786 -16230 21821 -16196
rect 21619 -16286 21821 -16230
rect 20331 -16353 20533 -16320
rect 21619 -16320 21651 -16286
rect 21685 -16320 21752 -16286
rect 21786 -16320 21821 -16286
rect 22907 -15330 22939 -15296
rect 22973 -15330 23040 -15296
rect 23074 -15330 23109 -15296
rect 24195 -15296 24397 -15267
rect 22907 -15386 23109 -15330
rect 22907 -15420 22939 -15386
rect 22973 -15420 23040 -15386
rect 23074 -15420 23109 -15386
rect 22907 -15476 23109 -15420
rect 22907 -15510 22939 -15476
rect 22973 -15510 23040 -15476
rect 23074 -15510 23109 -15476
rect 22907 -15566 23109 -15510
rect 22907 -15600 22939 -15566
rect 22973 -15600 23040 -15566
rect 23074 -15600 23109 -15566
rect 22907 -15656 23109 -15600
rect 22907 -15690 22939 -15656
rect 22973 -15690 23040 -15656
rect 23074 -15690 23109 -15656
rect 22907 -15746 23109 -15690
rect 22907 -15780 22939 -15746
rect 22973 -15780 23040 -15746
rect 23074 -15780 23109 -15746
rect 22907 -15836 23109 -15780
rect 22907 -15870 22939 -15836
rect 22973 -15870 23040 -15836
rect 23074 -15870 23109 -15836
rect 22907 -15926 23109 -15870
rect 22907 -15960 22939 -15926
rect 22973 -15960 23040 -15926
rect 23074 -15960 23109 -15926
rect 22907 -16016 23109 -15960
rect 22907 -16050 22939 -16016
rect 22973 -16050 23040 -16016
rect 23074 -16050 23109 -16016
rect 22907 -16106 23109 -16050
rect 22907 -16140 22939 -16106
rect 22973 -16140 23040 -16106
rect 23074 -16140 23109 -16106
rect 22907 -16196 23109 -16140
rect 22907 -16230 22939 -16196
rect 22973 -16230 23040 -16196
rect 23074 -16230 23109 -16196
rect 22907 -16286 23109 -16230
rect 21619 -16353 21821 -16320
rect 22907 -16320 22939 -16286
rect 22973 -16320 23040 -16286
rect 23074 -16320 23109 -16286
rect 24195 -15330 24227 -15296
rect 24261 -15330 24328 -15296
rect 24362 -15330 24397 -15296
rect 25483 -15296 25685 -15267
rect 24195 -15386 24397 -15330
rect 24195 -15420 24227 -15386
rect 24261 -15420 24328 -15386
rect 24362 -15420 24397 -15386
rect 24195 -15476 24397 -15420
rect 24195 -15510 24227 -15476
rect 24261 -15510 24328 -15476
rect 24362 -15510 24397 -15476
rect 24195 -15566 24397 -15510
rect 24195 -15600 24227 -15566
rect 24261 -15600 24328 -15566
rect 24362 -15600 24397 -15566
rect 24195 -15656 24397 -15600
rect 24195 -15690 24227 -15656
rect 24261 -15690 24328 -15656
rect 24362 -15690 24397 -15656
rect 24195 -15746 24397 -15690
rect 24195 -15780 24227 -15746
rect 24261 -15780 24328 -15746
rect 24362 -15780 24397 -15746
rect 24195 -15836 24397 -15780
rect 24195 -15870 24227 -15836
rect 24261 -15870 24328 -15836
rect 24362 -15870 24397 -15836
rect 24195 -15926 24397 -15870
rect 24195 -15960 24227 -15926
rect 24261 -15960 24328 -15926
rect 24362 -15960 24397 -15926
rect 24195 -16016 24397 -15960
rect 24195 -16050 24227 -16016
rect 24261 -16050 24328 -16016
rect 24362 -16050 24397 -16016
rect 24195 -16106 24397 -16050
rect 24195 -16140 24227 -16106
rect 24261 -16140 24328 -16106
rect 24362 -16140 24397 -16106
rect 24195 -16196 24397 -16140
rect 24195 -16230 24227 -16196
rect 24261 -16230 24328 -16196
rect 24362 -16230 24397 -16196
rect 24195 -16286 24397 -16230
rect 22907 -16353 23109 -16320
rect 24195 -16320 24227 -16286
rect 24261 -16320 24328 -16286
rect 24362 -16320 24397 -16286
rect 25483 -15330 25515 -15296
rect 25549 -15330 25616 -15296
rect 25650 -15330 25685 -15296
rect 26771 -15296 26872 -15267
rect 25483 -15386 25685 -15330
rect 25483 -15420 25515 -15386
rect 25549 -15420 25616 -15386
rect 25650 -15420 25685 -15386
rect 25483 -15476 25685 -15420
rect 25483 -15510 25515 -15476
rect 25549 -15510 25616 -15476
rect 25650 -15510 25685 -15476
rect 25483 -15566 25685 -15510
rect 25483 -15600 25515 -15566
rect 25549 -15600 25616 -15566
rect 25650 -15600 25685 -15566
rect 25483 -15656 25685 -15600
rect 25483 -15690 25515 -15656
rect 25549 -15690 25616 -15656
rect 25650 -15690 25685 -15656
rect 25483 -15746 25685 -15690
rect 25483 -15780 25515 -15746
rect 25549 -15780 25616 -15746
rect 25650 -15780 25685 -15746
rect 25483 -15836 25685 -15780
rect 25483 -15870 25515 -15836
rect 25549 -15870 25616 -15836
rect 25650 -15870 25685 -15836
rect 25483 -15926 25685 -15870
rect 25483 -15960 25515 -15926
rect 25549 -15960 25616 -15926
rect 25650 -15960 25685 -15926
rect 25483 -16016 25685 -15960
rect 25483 -16050 25515 -16016
rect 25549 -16050 25616 -16016
rect 25650 -16050 25685 -16016
rect 25483 -16106 25685 -16050
rect 25483 -16140 25515 -16106
rect 25549 -16140 25616 -16106
rect 25650 -16140 25685 -16106
rect 25483 -16196 25685 -16140
rect 25483 -16230 25515 -16196
rect 25549 -16230 25616 -16196
rect 25650 -16230 25685 -16196
rect 25483 -16286 25685 -16230
rect 24195 -16353 24397 -16320
rect 25483 -16320 25515 -16286
rect 25549 -16320 25616 -16286
rect 25650 -16320 25685 -16286
rect 26771 -15330 26803 -15296
rect 26837 -15330 26872 -15296
rect 26771 -15386 26872 -15330
rect 26771 -15420 26803 -15386
rect 26837 -15420 26872 -15386
rect 26771 -15476 26872 -15420
rect 26771 -15510 26803 -15476
rect 26837 -15510 26872 -15476
rect 26771 -15566 26872 -15510
rect 26771 -15600 26803 -15566
rect 26837 -15600 26872 -15566
rect 26771 -15656 26872 -15600
rect 26771 -15690 26803 -15656
rect 26837 -15690 26872 -15656
rect 26771 -15746 26872 -15690
rect 26771 -15780 26803 -15746
rect 26837 -15780 26872 -15746
rect 26771 -15836 26872 -15780
rect 26771 -15870 26803 -15836
rect 26837 -15870 26872 -15836
rect 26771 -15926 26872 -15870
rect 26771 -15960 26803 -15926
rect 26837 -15960 26872 -15926
rect 26771 -16016 26872 -15960
rect 26771 -16050 26803 -16016
rect 26837 -16050 26872 -16016
rect 26771 -16106 26872 -16050
rect 26771 -16140 26803 -16106
rect 26837 -16140 26872 -16106
rect 26771 -16196 26872 -16140
rect 26771 -16230 26803 -16196
rect 26837 -16230 26872 -16196
rect 26771 -16286 26872 -16230
rect 25483 -16353 25685 -16320
rect 26771 -16320 26803 -16286
rect 26837 -16320 26872 -16286
rect 26771 -16353 26872 -16320
rect 16568 -16387 26872 -16353
rect 16568 -16421 16684 -16387
rect 16718 -16421 16774 -16387
rect 16808 -16421 16864 -16387
rect 16898 -16421 16954 -16387
rect 16988 -16421 17044 -16387
rect 17078 -16421 17134 -16387
rect 17168 -16421 17224 -16387
rect 17258 -16421 17314 -16387
rect 17348 -16421 17404 -16387
rect 17438 -16421 17494 -16387
rect 17528 -16421 17584 -16387
rect 17618 -16421 17674 -16387
rect 17708 -16421 17764 -16387
rect 17798 -16421 17972 -16387
rect 18006 -16421 18062 -16387
rect 18096 -16421 18152 -16387
rect 18186 -16421 18242 -16387
rect 18276 -16421 18332 -16387
rect 18366 -16421 18422 -16387
rect 18456 -16421 18512 -16387
rect 18546 -16421 18602 -16387
rect 18636 -16421 18692 -16387
rect 18726 -16421 18782 -16387
rect 18816 -16421 18872 -16387
rect 18906 -16421 18962 -16387
rect 18996 -16421 19052 -16387
rect 19086 -16421 19260 -16387
rect 19294 -16421 19350 -16387
rect 19384 -16421 19440 -16387
rect 19474 -16421 19530 -16387
rect 19564 -16421 19620 -16387
rect 19654 -16421 19710 -16387
rect 19744 -16421 19800 -16387
rect 19834 -16421 19890 -16387
rect 19924 -16421 19980 -16387
rect 20014 -16421 20070 -16387
rect 20104 -16421 20160 -16387
rect 20194 -16421 20250 -16387
rect 20284 -16421 20340 -16387
rect 20374 -16421 20548 -16387
rect 20582 -16421 20638 -16387
rect 20672 -16421 20728 -16387
rect 20762 -16421 20818 -16387
rect 20852 -16421 20908 -16387
rect 20942 -16421 20998 -16387
rect 21032 -16421 21088 -16387
rect 21122 -16421 21178 -16387
rect 21212 -16421 21268 -16387
rect 21302 -16421 21358 -16387
rect 21392 -16421 21448 -16387
rect 21482 -16421 21538 -16387
rect 21572 -16421 21628 -16387
rect 21662 -16421 21836 -16387
rect 21870 -16421 21926 -16387
rect 21960 -16421 22016 -16387
rect 22050 -16421 22106 -16387
rect 22140 -16421 22196 -16387
rect 22230 -16421 22286 -16387
rect 22320 -16421 22376 -16387
rect 22410 -16421 22466 -16387
rect 22500 -16421 22556 -16387
rect 22590 -16421 22646 -16387
rect 22680 -16421 22736 -16387
rect 22770 -16421 22826 -16387
rect 22860 -16421 22916 -16387
rect 22950 -16421 23124 -16387
rect 23158 -16421 23214 -16387
rect 23248 -16421 23304 -16387
rect 23338 -16421 23394 -16387
rect 23428 -16421 23484 -16387
rect 23518 -16421 23574 -16387
rect 23608 -16421 23664 -16387
rect 23698 -16421 23754 -16387
rect 23788 -16421 23844 -16387
rect 23878 -16421 23934 -16387
rect 23968 -16421 24024 -16387
rect 24058 -16421 24114 -16387
rect 24148 -16421 24204 -16387
rect 24238 -16421 24412 -16387
rect 24446 -16421 24502 -16387
rect 24536 -16421 24592 -16387
rect 24626 -16421 24682 -16387
rect 24716 -16421 24772 -16387
rect 24806 -16421 24862 -16387
rect 24896 -16421 24952 -16387
rect 24986 -16421 25042 -16387
rect 25076 -16421 25132 -16387
rect 25166 -16421 25222 -16387
rect 25256 -16421 25312 -16387
rect 25346 -16421 25402 -16387
rect 25436 -16421 25492 -16387
rect 25526 -16421 25700 -16387
rect 25734 -16421 25790 -16387
rect 25824 -16421 25880 -16387
rect 25914 -16421 25970 -16387
rect 26004 -16421 26060 -16387
rect 26094 -16421 26150 -16387
rect 26184 -16421 26240 -16387
rect 26274 -16421 26330 -16387
rect 26364 -16421 26420 -16387
rect 26454 -16421 26510 -16387
rect 26544 -16421 26600 -16387
rect 26634 -16421 26690 -16387
rect 26724 -16421 26780 -16387
rect 26814 -16421 26872 -16387
rect 7278 -16480 13630 -16456
rect 7278 -17050 7302 -16480
rect 13606 -17050 13630 -16480
rect 7278 -17074 13630 -17050
rect 16568 -16488 26872 -16421
rect 16568 -16522 16684 -16488
rect 16718 -16522 16774 -16488
rect 16808 -16522 16864 -16488
rect 16898 -16522 16954 -16488
rect 16988 -16522 17044 -16488
rect 17078 -16522 17134 -16488
rect 17168 -16522 17224 -16488
rect 17258 -16522 17314 -16488
rect 17348 -16522 17404 -16488
rect 17438 -16522 17494 -16488
rect 17528 -16522 17584 -16488
rect 17618 -16522 17674 -16488
rect 17708 -16522 17764 -16488
rect 17798 -16522 17972 -16488
rect 18006 -16522 18062 -16488
rect 18096 -16522 18152 -16488
rect 18186 -16522 18242 -16488
rect 18276 -16522 18332 -16488
rect 18366 -16522 18422 -16488
rect 18456 -16522 18512 -16488
rect 18546 -16522 18602 -16488
rect 18636 -16522 18692 -16488
rect 18726 -16522 18782 -16488
rect 18816 -16522 18872 -16488
rect 18906 -16522 18962 -16488
rect 18996 -16522 19052 -16488
rect 19086 -16522 19260 -16488
rect 19294 -16522 19350 -16488
rect 19384 -16522 19440 -16488
rect 19474 -16522 19530 -16488
rect 19564 -16522 19620 -16488
rect 19654 -16522 19710 -16488
rect 19744 -16522 19800 -16488
rect 19834 -16522 19890 -16488
rect 19924 -16522 19980 -16488
rect 20014 -16522 20070 -16488
rect 20104 -16522 20160 -16488
rect 20194 -16522 20250 -16488
rect 20284 -16522 20340 -16488
rect 20374 -16522 20548 -16488
rect 20582 -16522 20638 -16488
rect 20672 -16522 20728 -16488
rect 20762 -16522 20818 -16488
rect 20852 -16522 20908 -16488
rect 20942 -16522 20998 -16488
rect 21032 -16522 21088 -16488
rect 21122 -16522 21178 -16488
rect 21212 -16522 21268 -16488
rect 21302 -16522 21358 -16488
rect 21392 -16522 21448 -16488
rect 21482 -16522 21538 -16488
rect 21572 -16522 21628 -16488
rect 21662 -16522 21836 -16488
rect 21870 -16522 21926 -16488
rect 21960 -16522 22016 -16488
rect 22050 -16522 22106 -16488
rect 22140 -16522 22196 -16488
rect 22230 -16522 22286 -16488
rect 22320 -16522 22376 -16488
rect 22410 -16522 22466 -16488
rect 22500 -16522 22556 -16488
rect 22590 -16522 22646 -16488
rect 22680 -16522 22736 -16488
rect 22770 -16522 22826 -16488
rect 22860 -16522 22916 -16488
rect 22950 -16522 23124 -16488
rect 23158 -16522 23214 -16488
rect 23248 -16522 23304 -16488
rect 23338 -16522 23394 -16488
rect 23428 -16522 23484 -16488
rect 23518 -16522 23574 -16488
rect 23608 -16522 23664 -16488
rect 23698 -16522 23754 -16488
rect 23788 -16522 23844 -16488
rect 23878 -16522 23934 -16488
rect 23968 -16522 24024 -16488
rect 24058 -16522 24114 -16488
rect 24148 -16522 24204 -16488
rect 24238 -16522 24412 -16488
rect 24446 -16522 24502 -16488
rect 24536 -16522 24592 -16488
rect 24626 -16522 24682 -16488
rect 24716 -16522 24772 -16488
rect 24806 -16522 24862 -16488
rect 24896 -16522 24952 -16488
rect 24986 -16522 25042 -16488
rect 25076 -16522 25132 -16488
rect 25166 -16522 25222 -16488
rect 25256 -16522 25312 -16488
rect 25346 -16522 25402 -16488
rect 25436 -16522 25492 -16488
rect 25526 -16522 25700 -16488
rect 25734 -16522 25790 -16488
rect 25824 -16522 25880 -16488
rect 25914 -16522 25970 -16488
rect 26004 -16522 26060 -16488
rect 26094 -16522 26150 -16488
rect 26184 -16522 26240 -16488
rect 26274 -16522 26330 -16488
rect 26364 -16522 26420 -16488
rect 26454 -16522 26510 -16488
rect 26544 -16522 26600 -16488
rect 26634 -16522 26690 -16488
rect 26724 -16522 26780 -16488
rect 26814 -16522 26872 -16488
rect 16568 -16555 26872 -16522
rect 16568 -16584 16669 -16555
rect 16568 -16618 16600 -16584
rect 16634 -16618 16669 -16584
rect 17755 -16584 17957 -16555
rect 16568 -16674 16669 -16618
rect 16568 -16708 16600 -16674
rect 16634 -16708 16669 -16674
rect 16568 -16764 16669 -16708
rect 16568 -16798 16600 -16764
rect 16634 -16798 16669 -16764
rect 16568 -16854 16669 -16798
rect 16568 -16888 16600 -16854
rect 16634 -16888 16669 -16854
rect 16568 -16944 16669 -16888
rect 16568 -16978 16600 -16944
rect 16634 -16978 16669 -16944
rect 16568 -17034 16669 -16978
rect 16568 -17068 16600 -17034
rect 16634 -17068 16669 -17034
rect 16568 -17124 16669 -17068
rect 16568 -17158 16600 -17124
rect 16634 -17158 16669 -17124
rect 16568 -17214 16669 -17158
rect 16568 -17248 16600 -17214
rect 16634 -17248 16669 -17214
rect 16568 -17304 16669 -17248
rect 16568 -17338 16600 -17304
rect 16634 -17338 16669 -17304
rect 16568 -17394 16669 -17338
rect 16568 -17428 16600 -17394
rect 16634 -17428 16669 -17394
rect 16568 -17484 16669 -17428
rect 16568 -17518 16600 -17484
rect 16634 -17518 16669 -17484
rect 16568 -17574 16669 -17518
rect 16568 -17608 16600 -17574
rect 16634 -17608 16669 -17574
rect 17755 -16618 17787 -16584
rect 17821 -16618 17888 -16584
rect 17922 -16618 17957 -16584
rect 19043 -16584 19245 -16555
rect 17755 -16674 17957 -16618
rect 17755 -16708 17787 -16674
rect 17821 -16708 17888 -16674
rect 17922 -16708 17957 -16674
rect 17755 -16764 17957 -16708
rect 17755 -16798 17787 -16764
rect 17821 -16798 17888 -16764
rect 17922 -16798 17957 -16764
rect 17755 -16854 17957 -16798
rect 17755 -16888 17787 -16854
rect 17821 -16888 17888 -16854
rect 17922 -16888 17957 -16854
rect 17755 -16944 17957 -16888
rect 17755 -16978 17787 -16944
rect 17821 -16978 17888 -16944
rect 17922 -16978 17957 -16944
rect 17755 -17034 17957 -16978
rect 17755 -17068 17787 -17034
rect 17821 -17068 17888 -17034
rect 17922 -17068 17957 -17034
rect 17755 -17124 17957 -17068
rect 17755 -17158 17787 -17124
rect 17821 -17158 17888 -17124
rect 17922 -17158 17957 -17124
rect 17755 -17214 17957 -17158
rect 17755 -17248 17787 -17214
rect 17821 -17248 17888 -17214
rect 17922 -17248 17957 -17214
rect 17755 -17304 17957 -17248
rect 17755 -17338 17787 -17304
rect 17821 -17338 17888 -17304
rect 17922 -17338 17957 -17304
rect 17755 -17394 17957 -17338
rect 17755 -17428 17787 -17394
rect 17821 -17428 17888 -17394
rect 17922 -17428 17957 -17394
rect 17755 -17484 17957 -17428
rect 17755 -17518 17787 -17484
rect 17821 -17518 17888 -17484
rect 17922 -17518 17957 -17484
rect 17755 -17574 17957 -17518
rect 16568 -17641 16669 -17608
rect 17755 -17608 17787 -17574
rect 17821 -17608 17888 -17574
rect 17922 -17608 17957 -17574
rect 19043 -16618 19075 -16584
rect 19109 -16618 19176 -16584
rect 19210 -16618 19245 -16584
rect 20331 -16584 20533 -16555
rect 19043 -16674 19245 -16618
rect 19043 -16708 19075 -16674
rect 19109 -16708 19176 -16674
rect 19210 -16708 19245 -16674
rect 19043 -16764 19245 -16708
rect 19043 -16798 19075 -16764
rect 19109 -16798 19176 -16764
rect 19210 -16798 19245 -16764
rect 19043 -16854 19245 -16798
rect 19043 -16888 19075 -16854
rect 19109 -16888 19176 -16854
rect 19210 -16888 19245 -16854
rect 19043 -16944 19245 -16888
rect 19043 -16978 19075 -16944
rect 19109 -16978 19176 -16944
rect 19210 -16978 19245 -16944
rect 19043 -17034 19245 -16978
rect 19043 -17068 19075 -17034
rect 19109 -17068 19176 -17034
rect 19210 -17068 19245 -17034
rect 19043 -17124 19245 -17068
rect 19043 -17158 19075 -17124
rect 19109 -17158 19176 -17124
rect 19210 -17158 19245 -17124
rect 19043 -17214 19245 -17158
rect 19043 -17248 19075 -17214
rect 19109 -17248 19176 -17214
rect 19210 -17248 19245 -17214
rect 19043 -17304 19245 -17248
rect 19043 -17338 19075 -17304
rect 19109 -17338 19176 -17304
rect 19210 -17338 19245 -17304
rect 19043 -17394 19245 -17338
rect 19043 -17428 19075 -17394
rect 19109 -17428 19176 -17394
rect 19210 -17428 19245 -17394
rect 19043 -17484 19245 -17428
rect 19043 -17518 19075 -17484
rect 19109 -17518 19176 -17484
rect 19210 -17518 19245 -17484
rect 19043 -17574 19245 -17518
rect 17755 -17641 17957 -17608
rect 19043 -17608 19075 -17574
rect 19109 -17608 19176 -17574
rect 19210 -17608 19245 -17574
rect 20331 -16618 20363 -16584
rect 20397 -16618 20464 -16584
rect 20498 -16618 20533 -16584
rect 21619 -16584 21821 -16555
rect 20331 -16674 20533 -16618
rect 20331 -16708 20363 -16674
rect 20397 -16708 20464 -16674
rect 20498 -16708 20533 -16674
rect 20331 -16764 20533 -16708
rect 20331 -16798 20363 -16764
rect 20397 -16798 20464 -16764
rect 20498 -16798 20533 -16764
rect 20331 -16854 20533 -16798
rect 20331 -16888 20363 -16854
rect 20397 -16888 20464 -16854
rect 20498 -16888 20533 -16854
rect 20331 -16944 20533 -16888
rect 20331 -16978 20363 -16944
rect 20397 -16978 20464 -16944
rect 20498 -16978 20533 -16944
rect 20331 -17034 20533 -16978
rect 20331 -17068 20363 -17034
rect 20397 -17068 20464 -17034
rect 20498 -17068 20533 -17034
rect 20331 -17124 20533 -17068
rect 20331 -17158 20363 -17124
rect 20397 -17158 20464 -17124
rect 20498 -17158 20533 -17124
rect 20331 -17214 20533 -17158
rect 20331 -17248 20363 -17214
rect 20397 -17248 20464 -17214
rect 20498 -17248 20533 -17214
rect 20331 -17304 20533 -17248
rect 20331 -17338 20363 -17304
rect 20397 -17338 20464 -17304
rect 20498 -17338 20533 -17304
rect 20331 -17394 20533 -17338
rect 20331 -17428 20363 -17394
rect 20397 -17428 20464 -17394
rect 20498 -17428 20533 -17394
rect 20331 -17484 20533 -17428
rect 20331 -17518 20363 -17484
rect 20397 -17518 20464 -17484
rect 20498 -17518 20533 -17484
rect 20331 -17574 20533 -17518
rect 19043 -17641 19245 -17608
rect 20331 -17608 20363 -17574
rect 20397 -17608 20464 -17574
rect 20498 -17608 20533 -17574
rect 21619 -16618 21651 -16584
rect 21685 -16618 21752 -16584
rect 21786 -16618 21821 -16584
rect 22907 -16584 23109 -16555
rect 21619 -16674 21821 -16618
rect 21619 -16708 21651 -16674
rect 21685 -16708 21752 -16674
rect 21786 -16708 21821 -16674
rect 21619 -16764 21821 -16708
rect 21619 -16798 21651 -16764
rect 21685 -16798 21752 -16764
rect 21786 -16798 21821 -16764
rect 21619 -16854 21821 -16798
rect 21619 -16888 21651 -16854
rect 21685 -16888 21752 -16854
rect 21786 -16888 21821 -16854
rect 21619 -16944 21821 -16888
rect 21619 -16978 21651 -16944
rect 21685 -16978 21752 -16944
rect 21786 -16978 21821 -16944
rect 21619 -17034 21821 -16978
rect 21619 -17068 21651 -17034
rect 21685 -17068 21752 -17034
rect 21786 -17068 21821 -17034
rect 21619 -17124 21821 -17068
rect 21619 -17158 21651 -17124
rect 21685 -17158 21752 -17124
rect 21786 -17158 21821 -17124
rect 21619 -17214 21821 -17158
rect 21619 -17248 21651 -17214
rect 21685 -17248 21752 -17214
rect 21786 -17248 21821 -17214
rect 21619 -17304 21821 -17248
rect 21619 -17338 21651 -17304
rect 21685 -17338 21752 -17304
rect 21786 -17338 21821 -17304
rect 21619 -17394 21821 -17338
rect 21619 -17428 21651 -17394
rect 21685 -17428 21752 -17394
rect 21786 -17428 21821 -17394
rect 21619 -17484 21821 -17428
rect 21619 -17518 21651 -17484
rect 21685 -17518 21752 -17484
rect 21786 -17518 21821 -17484
rect 21619 -17574 21821 -17518
rect 20331 -17641 20533 -17608
rect 21619 -17608 21651 -17574
rect 21685 -17608 21752 -17574
rect 21786 -17608 21821 -17574
rect 22907 -16618 22939 -16584
rect 22973 -16618 23040 -16584
rect 23074 -16618 23109 -16584
rect 24195 -16584 24397 -16555
rect 22907 -16674 23109 -16618
rect 22907 -16708 22939 -16674
rect 22973 -16708 23040 -16674
rect 23074 -16708 23109 -16674
rect 22907 -16764 23109 -16708
rect 22907 -16798 22939 -16764
rect 22973 -16798 23040 -16764
rect 23074 -16798 23109 -16764
rect 22907 -16854 23109 -16798
rect 22907 -16888 22939 -16854
rect 22973 -16888 23040 -16854
rect 23074 -16888 23109 -16854
rect 22907 -16944 23109 -16888
rect 22907 -16978 22939 -16944
rect 22973 -16978 23040 -16944
rect 23074 -16978 23109 -16944
rect 22907 -17034 23109 -16978
rect 22907 -17068 22939 -17034
rect 22973 -17068 23040 -17034
rect 23074 -17068 23109 -17034
rect 22907 -17124 23109 -17068
rect 22907 -17158 22939 -17124
rect 22973 -17158 23040 -17124
rect 23074 -17158 23109 -17124
rect 22907 -17214 23109 -17158
rect 22907 -17248 22939 -17214
rect 22973 -17248 23040 -17214
rect 23074 -17248 23109 -17214
rect 22907 -17304 23109 -17248
rect 22907 -17338 22939 -17304
rect 22973 -17338 23040 -17304
rect 23074 -17338 23109 -17304
rect 22907 -17394 23109 -17338
rect 22907 -17428 22939 -17394
rect 22973 -17428 23040 -17394
rect 23074 -17428 23109 -17394
rect 22907 -17484 23109 -17428
rect 22907 -17518 22939 -17484
rect 22973 -17518 23040 -17484
rect 23074 -17518 23109 -17484
rect 22907 -17574 23109 -17518
rect 21619 -17641 21821 -17608
rect 22907 -17608 22939 -17574
rect 22973 -17608 23040 -17574
rect 23074 -17608 23109 -17574
rect 24195 -16618 24227 -16584
rect 24261 -16618 24328 -16584
rect 24362 -16618 24397 -16584
rect 25483 -16584 25685 -16555
rect 24195 -16674 24397 -16618
rect 24195 -16708 24227 -16674
rect 24261 -16708 24328 -16674
rect 24362 -16708 24397 -16674
rect 24195 -16764 24397 -16708
rect 24195 -16798 24227 -16764
rect 24261 -16798 24328 -16764
rect 24362 -16798 24397 -16764
rect 24195 -16854 24397 -16798
rect 24195 -16888 24227 -16854
rect 24261 -16888 24328 -16854
rect 24362 -16888 24397 -16854
rect 24195 -16944 24397 -16888
rect 24195 -16978 24227 -16944
rect 24261 -16978 24328 -16944
rect 24362 -16978 24397 -16944
rect 24195 -17034 24397 -16978
rect 24195 -17068 24227 -17034
rect 24261 -17068 24328 -17034
rect 24362 -17068 24397 -17034
rect 24195 -17124 24397 -17068
rect 24195 -17158 24227 -17124
rect 24261 -17158 24328 -17124
rect 24362 -17158 24397 -17124
rect 24195 -17214 24397 -17158
rect 24195 -17248 24227 -17214
rect 24261 -17248 24328 -17214
rect 24362 -17248 24397 -17214
rect 24195 -17304 24397 -17248
rect 24195 -17338 24227 -17304
rect 24261 -17338 24328 -17304
rect 24362 -17338 24397 -17304
rect 24195 -17394 24397 -17338
rect 24195 -17428 24227 -17394
rect 24261 -17428 24328 -17394
rect 24362 -17428 24397 -17394
rect 24195 -17484 24397 -17428
rect 24195 -17518 24227 -17484
rect 24261 -17518 24328 -17484
rect 24362 -17518 24397 -17484
rect 24195 -17574 24397 -17518
rect 22907 -17641 23109 -17608
rect 24195 -17608 24227 -17574
rect 24261 -17608 24328 -17574
rect 24362 -17608 24397 -17574
rect 25483 -16618 25515 -16584
rect 25549 -16618 25616 -16584
rect 25650 -16618 25685 -16584
rect 26771 -16584 26872 -16555
rect 25483 -16674 25685 -16618
rect 25483 -16708 25515 -16674
rect 25549 -16708 25616 -16674
rect 25650 -16708 25685 -16674
rect 25483 -16764 25685 -16708
rect 25483 -16798 25515 -16764
rect 25549 -16798 25616 -16764
rect 25650 -16798 25685 -16764
rect 25483 -16854 25685 -16798
rect 25483 -16888 25515 -16854
rect 25549 -16888 25616 -16854
rect 25650 -16888 25685 -16854
rect 25483 -16944 25685 -16888
rect 25483 -16978 25515 -16944
rect 25549 -16978 25616 -16944
rect 25650 -16978 25685 -16944
rect 25483 -17034 25685 -16978
rect 25483 -17068 25515 -17034
rect 25549 -17068 25616 -17034
rect 25650 -17068 25685 -17034
rect 25483 -17124 25685 -17068
rect 25483 -17158 25515 -17124
rect 25549 -17158 25616 -17124
rect 25650 -17158 25685 -17124
rect 25483 -17214 25685 -17158
rect 25483 -17248 25515 -17214
rect 25549 -17248 25616 -17214
rect 25650 -17248 25685 -17214
rect 25483 -17304 25685 -17248
rect 25483 -17338 25515 -17304
rect 25549 -17338 25616 -17304
rect 25650 -17338 25685 -17304
rect 25483 -17394 25685 -17338
rect 25483 -17428 25515 -17394
rect 25549 -17428 25616 -17394
rect 25650 -17428 25685 -17394
rect 25483 -17484 25685 -17428
rect 25483 -17518 25515 -17484
rect 25549 -17518 25616 -17484
rect 25650 -17518 25685 -17484
rect 25483 -17574 25685 -17518
rect 24195 -17641 24397 -17608
rect 25483 -17608 25515 -17574
rect 25549 -17608 25616 -17574
rect 25650 -17608 25685 -17574
rect 26771 -16618 26803 -16584
rect 26837 -16618 26872 -16584
rect 26771 -16674 26872 -16618
rect 26771 -16708 26803 -16674
rect 26837 -16708 26872 -16674
rect 26771 -16764 26872 -16708
rect 26771 -16798 26803 -16764
rect 26837 -16798 26872 -16764
rect 26771 -16854 26872 -16798
rect 26771 -16888 26803 -16854
rect 26837 -16888 26872 -16854
rect 26771 -16944 26872 -16888
rect 26771 -16978 26803 -16944
rect 26837 -16978 26872 -16944
rect 26771 -17034 26872 -16978
rect 26771 -17068 26803 -17034
rect 26837 -17068 26872 -17034
rect 26771 -17124 26872 -17068
rect 26771 -17158 26803 -17124
rect 26837 -17158 26872 -17124
rect 26771 -17214 26872 -17158
rect 26771 -17248 26803 -17214
rect 26837 -17248 26872 -17214
rect 26771 -17304 26872 -17248
rect 26771 -17338 26803 -17304
rect 26837 -17338 26872 -17304
rect 26771 -17394 26872 -17338
rect 26771 -17428 26803 -17394
rect 26837 -17428 26872 -17394
rect 26771 -17484 26872 -17428
rect 26771 -17518 26803 -17484
rect 26837 -17518 26872 -17484
rect 26771 -17574 26872 -17518
rect 25483 -17641 25685 -17608
rect 26771 -17608 26803 -17574
rect 26837 -17608 26872 -17574
rect 26771 -17641 26872 -17608
rect 16568 -17675 26872 -17641
rect 16568 -17709 16684 -17675
rect 16718 -17709 16774 -17675
rect 16808 -17709 16864 -17675
rect 16898 -17709 16954 -17675
rect 16988 -17709 17044 -17675
rect 17078 -17709 17134 -17675
rect 17168 -17709 17224 -17675
rect 17258 -17709 17314 -17675
rect 17348 -17709 17404 -17675
rect 17438 -17709 17494 -17675
rect 17528 -17709 17584 -17675
rect 17618 -17709 17674 -17675
rect 17708 -17709 17764 -17675
rect 17798 -17709 17972 -17675
rect 18006 -17709 18062 -17675
rect 18096 -17709 18152 -17675
rect 18186 -17709 18242 -17675
rect 18276 -17709 18332 -17675
rect 18366 -17709 18422 -17675
rect 18456 -17709 18512 -17675
rect 18546 -17709 18602 -17675
rect 18636 -17709 18692 -17675
rect 18726 -17709 18782 -17675
rect 18816 -17709 18872 -17675
rect 18906 -17709 18962 -17675
rect 18996 -17709 19052 -17675
rect 19086 -17709 19260 -17675
rect 19294 -17709 19350 -17675
rect 19384 -17709 19440 -17675
rect 19474 -17709 19530 -17675
rect 19564 -17709 19620 -17675
rect 19654 -17709 19710 -17675
rect 19744 -17709 19800 -17675
rect 19834 -17709 19890 -17675
rect 19924 -17709 19980 -17675
rect 20014 -17709 20070 -17675
rect 20104 -17709 20160 -17675
rect 20194 -17709 20250 -17675
rect 20284 -17709 20340 -17675
rect 20374 -17709 20548 -17675
rect 20582 -17709 20638 -17675
rect 20672 -17709 20728 -17675
rect 20762 -17709 20818 -17675
rect 20852 -17709 20908 -17675
rect 20942 -17709 20998 -17675
rect 21032 -17709 21088 -17675
rect 21122 -17709 21178 -17675
rect 21212 -17709 21268 -17675
rect 21302 -17709 21358 -17675
rect 21392 -17709 21448 -17675
rect 21482 -17709 21538 -17675
rect 21572 -17709 21628 -17675
rect 21662 -17709 21836 -17675
rect 21870 -17709 21926 -17675
rect 21960 -17709 22016 -17675
rect 22050 -17709 22106 -17675
rect 22140 -17709 22196 -17675
rect 22230 -17709 22286 -17675
rect 22320 -17709 22376 -17675
rect 22410 -17709 22466 -17675
rect 22500 -17709 22556 -17675
rect 22590 -17709 22646 -17675
rect 22680 -17709 22736 -17675
rect 22770 -17709 22826 -17675
rect 22860 -17709 22916 -17675
rect 22950 -17709 23124 -17675
rect 23158 -17709 23214 -17675
rect 23248 -17709 23304 -17675
rect 23338 -17709 23394 -17675
rect 23428 -17709 23484 -17675
rect 23518 -17709 23574 -17675
rect 23608 -17709 23664 -17675
rect 23698 -17709 23754 -17675
rect 23788 -17709 23844 -17675
rect 23878 -17709 23934 -17675
rect 23968 -17709 24024 -17675
rect 24058 -17709 24114 -17675
rect 24148 -17709 24204 -17675
rect 24238 -17709 24412 -17675
rect 24446 -17709 24502 -17675
rect 24536 -17709 24592 -17675
rect 24626 -17709 24682 -17675
rect 24716 -17709 24772 -17675
rect 24806 -17709 24862 -17675
rect 24896 -17709 24952 -17675
rect 24986 -17709 25042 -17675
rect 25076 -17709 25132 -17675
rect 25166 -17709 25222 -17675
rect 25256 -17709 25312 -17675
rect 25346 -17709 25402 -17675
rect 25436 -17709 25492 -17675
rect 25526 -17709 25700 -17675
rect 25734 -17709 25790 -17675
rect 25824 -17709 25880 -17675
rect 25914 -17709 25970 -17675
rect 26004 -17709 26060 -17675
rect 26094 -17709 26150 -17675
rect 26184 -17709 26240 -17675
rect 26274 -17709 26330 -17675
rect 26364 -17709 26420 -17675
rect 26454 -17709 26510 -17675
rect 26544 -17709 26600 -17675
rect 26634 -17709 26690 -17675
rect 26724 -17709 26780 -17675
rect 26814 -17709 26872 -17675
rect 16568 -17742 26872 -17709
rect 7278 -31168 13630 -31144
rect 7278 -31738 7302 -31168
rect 13606 -31738 13630 -31168
rect 7278 -31762 13630 -31738
rect 7278 -36128 13630 -36104
rect 7278 -36698 7302 -36128
rect 13606 -36698 13630 -36128
rect 7278 -36722 13630 -36698
rect 7278 -39372 13630 -39348
rect 7278 -39942 7302 -39372
rect 13606 -39942 13630 -39372
rect 7278 -39966 13630 -39942
<< nsubdiff >>
rect 16731 -11484 17693 -11465
rect 16731 -11518 16863 -11484
rect 16897 -11518 16953 -11484
rect 16987 -11518 17043 -11484
rect 17077 -11518 17133 -11484
rect 17167 -11518 17223 -11484
rect 17257 -11518 17313 -11484
rect 17347 -11518 17403 -11484
rect 17437 -11518 17493 -11484
rect 17527 -11518 17583 -11484
rect 17617 -11518 17693 -11484
rect 16731 -11537 17693 -11518
rect 16731 -11562 16803 -11537
rect 16731 -11596 16750 -11562
rect 16784 -11596 16803 -11562
rect 16731 -11652 16803 -11596
rect 17621 -11596 17693 -11537
rect 16731 -11686 16750 -11652
rect 16784 -11686 16803 -11652
rect 16731 -11742 16803 -11686
rect 16731 -11776 16750 -11742
rect 16784 -11776 16803 -11742
rect 16731 -11832 16803 -11776
rect 16731 -11866 16750 -11832
rect 16784 -11866 16803 -11832
rect 16731 -11922 16803 -11866
rect 16731 -11956 16750 -11922
rect 16784 -11956 16803 -11922
rect 16731 -12012 16803 -11956
rect 16731 -12046 16750 -12012
rect 16784 -12046 16803 -12012
rect 16731 -12102 16803 -12046
rect 16731 -12136 16750 -12102
rect 16784 -12136 16803 -12102
rect 16731 -12192 16803 -12136
rect 16731 -12226 16750 -12192
rect 16784 -12226 16803 -12192
rect 16731 -12282 16803 -12226
rect 16731 -12316 16750 -12282
rect 16784 -12316 16803 -12282
rect 17621 -11630 17640 -11596
rect 17674 -11630 17693 -11596
rect 17621 -11686 17693 -11630
rect 17621 -11720 17640 -11686
rect 17674 -11720 17693 -11686
rect 17621 -11776 17693 -11720
rect 17621 -11810 17640 -11776
rect 17674 -11810 17693 -11776
rect 17621 -11866 17693 -11810
rect 17621 -11900 17640 -11866
rect 17674 -11900 17693 -11866
rect 17621 -11956 17693 -11900
rect 17621 -11990 17640 -11956
rect 17674 -11990 17693 -11956
rect 17621 -12046 17693 -11990
rect 17621 -12080 17640 -12046
rect 17674 -12080 17693 -12046
rect 17621 -12136 17693 -12080
rect 17621 -12170 17640 -12136
rect 17674 -12170 17693 -12136
rect 17621 -12226 17693 -12170
rect 17621 -12260 17640 -12226
rect 17674 -12260 17693 -12226
rect 16731 -12355 16803 -12316
rect 17621 -12316 17693 -12260
rect 17621 -12350 17640 -12316
rect 17674 -12350 17693 -12316
rect 17621 -12355 17693 -12350
rect 16731 -12374 17693 -12355
rect 16731 -12408 16844 -12374
rect 16878 -12408 16934 -12374
rect 16968 -12408 17024 -12374
rect 17058 -12408 17114 -12374
rect 17148 -12408 17204 -12374
rect 17238 -12408 17294 -12374
rect 17328 -12408 17384 -12374
rect 17418 -12408 17474 -12374
rect 17508 -12408 17564 -12374
rect 17598 -12408 17693 -12374
rect 16731 -12427 17693 -12408
rect 18019 -11484 18981 -11465
rect 18019 -11518 18151 -11484
rect 18185 -11518 18241 -11484
rect 18275 -11518 18331 -11484
rect 18365 -11518 18421 -11484
rect 18455 -11518 18511 -11484
rect 18545 -11518 18601 -11484
rect 18635 -11518 18691 -11484
rect 18725 -11518 18781 -11484
rect 18815 -11518 18871 -11484
rect 18905 -11518 18981 -11484
rect 18019 -11537 18981 -11518
rect 18019 -11562 18091 -11537
rect 18019 -11596 18038 -11562
rect 18072 -11596 18091 -11562
rect 18019 -11652 18091 -11596
rect 18909 -11596 18981 -11537
rect 18019 -11686 18038 -11652
rect 18072 -11686 18091 -11652
rect 18019 -11742 18091 -11686
rect 18019 -11776 18038 -11742
rect 18072 -11776 18091 -11742
rect 18019 -11832 18091 -11776
rect 18019 -11866 18038 -11832
rect 18072 -11866 18091 -11832
rect 18019 -11922 18091 -11866
rect 18019 -11956 18038 -11922
rect 18072 -11956 18091 -11922
rect 18019 -12012 18091 -11956
rect 18019 -12046 18038 -12012
rect 18072 -12046 18091 -12012
rect 18019 -12102 18091 -12046
rect 18019 -12136 18038 -12102
rect 18072 -12136 18091 -12102
rect 18019 -12192 18091 -12136
rect 18019 -12226 18038 -12192
rect 18072 -12226 18091 -12192
rect 18019 -12282 18091 -12226
rect 18019 -12316 18038 -12282
rect 18072 -12316 18091 -12282
rect 18909 -11630 18928 -11596
rect 18962 -11630 18981 -11596
rect 18909 -11686 18981 -11630
rect 18909 -11720 18928 -11686
rect 18962 -11720 18981 -11686
rect 18909 -11776 18981 -11720
rect 18909 -11810 18928 -11776
rect 18962 -11810 18981 -11776
rect 18909 -11866 18981 -11810
rect 18909 -11900 18928 -11866
rect 18962 -11900 18981 -11866
rect 18909 -11956 18981 -11900
rect 18909 -11990 18928 -11956
rect 18962 -11990 18981 -11956
rect 18909 -12046 18981 -11990
rect 18909 -12080 18928 -12046
rect 18962 -12080 18981 -12046
rect 18909 -12136 18981 -12080
rect 18909 -12170 18928 -12136
rect 18962 -12170 18981 -12136
rect 18909 -12226 18981 -12170
rect 18909 -12260 18928 -12226
rect 18962 -12260 18981 -12226
rect 18019 -12355 18091 -12316
rect 18909 -12316 18981 -12260
rect 18909 -12350 18928 -12316
rect 18962 -12350 18981 -12316
rect 18909 -12355 18981 -12350
rect 18019 -12374 18981 -12355
rect 18019 -12408 18132 -12374
rect 18166 -12408 18222 -12374
rect 18256 -12408 18312 -12374
rect 18346 -12408 18402 -12374
rect 18436 -12408 18492 -12374
rect 18526 -12408 18582 -12374
rect 18616 -12408 18672 -12374
rect 18706 -12408 18762 -12374
rect 18796 -12408 18852 -12374
rect 18886 -12408 18981 -12374
rect 18019 -12427 18981 -12408
rect 19307 -11484 20269 -11465
rect 19307 -11518 19439 -11484
rect 19473 -11518 19529 -11484
rect 19563 -11518 19619 -11484
rect 19653 -11518 19709 -11484
rect 19743 -11518 19799 -11484
rect 19833 -11518 19889 -11484
rect 19923 -11518 19979 -11484
rect 20013 -11518 20069 -11484
rect 20103 -11518 20159 -11484
rect 20193 -11518 20269 -11484
rect 19307 -11537 20269 -11518
rect 19307 -11562 19379 -11537
rect 19307 -11596 19326 -11562
rect 19360 -11596 19379 -11562
rect 19307 -11652 19379 -11596
rect 20197 -11596 20269 -11537
rect 19307 -11686 19326 -11652
rect 19360 -11686 19379 -11652
rect 19307 -11742 19379 -11686
rect 19307 -11776 19326 -11742
rect 19360 -11776 19379 -11742
rect 19307 -11832 19379 -11776
rect 19307 -11866 19326 -11832
rect 19360 -11866 19379 -11832
rect 19307 -11922 19379 -11866
rect 19307 -11956 19326 -11922
rect 19360 -11956 19379 -11922
rect 19307 -12012 19379 -11956
rect 19307 -12046 19326 -12012
rect 19360 -12046 19379 -12012
rect 19307 -12102 19379 -12046
rect 19307 -12136 19326 -12102
rect 19360 -12136 19379 -12102
rect 19307 -12192 19379 -12136
rect 19307 -12226 19326 -12192
rect 19360 -12226 19379 -12192
rect 19307 -12282 19379 -12226
rect 19307 -12316 19326 -12282
rect 19360 -12316 19379 -12282
rect 20197 -11630 20216 -11596
rect 20250 -11630 20269 -11596
rect 20197 -11686 20269 -11630
rect 20197 -11720 20216 -11686
rect 20250 -11720 20269 -11686
rect 20197 -11776 20269 -11720
rect 20197 -11810 20216 -11776
rect 20250 -11810 20269 -11776
rect 20197 -11866 20269 -11810
rect 20197 -11900 20216 -11866
rect 20250 -11900 20269 -11866
rect 20197 -11956 20269 -11900
rect 20197 -11990 20216 -11956
rect 20250 -11990 20269 -11956
rect 20197 -12046 20269 -11990
rect 20197 -12080 20216 -12046
rect 20250 -12080 20269 -12046
rect 20197 -12136 20269 -12080
rect 20197 -12170 20216 -12136
rect 20250 -12170 20269 -12136
rect 20197 -12226 20269 -12170
rect 20197 -12260 20216 -12226
rect 20250 -12260 20269 -12226
rect 19307 -12355 19379 -12316
rect 20197 -12316 20269 -12260
rect 20197 -12350 20216 -12316
rect 20250 -12350 20269 -12316
rect 20197 -12355 20269 -12350
rect 19307 -12374 20269 -12355
rect 19307 -12408 19420 -12374
rect 19454 -12408 19510 -12374
rect 19544 -12408 19600 -12374
rect 19634 -12408 19690 -12374
rect 19724 -12408 19780 -12374
rect 19814 -12408 19870 -12374
rect 19904 -12408 19960 -12374
rect 19994 -12408 20050 -12374
rect 20084 -12408 20140 -12374
rect 20174 -12408 20269 -12374
rect 19307 -12427 20269 -12408
rect 20595 -11484 21557 -11465
rect 20595 -11518 20727 -11484
rect 20761 -11518 20817 -11484
rect 20851 -11518 20907 -11484
rect 20941 -11518 20997 -11484
rect 21031 -11518 21087 -11484
rect 21121 -11518 21177 -11484
rect 21211 -11518 21267 -11484
rect 21301 -11518 21357 -11484
rect 21391 -11518 21447 -11484
rect 21481 -11518 21557 -11484
rect 20595 -11537 21557 -11518
rect 20595 -11562 20667 -11537
rect 20595 -11596 20614 -11562
rect 20648 -11596 20667 -11562
rect 20595 -11652 20667 -11596
rect 21485 -11596 21557 -11537
rect 20595 -11686 20614 -11652
rect 20648 -11686 20667 -11652
rect 20595 -11742 20667 -11686
rect 20595 -11776 20614 -11742
rect 20648 -11776 20667 -11742
rect 20595 -11832 20667 -11776
rect 20595 -11866 20614 -11832
rect 20648 -11866 20667 -11832
rect 20595 -11922 20667 -11866
rect 20595 -11956 20614 -11922
rect 20648 -11956 20667 -11922
rect 20595 -12012 20667 -11956
rect 20595 -12046 20614 -12012
rect 20648 -12046 20667 -12012
rect 20595 -12102 20667 -12046
rect 20595 -12136 20614 -12102
rect 20648 -12136 20667 -12102
rect 20595 -12192 20667 -12136
rect 20595 -12226 20614 -12192
rect 20648 -12226 20667 -12192
rect 20595 -12282 20667 -12226
rect 20595 -12316 20614 -12282
rect 20648 -12316 20667 -12282
rect 21485 -11630 21504 -11596
rect 21538 -11630 21557 -11596
rect 21485 -11686 21557 -11630
rect 21485 -11720 21504 -11686
rect 21538 -11720 21557 -11686
rect 21485 -11776 21557 -11720
rect 21485 -11810 21504 -11776
rect 21538 -11810 21557 -11776
rect 21485 -11866 21557 -11810
rect 21485 -11900 21504 -11866
rect 21538 -11900 21557 -11866
rect 21485 -11956 21557 -11900
rect 21485 -11990 21504 -11956
rect 21538 -11990 21557 -11956
rect 21485 -12046 21557 -11990
rect 21485 -12080 21504 -12046
rect 21538 -12080 21557 -12046
rect 21485 -12136 21557 -12080
rect 21485 -12170 21504 -12136
rect 21538 -12170 21557 -12136
rect 21485 -12226 21557 -12170
rect 21485 -12260 21504 -12226
rect 21538 -12260 21557 -12226
rect 20595 -12355 20667 -12316
rect 21485 -12316 21557 -12260
rect 21485 -12350 21504 -12316
rect 21538 -12350 21557 -12316
rect 21485 -12355 21557 -12350
rect 20595 -12374 21557 -12355
rect 20595 -12408 20708 -12374
rect 20742 -12408 20798 -12374
rect 20832 -12408 20888 -12374
rect 20922 -12408 20978 -12374
rect 21012 -12408 21068 -12374
rect 21102 -12408 21158 -12374
rect 21192 -12408 21248 -12374
rect 21282 -12408 21338 -12374
rect 21372 -12408 21428 -12374
rect 21462 -12408 21557 -12374
rect 20595 -12427 21557 -12408
rect 21883 -11484 22845 -11465
rect 21883 -11518 22015 -11484
rect 22049 -11518 22105 -11484
rect 22139 -11518 22195 -11484
rect 22229 -11518 22285 -11484
rect 22319 -11518 22375 -11484
rect 22409 -11518 22465 -11484
rect 22499 -11518 22555 -11484
rect 22589 -11518 22645 -11484
rect 22679 -11518 22735 -11484
rect 22769 -11518 22845 -11484
rect 21883 -11537 22845 -11518
rect 21883 -11562 21955 -11537
rect 21883 -11596 21902 -11562
rect 21936 -11596 21955 -11562
rect 21883 -11652 21955 -11596
rect 22773 -11596 22845 -11537
rect 21883 -11686 21902 -11652
rect 21936 -11686 21955 -11652
rect 21883 -11742 21955 -11686
rect 21883 -11776 21902 -11742
rect 21936 -11776 21955 -11742
rect 21883 -11832 21955 -11776
rect 21883 -11866 21902 -11832
rect 21936 -11866 21955 -11832
rect 21883 -11922 21955 -11866
rect 21883 -11956 21902 -11922
rect 21936 -11956 21955 -11922
rect 21883 -12012 21955 -11956
rect 21883 -12046 21902 -12012
rect 21936 -12046 21955 -12012
rect 21883 -12102 21955 -12046
rect 21883 -12136 21902 -12102
rect 21936 -12136 21955 -12102
rect 21883 -12192 21955 -12136
rect 21883 -12226 21902 -12192
rect 21936 -12226 21955 -12192
rect 21883 -12282 21955 -12226
rect 21883 -12316 21902 -12282
rect 21936 -12316 21955 -12282
rect 22773 -11630 22792 -11596
rect 22826 -11630 22845 -11596
rect 22773 -11686 22845 -11630
rect 22773 -11720 22792 -11686
rect 22826 -11720 22845 -11686
rect 22773 -11776 22845 -11720
rect 22773 -11810 22792 -11776
rect 22826 -11810 22845 -11776
rect 22773 -11866 22845 -11810
rect 22773 -11900 22792 -11866
rect 22826 -11900 22845 -11866
rect 22773 -11956 22845 -11900
rect 22773 -11990 22792 -11956
rect 22826 -11990 22845 -11956
rect 22773 -12046 22845 -11990
rect 22773 -12080 22792 -12046
rect 22826 -12080 22845 -12046
rect 22773 -12136 22845 -12080
rect 22773 -12170 22792 -12136
rect 22826 -12170 22845 -12136
rect 22773 -12226 22845 -12170
rect 22773 -12260 22792 -12226
rect 22826 -12260 22845 -12226
rect 21883 -12355 21955 -12316
rect 22773 -12316 22845 -12260
rect 22773 -12350 22792 -12316
rect 22826 -12350 22845 -12316
rect 22773 -12355 22845 -12350
rect 21883 -12374 22845 -12355
rect 21883 -12408 21996 -12374
rect 22030 -12408 22086 -12374
rect 22120 -12408 22176 -12374
rect 22210 -12408 22266 -12374
rect 22300 -12408 22356 -12374
rect 22390 -12408 22446 -12374
rect 22480 -12408 22536 -12374
rect 22570 -12408 22626 -12374
rect 22660 -12408 22716 -12374
rect 22750 -12408 22845 -12374
rect 21883 -12427 22845 -12408
rect 23171 -11484 24133 -11465
rect 23171 -11518 23303 -11484
rect 23337 -11518 23393 -11484
rect 23427 -11518 23483 -11484
rect 23517 -11518 23573 -11484
rect 23607 -11518 23663 -11484
rect 23697 -11518 23753 -11484
rect 23787 -11518 23843 -11484
rect 23877 -11518 23933 -11484
rect 23967 -11518 24023 -11484
rect 24057 -11518 24133 -11484
rect 23171 -11537 24133 -11518
rect 23171 -11562 23243 -11537
rect 23171 -11596 23190 -11562
rect 23224 -11596 23243 -11562
rect 23171 -11652 23243 -11596
rect 24061 -11596 24133 -11537
rect 23171 -11686 23190 -11652
rect 23224 -11686 23243 -11652
rect 23171 -11742 23243 -11686
rect 23171 -11776 23190 -11742
rect 23224 -11776 23243 -11742
rect 23171 -11832 23243 -11776
rect 23171 -11866 23190 -11832
rect 23224 -11866 23243 -11832
rect 23171 -11922 23243 -11866
rect 23171 -11956 23190 -11922
rect 23224 -11956 23243 -11922
rect 23171 -12012 23243 -11956
rect 23171 -12046 23190 -12012
rect 23224 -12046 23243 -12012
rect 23171 -12102 23243 -12046
rect 23171 -12136 23190 -12102
rect 23224 -12136 23243 -12102
rect 23171 -12192 23243 -12136
rect 23171 -12226 23190 -12192
rect 23224 -12226 23243 -12192
rect 23171 -12282 23243 -12226
rect 23171 -12316 23190 -12282
rect 23224 -12316 23243 -12282
rect 24061 -11630 24080 -11596
rect 24114 -11630 24133 -11596
rect 24061 -11686 24133 -11630
rect 24061 -11720 24080 -11686
rect 24114 -11720 24133 -11686
rect 24061 -11776 24133 -11720
rect 24061 -11810 24080 -11776
rect 24114 -11810 24133 -11776
rect 24061 -11866 24133 -11810
rect 24061 -11900 24080 -11866
rect 24114 -11900 24133 -11866
rect 24061 -11956 24133 -11900
rect 24061 -11990 24080 -11956
rect 24114 -11990 24133 -11956
rect 24061 -12046 24133 -11990
rect 24061 -12080 24080 -12046
rect 24114 -12080 24133 -12046
rect 24061 -12136 24133 -12080
rect 24061 -12170 24080 -12136
rect 24114 -12170 24133 -12136
rect 24061 -12226 24133 -12170
rect 24061 -12260 24080 -12226
rect 24114 -12260 24133 -12226
rect 23171 -12355 23243 -12316
rect 24061 -12316 24133 -12260
rect 24061 -12350 24080 -12316
rect 24114 -12350 24133 -12316
rect 24061 -12355 24133 -12350
rect 23171 -12374 24133 -12355
rect 23171 -12408 23284 -12374
rect 23318 -12408 23374 -12374
rect 23408 -12408 23464 -12374
rect 23498 -12408 23554 -12374
rect 23588 -12408 23644 -12374
rect 23678 -12408 23734 -12374
rect 23768 -12408 23824 -12374
rect 23858 -12408 23914 -12374
rect 23948 -12408 24004 -12374
rect 24038 -12408 24133 -12374
rect 23171 -12427 24133 -12408
rect 24459 -11484 25421 -11465
rect 24459 -11518 24591 -11484
rect 24625 -11518 24681 -11484
rect 24715 -11518 24771 -11484
rect 24805 -11518 24861 -11484
rect 24895 -11518 24951 -11484
rect 24985 -11518 25041 -11484
rect 25075 -11518 25131 -11484
rect 25165 -11518 25221 -11484
rect 25255 -11518 25311 -11484
rect 25345 -11518 25421 -11484
rect 24459 -11537 25421 -11518
rect 24459 -11562 24531 -11537
rect 24459 -11596 24478 -11562
rect 24512 -11596 24531 -11562
rect 24459 -11652 24531 -11596
rect 25349 -11596 25421 -11537
rect 24459 -11686 24478 -11652
rect 24512 -11686 24531 -11652
rect 24459 -11742 24531 -11686
rect 24459 -11776 24478 -11742
rect 24512 -11776 24531 -11742
rect 24459 -11832 24531 -11776
rect 24459 -11866 24478 -11832
rect 24512 -11866 24531 -11832
rect 24459 -11922 24531 -11866
rect 24459 -11956 24478 -11922
rect 24512 -11956 24531 -11922
rect 24459 -12012 24531 -11956
rect 24459 -12046 24478 -12012
rect 24512 -12046 24531 -12012
rect 24459 -12102 24531 -12046
rect 24459 -12136 24478 -12102
rect 24512 -12136 24531 -12102
rect 24459 -12192 24531 -12136
rect 24459 -12226 24478 -12192
rect 24512 -12226 24531 -12192
rect 24459 -12282 24531 -12226
rect 24459 -12316 24478 -12282
rect 24512 -12316 24531 -12282
rect 25349 -11630 25368 -11596
rect 25402 -11630 25421 -11596
rect 25349 -11686 25421 -11630
rect 25349 -11720 25368 -11686
rect 25402 -11720 25421 -11686
rect 25349 -11776 25421 -11720
rect 25349 -11810 25368 -11776
rect 25402 -11810 25421 -11776
rect 25349 -11866 25421 -11810
rect 25349 -11900 25368 -11866
rect 25402 -11900 25421 -11866
rect 25349 -11956 25421 -11900
rect 25349 -11990 25368 -11956
rect 25402 -11990 25421 -11956
rect 25349 -12046 25421 -11990
rect 25349 -12080 25368 -12046
rect 25402 -12080 25421 -12046
rect 25349 -12136 25421 -12080
rect 25349 -12170 25368 -12136
rect 25402 -12170 25421 -12136
rect 25349 -12226 25421 -12170
rect 25349 -12260 25368 -12226
rect 25402 -12260 25421 -12226
rect 24459 -12355 24531 -12316
rect 25349 -12316 25421 -12260
rect 25349 -12350 25368 -12316
rect 25402 -12350 25421 -12316
rect 25349 -12355 25421 -12350
rect 24459 -12374 25421 -12355
rect 24459 -12408 24572 -12374
rect 24606 -12408 24662 -12374
rect 24696 -12408 24752 -12374
rect 24786 -12408 24842 -12374
rect 24876 -12408 24932 -12374
rect 24966 -12408 25022 -12374
rect 25056 -12408 25112 -12374
rect 25146 -12408 25202 -12374
rect 25236 -12408 25292 -12374
rect 25326 -12408 25421 -12374
rect 24459 -12427 25421 -12408
rect 25747 -11484 26709 -11465
rect 25747 -11518 25879 -11484
rect 25913 -11518 25969 -11484
rect 26003 -11518 26059 -11484
rect 26093 -11518 26149 -11484
rect 26183 -11518 26239 -11484
rect 26273 -11518 26329 -11484
rect 26363 -11518 26419 -11484
rect 26453 -11518 26509 -11484
rect 26543 -11518 26599 -11484
rect 26633 -11518 26709 -11484
rect 25747 -11537 26709 -11518
rect 25747 -11562 25819 -11537
rect 25747 -11596 25766 -11562
rect 25800 -11596 25819 -11562
rect 25747 -11652 25819 -11596
rect 26637 -11596 26709 -11537
rect 25747 -11686 25766 -11652
rect 25800 -11686 25819 -11652
rect 25747 -11742 25819 -11686
rect 25747 -11776 25766 -11742
rect 25800 -11776 25819 -11742
rect 25747 -11832 25819 -11776
rect 25747 -11866 25766 -11832
rect 25800 -11866 25819 -11832
rect 25747 -11922 25819 -11866
rect 25747 -11956 25766 -11922
rect 25800 -11956 25819 -11922
rect 25747 -12012 25819 -11956
rect 25747 -12046 25766 -12012
rect 25800 -12046 25819 -12012
rect 25747 -12102 25819 -12046
rect 25747 -12136 25766 -12102
rect 25800 -12136 25819 -12102
rect 25747 -12192 25819 -12136
rect 25747 -12226 25766 -12192
rect 25800 -12226 25819 -12192
rect 25747 -12282 25819 -12226
rect 25747 -12316 25766 -12282
rect 25800 -12316 25819 -12282
rect 26637 -11630 26656 -11596
rect 26690 -11630 26709 -11596
rect 26637 -11686 26709 -11630
rect 26637 -11720 26656 -11686
rect 26690 -11720 26709 -11686
rect 26637 -11776 26709 -11720
rect 26637 -11810 26656 -11776
rect 26690 -11810 26709 -11776
rect 26637 -11866 26709 -11810
rect 26637 -11900 26656 -11866
rect 26690 -11900 26709 -11866
rect 26637 -11956 26709 -11900
rect 26637 -11990 26656 -11956
rect 26690 -11990 26709 -11956
rect 26637 -12046 26709 -11990
rect 26637 -12080 26656 -12046
rect 26690 -12080 26709 -12046
rect 26637 -12136 26709 -12080
rect 26637 -12170 26656 -12136
rect 26690 -12170 26709 -12136
rect 26637 -12226 26709 -12170
rect 26637 -12260 26656 -12226
rect 26690 -12260 26709 -12226
rect 25747 -12355 25819 -12316
rect 26637 -12316 26709 -12260
rect 26637 -12350 26656 -12316
rect 26690 -12350 26709 -12316
rect 26637 -12355 26709 -12350
rect 25747 -12374 26709 -12355
rect 25747 -12408 25860 -12374
rect 25894 -12408 25950 -12374
rect 25984 -12408 26040 -12374
rect 26074 -12408 26130 -12374
rect 26164 -12408 26220 -12374
rect 26254 -12408 26310 -12374
rect 26344 -12408 26400 -12374
rect 26434 -12408 26490 -12374
rect 26524 -12408 26580 -12374
rect 26614 -12408 26709 -12374
rect 25747 -12427 26709 -12408
rect 16731 -12772 17693 -12753
rect 16731 -12806 16863 -12772
rect 16897 -12806 16953 -12772
rect 16987 -12806 17043 -12772
rect 17077 -12806 17133 -12772
rect 17167 -12806 17223 -12772
rect 17257 -12806 17313 -12772
rect 17347 -12806 17403 -12772
rect 17437 -12806 17493 -12772
rect 17527 -12806 17583 -12772
rect 17617 -12806 17693 -12772
rect 16731 -12825 17693 -12806
rect 16731 -12850 16803 -12825
rect 16731 -12884 16750 -12850
rect 16784 -12884 16803 -12850
rect 16731 -12940 16803 -12884
rect 17621 -12884 17693 -12825
rect 16731 -12974 16750 -12940
rect 16784 -12974 16803 -12940
rect 16731 -13030 16803 -12974
rect 16731 -13064 16750 -13030
rect 16784 -13064 16803 -13030
rect 16731 -13120 16803 -13064
rect 16731 -13154 16750 -13120
rect 16784 -13154 16803 -13120
rect 16731 -13210 16803 -13154
rect 16731 -13244 16750 -13210
rect 16784 -13244 16803 -13210
rect 16731 -13300 16803 -13244
rect 16731 -13334 16750 -13300
rect 16784 -13334 16803 -13300
rect 16731 -13390 16803 -13334
rect 16731 -13424 16750 -13390
rect 16784 -13424 16803 -13390
rect 16731 -13480 16803 -13424
rect 16731 -13514 16750 -13480
rect 16784 -13514 16803 -13480
rect 16731 -13570 16803 -13514
rect 16731 -13604 16750 -13570
rect 16784 -13604 16803 -13570
rect 17621 -12918 17640 -12884
rect 17674 -12918 17693 -12884
rect 17621 -12974 17693 -12918
rect 17621 -13008 17640 -12974
rect 17674 -13008 17693 -12974
rect 17621 -13064 17693 -13008
rect 17621 -13098 17640 -13064
rect 17674 -13098 17693 -13064
rect 17621 -13154 17693 -13098
rect 17621 -13188 17640 -13154
rect 17674 -13188 17693 -13154
rect 17621 -13244 17693 -13188
rect 17621 -13278 17640 -13244
rect 17674 -13278 17693 -13244
rect 17621 -13334 17693 -13278
rect 17621 -13368 17640 -13334
rect 17674 -13368 17693 -13334
rect 17621 -13424 17693 -13368
rect 17621 -13458 17640 -13424
rect 17674 -13458 17693 -13424
rect 17621 -13514 17693 -13458
rect 17621 -13548 17640 -13514
rect 17674 -13548 17693 -13514
rect 16731 -13643 16803 -13604
rect 17621 -13604 17693 -13548
rect 17621 -13638 17640 -13604
rect 17674 -13638 17693 -13604
rect 17621 -13643 17693 -13638
rect 16731 -13662 17693 -13643
rect 16731 -13696 16844 -13662
rect 16878 -13696 16934 -13662
rect 16968 -13696 17024 -13662
rect 17058 -13696 17114 -13662
rect 17148 -13696 17204 -13662
rect 17238 -13696 17294 -13662
rect 17328 -13696 17384 -13662
rect 17418 -13696 17474 -13662
rect 17508 -13696 17564 -13662
rect 17598 -13696 17693 -13662
rect 16731 -13715 17693 -13696
rect 18019 -12772 18981 -12753
rect 18019 -12806 18151 -12772
rect 18185 -12806 18241 -12772
rect 18275 -12806 18331 -12772
rect 18365 -12806 18421 -12772
rect 18455 -12806 18511 -12772
rect 18545 -12806 18601 -12772
rect 18635 -12806 18691 -12772
rect 18725 -12806 18781 -12772
rect 18815 -12806 18871 -12772
rect 18905 -12806 18981 -12772
rect 18019 -12825 18981 -12806
rect 18019 -12850 18091 -12825
rect 18019 -12884 18038 -12850
rect 18072 -12884 18091 -12850
rect 18019 -12940 18091 -12884
rect 18909 -12884 18981 -12825
rect 18019 -12974 18038 -12940
rect 18072 -12974 18091 -12940
rect 18019 -13030 18091 -12974
rect 18019 -13064 18038 -13030
rect 18072 -13064 18091 -13030
rect 18019 -13120 18091 -13064
rect 18019 -13154 18038 -13120
rect 18072 -13154 18091 -13120
rect 18019 -13210 18091 -13154
rect 18019 -13244 18038 -13210
rect 18072 -13244 18091 -13210
rect 18019 -13300 18091 -13244
rect 18019 -13334 18038 -13300
rect 18072 -13334 18091 -13300
rect 18019 -13390 18091 -13334
rect 18019 -13424 18038 -13390
rect 18072 -13424 18091 -13390
rect 18019 -13480 18091 -13424
rect 18019 -13514 18038 -13480
rect 18072 -13514 18091 -13480
rect 18019 -13570 18091 -13514
rect 18019 -13604 18038 -13570
rect 18072 -13604 18091 -13570
rect 18909 -12918 18928 -12884
rect 18962 -12918 18981 -12884
rect 18909 -12974 18981 -12918
rect 18909 -13008 18928 -12974
rect 18962 -13008 18981 -12974
rect 18909 -13064 18981 -13008
rect 18909 -13098 18928 -13064
rect 18962 -13098 18981 -13064
rect 18909 -13154 18981 -13098
rect 18909 -13188 18928 -13154
rect 18962 -13188 18981 -13154
rect 18909 -13244 18981 -13188
rect 18909 -13278 18928 -13244
rect 18962 -13278 18981 -13244
rect 18909 -13334 18981 -13278
rect 18909 -13368 18928 -13334
rect 18962 -13368 18981 -13334
rect 18909 -13424 18981 -13368
rect 18909 -13458 18928 -13424
rect 18962 -13458 18981 -13424
rect 18909 -13514 18981 -13458
rect 18909 -13548 18928 -13514
rect 18962 -13548 18981 -13514
rect 18019 -13643 18091 -13604
rect 18909 -13604 18981 -13548
rect 18909 -13638 18928 -13604
rect 18962 -13638 18981 -13604
rect 18909 -13643 18981 -13638
rect 18019 -13662 18981 -13643
rect 18019 -13696 18132 -13662
rect 18166 -13696 18222 -13662
rect 18256 -13696 18312 -13662
rect 18346 -13696 18402 -13662
rect 18436 -13696 18492 -13662
rect 18526 -13696 18582 -13662
rect 18616 -13696 18672 -13662
rect 18706 -13696 18762 -13662
rect 18796 -13696 18852 -13662
rect 18886 -13696 18981 -13662
rect 18019 -13715 18981 -13696
rect 19307 -12772 20269 -12753
rect 19307 -12806 19439 -12772
rect 19473 -12806 19529 -12772
rect 19563 -12806 19619 -12772
rect 19653 -12806 19709 -12772
rect 19743 -12806 19799 -12772
rect 19833 -12806 19889 -12772
rect 19923 -12806 19979 -12772
rect 20013 -12806 20069 -12772
rect 20103 -12806 20159 -12772
rect 20193 -12806 20269 -12772
rect 19307 -12825 20269 -12806
rect 19307 -12850 19379 -12825
rect 19307 -12884 19326 -12850
rect 19360 -12884 19379 -12850
rect 19307 -12940 19379 -12884
rect 20197 -12884 20269 -12825
rect 19307 -12974 19326 -12940
rect 19360 -12974 19379 -12940
rect 19307 -13030 19379 -12974
rect 19307 -13064 19326 -13030
rect 19360 -13064 19379 -13030
rect 19307 -13120 19379 -13064
rect 19307 -13154 19326 -13120
rect 19360 -13154 19379 -13120
rect 19307 -13210 19379 -13154
rect 19307 -13244 19326 -13210
rect 19360 -13244 19379 -13210
rect 19307 -13300 19379 -13244
rect 19307 -13334 19326 -13300
rect 19360 -13334 19379 -13300
rect 19307 -13390 19379 -13334
rect 19307 -13424 19326 -13390
rect 19360 -13424 19379 -13390
rect 19307 -13480 19379 -13424
rect 19307 -13514 19326 -13480
rect 19360 -13514 19379 -13480
rect 19307 -13570 19379 -13514
rect 19307 -13604 19326 -13570
rect 19360 -13604 19379 -13570
rect 20197 -12918 20216 -12884
rect 20250 -12918 20269 -12884
rect 20197 -12974 20269 -12918
rect 20197 -13008 20216 -12974
rect 20250 -13008 20269 -12974
rect 20197 -13064 20269 -13008
rect 20197 -13098 20216 -13064
rect 20250 -13098 20269 -13064
rect 20197 -13154 20269 -13098
rect 20197 -13188 20216 -13154
rect 20250 -13188 20269 -13154
rect 20197 -13244 20269 -13188
rect 20197 -13278 20216 -13244
rect 20250 -13278 20269 -13244
rect 20197 -13334 20269 -13278
rect 20197 -13368 20216 -13334
rect 20250 -13368 20269 -13334
rect 20197 -13424 20269 -13368
rect 20197 -13458 20216 -13424
rect 20250 -13458 20269 -13424
rect 20197 -13514 20269 -13458
rect 20197 -13548 20216 -13514
rect 20250 -13548 20269 -13514
rect 19307 -13643 19379 -13604
rect 20197 -13604 20269 -13548
rect 20197 -13638 20216 -13604
rect 20250 -13638 20269 -13604
rect 20197 -13643 20269 -13638
rect 19307 -13662 20269 -13643
rect 19307 -13696 19420 -13662
rect 19454 -13696 19510 -13662
rect 19544 -13696 19600 -13662
rect 19634 -13696 19690 -13662
rect 19724 -13696 19780 -13662
rect 19814 -13696 19870 -13662
rect 19904 -13696 19960 -13662
rect 19994 -13696 20050 -13662
rect 20084 -13696 20140 -13662
rect 20174 -13696 20269 -13662
rect 19307 -13715 20269 -13696
rect 20595 -12772 21557 -12753
rect 20595 -12806 20727 -12772
rect 20761 -12806 20817 -12772
rect 20851 -12806 20907 -12772
rect 20941 -12806 20997 -12772
rect 21031 -12806 21087 -12772
rect 21121 -12806 21177 -12772
rect 21211 -12806 21267 -12772
rect 21301 -12806 21357 -12772
rect 21391 -12806 21447 -12772
rect 21481 -12806 21557 -12772
rect 20595 -12825 21557 -12806
rect 20595 -12850 20667 -12825
rect 20595 -12884 20614 -12850
rect 20648 -12884 20667 -12850
rect 20595 -12940 20667 -12884
rect 21485 -12884 21557 -12825
rect 20595 -12974 20614 -12940
rect 20648 -12974 20667 -12940
rect 20595 -13030 20667 -12974
rect 20595 -13064 20614 -13030
rect 20648 -13064 20667 -13030
rect 20595 -13120 20667 -13064
rect 20595 -13154 20614 -13120
rect 20648 -13154 20667 -13120
rect 20595 -13210 20667 -13154
rect 20595 -13244 20614 -13210
rect 20648 -13244 20667 -13210
rect 20595 -13300 20667 -13244
rect 20595 -13334 20614 -13300
rect 20648 -13334 20667 -13300
rect 20595 -13390 20667 -13334
rect 20595 -13424 20614 -13390
rect 20648 -13424 20667 -13390
rect 20595 -13480 20667 -13424
rect 20595 -13514 20614 -13480
rect 20648 -13514 20667 -13480
rect 20595 -13570 20667 -13514
rect 20595 -13604 20614 -13570
rect 20648 -13604 20667 -13570
rect 21485 -12918 21504 -12884
rect 21538 -12918 21557 -12884
rect 21485 -12974 21557 -12918
rect 21485 -13008 21504 -12974
rect 21538 -13008 21557 -12974
rect 21485 -13064 21557 -13008
rect 21485 -13098 21504 -13064
rect 21538 -13098 21557 -13064
rect 21485 -13154 21557 -13098
rect 21485 -13188 21504 -13154
rect 21538 -13188 21557 -13154
rect 21485 -13244 21557 -13188
rect 21485 -13278 21504 -13244
rect 21538 -13278 21557 -13244
rect 21485 -13334 21557 -13278
rect 21485 -13368 21504 -13334
rect 21538 -13368 21557 -13334
rect 21485 -13424 21557 -13368
rect 21485 -13458 21504 -13424
rect 21538 -13458 21557 -13424
rect 21485 -13514 21557 -13458
rect 21485 -13548 21504 -13514
rect 21538 -13548 21557 -13514
rect 20595 -13643 20667 -13604
rect 21485 -13604 21557 -13548
rect 21485 -13638 21504 -13604
rect 21538 -13638 21557 -13604
rect 21485 -13643 21557 -13638
rect 20595 -13662 21557 -13643
rect 20595 -13696 20708 -13662
rect 20742 -13696 20798 -13662
rect 20832 -13696 20888 -13662
rect 20922 -13696 20978 -13662
rect 21012 -13696 21068 -13662
rect 21102 -13696 21158 -13662
rect 21192 -13696 21248 -13662
rect 21282 -13696 21338 -13662
rect 21372 -13696 21428 -13662
rect 21462 -13696 21557 -13662
rect 20595 -13715 21557 -13696
rect 21883 -12772 22845 -12753
rect 21883 -12806 22015 -12772
rect 22049 -12806 22105 -12772
rect 22139 -12806 22195 -12772
rect 22229 -12806 22285 -12772
rect 22319 -12806 22375 -12772
rect 22409 -12806 22465 -12772
rect 22499 -12806 22555 -12772
rect 22589 -12806 22645 -12772
rect 22679 -12806 22735 -12772
rect 22769 -12806 22845 -12772
rect 21883 -12825 22845 -12806
rect 21883 -12850 21955 -12825
rect 21883 -12884 21902 -12850
rect 21936 -12884 21955 -12850
rect 21883 -12940 21955 -12884
rect 22773 -12884 22845 -12825
rect 21883 -12974 21902 -12940
rect 21936 -12974 21955 -12940
rect 21883 -13030 21955 -12974
rect 21883 -13064 21902 -13030
rect 21936 -13064 21955 -13030
rect 21883 -13120 21955 -13064
rect 21883 -13154 21902 -13120
rect 21936 -13154 21955 -13120
rect 21883 -13210 21955 -13154
rect 21883 -13244 21902 -13210
rect 21936 -13244 21955 -13210
rect 21883 -13300 21955 -13244
rect 21883 -13334 21902 -13300
rect 21936 -13334 21955 -13300
rect 21883 -13390 21955 -13334
rect 21883 -13424 21902 -13390
rect 21936 -13424 21955 -13390
rect 21883 -13480 21955 -13424
rect 21883 -13514 21902 -13480
rect 21936 -13514 21955 -13480
rect 21883 -13570 21955 -13514
rect 21883 -13604 21902 -13570
rect 21936 -13604 21955 -13570
rect 22773 -12918 22792 -12884
rect 22826 -12918 22845 -12884
rect 22773 -12974 22845 -12918
rect 22773 -13008 22792 -12974
rect 22826 -13008 22845 -12974
rect 22773 -13064 22845 -13008
rect 22773 -13098 22792 -13064
rect 22826 -13098 22845 -13064
rect 22773 -13154 22845 -13098
rect 22773 -13188 22792 -13154
rect 22826 -13188 22845 -13154
rect 22773 -13244 22845 -13188
rect 22773 -13278 22792 -13244
rect 22826 -13278 22845 -13244
rect 22773 -13334 22845 -13278
rect 22773 -13368 22792 -13334
rect 22826 -13368 22845 -13334
rect 22773 -13424 22845 -13368
rect 22773 -13458 22792 -13424
rect 22826 -13458 22845 -13424
rect 22773 -13514 22845 -13458
rect 22773 -13548 22792 -13514
rect 22826 -13548 22845 -13514
rect 21883 -13643 21955 -13604
rect 22773 -13604 22845 -13548
rect 22773 -13638 22792 -13604
rect 22826 -13638 22845 -13604
rect 22773 -13643 22845 -13638
rect 21883 -13662 22845 -13643
rect 21883 -13696 21996 -13662
rect 22030 -13696 22086 -13662
rect 22120 -13696 22176 -13662
rect 22210 -13696 22266 -13662
rect 22300 -13696 22356 -13662
rect 22390 -13696 22446 -13662
rect 22480 -13696 22536 -13662
rect 22570 -13696 22626 -13662
rect 22660 -13696 22716 -13662
rect 22750 -13696 22845 -13662
rect 21883 -13715 22845 -13696
rect 23171 -12772 24133 -12753
rect 23171 -12806 23303 -12772
rect 23337 -12806 23393 -12772
rect 23427 -12806 23483 -12772
rect 23517 -12806 23573 -12772
rect 23607 -12806 23663 -12772
rect 23697 -12806 23753 -12772
rect 23787 -12806 23843 -12772
rect 23877 -12806 23933 -12772
rect 23967 -12806 24023 -12772
rect 24057 -12806 24133 -12772
rect 23171 -12825 24133 -12806
rect 23171 -12850 23243 -12825
rect 23171 -12884 23190 -12850
rect 23224 -12884 23243 -12850
rect 23171 -12940 23243 -12884
rect 24061 -12884 24133 -12825
rect 23171 -12974 23190 -12940
rect 23224 -12974 23243 -12940
rect 23171 -13030 23243 -12974
rect 23171 -13064 23190 -13030
rect 23224 -13064 23243 -13030
rect 23171 -13120 23243 -13064
rect 23171 -13154 23190 -13120
rect 23224 -13154 23243 -13120
rect 23171 -13210 23243 -13154
rect 23171 -13244 23190 -13210
rect 23224 -13244 23243 -13210
rect 23171 -13300 23243 -13244
rect 23171 -13334 23190 -13300
rect 23224 -13334 23243 -13300
rect 23171 -13390 23243 -13334
rect 23171 -13424 23190 -13390
rect 23224 -13424 23243 -13390
rect 23171 -13480 23243 -13424
rect 23171 -13514 23190 -13480
rect 23224 -13514 23243 -13480
rect 23171 -13570 23243 -13514
rect 23171 -13604 23190 -13570
rect 23224 -13604 23243 -13570
rect 24061 -12918 24080 -12884
rect 24114 -12918 24133 -12884
rect 24061 -12974 24133 -12918
rect 24061 -13008 24080 -12974
rect 24114 -13008 24133 -12974
rect 24061 -13064 24133 -13008
rect 24061 -13098 24080 -13064
rect 24114 -13098 24133 -13064
rect 24061 -13154 24133 -13098
rect 24061 -13188 24080 -13154
rect 24114 -13188 24133 -13154
rect 24061 -13244 24133 -13188
rect 24061 -13278 24080 -13244
rect 24114 -13278 24133 -13244
rect 24061 -13334 24133 -13278
rect 24061 -13368 24080 -13334
rect 24114 -13368 24133 -13334
rect 24061 -13424 24133 -13368
rect 24061 -13458 24080 -13424
rect 24114 -13458 24133 -13424
rect 24061 -13514 24133 -13458
rect 24061 -13548 24080 -13514
rect 24114 -13548 24133 -13514
rect 23171 -13643 23243 -13604
rect 24061 -13604 24133 -13548
rect 24061 -13638 24080 -13604
rect 24114 -13638 24133 -13604
rect 24061 -13643 24133 -13638
rect 23171 -13662 24133 -13643
rect 23171 -13696 23284 -13662
rect 23318 -13696 23374 -13662
rect 23408 -13696 23464 -13662
rect 23498 -13696 23554 -13662
rect 23588 -13696 23644 -13662
rect 23678 -13696 23734 -13662
rect 23768 -13696 23824 -13662
rect 23858 -13696 23914 -13662
rect 23948 -13696 24004 -13662
rect 24038 -13696 24133 -13662
rect 23171 -13715 24133 -13696
rect 24459 -12772 25421 -12753
rect 24459 -12806 24591 -12772
rect 24625 -12806 24681 -12772
rect 24715 -12806 24771 -12772
rect 24805 -12806 24861 -12772
rect 24895 -12806 24951 -12772
rect 24985 -12806 25041 -12772
rect 25075 -12806 25131 -12772
rect 25165 -12806 25221 -12772
rect 25255 -12806 25311 -12772
rect 25345 -12806 25421 -12772
rect 24459 -12825 25421 -12806
rect 24459 -12850 24531 -12825
rect 24459 -12884 24478 -12850
rect 24512 -12884 24531 -12850
rect 24459 -12940 24531 -12884
rect 25349 -12884 25421 -12825
rect 24459 -12974 24478 -12940
rect 24512 -12974 24531 -12940
rect 24459 -13030 24531 -12974
rect 24459 -13064 24478 -13030
rect 24512 -13064 24531 -13030
rect 24459 -13120 24531 -13064
rect 24459 -13154 24478 -13120
rect 24512 -13154 24531 -13120
rect 24459 -13210 24531 -13154
rect 24459 -13244 24478 -13210
rect 24512 -13244 24531 -13210
rect 24459 -13300 24531 -13244
rect 24459 -13334 24478 -13300
rect 24512 -13334 24531 -13300
rect 24459 -13390 24531 -13334
rect 24459 -13424 24478 -13390
rect 24512 -13424 24531 -13390
rect 24459 -13480 24531 -13424
rect 24459 -13514 24478 -13480
rect 24512 -13514 24531 -13480
rect 24459 -13570 24531 -13514
rect 24459 -13604 24478 -13570
rect 24512 -13604 24531 -13570
rect 25349 -12918 25368 -12884
rect 25402 -12918 25421 -12884
rect 25349 -12974 25421 -12918
rect 25349 -13008 25368 -12974
rect 25402 -13008 25421 -12974
rect 25349 -13064 25421 -13008
rect 25349 -13098 25368 -13064
rect 25402 -13098 25421 -13064
rect 25349 -13154 25421 -13098
rect 25349 -13188 25368 -13154
rect 25402 -13188 25421 -13154
rect 25349 -13244 25421 -13188
rect 25349 -13278 25368 -13244
rect 25402 -13278 25421 -13244
rect 25349 -13334 25421 -13278
rect 25349 -13368 25368 -13334
rect 25402 -13368 25421 -13334
rect 25349 -13424 25421 -13368
rect 25349 -13458 25368 -13424
rect 25402 -13458 25421 -13424
rect 25349 -13514 25421 -13458
rect 25349 -13548 25368 -13514
rect 25402 -13548 25421 -13514
rect 24459 -13643 24531 -13604
rect 25349 -13604 25421 -13548
rect 25349 -13638 25368 -13604
rect 25402 -13638 25421 -13604
rect 25349 -13643 25421 -13638
rect 24459 -13662 25421 -13643
rect 24459 -13696 24572 -13662
rect 24606 -13696 24662 -13662
rect 24696 -13696 24752 -13662
rect 24786 -13696 24842 -13662
rect 24876 -13696 24932 -13662
rect 24966 -13696 25022 -13662
rect 25056 -13696 25112 -13662
rect 25146 -13696 25202 -13662
rect 25236 -13696 25292 -13662
rect 25326 -13696 25421 -13662
rect 24459 -13715 25421 -13696
rect 25747 -12772 26709 -12753
rect 25747 -12806 25879 -12772
rect 25913 -12806 25969 -12772
rect 26003 -12806 26059 -12772
rect 26093 -12806 26149 -12772
rect 26183 -12806 26239 -12772
rect 26273 -12806 26329 -12772
rect 26363 -12806 26419 -12772
rect 26453 -12806 26509 -12772
rect 26543 -12806 26599 -12772
rect 26633 -12806 26709 -12772
rect 25747 -12825 26709 -12806
rect 25747 -12850 25819 -12825
rect 25747 -12884 25766 -12850
rect 25800 -12884 25819 -12850
rect 25747 -12940 25819 -12884
rect 26637 -12884 26709 -12825
rect 25747 -12974 25766 -12940
rect 25800 -12974 25819 -12940
rect 25747 -13030 25819 -12974
rect 25747 -13064 25766 -13030
rect 25800 -13064 25819 -13030
rect 25747 -13120 25819 -13064
rect 25747 -13154 25766 -13120
rect 25800 -13154 25819 -13120
rect 25747 -13210 25819 -13154
rect 25747 -13244 25766 -13210
rect 25800 -13244 25819 -13210
rect 25747 -13300 25819 -13244
rect 25747 -13334 25766 -13300
rect 25800 -13334 25819 -13300
rect 25747 -13390 25819 -13334
rect 25747 -13424 25766 -13390
rect 25800 -13424 25819 -13390
rect 25747 -13480 25819 -13424
rect 25747 -13514 25766 -13480
rect 25800 -13514 25819 -13480
rect 25747 -13570 25819 -13514
rect 25747 -13604 25766 -13570
rect 25800 -13604 25819 -13570
rect 26637 -12918 26656 -12884
rect 26690 -12918 26709 -12884
rect 26637 -12974 26709 -12918
rect 26637 -13008 26656 -12974
rect 26690 -13008 26709 -12974
rect 26637 -13064 26709 -13008
rect 26637 -13098 26656 -13064
rect 26690 -13098 26709 -13064
rect 26637 -13154 26709 -13098
rect 26637 -13188 26656 -13154
rect 26690 -13188 26709 -13154
rect 26637 -13244 26709 -13188
rect 26637 -13278 26656 -13244
rect 26690 -13278 26709 -13244
rect 26637 -13334 26709 -13278
rect 26637 -13368 26656 -13334
rect 26690 -13368 26709 -13334
rect 26637 -13424 26709 -13368
rect 26637 -13458 26656 -13424
rect 26690 -13458 26709 -13424
rect 26637 -13514 26709 -13458
rect 26637 -13548 26656 -13514
rect 26690 -13548 26709 -13514
rect 25747 -13643 25819 -13604
rect 26637 -13604 26709 -13548
rect 26637 -13638 26656 -13604
rect 26690 -13638 26709 -13604
rect 26637 -13643 26709 -13638
rect 25747 -13662 26709 -13643
rect 25747 -13696 25860 -13662
rect 25894 -13696 25950 -13662
rect 25984 -13696 26040 -13662
rect 26074 -13696 26130 -13662
rect 26164 -13696 26220 -13662
rect 26254 -13696 26310 -13662
rect 26344 -13696 26400 -13662
rect 26434 -13696 26490 -13662
rect 26524 -13696 26580 -13662
rect 26614 -13696 26709 -13662
rect 25747 -13715 26709 -13696
rect 16731 -14060 17693 -14041
rect 16731 -14094 16863 -14060
rect 16897 -14094 16953 -14060
rect 16987 -14094 17043 -14060
rect 17077 -14094 17133 -14060
rect 17167 -14094 17223 -14060
rect 17257 -14094 17313 -14060
rect 17347 -14094 17403 -14060
rect 17437 -14094 17493 -14060
rect 17527 -14094 17583 -14060
rect 17617 -14094 17693 -14060
rect 16731 -14113 17693 -14094
rect 16731 -14138 16803 -14113
rect 16731 -14172 16750 -14138
rect 16784 -14172 16803 -14138
rect 16731 -14228 16803 -14172
rect 17621 -14172 17693 -14113
rect 16731 -14262 16750 -14228
rect 16784 -14262 16803 -14228
rect 16731 -14318 16803 -14262
rect 16731 -14352 16750 -14318
rect 16784 -14352 16803 -14318
rect 16731 -14408 16803 -14352
rect 16731 -14442 16750 -14408
rect 16784 -14442 16803 -14408
rect 16731 -14498 16803 -14442
rect 16731 -14532 16750 -14498
rect 16784 -14532 16803 -14498
rect 16731 -14588 16803 -14532
rect 16731 -14622 16750 -14588
rect 16784 -14622 16803 -14588
rect 16731 -14678 16803 -14622
rect 16731 -14712 16750 -14678
rect 16784 -14712 16803 -14678
rect 16731 -14768 16803 -14712
rect 16731 -14802 16750 -14768
rect 16784 -14802 16803 -14768
rect 16731 -14858 16803 -14802
rect 16731 -14892 16750 -14858
rect 16784 -14892 16803 -14858
rect 17621 -14206 17640 -14172
rect 17674 -14206 17693 -14172
rect 17621 -14262 17693 -14206
rect 17621 -14296 17640 -14262
rect 17674 -14296 17693 -14262
rect 17621 -14352 17693 -14296
rect 17621 -14386 17640 -14352
rect 17674 -14386 17693 -14352
rect 17621 -14442 17693 -14386
rect 17621 -14476 17640 -14442
rect 17674 -14476 17693 -14442
rect 17621 -14532 17693 -14476
rect 17621 -14566 17640 -14532
rect 17674 -14566 17693 -14532
rect 17621 -14622 17693 -14566
rect 17621 -14656 17640 -14622
rect 17674 -14656 17693 -14622
rect 17621 -14712 17693 -14656
rect 17621 -14746 17640 -14712
rect 17674 -14746 17693 -14712
rect 17621 -14802 17693 -14746
rect 17621 -14836 17640 -14802
rect 17674 -14836 17693 -14802
rect 16731 -14931 16803 -14892
rect 17621 -14892 17693 -14836
rect 17621 -14926 17640 -14892
rect 17674 -14926 17693 -14892
rect 17621 -14931 17693 -14926
rect 16731 -14950 17693 -14931
rect 16731 -14984 16844 -14950
rect 16878 -14984 16934 -14950
rect 16968 -14984 17024 -14950
rect 17058 -14984 17114 -14950
rect 17148 -14984 17204 -14950
rect 17238 -14984 17294 -14950
rect 17328 -14984 17384 -14950
rect 17418 -14984 17474 -14950
rect 17508 -14984 17564 -14950
rect 17598 -14984 17693 -14950
rect 16731 -15003 17693 -14984
rect 18019 -14060 18981 -14041
rect 18019 -14094 18151 -14060
rect 18185 -14094 18241 -14060
rect 18275 -14094 18331 -14060
rect 18365 -14094 18421 -14060
rect 18455 -14094 18511 -14060
rect 18545 -14094 18601 -14060
rect 18635 -14094 18691 -14060
rect 18725 -14094 18781 -14060
rect 18815 -14094 18871 -14060
rect 18905 -14094 18981 -14060
rect 18019 -14113 18981 -14094
rect 18019 -14138 18091 -14113
rect 18019 -14172 18038 -14138
rect 18072 -14172 18091 -14138
rect 18019 -14228 18091 -14172
rect 18909 -14172 18981 -14113
rect 18019 -14262 18038 -14228
rect 18072 -14262 18091 -14228
rect 18019 -14318 18091 -14262
rect 18019 -14352 18038 -14318
rect 18072 -14352 18091 -14318
rect 18019 -14408 18091 -14352
rect 18019 -14442 18038 -14408
rect 18072 -14442 18091 -14408
rect 18019 -14498 18091 -14442
rect 18019 -14532 18038 -14498
rect 18072 -14532 18091 -14498
rect 18019 -14588 18091 -14532
rect 18019 -14622 18038 -14588
rect 18072 -14622 18091 -14588
rect 18019 -14678 18091 -14622
rect 18019 -14712 18038 -14678
rect 18072 -14712 18091 -14678
rect 18019 -14768 18091 -14712
rect 18019 -14802 18038 -14768
rect 18072 -14802 18091 -14768
rect 18019 -14858 18091 -14802
rect 18019 -14892 18038 -14858
rect 18072 -14892 18091 -14858
rect 18909 -14206 18928 -14172
rect 18962 -14206 18981 -14172
rect 18909 -14262 18981 -14206
rect 18909 -14296 18928 -14262
rect 18962 -14296 18981 -14262
rect 18909 -14352 18981 -14296
rect 18909 -14386 18928 -14352
rect 18962 -14386 18981 -14352
rect 18909 -14442 18981 -14386
rect 18909 -14476 18928 -14442
rect 18962 -14476 18981 -14442
rect 18909 -14532 18981 -14476
rect 18909 -14566 18928 -14532
rect 18962 -14566 18981 -14532
rect 18909 -14622 18981 -14566
rect 18909 -14656 18928 -14622
rect 18962 -14656 18981 -14622
rect 18909 -14712 18981 -14656
rect 18909 -14746 18928 -14712
rect 18962 -14746 18981 -14712
rect 18909 -14802 18981 -14746
rect 18909 -14836 18928 -14802
rect 18962 -14836 18981 -14802
rect 18019 -14931 18091 -14892
rect 18909 -14892 18981 -14836
rect 18909 -14926 18928 -14892
rect 18962 -14926 18981 -14892
rect 18909 -14931 18981 -14926
rect 18019 -14950 18981 -14931
rect 18019 -14984 18132 -14950
rect 18166 -14984 18222 -14950
rect 18256 -14984 18312 -14950
rect 18346 -14984 18402 -14950
rect 18436 -14984 18492 -14950
rect 18526 -14984 18582 -14950
rect 18616 -14984 18672 -14950
rect 18706 -14984 18762 -14950
rect 18796 -14984 18852 -14950
rect 18886 -14984 18981 -14950
rect 18019 -15003 18981 -14984
rect 19307 -14060 20269 -14041
rect 19307 -14094 19439 -14060
rect 19473 -14094 19529 -14060
rect 19563 -14094 19619 -14060
rect 19653 -14094 19709 -14060
rect 19743 -14094 19799 -14060
rect 19833 -14094 19889 -14060
rect 19923 -14094 19979 -14060
rect 20013 -14094 20069 -14060
rect 20103 -14094 20159 -14060
rect 20193 -14094 20269 -14060
rect 19307 -14113 20269 -14094
rect 19307 -14138 19379 -14113
rect 19307 -14172 19326 -14138
rect 19360 -14172 19379 -14138
rect 19307 -14228 19379 -14172
rect 20197 -14172 20269 -14113
rect 19307 -14262 19326 -14228
rect 19360 -14262 19379 -14228
rect 19307 -14318 19379 -14262
rect 19307 -14352 19326 -14318
rect 19360 -14352 19379 -14318
rect 19307 -14408 19379 -14352
rect 19307 -14442 19326 -14408
rect 19360 -14442 19379 -14408
rect 19307 -14498 19379 -14442
rect 19307 -14532 19326 -14498
rect 19360 -14532 19379 -14498
rect 19307 -14588 19379 -14532
rect 19307 -14622 19326 -14588
rect 19360 -14622 19379 -14588
rect 19307 -14678 19379 -14622
rect 19307 -14712 19326 -14678
rect 19360 -14712 19379 -14678
rect 19307 -14768 19379 -14712
rect 19307 -14802 19326 -14768
rect 19360 -14802 19379 -14768
rect 19307 -14858 19379 -14802
rect 19307 -14892 19326 -14858
rect 19360 -14892 19379 -14858
rect 20197 -14206 20216 -14172
rect 20250 -14206 20269 -14172
rect 20197 -14262 20269 -14206
rect 20197 -14296 20216 -14262
rect 20250 -14296 20269 -14262
rect 20197 -14352 20269 -14296
rect 20197 -14386 20216 -14352
rect 20250 -14386 20269 -14352
rect 20197 -14442 20269 -14386
rect 20197 -14476 20216 -14442
rect 20250 -14476 20269 -14442
rect 20197 -14532 20269 -14476
rect 20197 -14566 20216 -14532
rect 20250 -14566 20269 -14532
rect 20197 -14622 20269 -14566
rect 20197 -14656 20216 -14622
rect 20250 -14656 20269 -14622
rect 20197 -14712 20269 -14656
rect 20197 -14746 20216 -14712
rect 20250 -14746 20269 -14712
rect 20197 -14802 20269 -14746
rect 20197 -14836 20216 -14802
rect 20250 -14836 20269 -14802
rect 19307 -14931 19379 -14892
rect 20197 -14892 20269 -14836
rect 20197 -14926 20216 -14892
rect 20250 -14926 20269 -14892
rect 20197 -14931 20269 -14926
rect 19307 -14950 20269 -14931
rect 19307 -14984 19420 -14950
rect 19454 -14984 19510 -14950
rect 19544 -14984 19600 -14950
rect 19634 -14984 19690 -14950
rect 19724 -14984 19780 -14950
rect 19814 -14984 19870 -14950
rect 19904 -14984 19960 -14950
rect 19994 -14984 20050 -14950
rect 20084 -14984 20140 -14950
rect 20174 -14984 20269 -14950
rect 19307 -15003 20269 -14984
rect 20595 -14060 21557 -14041
rect 20595 -14094 20727 -14060
rect 20761 -14094 20817 -14060
rect 20851 -14094 20907 -14060
rect 20941 -14094 20997 -14060
rect 21031 -14094 21087 -14060
rect 21121 -14094 21177 -14060
rect 21211 -14094 21267 -14060
rect 21301 -14094 21357 -14060
rect 21391 -14094 21447 -14060
rect 21481 -14094 21557 -14060
rect 20595 -14113 21557 -14094
rect 20595 -14138 20667 -14113
rect 20595 -14172 20614 -14138
rect 20648 -14172 20667 -14138
rect 20595 -14228 20667 -14172
rect 21485 -14172 21557 -14113
rect 20595 -14262 20614 -14228
rect 20648 -14262 20667 -14228
rect 20595 -14318 20667 -14262
rect 20595 -14352 20614 -14318
rect 20648 -14352 20667 -14318
rect 20595 -14408 20667 -14352
rect 20595 -14442 20614 -14408
rect 20648 -14442 20667 -14408
rect 20595 -14498 20667 -14442
rect 20595 -14532 20614 -14498
rect 20648 -14532 20667 -14498
rect 20595 -14588 20667 -14532
rect 20595 -14622 20614 -14588
rect 20648 -14622 20667 -14588
rect 20595 -14678 20667 -14622
rect 20595 -14712 20614 -14678
rect 20648 -14712 20667 -14678
rect 20595 -14768 20667 -14712
rect 20595 -14802 20614 -14768
rect 20648 -14802 20667 -14768
rect 20595 -14858 20667 -14802
rect 20595 -14892 20614 -14858
rect 20648 -14892 20667 -14858
rect 21485 -14206 21504 -14172
rect 21538 -14206 21557 -14172
rect 21485 -14262 21557 -14206
rect 21485 -14296 21504 -14262
rect 21538 -14296 21557 -14262
rect 21485 -14352 21557 -14296
rect 21485 -14386 21504 -14352
rect 21538 -14386 21557 -14352
rect 21485 -14442 21557 -14386
rect 21485 -14476 21504 -14442
rect 21538 -14476 21557 -14442
rect 21485 -14532 21557 -14476
rect 21485 -14566 21504 -14532
rect 21538 -14566 21557 -14532
rect 21485 -14622 21557 -14566
rect 21485 -14656 21504 -14622
rect 21538 -14656 21557 -14622
rect 21485 -14712 21557 -14656
rect 21485 -14746 21504 -14712
rect 21538 -14746 21557 -14712
rect 21485 -14802 21557 -14746
rect 21485 -14836 21504 -14802
rect 21538 -14836 21557 -14802
rect 20595 -14931 20667 -14892
rect 21485 -14892 21557 -14836
rect 21485 -14926 21504 -14892
rect 21538 -14926 21557 -14892
rect 21485 -14931 21557 -14926
rect 20595 -14950 21557 -14931
rect 20595 -14984 20708 -14950
rect 20742 -14984 20798 -14950
rect 20832 -14984 20888 -14950
rect 20922 -14984 20978 -14950
rect 21012 -14984 21068 -14950
rect 21102 -14984 21158 -14950
rect 21192 -14984 21248 -14950
rect 21282 -14984 21338 -14950
rect 21372 -14984 21428 -14950
rect 21462 -14984 21557 -14950
rect 20595 -15003 21557 -14984
rect 21883 -14060 22845 -14041
rect 21883 -14094 22015 -14060
rect 22049 -14094 22105 -14060
rect 22139 -14094 22195 -14060
rect 22229 -14094 22285 -14060
rect 22319 -14094 22375 -14060
rect 22409 -14094 22465 -14060
rect 22499 -14094 22555 -14060
rect 22589 -14094 22645 -14060
rect 22679 -14094 22735 -14060
rect 22769 -14094 22845 -14060
rect 21883 -14113 22845 -14094
rect 21883 -14138 21955 -14113
rect 21883 -14172 21902 -14138
rect 21936 -14172 21955 -14138
rect 21883 -14228 21955 -14172
rect 22773 -14172 22845 -14113
rect 21883 -14262 21902 -14228
rect 21936 -14262 21955 -14228
rect 21883 -14318 21955 -14262
rect 21883 -14352 21902 -14318
rect 21936 -14352 21955 -14318
rect 21883 -14408 21955 -14352
rect 21883 -14442 21902 -14408
rect 21936 -14442 21955 -14408
rect 21883 -14498 21955 -14442
rect 21883 -14532 21902 -14498
rect 21936 -14532 21955 -14498
rect 21883 -14588 21955 -14532
rect 21883 -14622 21902 -14588
rect 21936 -14622 21955 -14588
rect 21883 -14678 21955 -14622
rect 21883 -14712 21902 -14678
rect 21936 -14712 21955 -14678
rect 21883 -14768 21955 -14712
rect 21883 -14802 21902 -14768
rect 21936 -14802 21955 -14768
rect 21883 -14858 21955 -14802
rect 21883 -14892 21902 -14858
rect 21936 -14892 21955 -14858
rect 22773 -14206 22792 -14172
rect 22826 -14206 22845 -14172
rect 22773 -14262 22845 -14206
rect 22773 -14296 22792 -14262
rect 22826 -14296 22845 -14262
rect 22773 -14352 22845 -14296
rect 22773 -14386 22792 -14352
rect 22826 -14386 22845 -14352
rect 22773 -14442 22845 -14386
rect 22773 -14476 22792 -14442
rect 22826 -14476 22845 -14442
rect 22773 -14532 22845 -14476
rect 22773 -14566 22792 -14532
rect 22826 -14566 22845 -14532
rect 22773 -14622 22845 -14566
rect 22773 -14656 22792 -14622
rect 22826 -14656 22845 -14622
rect 22773 -14712 22845 -14656
rect 22773 -14746 22792 -14712
rect 22826 -14746 22845 -14712
rect 22773 -14802 22845 -14746
rect 22773 -14836 22792 -14802
rect 22826 -14836 22845 -14802
rect 21883 -14931 21955 -14892
rect 22773 -14892 22845 -14836
rect 22773 -14926 22792 -14892
rect 22826 -14926 22845 -14892
rect 22773 -14931 22845 -14926
rect 21883 -14950 22845 -14931
rect 21883 -14984 21996 -14950
rect 22030 -14984 22086 -14950
rect 22120 -14984 22176 -14950
rect 22210 -14984 22266 -14950
rect 22300 -14984 22356 -14950
rect 22390 -14984 22446 -14950
rect 22480 -14984 22536 -14950
rect 22570 -14984 22626 -14950
rect 22660 -14984 22716 -14950
rect 22750 -14984 22845 -14950
rect 21883 -15003 22845 -14984
rect 23171 -14060 24133 -14041
rect 23171 -14094 23303 -14060
rect 23337 -14094 23393 -14060
rect 23427 -14094 23483 -14060
rect 23517 -14094 23573 -14060
rect 23607 -14094 23663 -14060
rect 23697 -14094 23753 -14060
rect 23787 -14094 23843 -14060
rect 23877 -14094 23933 -14060
rect 23967 -14094 24023 -14060
rect 24057 -14094 24133 -14060
rect 23171 -14113 24133 -14094
rect 23171 -14138 23243 -14113
rect 23171 -14172 23190 -14138
rect 23224 -14172 23243 -14138
rect 23171 -14228 23243 -14172
rect 24061 -14172 24133 -14113
rect 23171 -14262 23190 -14228
rect 23224 -14262 23243 -14228
rect 23171 -14318 23243 -14262
rect 23171 -14352 23190 -14318
rect 23224 -14352 23243 -14318
rect 23171 -14408 23243 -14352
rect 23171 -14442 23190 -14408
rect 23224 -14442 23243 -14408
rect 23171 -14498 23243 -14442
rect 23171 -14532 23190 -14498
rect 23224 -14532 23243 -14498
rect 23171 -14588 23243 -14532
rect 23171 -14622 23190 -14588
rect 23224 -14622 23243 -14588
rect 23171 -14678 23243 -14622
rect 23171 -14712 23190 -14678
rect 23224 -14712 23243 -14678
rect 23171 -14768 23243 -14712
rect 23171 -14802 23190 -14768
rect 23224 -14802 23243 -14768
rect 23171 -14858 23243 -14802
rect 23171 -14892 23190 -14858
rect 23224 -14892 23243 -14858
rect 24061 -14206 24080 -14172
rect 24114 -14206 24133 -14172
rect 24061 -14262 24133 -14206
rect 24061 -14296 24080 -14262
rect 24114 -14296 24133 -14262
rect 24061 -14352 24133 -14296
rect 24061 -14386 24080 -14352
rect 24114 -14386 24133 -14352
rect 24061 -14442 24133 -14386
rect 24061 -14476 24080 -14442
rect 24114 -14476 24133 -14442
rect 24061 -14532 24133 -14476
rect 24061 -14566 24080 -14532
rect 24114 -14566 24133 -14532
rect 24061 -14622 24133 -14566
rect 24061 -14656 24080 -14622
rect 24114 -14656 24133 -14622
rect 24061 -14712 24133 -14656
rect 24061 -14746 24080 -14712
rect 24114 -14746 24133 -14712
rect 24061 -14802 24133 -14746
rect 24061 -14836 24080 -14802
rect 24114 -14836 24133 -14802
rect 23171 -14931 23243 -14892
rect 24061 -14892 24133 -14836
rect 24061 -14926 24080 -14892
rect 24114 -14926 24133 -14892
rect 24061 -14931 24133 -14926
rect 23171 -14950 24133 -14931
rect 23171 -14984 23284 -14950
rect 23318 -14984 23374 -14950
rect 23408 -14984 23464 -14950
rect 23498 -14984 23554 -14950
rect 23588 -14984 23644 -14950
rect 23678 -14984 23734 -14950
rect 23768 -14984 23824 -14950
rect 23858 -14984 23914 -14950
rect 23948 -14984 24004 -14950
rect 24038 -14984 24133 -14950
rect 23171 -15003 24133 -14984
rect 24459 -14060 25421 -14041
rect 24459 -14094 24591 -14060
rect 24625 -14094 24681 -14060
rect 24715 -14094 24771 -14060
rect 24805 -14094 24861 -14060
rect 24895 -14094 24951 -14060
rect 24985 -14094 25041 -14060
rect 25075 -14094 25131 -14060
rect 25165 -14094 25221 -14060
rect 25255 -14094 25311 -14060
rect 25345 -14094 25421 -14060
rect 24459 -14113 25421 -14094
rect 24459 -14138 24531 -14113
rect 24459 -14172 24478 -14138
rect 24512 -14172 24531 -14138
rect 24459 -14228 24531 -14172
rect 25349 -14172 25421 -14113
rect 24459 -14262 24478 -14228
rect 24512 -14262 24531 -14228
rect 24459 -14318 24531 -14262
rect 24459 -14352 24478 -14318
rect 24512 -14352 24531 -14318
rect 24459 -14408 24531 -14352
rect 24459 -14442 24478 -14408
rect 24512 -14442 24531 -14408
rect 24459 -14498 24531 -14442
rect 24459 -14532 24478 -14498
rect 24512 -14532 24531 -14498
rect 24459 -14588 24531 -14532
rect 24459 -14622 24478 -14588
rect 24512 -14622 24531 -14588
rect 24459 -14678 24531 -14622
rect 24459 -14712 24478 -14678
rect 24512 -14712 24531 -14678
rect 24459 -14768 24531 -14712
rect 24459 -14802 24478 -14768
rect 24512 -14802 24531 -14768
rect 24459 -14858 24531 -14802
rect 24459 -14892 24478 -14858
rect 24512 -14892 24531 -14858
rect 25349 -14206 25368 -14172
rect 25402 -14206 25421 -14172
rect 25349 -14262 25421 -14206
rect 25349 -14296 25368 -14262
rect 25402 -14296 25421 -14262
rect 25349 -14352 25421 -14296
rect 25349 -14386 25368 -14352
rect 25402 -14386 25421 -14352
rect 25349 -14442 25421 -14386
rect 25349 -14476 25368 -14442
rect 25402 -14476 25421 -14442
rect 25349 -14532 25421 -14476
rect 25349 -14566 25368 -14532
rect 25402 -14566 25421 -14532
rect 25349 -14622 25421 -14566
rect 25349 -14656 25368 -14622
rect 25402 -14656 25421 -14622
rect 25349 -14712 25421 -14656
rect 25349 -14746 25368 -14712
rect 25402 -14746 25421 -14712
rect 25349 -14802 25421 -14746
rect 25349 -14836 25368 -14802
rect 25402 -14836 25421 -14802
rect 24459 -14931 24531 -14892
rect 25349 -14892 25421 -14836
rect 25349 -14926 25368 -14892
rect 25402 -14926 25421 -14892
rect 25349 -14931 25421 -14926
rect 24459 -14950 25421 -14931
rect 24459 -14984 24572 -14950
rect 24606 -14984 24662 -14950
rect 24696 -14984 24752 -14950
rect 24786 -14984 24842 -14950
rect 24876 -14984 24932 -14950
rect 24966 -14984 25022 -14950
rect 25056 -14984 25112 -14950
rect 25146 -14984 25202 -14950
rect 25236 -14984 25292 -14950
rect 25326 -14984 25421 -14950
rect 24459 -15003 25421 -14984
rect 25747 -14060 26709 -14041
rect 25747 -14094 25879 -14060
rect 25913 -14094 25969 -14060
rect 26003 -14094 26059 -14060
rect 26093 -14094 26149 -14060
rect 26183 -14094 26239 -14060
rect 26273 -14094 26329 -14060
rect 26363 -14094 26419 -14060
rect 26453 -14094 26509 -14060
rect 26543 -14094 26599 -14060
rect 26633 -14094 26709 -14060
rect 25747 -14113 26709 -14094
rect 25747 -14138 25819 -14113
rect 25747 -14172 25766 -14138
rect 25800 -14172 25819 -14138
rect 25747 -14228 25819 -14172
rect 26637 -14172 26709 -14113
rect 25747 -14262 25766 -14228
rect 25800 -14262 25819 -14228
rect 25747 -14318 25819 -14262
rect 25747 -14352 25766 -14318
rect 25800 -14352 25819 -14318
rect 25747 -14408 25819 -14352
rect 25747 -14442 25766 -14408
rect 25800 -14442 25819 -14408
rect 25747 -14498 25819 -14442
rect 25747 -14532 25766 -14498
rect 25800 -14532 25819 -14498
rect 25747 -14588 25819 -14532
rect 25747 -14622 25766 -14588
rect 25800 -14622 25819 -14588
rect 25747 -14678 25819 -14622
rect 25747 -14712 25766 -14678
rect 25800 -14712 25819 -14678
rect 25747 -14768 25819 -14712
rect 25747 -14802 25766 -14768
rect 25800 -14802 25819 -14768
rect 25747 -14858 25819 -14802
rect 25747 -14892 25766 -14858
rect 25800 -14892 25819 -14858
rect 26637 -14206 26656 -14172
rect 26690 -14206 26709 -14172
rect 26637 -14262 26709 -14206
rect 26637 -14296 26656 -14262
rect 26690 -14296 26709 -14262
rect 26637 -14352 26709 -14296
rect 26637 -14386 26656 -14352
rect 26690 -14386 26709 -14352
rect 26637 -14442 26709 -14386
rect 26637 -14476 26656 -14442
rect 26690 -14476 26709 -14442
rect 26637 -14532 26709 -14476
rect 26637 -14566 26656 -14532
rect 26690 -14566 26709 -14532
rect 26637 -14622 26709 -14566
rect 26637 -14656 26656 -14622
rect 26690 -14656 26709 -14622
rect 26637 -14712 26709 -14656
rect 26637 -14746 26656 -14712
rect 26690 -14746 26709 -14712
rect 26637 -14802 26709 -14746
rect 26637 -14836 26656 -14802
rect 26690 -14836 26709 -14802
rect 25747 -14931 25819 -14892
rect 26637 -14892 26709 -14836
rect 26637 -14926 26656 -14892
rect 26690 -14926 26709 -14892
rect 26637 -14931 26709 -14926
rect 25747 -14950 26709 -14931
rect 25747 -14984 25860 -14950
rect 25894 -14984 25950 -14950
rect 25984 -14984 26040 -14950
rect 26074 -14984 26130 -14950
rect 26164 -14984 26220 -14950
rect 26254 -14984 26310 -14950
rect 26344 -14984 26400 -14950
rect 26434 -14984 26490 -14950
rect 26524 -14984 26580 -14950
rect 26614 -14984 26709 -14950
rect 25747 -15003 26709 -14984
rect 16731 -15348 17693 -15329
rect 16731 -15382 16863 -15348
rect 16897 -15382 16953 -15348
rect 16987 -15382 17043 -15348
rect 17077 -15382 17133 -15348
rect 17167 -15382 17223 -15348
rect 17257 -15382 17313 -15348
rect 17347 -15382 17403 -15348
rect 17437 -15382 17493 -15348
rect 17527 -15382 17583 -15348
rect 17617 -15382 17693 -15348
rect 16731 -15401 17693 -15382
rect 16731 -15426 16803 -15401
rect 16731 -15460 16750 -15426
rect 16784 -15460 16803 -15426
rect 16731 -15516 16803 -15460
rect 17621 -15460 17693 -15401
rect 16731 -15550 16750 -15516
rect 16784 -15550 16803 -15516
rect 16731 -15606 16803 -15550
rect 16731 -15640 16750 -15606
rect 16784 -15640 16803 -15606
rect 16731 -15696 16803 -15640
rect 16731 -15730 16750 -15696
rect 16784 -15730 16803 -15696
rect 16731 -15786 16803 -15730
rect 16731 -15820 16750 -15786
rect 16784 -15820 16803 -15786
rect 16731 -15876 16803 -15820
rect 16731 -15910 16750 -15876
rect 16784 -15910 16803 -15876
rect 16731 -15966 16803 -15910
rect 16731 -16000 16750 -15966
rect 16784 -16000 16803 -15966
rect 16731 -16056 16803 -16000
rect 16731 -16090 16750 -16056
rect 16784 -16090 16803 -16056
rect 16731 -16146 16803 -16090
rect 16731 -16180 16750 -16146
rect 16784 -16180 16803 -16146
rect 17621 -15494 17640 -15460
rect 17674 -15494 17693 -15460
rect 17621 -15550 17693 -15494
rect 17621 -15584 17640 -15550
rect 17674 -15584 17693 -15550
rect 17621 -15640 17693 -15584
rect 17621 -15674 17640 -15640
rect 17674 -15674 17693 -15640
rect 17621 -15730 17693 -15674
rect 17621 -15764 17640 -15730
rect 17674 -15764 17693 -15730
rect 17621 -15820 17693 -15764
rect 17621 -15854 17640 -15820
rect 17674 -15854 17693 -15820
rect 17621 -15910 17693 -15854
rect 17621 -15944 17640 -15910
rect 17674 -15944 17693 -15910
rect 17621 -16000 17693 -15944
rect 17621 -16034 17640 -16000
rect 17674 -16034 17693 -16000
rect 17621 -16090 17693 -16034
rect 17621 -16124 17640 -16090
rect 17674 -16124 17693 -16090
rect 16731 -16219 16803 -16180
rect 17621 -16180 17693 -16124
rect 17621 -16214 17640 -16180
rect 17674 -16214 17693 -16180
rect 17621 -16219 17693 -16214
rect 16731 -16238 17693 -16219
rect 16731 -16272 16844 -16238
rect 16878 -16272 16934 -16238
rect 16968 -16272 17024 -16238
rect 17058 -16272 17114 -16238
rect 17148 -16272 17204 -16238
rect 17238 -16272 17294 -16238
rect 17328 -16272 17384 -16238
rect 17418 -16272 17474 -16238
rect 17508 -16272 17564 -16238
rect 17598 -16272 17693 -16238
rect 16731 -16291 17693 -16272
rect 18019 -15348 18981 -15329
rect 18019 -15382 18151 -15348
rect 18185 -15382 18241 -15348
rect 18275 -15382 18331 -15348
rect 18365 -15382 18421 -15348
rect 18455 -15382 18511 -15348
rect 18545 -15382 18601 -15348
rect 18635 -15382 18691 -15348
rect 18725 -15382 18781 -15348
rect 18815 -15382 18871 -15348
rect 18905 -15382 18981 -15348
rect 18019 -15401 18981 -15382
rect 18019 -15426 18091 -15401
rect 18019 -15460 18038 -15426
rect 18072 -15460 18091 -15426
rect 18019 -15516 18091 -15460
rect 18909 -15460 18981 -15401
rect 18019 -15550 18038 -15516
rect 18072 -15550 18091 -15516
rect 18019 -15606 18091 -15550
rect 18019 -15640 18038 -15606
rect 18072 -15640 18091 -15606
rect 18019 -15696 18091 -15640
rect 18019 -15730 18038 -15696
rect 18072 -15730 18091 -15696
rect 18019 -15786 18091 -15730
rect 18019 -15820 18038 -15786
rect 18072 -15820 18091 -15786
rect 18019 -15876 18091 -15820
rect 18019 -15910 18038 -15876
rect 18072 -15910 18091 -15876
rect 18019 -15966 18091 -15910
rect 18019 -16000 18038 -15966
rect 18072 -16000 18091 -15966
rect 18019 -16056 18091 -16000
rect 18019 -16090 18038 -16056
rect 18072 -16090 18091 -16056
rect 18019 -16146 18091 -16090
rect 18019 -16180 18038 -16146
rect 18072 -16180 18091 -16146
rect 18909 -15494 18928 -15460
rect 18962 -15494 18981 -15460
rect 18909 -15550 18981 -15494
rect 18909 -15584 18928 -15550
rect 18962 -15584 18981 -15550
rect 18909 -15640 18981 -15584
rect 18909 -15674 18928 -15640
rect 18962 -15674 18981 -15640
rect 18909 -15730 18981 -15674
rect 18909 -15764 18928 -15730
rect 18962 -15764 18981 -15730
rect 18909 -15820 18981 -15764
rect 18909 -15854 18928 -15820
rect 18962 -15854 18981 -15820
rect 18909 -15910 18981 -15854
rect 18909 -15944 18928 -15910
rect 18962 -15944 18981 -15910
rect 18909 -16000 18981 -15944
rect 18909 -16034 18928 -16000
rect 18962 -16034 18981 -16000
rect 18909 -16090 18981 -16034
rect 18909 -16124 18928 -16090
rect 18962 -16124 18981 -16090
rect 18019 -16219 18091 -16180
rect 18909 -16180 18981 -16124
rect 18909 -16214 18928 -16180
rect 18962 -16214 18981 -16180
rect 18909 -16219 18981 -16214
rect 18019 -16238 18981 -16219
rect 18019 -16272 18132 -16238
rect 18166 -16272 18222 -16238
rect 18256 -16272 18312 -16238
rect 18346 -16272 18402 -16238
rect 18436 -16272 18492 -16238
rect 18526 -16272 18582 -16238
rect 18616 -16272 18672 -16238
rect 18706 -16272 18762 -16238
rect 18796 -16272 18852 -16238
rect 18886 -16272 18981 -16238
rect 18019 -16291 18981 -16272
rect 19307 -15348 20269 -15329
rect 19307 -15382 19439 -15348
rect 19473 -15382 19529 -15348
rect 19563 -15382 19619 -15348
rect 19653 -15382 19709 -15348
rect 19743 -15382 19799 -15348
rect 19833 -15382 19889 -15348
rect 19923 -15382 19979 -15348
rect 20013 -15382 20069 -15348
rect 20103 -15382 20159 -15348
rect 20193 -15382 20269 -15348
rect 19307 -15401 20269 -15382
rect 19307 -15426 19379 -15401
rect 19307 -15460 19326 -15426
rect 19360 -15460 19379 -15426
rect 19307 -15516 19379 -15460
rect 20197 -15460 20269 -15401
rect 19307 -15550 19326 -15516
rect 19360 -15550 19379 -15516
rect 19307 -15606 19379 -15550
rect 19307 -15640 19326 -15606
rect 19360 -15640 19379 -15606
rect 19307 -15696 19379 -15640
rect 19307 -15730 19326 -15696
rect 19360 -15730 19379 -15696
rect 19307 -15786 19379 -15730
rect 19307 -15820 19326 -15786
rect 19360 -15820 19379 -15786
rect 19307 -15876 19379 -15820
rect 19307 -15910 19326 -15876
rect 19360 -15910 19379 -15876
rect 19307 -15966 19379 -15910
rect 19307 -16000 19326 -15966
rect 19360 -16000 19379 -15966
rect 19307 -16056 19379 -16000
rect 19307 -16090 19326 -16056
rect 19360 -16090 19379 -16056
rect 19307 -16146 19379 -16090
rect 19307 -16180 19326 -16146
rect 19360 -16180 19379 -16146
rect 20197 -15494 20216 -15460
rect 20250 -15494 20269 -15460
rect 20197 -15550 20269 -15494
rect 20197 -15584 20216 -15550
rect 20250 -15584 20269 -15550
rect 20197 -15640 20269 -15584
rect 20197 -15674 20216 -15640
rect 20250 -15674 20269 -15640
rect 20197 -15730 20269 -15674
rect 20197 -15764 20216 -15730
rect 20250 -15764 20269 -15730
rect 20197 -15820 20269 -15764
rect 20197 -15854 20216 -15820
rect 20250 -15854 20269 -15820
rect 20197 -15910 20269 -15854
rect 20197 -15944 20216 -15910
rect 20250 -15944 20269 -15910
rect 20197 -16000 20269 -15944
rect 20197 -16034 20216 -16000
rect 20250 -16034 20269 -16000
rect 20197 -16090 20269 -16034
rect 20197 -16124 20216 -16090
rect 20250 -16124 20269 -16090
rect 19307 -16219 19379 -16180
rect 20197 -16180 20269 -16124
rect 20197 -16214 20216 -16180
rect 20250 -16214 20269 -16180
rect 20197 -16219 20269 -16214
rect 19307 -16238 20269 -16219
rect 19307 -16272 19420 -16238
rect 19454 -16272 19510 -16238
rect 19544 -16272 19600 -16238
rect 19634 -16272 19690 -16238
rect 19724 -16272 19780 -16238
rect 19814 -16272 19870 -16238
rect 19904 -16272 19960 -16238
rect 19994 -16272 20050 -16238
rect 20084 -16272 20140 -16238
rect 20174 -16272 20269 -16238
rect 19307 -16291 20269 -16272
rect 20595 -15348 21557 -15329
rect 20595 -15382 20727 -15348
rect 20761 -15382 20817 -15348
rect 20851 -15382 20907 -15348
rect 20941 -15382 20997 -15348
rect 21031 -15382 21087 -15348
rect 21121 -15382 21177 -15348
rect 21211 -15382 21267 -15348
rect 21301 -15382 21357 -15348
rect 21391 -15382 21447 -15348
rect 21481 -15382 21557 -15348
rect 20595 -15401 21557 -15382
rect 20595 -15426 20667 -15401
rect 20595 -15460 20614 -15426
rect 20648 -15460 20667 -15426
rect 20595 -15516 20667 -15460
rect 21485 -15460 21557 -15401
rect 20595 -15550 20614 -15516
rect 20648 -15550 20667 -15516
rect 20595 -15606 20667 -15550
rect 20595 -15640 20614 -15606
rect 20648 -15640 20667 -15606
rect 20595 -15696 20667 -15640
rect 20595 -15730 20614 -15696
rect 20648 -15730 20667 -15696
rect 20595 -15786 20667 -15730
rect 20595 -15820 20614 -15786
rect 20648 -15820 20667 -15786
rect 20595 -15876 20667 -15820
rect 20595 -15910 20614 -15876
rect 20648 -15910 20667 -15876
rect 20595 -15966 20667 -15910
rect 20595 -16000 20614 -15966
rect 20648 -16000 20667 -15966
rect 20595 -16056 20667 -16000
rect 20595 -16090 20614 -16056
rect 20648 -16090 20667 -16056
rect 20595 -16146 20667 -16090
rect 20595 -16180 20614 -16146
rect 20648 -16180 20667 -16146
rect 21485 -15494 21504 -15460
rect 21538 -15494 21557 -15460
rect 21485 -15550 21557 -15494
rect 21485 -15584 21504 -15550
rect 21538 -15584 21557 -15550
rect 21485 -15640 21557 -15584
rect 21485 -15674 21504 -15640
rect 21538 -15674 21557 -15640
rect 21485 -15730 21557 -15674
rect 21485 -15764 21504 -15730
rect 21538 -15764 21557 -15730
rect 21485 -15820 21557 -15764
rect 21485 -15854 21504 -15820
rect 21538 -15854 21557 -15820
rect 21485 -15910 21557 -15854
rect 21485 -15944 21504 -15910
rect 21538 -15944 21557 -15910
rect 21485 -16000 21557 -15944
rect 21485 -16034 21504 -16000
rect 21538 -16034 21557 -16000
rect 21485 -16090 21557 -16034
rect 21485 -16124 21504 -16090
rect 21538 -16124 21557 -16090
rect 20595 -16219 20667 -16180
rect 21485 -16180 21557 -16124
rect 21485 -16214 21504 -16180
rect 21538 -16214 21557 -16180
rect 21485 -16219 21557 -16214
rect 20595 -16238 21557 -16219
rect 20595 -16272 20708 -16238
rect 20742 -16272 20798 -16238
rect 20832 -16272 20888 -16238
rect 20922 -16272 20978 -16238
rect 21012 -16272 21068 -16238
rect 21102 -16272 21158 -16238
rect 21192 -16272 21248 -16238
rect 21282 -16272 21338 -16238
rect 21372 -16272 21428 -16238
rect 21462 -16272 21557 -16238
rect 20595 -16291 21557 -16272
rect 21883 -15348 22845 -15329
rect 21883 -15382 22015 -15348
rect 22049 -15382 22105 -15348
rect 22139 -15382 22195 -15348
rect 22229 -15382 22285 -15348
rect 22319 -15382 22375 -15348
rect 22409 -15382 22465 -15348
rect 22499 -15382 22555 -15348
rect 22589 -15382 22645 -15348
rect 22679 -15382 22735 -15348
rect 22769 -15382 22845 -15348
rect 21883 -15401 22845 -15382
rect 21883 -15426 21955 -15401
rect 21883 -15460 21902 -15426
rect 21936 -15460 21955 -15426
rect 21883 -15516 21955 -15460
rect 22773 -15460 22845 -15401
rect 21883 -15550 21902 -15516
rect 21936 -15550 21955 -15516
rect 21883 -15606 21955 -15550
rect 21883 -15640 21902 -15606
rect 21936 -15640 21955 -15606
rect 21883 -15696 21955 -15640
rect 21883 -15730 21902 -15696
rect 21936 -15730 21955 -15696
rect 21883 -15786 21955 -15730
rect 21883 -15820 21902 -15786
rect 21936 -15820 21955 -15786
rect 21883 -15876 21955 -15820
rect 21883 -15910 21902 -15876
rect 21936 -15910 21955 -15876
rect 21883 -15966 21955 -15910
rect 21883 -16000 21902 -15966
rect 21936 -16000 21955 -15966
rect 21883 -16056 21955 -16000
rect 21883 -16090 21902 -16056
rect 21936 -16090 21955 -16056
rect 21883 -16146 21955 -16090
rect 21883 -16180 21902 -16146
rect 21936 -16180 21955 -16146
rect 22773 -15494 22792 -15460
rect 22826 -15494 22845 -15460
rect 22773 -15550 22845 -15494
rect 22773 -15584 22792 -15550
rect 22826 -15584 22845 -15550
rect 22773 -15640 22845 -15584
rect 22773 -15674 22792 -15640
rect 22826 -15674 22845 -15640
rect 22773 -15730 22845 -15674
rect 22773 -15764 22792 -15730
rect 22826 -15764 22845 -15730
rect 22773 -15820 22845 -15764
rect 22773 -15854 22792 -15820
rect 22826 -15854 22845 -15820
rect 22773 -15910 22845 -15854
rect 22773 -15944 22792 -15910
rect 22826 -15944 22845 -15910
rect 22773 -16000 22845 -15944
rect 22773 -16034 22792 -16000
rect 22826 -16034 22845 -16000
rect 22773 -16090 22845 -16034
rect 22773 -16124 22792 -16090
rect 22826 -16124 22845 -16090
rect 21883 -16219 21955 -16180
rect 22773 -16180 22845 -16124
rect 22773 -16214 22792 -16180
rect 22826 -16214 22845 -16180
rect 22773 -16219 22845 -16214
rect 21883 -16238 22845 -16219
rect 21883 -16272 21996 -16238
rect 22030 -16272 22086 -16238
rect 22120 -16272 22176 -16238
rect 22210 -16272 22266 -16238
rect 22300 -16272 22356 -16238
rect 22390 -16272 22446 -16238
rect 22480 -16272 22536 -16238
rect 22570 -16272 22626 -16238
rect 22660 -16272 22716 -16238
rect 22750 -16272 22845 -16238
rect 21883 -16291 22845 -16272
rect 23171 -15348 24133 -15329
rect 23171 -15382 23303 -15348
rect 23337 -15382 23393 -15348
rect 23427 -15382 23483 -15348
rect 23517 -15382 23573 -15348
rect 23607 -15382 23663 -15348
rect 23697 -15382 23753 -15348
rect 23787 -15382 23843 -15348
rect 23877 -15382 23933 -15348
rect 23967 -15382 24023 -15348
rect 24057 -15382 24133 -15348
rect 23171 -15401 24133 -15382
rect 23171 -15426 23243 -15401
rect 23171 -15460 23190 -15426
rect 23224 -15460 23243 -15426
rect 23171 -15516 23243 -15460
rect 24061 -15460 24133 -15401
rect 23171 -15550 23190 -15516
rect 23224 -15550 23243 -15516
rect 23171 -15606 23243 -15550
rect 23171 -15640 23190 -15606
rect 23224 -15640 23243 -15606
rect 23171 -15696 23243 -15640
rect 23171 -15730 23190 -15696
rect 23224 -15730 23243 -15696
rect 23171 -15786 23243 -15730
rect 23171 -15820 23190 -15786
rect 23224 -15820 23243 -15786
rect 23171 -15876 23243 -15820
rect 23171 -15910 23190 -15876
rect 23224 -15910 23243 -15876
rect 23171 -15966 23243 -15910
rect 23171 -16000 23190 -15966
rect 23224 -16000 23243 -15966
rect 23171 -16056 23243 -16000
rect 23171 -16090 23190 -16056
rect 23224 -16090 23243 -16056
rect 23171 -16146 23243 -16090
rect 23171 -16180 23190 -16146
rect 23224 -16180 23243 -16146
rect 24061 -15494 24080 -15460
rect 24114 -15494 24133 -15460
rect 24061 -15550 24133 -15494
rect 24061 -15584 24080 -15550
rect 24114 -15584 24133 -15550
rect 24061 -15640 24133 -15584
rect 24061 -15674 24080 -15640
rect 24114 -15674 24133 -15640
rect 24061 -15730 24133 -15674
rect 24061 -15764 24080 -15730
rect 24114 -15764 24133 -15730
rect 24061 -15820 24133 -15764
rect 24061 -15854 24080 -15820
rect 24114 -15854 24133 -15820
rect 24061 -15910 24133 -15854
rect 24061 -15944 24080 -15910
rect 24114 -15944 24133 -15910
rect 24061 -16000 24133 -15944
rect 24061 -16034 24080 -16000
rect 24114 -16034 24133 -16000
rect 24061 -16090 24133 -16034
rect 24061 -16124 24080 -16090
rect 24114 -16124 24133 -16090
rect 23171 -16219 23243 -16180
rect 24061 -16180 24133 -16124
rect 24061 -16214 24080 -16180
rect 24114 -16214 24133 -16180
rect 24061 -16219 24133 -16214
rect 23171 -16238 24133 -16219
rect 23171 -16272 23284 -16238
rect 23318 -16272 23374 -16238
rect 23408 -16272 23464 -16238
rect 23498 -16272 23554 -16238
rect 23588 -16272 23644 -16238
rect 23678 -16272 23734 -16238
rect 23768 -16272 23824 -16238
rect 23858 -16272 23914 -16238
rect 23948 -16272 24004 -16238
rect 24038 -16272 24133 -16238
rect 23171 -16291 24133 -16272
rect 24459 -15348 25421 -15329
rect 24459 -15382 24591 -15348
rect 24625 -15382 24681 -15348
rect 24715 -15382 24771 -15348
rect 24805 -15382 24861 -15348
rect 24895 -15382 24951 -15348
rect 24985 -15382 25041 -15348
rect 25075 -15382 25131 -15348
rect 25165 -15382 25221 -15348
rect 25255 -15382 25311 -15348
rect 25345 -15382 25421 -15348
rect 24459 -15401 25421 -15382
rect 24459 -15426 24531 -15401
rect 24459 -15460 24478 -15426
rect 24512 -15460 24531 -15426
rect 24459 -15516 24531 -15460
rect 25349 -15460 25421 -15401
rect 24459 -15550 24478 -15516
rect 24512 -15550 24531 -15516
rect 24459 -15606 24531 -15550
rect 24459 -15640 24478 -15606
rect 24512 -15640 24531 -15606
rect 24459 -15696 24531 -15640
rect 24459 -15730 24478 -15696
rect 24512 -15730 24531 -15696
rect 24459 -15786 24531 -15730
rect 24459 -15820 24478 -15786
rect 24512 -15820 24531 -15786
rect 24459 -15876 24531 -15820
rect 24459 -15910 24478 -15876
rect 24512 -15910 24531 -15876
rect 24459 -15966 24531 -15910
rect 24459 -16000 24478 -15966
rect 24512 -16000 24531 -15966
rect 24459 -16056 24531 -16000
rect 24459 -16090 24478 -16056
rect 24512 -16090 24531 -16056
rect 24459 -16146 24531 -16090
rect 24459 -16180 24478 -16146
rect 24512 -16180 24531 -16146
rect 25349 -15494 25368 -15460
rect 25402 -15494 25421 -15460
rect 25349 -15550 25421 -15494
rect 25349 -15584 25368 -15550
rect 25402 -15584 25421 -15550
rect 25349 -15640 25421 -15584
rect 25349 -15674 25368 -15640
rect 25402 -15674 25421 -15640
rect 25349 -15730 25421 -15674
rect 25349 -15764 25368 -15730
rect 25402 -15764 25421 -15730
rect 25349 -15820 25421 -15764
rect 25349 -15854 25368 -15820
rect 25402 -15854 25421 -15820
rect 25349 -15910 25421 -15854
rect 25349 -15944 25368 -15910
rect 25402 -15944 25421 -15910
rect 25349 -16000 25421 -15944
rect 25349 -16034 25368 -16000
rect 25402 -16034 25421 -16000
rect 25349 -16090 25421 -16034
rect 25349 -16124 25368 -16090
rect 25402 -16124 25421 -16090
rect 24459 -16219 24531 -16180
rect 25349 -16180 25421 -16124
rect 25349 -16214 25368 -16180
rect 25402 -16214 25421 -16180
rect 25349 -16219 25421 -16214
rect 24459 -16238 25421 -16219
rect 24459 -16272 24572 -16238
rect 24606 -16272 24662 -16238
rect 24696 -16272 24752 -16238
rect 24786 -16272 24842 -16238
rect 24876 -16272 24932 -16238
rect 24966 -16272 25022 -16238
rect 25056 -16272 25112 -16238
rect 25146 -16272 25202 -16238
rect 25236 -16272 25292 -16238
rect 25326 -16272 25421 -16238
rect 24459 -16291 25421 -16272
rect 25747 -15348 26709 -15329
rect 25747 -15382 25879 -15348
rect 25913 -15382 25969 -15348
rect 26003 -15382 26059 -15348
rect 26093 -15382 26149 -15348
rect 26183 -15382 26239 -15348
rect 26273 -15382 26329 -15348
rect 26363 -15382 26419 -15348
rect 26453 -15382 26509 -15348
rect 26543 -15382 26599 -15348
rect 26633 -15382 26709 -15348
rect 25747 -15401 26709 -15382
rect 25747 -15426 25819 -15401
rect 25747 -15460 25766 -15426
rect 25800 -15460 25819 -15426
rect 25747 -15516 25819 -15460
rect 26637 -15460 26709 -15401
rect 25747 -15550 25766 -15516
rect 25800 -15550 25819 -15516
rect 25747 -15606 25819 -15550
rect 25747 -15640 25766 -15606
rect 25800 -15640 25819 -15606
rect 25747 -15696 25819 -15640
rect 25747 -15730 25766 -15696
rect 25800 -15730 25819 -15696
rect 25747 -15786 25819 -15730
rect 25747 -15820 25766 -15786
rect 25800 -15820 25819 -15786
rect 25747 -15876 25819 -15820
rect 25747 -15910 25766 -15876
rect 25800 -15910 25819 -15876
rect 25747 -15966 25819 -15910
rect 25747 -16000 25766 -15966
rect 25800 -16000 25819 -15966
rect 25747 -16056 25819 -16000
rect 25747 -16090 25766 -16056
rect 25800 -16090 25819 -16056
rect 25747 -16146 25819 -16090
rect 25747 -16180 25766 -16146
rect 25800 -16180 25819 -16146
rect 26637 -15494 26656 -15460
rect 26690 -15494 26709 -15460
rect 26637 -15550 26709 -15494
rect 26637 -15584 26656 -15550
rect 26690 -15584 26709 -15550
rect 26637 -15640 26709 -15584
rect 26637 -15674 26656 -15640
rect 26690 -15674 26709 -15640
rect 26637 -15730 26709 -15674
rect 26637 -15764 26656 -15730
rect 26690 -15764 26709 -15730
rect 26637 -15820 26709 -15764
rect 26637 -15854 26656 -15820
rect 26690 -15854 26709 -15820
rect 26637 -15910 26709 -15854
rect 26637 -15944 26656 -15910
rect 26690 -15944 26709 -15910
rect 26637 -16000 26709 -15944
rect 26637 -16034 26656 -16000
rect 26690 -16034 26709 -16000
rect 26637 -16090 26709 -16034
rect 26637 -16124 26656 -16090
rect 26690 -16124 26709 -16090
rect 25747 -16219 25819 -16180
rect 26637 -16180 26709 -16124
rect 26637 -16214 26656 -16180
rect 26690 -16214 26709 -16180
rect 26637 -16219 26709 -16214
rect 25747 -16238 26709 -16219
rect 25747 -16272 25860 -16238
rect 25894 -16272 25950 -16238
rect 25984 -16272 26040 -16238
rect 26074 -16272 26130 -16238
rect 26164 -16272 26220 -16238
rect 26254 -16272 26310 -16238
rect 26344 -16272 26400 -16238
rect 26434 -16272 26490 -16238
rect 26524 -16272 26580 -16238
rect 26614 -16272 26709 -16238
rect 25747 -16291 26709 -16272
rect 16731 -16636 17693 -16617
rect 16731 -16670 16863 -16636
rect 16897 -16670 16953 -16636
rect 16987 -16670 17043 -16636
rect 17077 -16670 17133 -16636
rect 17167 -16670 17223 -16636
rect 17257 -16670 17313 -16636
rect 17347 -16670 17403 -16636
rect 17437 -16670 17493 -16636
rect 17527 -16670 17583 -16636
rect 17617 -16670 17693 -16636
rect 16731 -16689 17693 -16670
rect 16731 -16714 16803 -16689
rect 16731 -16748 16750 -16714
rect 16784 -16748 16803 -16714
rect 16731 -16804 16803 -16748
rect 17621 -16748 17693 -16689
rect 16731 -16838 16750 -16804
rect 16784 -16838 16803 -16804
rect 16731 -16894 16803 -16838
rect 16731 -16928 16750 -16894
rect 16784 -16928 16803 -16894
rect 16731 -16984 16803 -16928
rect 16731 -17018 16750 -16984
rect 16784 -17018 16803 -16984
rect 16731 -17074 16803 -17018
rect 16731 -17108 16750 -17074
rect 16784 -17108 16803 -17074
rect 16731 -17164 16803 -17108
rect 16731 -17198 16750 -17164
rect 16784 -17198 16803 -17164
rect 16731 -17254 16803 -17198
rect 16731 -17288 16750 -17254
rect 16784 -17288 16803 -17254
rect 16731 -17344 16803 -17288
rect 16731 -17378 16750 -17344
rect 16784 -17378 16803 -17344
rect 16731 -17434 16803 -17378
rect 16731 -17468 16750 -17434
rect 16784 -17468 16803 -17434
rect 17621 -16782 17640 -16748
rect 17674 -16782 17693 -16748
rect 17621 -16838 17693 -16782
rect 17621 -16872 17640 -16838
rect 17674 -16872 17693 -16838
rect 17621 -16928 17693 -16872
rect 17621 -16962 17640 -16928
rect 17674 -16962 17693 -16928
rect 17621 -17018 17693 -16962
rect 17621 -17052 17640 -17018
rect 17674 -17052 17693 -17018
rect 17621 -17108 17693 -17052
rect 17621 -17142 17640 -17108
rect 17674 -17142 17693 -17108
rect 17621 -17198 17693 -17142
rect 17621 -17232 17640 -17198
rect 17674 -17232 17693 -17198
rect 17621 -17288 17693 -17232
rect 17621 -17322 17640 -17288
rect 17674 -17322 17693 -17288
rect 17621 -17378 17693 -17322
rect 17621 -17412 17640 -17378
rect 17674 -17412 17693 -17378
rect 16731 -17507 16803 -17468
rect 17621 -17468 17693 -17412
rect 17621 -17502 17640 -17468
rect 17674 -17502 17693 -17468
rect 17621 -17507 17693 -17502
rect 16731 -17526 17693 -17507
rect 16731 -17560 16844 -17526
rect 16878 -17560 16934 -17526
rect 16968 -17560 17024 -17526
rect 17058 -17560 17114 -17526
rect 17148 -17560 17204 -17526
rect 17238 -17560 17294 -17526
rect 17328 -17560 17384 -17526
rect 17418 -17560 17474 -17526
rect 17508 -17560 17564 -17526
rect 17598 -17560 17693 -17526
rect 16731 -17579 17693 -17560
rect 18019 -16636 18981 -16617
rect 18019 -16670 18151 -16636
rect 18185 -16670 18241 -16636
rect 18275 -16670 18331 -16636
rect 18365 -16670 18421 -16636
rect 18455 -16670 18511 -16636
rect 18545 -16670 18601 -16636
rect 18635 -16670 18691 -16636
rect 18725 -16670 18781 -16636
rect 18815 -16670 18871 -16636
rect 18905 -16670 18981 -16636
rect 18019 -16689 18981 -16670
rect 18019 -16714 18091 -16689
rect 18019 -16748 18038 -16714
rect 18072 -16748 18091 -16714
rect 18019 -16804 18091 -16748
rect 18909 -16748 18981 -16689
rect 18019 -16838 18038 -16804
rect 18072 -16838 18091 -16804
rect 18019 -16894 18091 -16838
rect 18019 -16928 18038 -16894
rect 18072 -16928 18091 -16894
rect 18019 -16984 18091 -16928
rect 18019 -17018 18038 -16984
rect 18072 -17018 18091 -16984
rect 18019 -17074 18091 -17018
rect 18019 -17108 18038 -17074
rect 18072 -17108 18091 -17074
rect 18019 -17164 18091 -17108
rect 18019 -17198 18038 -17164
rect 18072 -17198 18091 -17164
rect 18019 -17254 18091 -17198
rect 18019 -17288 18038 -17254
rect 18072 -17288 18091 -17254
rect 18019 -17344 18091 -17288
rect 18019 -17378 18038 -17344
rect 18072 -17378 18091 -17344
rect 18019 -17434 18091 -17378
rect 18019 -17468 18038 -17434
rect 18072 -17468 18091 -17434
rect 18909 -16782 18928 -16748
rect 18962 -16782 18981 -16748
rect 18909 -16838 18981 -16782
rect 18909 -16872 18928 -16838
rect 18962 -16872 18981 -16838
rect 18909 -16928 18981 -16872
rect 18909 -16962 18928 -16928
rect 18962 -16962 18981 -16928
rect 18909 -17018 18981 -16962
rect 18909 -17052 18928 -17018
rect 18962 -17052 18981 -17018
rect 18909 -17108 18981 -17052
rect 18909 -17142 18928 -17108
rect 18962 -17142 18981 -17108
rect 18909 -17198 18981 -17142
rect 18909 -17232 18928 -17198
rect 18962 -17232 18981 -17198
rect 18909 -17288 18981 -17232
rect 18909 -17322 18928 -17288
rect 18962 -17322 18981 -17288
rect 18909 -17378 18981 -17322
rect 18909 -17412 18928 -17378
rect 18962 -17412 18981 -17378
rect 18019 -17507 18091 -17468
rect 18909 -17468 18981 -17412
rect 18909 -17502 18928 -17468
rect 18962 -17502 18981 -17468
rect 18909 -17507 18981 -17502
rect 18019 -17526 18981 -17507
rect 18019 -17560 18132 -17526
rect 18166 -17560 18222 -17526
rect 18256 -17560 18312 -17526
rect 18346 -17560 18402 -17526
rect 18436 -17560 18492 -17526
rect 18526 -17560 18582 -17526
rect 18616 -17560 18672 -17526
rect 18706 -17560 18762 -17526
rect 18796 -17560 18852 -17526
rect 18886 -17560 18981 -17526
rect 18019 -17579 18981 -17560
rect 19307 -16636 20269 -16617
rect 19307 -16670 19439 -16636
rect 19473 -16670 19529 -16636
rect 19563 -16670 19619 -16636
rect 19653 -16670 19709 -16636
rect 19743 -16670 19799 -16636
rect 19833 -16670 19889 -16636
rect 19923 -16670 19979 -16636
rect 20013 -16670 20069 -16636
rect 20103 -16670 20159 -16636
rect 20193 -16670 20269 -16636
rect 19307 -16689 20269 -16670
rect 19307 -16714 19379 -16689
rect 19307 -16748 19326 -16714
rect 19360 -16748 19379 -16714
rect 19307 -16804 19379 -16748
rect 20197 -16748 20269 -16689
rect 19307 -16838 19326 -16804
rect 19360 -16838 19379 -16804
rect 19307 -16894 19379 -16838
rect 19307 -16928 19326 -16894
rect 19360 -16928 19379 -16894
rect 19307 -16984 19379 -16928
rect 19307 -17018 19326 -16984
rect 19360 -17018 19379 -16984
rect 19307 -17074 19379 -17018
rect 19307 -17108 19326 -17074
rect 19360 -17108 19379 -17074
rect 19307 -17164 19379 -17108
rect 19307 -17198 19326 -17164
rect 19360 -17198 19379 -17164
rect 19307 -17254 19379 -17198
rect 19307 -17288 19326 -17254
rect 19360 -17288 19379 -17254
rect 19307 -17344 19379 -17288
rect 19307 -17378 19326 -17344
rect 19360 -17378 19379 -17344
rect 19307 -17434 19379 -17378
rect 19307 -17468 19326 -17434
rect 19360 -17468 19379 -17434
rect 20197 -16782 20216 -16748
rect 20250 -16782 20269 -16748
rect 20197 -16838 20269 -16782
rect 20197 -16872 20216 -16838
rect 20250 -16872 20269 -16838
rect 20197 -16928 20269 -16872
rect 20197 -16962 20216 -16928
rect 20250 -16962 20269 -16928
rect 20197 -17018 20269 -16962
rect 20197 -17052 20216 -17018
rect 20250 -17052 20269 -17018
rect 20197 -17108 20269 -17052
rect 20197 -17142 20216 -17108
rect 20250 -17142 20269 -17108
rect 20197 -17198 20269 -17142
rect 20197 -17232 20216 -17198
rect 20250 -17232 20269 -17198
rect 20197 -17288 20269 -17232
rect 20197 -17322 20216 -17288
rect 20250 -17322 20269 -17288
rect 20197 -17378 20269 -17322
rect 20197 -17412 20216 -17378
rect 20250 -17412 20269 -17378
rect 19307 -17507 19379 -17468
rect 20197 -17468 20269 -17412
rect 20197 -17502 20216 -17468
rect 20250 -17502 20269 -17468
rect 20197 -17507 20269 -17502
rect 19307 -17526 20269 -17507
rect 19307 -17560 19420 -17526
rect 19454 -17560 19510 -17526
rect 19544 -17560 19600 -17526
rect 19634 -17560 19690 -17526
rect 19724 -17560 19780 -17526
rect 19814 -17560 19870 -17526
rect 19904 -17560 19960 -17526
rect 19994 -17560 20050 -17526
rect 20084 -17560 20140 -17526
rect 20174 -17560 20269 -17526
rect 19307 -17579 20269 -17560
rect 20595 -16636 21557 -16617
rect 20595 -16670 20727 -16636
rect 20761 -16670 20817 -16636
rect 20851 -16670 20907 -16636
rect 20941 -16670 20997 -16636
rect 21031 -16670 21087 -16636
rect 21121 -16670 21177 -16636
rect 21211 -16670 21267 -16636
rect 21301 -16670 21357 -16636
rect 21391 -16670 21447 -16636
rect 21481 -16670 21557 -16636
rect 20595 -16689 21557 -16670
rect 20595 -16714 20667 -16689
rect 20595 -16748 20614 -16714
rect 20648 -16748 20667 -16714
rect 20595 -16804 20667 -16748
rect 21485 -16748 21557 -16689
rect 20595 -16838 20614 -16804
rect 20648 -16838 20667 -16804
rect 20595 -16894 20667 -16838
rect 20595 -16928 20614 -16894
rect 20648 -16928 20667 -16894
rect 20595 -16984 20667 -16928
rect 20595 -17018 20614 -16984
rect 20648 -17018 20667 -16984
rect 20595 -17074 20667 -17018
rect 20595 -17108 20614 -17074
rect 20648 -17108 20667 -17074
rect 20595 -17164 20667 -17108
rect 20595 -17198 20614 -17164
rect 20648 -17198 20667 -17164
rect 20595 -17254 20667 -17198
rect 20595 -17288 20614 -17254
rect 20648 -17288 20667 -17254
rect 20595 -17344 20667 -17288
rect 20595 -17378 20614 -17344
rect 20648 -17378 20667 -17344
rect 20595 -17434 20667 -17378
rect 20595 -17468 20614 -17434
rect 20648 -17468 20667 -17434
rect 21485 -16782 21504 -16748
rect 21538 -16782 21557 -16748
rect 21485 -16838 21557 -16782
rect 21485 -16872 21504 -16838
rect 21538 -16872 21557 -16838
rect 21485 -16928 21557 -16872
rect 21485 -16962 21504 -16928
rect 21538 -16962 21557 -16928
rect 21485 -17018 21557 -16962
rect 21485 -17052 21504 -17018
rect 21538 -17052 21557 -17018
rect 21485 -17108 21557 -17052
rect 21485 -17142 21504 -17108
rect 21538 -17142 21557 -17108
rect 21485 -17198 21557 -17142
rect 21485 -17232 21504 -17198
rect 21538 -17232 21557 -17198
rect 21485 -17288 21557 -17232
rect 21485 -17322 21504 -17288
rect 21538 -17322 21557 -17288
rect 21485 -17378 21557 -17322
rect 21485 -17412 21504 -17378
rect 21538 -17412 21557 -17378
rect 20595 -17507 20667 -17468
rect 21485 -17468 21557 -17412
rect 21485 -17502 21504 -17468
rect 21538 -17502 21557 -17468
rect 21485 -17507 21557 -17502
rect 20595 -17526 21557 -17507
rect 20595 -17560 20708 -17526
rect 20742 -17560 20798 -17526
rect 20832 -17560 20888 -17526
rect 20922 -17560 20978 -17526
rect 21012 -17560 21068 -17526
rect 21102 -17560 21158 -17526
rect 21192 -17560 21248 -17526
rect 21282 -17560 21338 -17526
rect 21372 -17560 21428 -17526
rect 21462 -17560 21557 -17526
rect 20595 -17579 21557 -17560
rect 21883 -16636 22845 -16617
rect 21883 -16670 22015 -16636
rect 22049 -16670 22105 -16636
rect 22139 -16670 22195 -16636
rect 22229 -16670 22285 -16636
rect 22319 -16670 22375 -16636
rect 22409 -16670 22465 -16636
rect 22499 -16670 22555 -16636
rect 22589 -16670 22645 -16636
rect 22679 -16670 22735 -16636
rect 22769 -16670 22845 -16636
rect 21883 -16689 22845 -16670
rect 21883 -16714 21955 -16689
rect 21883 -16748 21902 -16714
rect 21936 -16748 21955 -16714
rect 21883 -16804 21955 -16748
rect 22773 -16748 22845 -16689
rect 21883 -16838 21902 -16804
rect 21936 -16838 21955 -16804
rect 21883 -16894 21955 -16838
rect 21883 -16928 21902 -16894
rect 21936 -16928 21955 -16894
rect 21883 -16984 21955 -16928
rect 21883 -17018 21902 -16984
rect 21936 -17018 21955 -16984
rect 21883 -17074 21955 -17018
rect 21883 -17108 21902 -17074
rect 21936 -17108 21955 -17074
rect 21883 -17164 21955 -17108
rect 21883 -17198 21902 -17164
rect 21936 -17198 21955 -17164
rect 21883 -17254 21955 -17198
rect 21883 -17288 21902 -17254
rect 21936 -17288 21955 -17254
rect 21883 -17344 21955 -17288
rect 21883 -17378 21902 -17344
rect 21936 -17378 21955 -17344
rect 21883 -17434 21955 -17378
rect 21883 -17468 21902 -17434
rect 21936 -17468 21955 -17434
rect 22773 -16782 22792 -16748
rect 22826 -16782 22845 -16748
rect 22773 -16838 22845 -16782
rect 22773 -16872 22792 -16838
rect 22826 -16872 22845 -16838
rect 22773 -16928 22845 -16872
rect 22773 -16962 22792 -16928
rect 22826 -16962 22845 -16928
rect 22773 -17018 22845 -16962
rect 22773 -17052 22792 -17018
rect 22826 -17052 22845 -17018
rect 22773 -17108 22845 -17052
rect 22773 -17142 22792 -17108
rect 22826 -17142 22845 -17108
rect 22773 -17198 22845 -17142
rect 22773 -17232 22792 -17198
rect 22826 -17232 22845 -17198
rect 22773 -17288 22845 -17232
rect 22773 -17322 22792 -17288
rect 22826 -17322 22845 -17288
rect 22773 -17378 22845 -17322
rect 22773 -17412 22792 -17378
rect 22826 -17412 22845 -17378
rect 21883 -17507 21955 -17468
rect 22773 -17468 22845 -17412
rect 22773 -17502 22792 -17468
rect 22826 -17502 22845 -17468
rect 22773 -17507 22845 -17502
rect 21883 -17526 22845 -17507
rect 21883 -17560 21996 -17526
rect 22030 -17560 22086 -17526
rect 22120 -17560 22176 -17526
rect 22210 -17560 22266 -17526
rect 22300 -17560 22356 -17526
rect 22390 -17560 22446 -17526
rect 22480 -17560 22536 -17526
rect 22570 -17560 22626 -17526
rect 22660 -17560 22716 -17526
rect 22750 -17560 22845 -17526
rect 21883 -17579 22845 -17560
rect 23171 -16636 24133 -16617
rect 23171 -16670 23303 -16636
rect 23337 -16670 23393 -16636
rect 23427 -16670 23483 -16636
rect 23517 -16670 23573 -16636
rect 23607 -16670 23663 -16636
rect 23697 -16670 23753 -16636
rect 23787 -16670 23843 -16636
rect 23877 -16670 23933 -16636
rect 23967 -16670 24023 -16636
rect 24057 -16670 24133 -16636
rect 23171 -16689 24133 -16670
rect 23171 -16714 23243 -16689
rect 23171 -16748 23190 -16714
rect 23224 -16748 23243 -16714
rect 23171 -16804 23243 -16748
rect 24061 -16748 24133 -16689
rect 23171 -16838 23190 -16804
rect 23224 -16838 23243 -16804
rect 23171 -16894 23243 -16838
rect 23171 -16928 23190 -16894
rect 23224 -16928 23243 -16894
rect 23171 -16984 23243 -16928
rect 23171 -17018 23190 -16984
rect 23224 -17018 23243 -16984
rect 23171 -17074 23243 -17018
rect 23171 -17108 23190 -17074
rect 23224 -17108 23243 -17074
rect 23171 -17164 23243 -17108
rect 23171 -17198 23190 -17164
rect 23224 -17198 23243 -17164
rect 23171 -17254 23243 -17198
rect 23171 -17288 23190 -17254
rect 23224 -17288 23243 -17254
rect 23171 -17344 23243 -17288
rect 23171 -17378 23190 -17344
rect 23224 -17378 23243 -17344
rect 23171 -17434 23243 -17378
rect 23171 -17468 23190 -17434
rect 23224 -17468 23243 -17434
rect 24061 -16782 24080 -16748
rect 24114 -16782 24133 -16748
rect 24061 -16838 24133 -16782
rect 24061 -16872 24080 -16838
rect 24114 -16872 24133 -16838
rect 24061 -16928 24133 -16872
rect 24061 -16962 24080 -16928
rect 24114 -16962 24133 -16928
rect 24061 -17018 24133 -16962
rect 24061 -17052 24080 -17018
rect 24114 -17052 24133 -17018
rect 24061 -17108 24133 -17052
rect 24061 -17142 24080 -17108
rect 24114 -17142 24133 -17108
rect 24061 -17198 24133 -17142
rect 24061 -17232 24080 -17198
rect 24114 -17232 24133 -17198
rect 24061 -17288 24133 -17232
rect 24061 -17322 24080 -17288
rect 24114 -17322 24133 -17288
rect 24061 -17378 24133 -17322
rect 24061 -17412 24080 -17378
rect 24114 -17412 24133 -17378
rect 23171 -17507 23243 -17468
rect 24061 -17468 24133 -17412
rect 24061 -17502 24080 -17468
rect 24114 -17502 24133 -17468
rect 24061 -17507 24133 -17502
rect 23171 -17526 24133 -17507
rect 23171 -17560 23284 -17526
rect 23318 -17560 23374 -17526
rect 23408 -17560 23464 -17526
rect 23498 -17560 23554 -17526
rect 23588 -17560 23644 -17526
rect 23678 -17560 23734 -17526
rect 23768 -17560 23824 -17526
rect 23858 -17560 23914 -17526
rect 23948 -17560 24004 -17526
rect 24038 -17560 24133 -17526
rect 23171 -17579 24133 -17560
rect 24459 -16636 25421 -16617
rect 24459 -16670 24591 -16636
rect 24625 -16670 24681 -16636
rect 24715 -16670 24771 -16636
rect 24805 -16670 24861 -16636
rect 24895 -16670 24951 -16636
rect 24985 -16670 25041 -16636
rect 25075 -16670 25131 -16636
rect 25165 -16670 25221 -16636
rect 25255 -16670 25311 -16636
rect 25345 -16670 25421 -16636
rect 24459 -16689 25421 -16670
rect 24459 -16714 24531 -16689
rect 24459 -16748 24478 -16714
rect 24512 -16748 24531 -16714
rect 24459 -16804 24531 -16748
rect 25349 -16748 25421 -16689
rect 24459 -16838 24478 -16804
rect 24512 -16838 24531 -16804
rect 24459 -16894 24531 -16838
rect 24459 -16928 24478 -16894
rect 24512 -16928 24531 -16894
rect 24459 -16984 24531 -16928
rect 24459 -17018 24478 -16984
rect 24512 -17018 24531 -16984
rect 24459 -17074 24531 -17018
rect 24459 -17108 24478 -17074
rect 24512 -17108 24531 -17074
rect 24459 -17164 24531 -17108
rect 24459 -17198 24478 -17164
rect 24512 -17198 24531 -17164
rect 24459 -17254 24531 -17198
rect 24459 -17288 24478 -17254
rect 24512 -17288 24531 -17254
rect 24459 -17344 24531 -17288
rect 24459 -17378 24478 -17344
rect 24512 -17378 24531 -17344
rect 24459 -17434 24531 -17378
rect 24459 -17468 24478 -17434
rect 24512 -17468 24531 -17434
rect 25349 -16782 25368 -16748
rect 25402 -16782 25421 -16748
rect 25349 -16838 25421 -16782
rect 25349 -16872 25368 -16838
rect 25402 -16872 25421 -16838
rect 25349 -16928 25421 -16872
rect 25349 -16962 25368 -16928
rect 25402 -16962 25421 -16928
rect 25349 -17018 25421 -16962
rect 25349 -17052 25368 -17018
rect 25402 -17052 25421 -17018
rect 25349 -17108 25421 -17052
rect 25349 -17142 25368 -17108
rect 25402 -17142 25421 -17108
rect 25349 -17198 25421 -17142
rect 25349 -17232 25368 -17198
rect 25402 -17232 25421 -17198
rect 25349 -17288 25421 -17232
rect 25349 -17322 25368 -17288
rect 25402 -17322 25421 -17288
rect 25349 -17378 25421 -17322
rect 25349 -17412 25368 -17378
rect 25402 -17412 25421 -17378
rect 24459 -17507 24531 -17468
rect 25349 -17468 25421 -17412
rect 25349 -17502 25368 -17468
rect 25402 -17502 25421 -17468
rect 25349 -17507 25421 -17502
rect 24459 -17526 25421 -17507
rect 24459 -17560 24572 -17526
rect 24606 -17560 24662 -17526
rect 24696 -17560 24752 -17526
rect 24786 -17560 24842 -17526
rect 24876 -17560 24932 -17526
rect 24966 -17560 25022 -17526
rect 25056 -17560 25112 -17526
rect 25146 -17560 25202 -17526
rect 25236 -17560 25292 -17526
rect 25326 -17560 25421 -17526
rect 24459 -17579 25421 -17560
rect 25747 -16636 26709 -16617
rect 25747 -16670 25879 -16636
rect 25913 -16670 25969 -16636
rect 26003 -16670 26059 -16636
rect 26093 -16670 26149 -16636
rect 26183 -16670 26239 -16636
rect 26273 -16670 26329 -16636
rect 26363 -16670 26419 -16636
rect 26453 -16670 26509 -16636
rect 26543 -16670 26599 -16636
rect 26633 -16670 26709 -16636
rect 25747 -16689 26709 -16670
rect 25747 -16714 25819 -16689
rect 25747 -16748 25766 -16714
rect 25800 -16748 25819 -16714
rect 25747 -16804 25819 -16748
rect 26637 -16748 26709 -16689
rect 25747 -16838 25766 -16804
rect 25800 -16838 25819 -16804
rect 25747 -16894 25819 -16838
rect 25747 -16928 25766 -16894
rect 25800 -16928 25819 -16894
rect 25747 -16984 25819 -16928
rect 25747 -17018 25766 -16984
rect 25800 -17018 25819 -16984
rect 25747 -17074 25819 -17018
rect 25747 -17108 25766 -17074
rect 25800 -17108 25819 -17074
rect 25747 -17164 25819 -17108
rect 25747 -17198 25766 -17164
rect 25800 -17198 25819 -17164
rect 25747 -17254 25819 -17198
rect 25747 -17288 25766 -17254
rect 25800 -17288 25819 -17254
rect 25747 -17344 25819 -17288
rect 25747 -17378 25766 -17344
rect 25800 -17378 25819 -17344
rect 25747 -17434 25819 -17378
rect 25747 -17468 25766 -17434
rect 25800 -17468 25819 -17434
rect 26637 -16782 26656 -16748
rect 26690 -16782 26709 -16748
rect 26637 -16838 26709 -16782
rect 26637 -16872 26656 -16838
rect 26690 -16872 26709 -16838
rect 26637 -16928 26709 -16872
rect 26637 -16962 26656 -16928
rect 26690 -16962 26709 -16928
rect 26637 -17018 26709 -16962
rect 26637 -17052 26656 -17018
rect 26690 -17052 26709 -17018
rect 26637 -17108 26709 -17052
rect 26637 -17142 26656 -17108
rect 26690 -17142 26709 -17108
rect 26637 -17198 26709 -17142
rect 26637 -17232 26656 -17198
rect 26690 -17232 26709 -17198
rect 26637 -17288 26709 -17232
rect 26637 -17322 26656 -17288
rect 26690 -17322 26709 -17288
rect 26637 -17378 26709 -17322
rect 26637 -17412 26656 -17378
rect 26690 -17412 26709 -17378
rect 25747 -17507 25819 -17468
rect 26637 -17468 26709 -17412
rect 26637 -17502 26656 -17468
rect 26690 -17502 26709 -17468
rect 26637 -17507 26709 -17502
rect 25747 -17526 26709 -17507
rect 25747 -17560 25860 -17526
rect 25894 -17560 25950 -17526
rect 25984 -17560 26040 -17526
rect 26074 -17560 26130 -17526
rect 26164 -17560 26220 -17526
rect 26254 -17560 26310 -17526
rect 26344 -17560 26400 -17526
rect 26434 -17560 26490 -17526
rect 26524 -17560 26580 -17526
rect 26614 -17560 26709 -17526
rect 25747 -17579 26709 -17560
<< psubdiffcont >>
rect 16684 -11370 16718 -11336
rect 16774 -11370 16808 -11336
rect 16864 -11370 16898 -11336
rect 16954 -11370 16988 -11336
rect 17044 -11370 17078 -11336
rect 17134 -11370 17168 -11336
rect 17224 -11370 17258 -11336
rect 17314 -11370 17348 -11336
rect 17404 -11370 17438 -11336
rect 17494 -11370 17528 -11336
rect 17584 -11370 17618 -11336
rect 17674 -11370 17708 -11336
rect 17764 -11370 17798 -11336
rect 17972 -11370 18006 -11336
rect 18062 -11370 18096 -11336
rect 18152 -11370 18186 -11336
rect 18242 -11370 18276 -11336
rect 18332 -11370 18366 -11336
rect 18422 -11370 18456 -11336
rect 18512 -11370 18546 -11336
rect 18602 -11370 18636 -11336
rect 18692 -11370 18726 -11336
rect 18782 -11370 18816 -11336
rect 18872 -11370 18906 -11336
rect 18962 -11370 18996 -11336
rect 19052 -11370 19086 -11336
rect 19260 -11370 19294 -11336
rect 19350 -11370 19384 -11336
rect 19440 -11370 19474 -11336
rect 19530 -11370 19564 -11336
rect 19620 -11370 19654 -11336
rect 19710 -11370 19744 -11336
rect 19800 -11370 19834 -11336
rect 19890 -11370 19924 -11336
rect 19980 -11370 20014 -11336
rect 20070 -11370 20104 -11336
rect 20160 -11370 20194 -11336
rect 20250 -11370 20284 -11336
rect 20340 -11370 20374 -11336
rect 20548 -11370 20582 -11336
rect 20638 -11370 20672 -11336
rect 20728 -11370 20762 -11336
rect 20818 -11370 20852 -11336
rect 20908 -11370 20942 -11336
rect 20998 -11370 21032 -11336
rect 21088 -11370 21122 -11336
rect 21178 -11370 21212 -11336
rect 21268 -11370 21302 -11336
rect 21358 -11370 21392 -11336
rect 21448 -11370 21482 -11336
rect 21538 -11370 21572 -11336
rect 21628 -11370 21662 -11336
rect 21836 -11370 21870 -11336
rect 21926 -11370 21960 -11336
rect 22016 -11370 22050 -11336
rect 22106 -11370 22140 -11336
rect 22196 -11370 22230 -11336
rect 22286 -11370 22320 -11336
rect 22376 -11370 22410 -11336
rect 22466 -11370 22500 -11336
rect 22556 -11370 22590 -11336
rect 22646 -11370 22680 -11336
rect 22736 -11370 22770 -11336
rect 22826 -11370 22860 -11336
rect 22916 -11370 22950 -11336
rect 23124 -11370 23158 -11336
rect 23214 -11370 23248 -11336
rect 23304 -11370 23338 -11336
rect 23394 -11370 23428 -11336
rect 23484 -11370 23518 -11336
rect 23574 -11370 23608 -11336
rect 23664 -11370 23698 -11336
rect 23754 -11370 23788 -11336
rect 23844 -11370 23878 -11336
rect 23934 -11370 23968 -11336
rect 24024 -11370 24058 -11336
rect 24114 -11370 24148 -11336
rect 24204 -11370 24238 -11336
rect 24412 -11370 24446 -11336
rect 24502 -11370 24536 -11336
rect 24592 -11370 24626 -11336
rect 24682 -11370 24716 -11336
rect 24772 -11370 24806 -11336
rect 24862 -11370 24896 -11336
rect 24952 -11370 24986 -11336
rect 25042 -11370 25076 -11336
rect 25132 -11370 25166 -11336
rect 25222 -11370 25256 -11336
rect 25312 -11370 25346 -11336
rect 25402 -11370 25436 -11336
rect 25492 -11370 25526 -11336
rect 25700 -11370 25734 -11336
rect 25790 -11370 25824 -11336
rect 25880 -11370 25914 -11336
rect 25970 -11370 26004 -11336
rect 26060 -11370 26094 -11336
rect 26150 -11370 26184 -11336
rect 26240 -11370 26274 -11336
rect 26330 -11370 26364 -11336
rect 26420 -11370 26454 -11336
rect 26510 -11370 26544 -11336
rect 26600 -11370 26634 -11336
rect 26690 -11370 26724 -11336
rect 26780 -11370 26814 -11336
rect 16600 -11466 16634 -11432
rect 16600 -11556 16634 -11522
rect 16600 -11646 16634 -11612
rect 16600 -11736 16634 -11702
rect 16600 -11826 16634 -11792
rect 16600 -11916 16634 -11882
rect 16600 -12006 16634 -11972
rect 16600 -12096 16634 -12062
rect 16600 -12186 16634 -12152
rect 16600 -12276 16634 -12242
rect 16600 -12366 16634 -12332
rect 16600 -12456 16634 -12422
rect 17787 -11466 17821 -11432
rect 17888 -11466 17922 -11432
rect 17787 -11556 17821 -11522
rect 17888 -11556 17922 -11522
rect 17787 -11646 17821 -11612
rect 17888 -11646 17922 -11612
rect 17787 -11736 17821 -11702
rect 17888 -11736 17922 -11702
rect 17787 -11826 17821 -11792
rect 17888 -11826 17922 -11792
rect 17787 -11916 17821 -11882
rect 17888 -11916 17922 -11882
rect 17787 -12006 17821 -11972
rect 17888 -12006 17922 -11972
rect 17787 -12096 17821 -12062
rect 17888 -12096 17922 -12062
rect 17787 -12186 17821 -12152
rect 17888 -12186 17922 -12152
rect 17787 -12276 17821 -12242
rect 17888 -12276 17922 -12242
rect 17787 -12366 17821 -12332
rect 17888 -12366 17922 -12332
rect 17787 -12456 17821 -12422
rect 17888 -12456 17922 -12422
rect 19075 -11466 19109 -11432
rect 19176 -11466 19210 -11432
rect 19075 -11556 19109 -11522
rect 19176 -11556 19210 -11522
rect 19075 -11646 19109 -11612
rect 19176 -11646 19210 -11612
rect 19075 -11736 19109 -11702
rect 19176 -11736 19210 -11702
rect 19075 -11826 19109 -11792
rect 19176 -11826 19210 -11792
rect 19075 -11916 19109 -11882
rect 19176 -11916 19210 -11882
rect 19075 -12006 19109 -11972
rect 19176 -12006 19210 -11972
rect 19075 -12096 19109 -12062
rect 19176 -12096 19210 -12062
rect 19075 -12186 19109 -12152
rect 19176 -12186 19210 -12152
rect 19075 -12276 19109 -12242
rect 19176 -12276 19210 -12242
rect 19075 -12366 19109 -12332
rect 19176 -12366 19210 -12332
rect 19075 -12456 19109 -12422
rect 19176 -12456 19210 -12422
rect 20363 -11466 20397 -11432
rect 20464 -11466 20498 -11432
rect 20363 -11556 20397 -11522
rect 20464 -11556 20498 -11522
rect 20363 -11646 20397 -11612
rect 20464 -11646 20498 -11612
rect 20363 -11736 20397 -11702
rect 20464 -11736 20498 -11702
rect 20363 -11826 20397 -11792
rect 20464 -11826 20498 -11792
rect 20363 -11916 20397 -11882
rect 20464 -11916 20498 -11882
rect 20363 -12006 20397 -11972
rect 20464 -12006 20498 -11972
rect 20363 -12096 20397 -12062
rect 20464 -12096 20498 -12062
rect 20363 -12186 20397 -12152
rect 20464 -12186 20498 -12152
rect 20363 -12276 20397 -12242
rect 20464 -12276 20498 -12242
rect 20363 -12366 20397 -12332
rect 20464 -12366 20498 -12332
rect 20363 -12456 20397 -12422
rect 20464 -12456 20498 -12422
rect 21651 -11466 21685 -11432
rect 21752 -11466 21786 -11432
rect 21651 -11556 21685 -11522
rect 21752 -11556 21786 -11522
rect 21651 -11646 21685 -11612
rect 21752 -11646 21786 -11612
rect 21651 -11736 21685 -11702
rect 21752 -11736 21786 -11702
rect 21651 -11826 21685 -11792
rect 21752 -11826 21786 -11792
rect 21651 -11916 21685 -11882
rect 21752 -11916 21786 -11882
rect 21651 -12006 21685 -11972
rect 21752 -12006 21786 -11972
rect 21651 -12096 21685 -12062
rect 21752 -12096 21786 -12062
rect 21651 -12186 21685 -12152
rect 21752 -12186 21786 -12152
rect 21651 -12276 21685 -12242
rect 21752 -12276 21786 -12242
rect 21651 -12366 21685 -12332
rect 21752 -12366 21786 -12332
rect 21651 -12456 21685 -12422
rect 21752 -12456 21786 -12422
rect 22939 -11466 22973 -11432
rect 23040 -11466 23074 -11432
rect 22939 -11556 22973 -11522
rect 23040 -11556 23074 -11522
rect 22939 -11646 22973 -11612
rect 23040 -11646 23074 -11612
rect 22939 -11736 22973 -11702
rect 23040 -11736 23074 -11702
rect 22939 -11826 22973 -11792
rect 23040 -11826 23074 -11792
rect 22939 -11916 22973 -11882
rect 23040 -11916 23074 -11882
rect 22939 -12006 22973 -11972
rect 23040 -12006 23074 -11972
rect 22939 -12096 22973 -12062
rect 23040 -12096 23074 -12062
rect 22939 -12186 22973 -12152
rect 23040 -12186 23074 -12152
rect 22939 -12276 22973 -12242
rect 23040 -12276 23074 -12242
rect 22939 -12366 22973 -12332
rect 23040 -12366 23074 -12332
rect 22939 -12456 22973 -12422
rect 23040 -12456 23074 -12422
rect 24227 -11466 24261 -11432
rect 24328 -11466 24362 -11432
rect 24227 -11556 24261 -11522
rect 24328 -11556 24362 -11522
rect 24227 -11646 24261 -11612
rect 24328 -11646 24362 -11612
rect 24227 -11736 24261 -11702
rect 24328 -11736 24362 -11702
rect 24227 -11826 24261 -11792
rect 24328 -11826 24362 -11792
rect 24227 -11916 24261 -11882
rect 24328 -11916 24362 -11882
rect 24227 -12006 24261 -11972
rect 24328 -12006 24362 -11972
rect 24227 -12096 24261 -12062
rect 24328 -12096 24362 -12062
rect 24227 -12186 24261 -12152
rect 24328 -12186 24362 -12152
rect 24227 -12276 24261 -12242
rect 24328 -12276 24362 -12242
rect 24227 -12366 24261 -12332
rect 24328 -12366 24362 -12332
rect 24227 -12456 24261 -12422
rect 24328 -12456 24362 -12422
rect 25515 -11466 25549 -11432
rect 25616 -11466 25650 -11432
rect 25515 -11556 25549 -11522
rect 25616 -11556 25650 -11522
rect 25515 -11646 25549 -11612
rect 25616 -11646 25650 -11612
rect 25515 -11736 25549 -11702
rect 25616 -11736 25650 -11702
rect 25515 -11826 25549 -11792
rect 25616 -11826 25650 -11792
rect 25515 -11916 25549 -11882
rect 25616 -11916 25650 -11882
rect 25515 -12006 25549 -11972
rect 25616 -12006 25650 -11972
rect 25515 -12096 25549 -12062
rect 25616 -12096 25650 -12062
rect 25515 -12186 25549 -12152
rect 25616 -12186 25650 -12152
rect 25515 -12276 25549 -12242
rect 25616 -12276 25650 -12242
rect 25515 -12366 25549 -12332
rect 25616 -12366 25650 -12332
rect 25515 -12456 25549 -12422
rect 25616 -12456 25650 -12422
rect 26803 -11466 26837 -11432
rect 26803 -11556 26837 -11522
rect 26803 -11646 26837 -11612
rect 26803 -11736 26837 -11702
rect 26803 -11826 26837 -11792
rect 26803 -11916 26837 -11882
rect 26803 -12006 26837 -11972
rect 26803 -12096 26837 -12062
rect 26803 -12186 26837 -12152
rect 26803 -12276 26837 -12242
rect 26803 -12366 26837 -12332
rect 26803 -12456 26837 -12422
rect 16684 -12557 16718 -12523
rect 16774 -12557 16808 -12523
rect 16864 -12557 16898 -12523
rect 16954 -12557 16988 -12523
rect 17044 -12557 17078 -12523
rect 17134 -12557 17168 -12523
rect 17224 -12557 17258 -12523
rect 17314 -12557 17348 -12523
rect 17404 -12557 17438 -12523
rect 17494 -12557 17528 -12523
rect 17584 -12557 17618 -12523
rect 17674 -12557 17708 -12523
rect 17764 -12557 17798 -12523
rect 17972 -12557 18006 -12523
rect 18062 -12557 18096 -12523
rect 18152 -12557 18186 -12523
rect 18242 -12557 18276 -12523
rect 18332 -12557 18366 -12523
rect 18422 -12557 18456 -12523
rect 18512 -12557 18546 -12523
rect 18602 -12557 18636 -12523
rect 18692 -12557 18726 -12523
rect 18782 -12557 18816 -12523
rect 18872 -12557 18906 -12523
rect 18962 -12557 18996 -12523
rect 19052 -12557 19086 -12523
rect 19260 -12557 19294 -12523
rect 19350 -12557 19384 -12523
rect 19440 -12557 19474 -12523
rect 19530 -12557 19564 -12523
rect 19620 -12557 19654 -12523
rect 19710 -12557 19744 -12523
rect 19800 -12557 19834 -12523
rect 19890 -12557 19924 -12523
rect 19980 -12557 20014 -12523
rect 20070 -12557 20104 -12523
rect 20160 -12557 20194 -12523
rect 20250 -12557 20284 -12523
rect 20340 -12557 20374 -12523
rect 20548 -12557 20582 -12523
rect 20638 -12557 20672 -12523
rect 20728 -12557 20762 -12523
rect 20818 -12557 20852 -12523
rect 20908 -12557 20942 -12523
rect 20998 -12557 21032 -12523
rect 21088 -12557 21122 -12523
rect 21178 -12557 21212 -12523
rect 21268 -12557 21302 -12523
rect 21358 -12557 21392 -12523
rect 21448 -12557 21482 -12523
rect 21538 -12557 21572 -12523
rect 21628 -12557 21662 -12523
rect 21836 -12557 21870 -12523
rect 21926 -12557 21960 -12523
rect 22016 -12557 22050 -12523
rect 22106 -12557 22140 -12523
rect 22196 -12557 22230 -12523
rect 22286 -12557 22320 -12523
rect 22376 -12557 22410 -12523
rect 22466 -12557 22500 -12523
rect 22556 -12557 22590 -12523
rect 22646 -12557 22680 -12523
rect 22736 -12557 22770 -12523
rect 22826 -12557 22860 -12523
rect 22916 -12557 22950 -12523
rect 23124 -12557 23158 -12523
rect 23214 -12557 23248 -12523
rect 23304 -12557 23338 -12523
rect 23394 -12557 23428 -12523
rect 23484 -12557 23518 -12523
rect 23574 -12557 23608 -12523
rect 23664 -12557 23698 -12523
rect 23754 -12557 23788 -12523
rect 23844 -12557 23878 -12523
rect 23934 -12557 23968 -12523
rect 24024 -12557 24058 -12523
rect 24114 -12557 24148 -12523
rect 24204 -12557 24238 -12523
rect 24412 -12557 24446 -12523
rect 24502 -12557 24536 -12523
rect 24592 -12557 24626 -12523
rect 24682 -12557 24716 -12523
rect 24772 -12557 24806 -12523
rect 24862 -12557 24896 -12523
rect 24952 -12557 24986 -12523
rect 25042 -12557 25076 -12523
rect 25132 -12557 25166 -12523
rect 25222 -12557 25256 -12523
rect 25312 -12557 25346 -12523
rect 25402 -12557 25436 -12523
rect 25492 -12557 25526 -12523
rect 25700 -12557 25734 -12523
rect 25790 -12557 25824 -12523
rect 25880 -12557 25914 -12523
rect 25970 -12557 26004 -12523
rect 26060 -12557 26094 -12523
rect 26150 -12557 26184 -12523
rect 26240 -12557 26274 -12523
rect 26330 -12557 26364 -12523
rect 26420 -12557 26454 -12523
rect 26510 -12557 26544 -12523
rect 26600 -12557 26634 -12523
rect 26690 -12557 26724 -12523
rect 26780 -12557 26814 -12523
rect 16684 -12658 16718 -12624
rect 16774 -12658 16808 -12624
rect 16864 -12658 16898 -12624
rect 16954 -12658 16988 -12624
rect 17044 -12658 17078 -12624
rect 17134 -12658 17168 -12624
rect 17224 -12658 17258 -12624
rect 17314 -12658 17348 -12624
rect 17404 -12658 17438 -12624
rect 17494 -12658 17528 -12624
rect 17584 -12658 17618 -12624
rect 17674 -12658 17708 -12624
rect 17764 -12658 17798 -12624
rect 17972 -12658 18006 -12624
rect 18062 -12658 18096 -12624
rect 18152 -12658 18186 -12624
rect 18242 -12658 18276 -12624
rect 18332 -12658 18366 -12624
rect 18422 -12658 18456 -12624
rect 18512 -12658 18546 -12624
rect 18602 -12658 18636 -12624
rect 18692 -12658 18726 -12624
rect 18782 -12658 18816 -12624
rect 18872 -12658 18906 -12624
rect 18962 -12658 18996 -12624
rect 19052 -12658 19086 -12624
rect 19260 -12658 19294 -12624
rect 19350 -12658 19384 -12624
rect 19440 -12658 19474 -12624
rect 19530 -12658 19564 -12624
rect 19620 -12658 19654 -12624
rect 19710 -12658 19744 -12624
rect 19800 -12658 19834 -12624
rect 19890 -12658 19924 -12624
rect 19980 -12658 20014 -12624
rect 20070 -12658 20104 -12624
rect 20160 -12658 20194 -12624
rect 20250 -12658 20284 -12624
rect 20340 -12658 20374 -12624
rect 20548 -12658 20582 -12624
rect 20638 -12658 20672 -12624
rect 20728 -12658 20762 -12624
rect 20818 -12658 20852 -12624
rect 20908 -12658 20942 -12624
rect 20998 -12658 21032 -12624
rect 21088 -12658 21122 -12624
rect 21178 -12658 21212 -12624
rect 21268 -12658 21302 -12624
rect 21358 -12658 21392 -12624
rect 21448 -12658 21482 -12624
rect 21538 -12658 21572 -12624
rect 21628 -12658 21662 -12624
rect 21836 -12658 21870 -12624
rect 21926 -12658 21960 -12624
rect 22016 -12658 22050 -12624
rect 22106 -12658 22140 -12624
rect 22196 -12658 22230 -12624
rect 22286 -12658 22320 -12624
rect 22376 -12658 22410 -12624
rect 22466 -12658 22500 -12624
rect 22556 -12658 22590 -12624
rect 22646 -12658 22680 -12624
rect 22736 -12658 22770 -12624
rect 22826 -12658 22860 -12624
rect 22916 -12658 22950 -12624
rect 23124 -12658 23158 -12624
rect 23214 -12658 23248 -12624
rect 23304 -12658 23338 -12624
rect 23394 -12658 23428 -12624
rect 23484 -12658 23518 -12624
rect 23574 -12658 23608 -12624
rect 23664 -12658 23698 -12624
rect 23754 -12658 23788 -12624
rect 23844 -12658 23878 -12624
rect 23934 -12658 23968 -12624
rect 24024 -12658 24058 -12624
rect 24114 -12658 24148 -12624
rect 24204 -12658 24238 -12624
rect 24412 -12658 24446 -12624
rect 24502 -12658 24536 -12624
rect 24592 -12658 24626 -12624
rect 24682 -12658 24716 -12624
rect 24772 -12658 24806 -12624
rect 24862 -12658 24896 -12624
rect 24952 -12658 24986 -12624
rect 25042 -12658 25076 -12624
rect 25132 -12658 25166 -12624
rect 25222 -12658 25256 -12624
rect 25312 -12658 25346 -12624
rect 25402 -12658 25436 -12624
rect 25492 -12658 25526 -12624
rect 25700 -12658 25734 -12624
rect 25790 -12658 25824 -12624
rect 25880 -12658 25914 -12624
rect 25970 -12658 26004 -12624
rect 26060 -12658 26094 -12624
rect 26150 -12658 26184 -12624
rect 26240 -12658 26274 -12624
rect 26330 -12658 26364 -12624
rect 26420 -12658 26454 -12624
rect 26510 -12658 26544 -12624
rect 26600 -12658 26634 -12624
rect 26690 -12658 26724 -12624
rect 26780 -12658 26814 -12624
rect 16600 -12754 16634 -12720
rect 16600 -12844 16634 -12810
rect 16600 -12934 16634 -12900
rect 16600 -13024 16634 -12990
rect 16600 -13114 16634 -13080
rect 16600 -13204 16634 -13170
rect 16600 -13294 16634 -13260
rect 16600 -13384 16634 -13350
rect 16600 -13474 16634 -13440
rect 16600 -13564 16634 -13530
rect 16600 -13654 16634 -13620
rect 16600 -13744 16634 -13710
rect 17787 -12754 17821 -12720
rect 17888 -12754 17922 -12720
rect 17787 -12844 17821 -12810
rect 17888 -12844 17922 -12810
rect 17787 -12934 17821 -12900
rect 17888 -12934 17922 -12900
rect 17787 -13024 17821 -12990
rect 17888 -13024 17922 -12990
rect 17787 -13114 17821 -13080
rect 17888 -13114 17922 -13080
rect 17787 -13204 17821 -13170
rect 17888 -13204 17922 -13170
rect 17787 -13294 17821 -13260
rect 17888 -13294 17922 -13260
rect 17787 -13384 17821 -13350
rect 17888 -13384 17922 -13350
rect 17787 -13474 17821 -13440
rect 17888 -13474 17922 -13440
rect 17787 -13564 17821 -13530
rect 17888 -13564 17922 -13530
rect 17787 -13654 17821 -13620
rect 17888 -13654 17922 -13620
rect 17787 -13744 17821 -13710
rect 17888 -13744 17922 -13710
rect 19075 -12754 19109 -12720
rect 19176 -12754 19210 -12720
rect 19075 -12844 19109 -12810
rect 19176 -12844 19210 -12810
rect 19075 -12934 19109 -12900
rect 19176 -12934 19210 -12900
rect 19075 -13024 19109 -12990
rect 19176 -13024 19210 -12990
rect 19075 -13114 19109 -13080
rect 19176 -13114 19210 -13080
rect 19075 -13204 19109 -13170
rect 19176 -13204 19210 -13170
rect 19075 -13294 19109 -13260
rect 19176 -13294 19210 -13260
rect 19075 -13384 19109 -13350
rect 19176 -13384 19210 -13350
rect 19075 -13474 19109 -13440
rect 19176 -13474 19210 -13440
rect 19075 -13564 19109 -13530
rect 19176 -13564 19210 -13530
rect 19075 -13654 19109 -13620
rect 19176 -13654 19210 -13620
rect 19075 -13744 19109 -13710
rect 19176 -13744 19210 -13710
rect 20363 -12754 20397 -12720
rect 20464 -12754 20498 -12720
rect 20363 -12844 20397 -12810
rect 20464 -12844 20498 -12810
rect 20363 -12934 20397 -12900
rect 20464 -12934 20498 -12900
rect 20363 -13024 20397 -12990
rect 20464 -13024 20498 -12990
rect 20363 -13114 20397 -13080
rect 20464 -13114 20498 -13080
rect 20363 -13204 20397 -13170
rect 20464 -13204 20498 -13170
rect 20363 -13294 20397 -13260
rect 20464 -13294 20498 -13260
rect 20363 -13384 20397 -13350
rect 20464 -13384 20498 -13350
rect 20363 -13474 20397 -13440
rect 20464 -13474 20498 -13440
rect 20363 -13564 20397 -13530
rect 20464 -13564 20498 -13530
rect 20363 -13654 20397 -13620
rect 20464 -13654 20498 -13620
rect 20363 -13744 20397 -13710
rect 20464 -13744 20498 -13710
rect 21651 -12754 21685 -12720
rect 21752 -12754 21786 -12720
rect 21651 -12844 21685 -12810
rect 21752 -12844 21786 -12810
rect 21651 -12934 21685 -12900
rect 21752 -12934 21786 -12900
rect 21651 -13024 21685 -12990
rect 21752 -13024 21786 -12990
rect 21651 -13114 21685 -13080
rect 21752 -13114 21786 -13080
rect 21651 -13204 21685 -13170
rect 21752 -13204 21786 -13170
rect 21651 -13294 21685 -13260
rect 21752 -13294 21786 -13260
rect 21651 -13384 21685 -13350
rect 21752 -13384 21786 -13350
rect 21651 -13474 21685 -13440
rect 21752 -13474 21786 -13440
rect 21651 -13564 21685 -13530
rect 21752 -13564 21786 -13530
rect 21651 -13654 21685 -13620
rect 21752 -13654 21786 -13620
rect 21651 -13744 21685 -13710
rect 21752 -13744 21786 -13710
rect 22939 -12754 22973 -12720
rect 23040 -12754 23074 -12720
rect 22939 -12844 22973 -12810
rect 23040 -12844 23074 -12810
rect 22939 -12934 22973 -12900
rect 23040 -12934 23074 -12900
rect 22939 -13024 22973 -12990
rect 23040 -13024 23074 -12990
rect 22939 -13114 22973 -13080
rect 23040 -13114 23074 -13080
rect 22939 -13204 22973 -13170
rect 23040 -13204 23074 -13170
rect 22939 -13294 22973 -13260
rect 23040 -13294 23074 -13260
rect 22939 -13384 22973 -13350
rect 23040 -13384 23074 -13350
rect 22939 -13474 22973 -13440
rect 23040 -13474 23074 -13440
rect 22939 -13564 22973 -13530
rect 23040 -13564 23074 -13530
rect 22939 -13654 22973 -13620
rect 23040 -13654 23074 -13620
rect 22939 -13744 22973 -13710
rect 23040 -13744 23074 -13710
rect 24227 -12754 24261 -12720
rect 24328 -12754 24362 -12720
rect 24227 -12844 24261 -12810
rect 24328 -12844 24362 -12810
rect 24227 -12934 24261 -12900
rect 24328 -12934 24362 -12900
rect 24227 -13024 24261 -12990
rect 24328 -13024 24362 -12990
rect 24227 -13114 24261 -13080
rect 24328 -13114 24362 -13080
rect 24227 -13204 24261 -13170
rect 24328 -13204 24362 -13170
rect 24227 -13294 24261 -13260
rect 24328 -13294 24362 -13260
rect 24227 -13384 24261 -13350
rect 24328 -13384 24362 -13350
rect 24227 -13474 24261 -13440
rect 24328 -13474 24362 -13440
rect 24227 -13564 24261 -13530
rect 24328 -13564 24362 -13530
rect 24227 -13654 24261 -13620
rect 24328 -13654 24362 -13620
rect 24227 -13744 24261 -13710
rect 24328 -13744 24362 -13710
rect 25515 -12754 25549 -12720
rect 25616 -12754 25650 -12720
rect 25515 -12844 25549 -12810
rect 25616 -12844 25650 -12810
rect 25515 -12934 25549 -12900
rect 25616 -12934 25650 -12900
rect 25515 -13024 25549 -12990
rect 25616 -13024 25650 -12990
rect 25515 -13114 25549 -13080
rect 25616 -13114 25650 -13080
rect 25515 -13204 25549 -13170
rect 25616 -13204 25650 -13170
rect 25515 -13294 25549 -13260
rect 25616 -13294 25650 -13260
rect 25515 -13384 25549 -13350
rect 25616 -13384 25650 -13350
rect 25515 -13474 25549 -13440
rect 25616 -13474 25650 -13440
rect 25515 -13564 25549 -13530
rect 25616 -13564 25650 -13530
rect 25515 -13654 25549 -13620
rect 25616 -13654 25650 -13620
rect 25515 -13744 25549 -13710
rect 25616 -13744 25650 -13710
rect 26803 -12754 26837 -12720
rect 26803 -12844 26837 -12810
rect 26803 -12934 26837 -12900
rect 26803 -13024 26837 -12990
rect 26803 -13114 26837 -13080
rect 26803 -13204 26837 -13170
rect 26803 -13294 26837 -13260
rect 26803 -13384 26837 -13350
rect 26803 -13474 26837 -13440
rect 26803 -13564 26837 -13530
rect 26803 -13654 26837 -13620
rect 26803 -13744 26837 -13710
rect 16684 -13845 16718 -13811
rect 16774 -13845 16808 -13811
rect 16864 -13845 16898 -13811
rect 16954 -13845 16988 -13811
rect 17044 -13845 17078 -13811
rect 17134 -13845 17168 -13811
rect 17224 -13845 17258 -13811
rect 17314 -13845 17348 -13811
rect 17404 -13845 17438 -13811
rect 17494 -13845 17528 -13811
rect 17584 -13845 17618 -13811
rect 17674 -13845 17708 -13811
rect 17764 -13845 17798 -13811
rect 17972 -13845 18006 -13811
rect 18062 -13845 18096 -13811
rect 18152 -13845 18186 -13811
rect 18242 -13845 18276 -13811
rect 18332 -13845 18366 -13811
rect 18422 -13845 18456 -13811
rect 18512 -13845 18546 -13811
rect 18602 -13845 18636 -13811
rect 18692 -13845 18726 -13811
rect 18782 -13845 18816 -13811
rect 18872 -13845 18906 -13811
rect 18962 -13845 18996 -13811
rect 19052 -13845 19086 -13811
rect 19260 -13845 19294 -13811
rect 19350 -13845 19384 -13811
rect 19440 -13845 19474 -13811
rect 19530 -13845 19564 -13811
rect 19620 -13845 19654 -13811
rect 19710 -13845 19744 -13811
rect 19800 -13845 19834 -13811
rect 19890 -13845 19924 -13811
rect 19980 -13845 20014 -13811
rect 20070 -13845 20104 -13811
rect 20160 -13845 20194 -13811
rect 20250 -13845 20284 -13811
rect 20340 -13845 20374 -13811
rect 20548 -13845 20582 -13811
rect 20638 -13845 20672 -13811
rect 20728 -13845 20762 -13811
rect 20818 -13845 20852 -13811
rect 20908 -13845 20942 -13811
rect 20998 -13845 21032 -13811
rect 21088 -13845 21122 -13811
rect 21178 -13845 21212 -13811
rect 21268 -13845 21302 -13811
rect 21358 -13845 21392 -13811
rect 21448 -13845 21482 -13811
rect 21538 -13845 21572 -13811
rect 21628 -13845 21662 -13811
rect 21836 -13845 21870 -13811
rect 21926 -13845 21960 -13811
rect 22016 -13845 22050 -13811
rect 22106 -13845 22140 -13811
rect 22196 -13845 22230 -13811
rect 22286 -13845 22320 -13811
rect 22376 -13845 22410 -13811
rect 22466 -13845 22500 -13811
rect 22556 -13845 22590 -13811
rect 22646 -13845 22680 -13811
rect 22736 -13845 22770 -13811
rect 22826 -13845 22860 -13811
rect 22916 -13845 22950 -13811
rect 23124 -13845 23158 -13811
rect 23214 -13845 23248 -13811
rect 23304 -13845 23338 -13811
rect 23394 -13845 23428 -13811
rect 23484 -13845 23518 -13811
rect 23574 -13845 23608 -13811
rect 23664 -13845 23698 -13811
rect 23754 -13845 23788 -13811
rect 23844 -13845 23878 -13811
rect 23934 -13845 23968 -13811
rect 24024 -13845 24058 -13811
rect 24114 -13845 24148 -13811
rect 24204 -13845 24238 -13811
rect 24412 -13845 24446 -13811
rect 24502 -13845 24536 -13811
rect 24592 -13845 24626 -13811
rect 24682 -13845 24716 -13811
rect 24772 -13845 24806 -13811
rect 24862 -13845 24896 -13811
rect 24952 -13845 24986 -13811
rect 25042 -13845 25076 -13811
rect 25132 -13845 25166 -13811
rect 25222 -13845 25256 -13811
rect 25312 -13845 25346 -13811
rect 25402 -13845 25436 -13811
rect 25492 -13845 25526 -13811
rect 25700 -13845 25734 -13811
rect 25790 -13845 25824 -13811
rect 25880 -13845 25914 -13811
rect 25970 -13845 26004 -13811
rect 26060 -13845 26094 -13811
rect 26150 -13845 26184 -13811
rect 26240 -13845 26274 -13811
rect 26330 -13845 26364 -13811
rect 26420 -13845 26454 -13811
rect 26510 -13845 26544 -13811
rect 26600 -13845 26634 -13811
rect 26690 -13845 26724 -13811
rect 26780 -13845 26814 -13811
rect 16684 -13946 16718 -13912
rect 16774 -13946 16808 -13912
rect 16864 -13946 16898 -13912
rect 16954 -13946 16988 -13912
rect 17044 -13946 17078 -13912
rect 17134 -13946 17168 -13912
rect 17224 -13946 17258 -13912
rect 17314 -13946 17348 -13912
rect 17404 -13946 17438 -13912
rect 17494 -13946 17528 -13912
rect 17584 -13946 17618 -13912
rect 17674 -13946 17708 -13912
rect 17764 -13946 17798 -13912
rect 17972 -13946 18006 -13912
rect 18062 -13946 18096 -13912
rect 18152 -13946 18186 -13912
rect 18242 -13946 18276 -13912
rect 18332 -13946 18366 -13912
rect 18422 -13946 18456 -13912
rect 18512 -13946 18546 -13912
rect 18602 -13946 18636 -13912
rect 18692 -13946 18726 -13912
rect 18782 -13946 18816 -13912
rect 18872 -13946 18906 -13912
rect 18962 -13946 18996 -13912
rect 19052 -13946 19086 -13912
rect 19260 -13946 19294 -13912
rect 19350 -13946 19384 -13912
rect 19440 -13946 19474 -13912
rect 19530 -13946 19564 -13912
rect 19620 -13946 19654 -13912
rect 19710 -13946 19744 -13912
rect 19800 -13946 19834 -13912
rect 19890 -13946 19924 -13912
rect 19980 -13946 20014 -13912
rect 20070 -13946 20104 -13912
rect 20160 -13946 20194 -13912
rect 20250 -13946 20284 -13912
rect 20340 -13946 20374 -13912
rect 20548 -13946 20582 -13912
rect 20638 -13946 20672 -13912
rect 20728 -13946 20762 -13912
rect 20818 -13946 20852 -13912
rect 20908 -13946 20942 -13912
rect 20998 -13946 21032 -13912
rect 21088 -13946 21122 -13912
rect 21178 -13946 21212 -13912
rect 21268 -13946 21302 -13912
rect 21358 -13946 21392 -13912
rect 21448 -13946 21482 -13912
rect 21538 -13946 21572 -13912
rect 21628 -13946 21662 -13912
rect 21836 -13946 21870 -13912
rect 21926 -13946 21960 -13912
rect 22016 -13946 22050 -13912
rect 22106 -13946 22140 -13912
rect 22196 -13946 22230 -13912
rect 22286 -13946 22320 -13912
rect 22376 -13946 22410 -13912
rect 22466 -13946 22500 -13912
rect 22556 -13946 22590 -13912
rect 22646 -13946 22680 -13912
rect 22736 -13946 22770 -13912
rect 22826 -13946 22860 -13912
rect 22916 -13946 22950 -13912
rect 23124 -13946 23158 -13912
rect 23214 -13946 23248 -13912
rect 23304 -13946 23338 -13912
rect 23394 -13946 23428 -13912
rect 23484 -13946 23518 -13912
rect 23574 -13946 23608 -13912
rect 23664 -13946 23698 -13912
rect 23754 -13946 23788 -13912
rect 23844 -13946 23878 -13912
rect 23934 -13946 23968 -13912
rect 24024 -13946 24058 -13912
rect 24114 -13946 24148 -13912
rect 24204 -13946 24238 -13912
rect 24412 -13946 24446 -13912
rect 24502 -13946 24536 -13912
rect 24592 -13946 24626 -13912
rect 24682 -13946 24716 -13912
rect 24772 -13946 24806 -13912
rect 24862 -13946 24896 -13912
rect 24952 -13946 24986 -13912
rect 25042 -13946 25076 -13912
rect 25132 -13946 25166 -13912
rect 25222 -13946 25256 -13912
rect 25312 -13946 25346 -13912
rect 25402 -13946 25436 -13912
rect 25492 -13946 25526 -13912
rect 25700 -13946 25734 -13912
rect 25790 -13946 25824 -13912
rect 25880 -13946 25914 -13912
rect 25970 -13946 26004 -13912
rect 26060 -13946 26094 -13912
rect 26150 -13946 26184 -13912
rect 26240 -13946 26274 -13912
rect 26330 -13946 26364 -13912
rect 26420 -13946 26454 -13912
rect 26510 -13946 26544 -13912
rect 26600 -13946 26634 -13912
rect 26690 -13946 26724 -13912
rect 26780 -13946 26814 -13912
rect 16600 -14042 16634 -14008
rect 16600 -14132 16634 -14098
rect 16600 -14222 16634 -14188
rect 16600 -14312 16634 -14278
rect 16600 -14402 16634 -14368
rect 16600 -14492 16634 -14458
rect 16600 -14582 16634 -14548
rect 16600 -14672 16634 -14638
rect 16600 -14762 16634 -14728
rect 16600 -14852 16634 -14818
rect 16600 -14942 16634 -14908
rect 16600 -15032 16634 -14998
rect 17787 -14042 17821 -14008
rect 17888 -14042 17922 -14008
rect 17787 -14132 17821 -14098
rect 17888 -14132 17922 -14098
rect 17787 -14222 17821 -14188
rect 17888 -14222 17922 -14188
rect 17787 -14312 17821 -14278
rect 17888 -14312 17922 -14278
rect 17787 -14402 17821 -14368
rect 17888 -14402 17922 -14368
rect 17787 -14492 17821 -14458
rect 17888 -14492 17922 -14458
rect 17787 -14582 17821 -14548
rect 17888 -14582 17922 -14548
rect 17787 -14672 17821 -14638
rect 17888 -14672 17922 -14638
rect 17787 -14762 17821 -14728
rect 17888 -14762 17922 -14728
rect 17787 -14852 17821 -14818
rect 17888 -14852 17922 -14818
rect 17787 -14942 17821 -14908
rect 17888 -14942 17922 -14908
rect 17787 -15032 17821 -14998
rect 17888 -15032 17922 -14998
rect 19075 -14042 19109 -14008
rect 19176 -14042 19210 -14008
rect 19075 -14132 19109 -14098
rect 19176 -14132 19210 -14098
rect 19075 -14222 19109 -14188
rect 19176 -14222 19210 -14188
rect 19075 -14312 19109 -14278
rect 19176 -14312 19210 -14278
rect 19075 -14402 19109 -14368
rect 19176 -14402 19210 -14368
rect 19075 -14492 19109 -14458
rect 19176 -14492 19210 -14458
rect 19075 -14582 19109 -14548
rect 19176 -14582 19210 -14548
rect 19075 -14672 19109 -14638
rect 19176 -14672 19210 -14638
rect 19075 -14762 19109 -14728
rect 19176 -14762 19210 -14728
rect 19075 -14852 19109 -14818
rect 19176 -14852 19210 -14818
rect 19075 -14942 19109 -14908
rect 19176 -14942 19210 -14908
rect 19075 -15032 19109 -14998
rect 19176 -15032 19210 -14998
rect 20363 -14042 20397 -14008
rect 20464 -14042 20498 -14008
rect 20363 -14132 20397 -14098
rect 20464 -14132 20498 -14098
rect 20363 -14222 20397 -14188
rect 20464 -14222 20498 -14188
rect 20363 -14312 20397 -14278
rect 20464 -14312 20498 -14278
rect 20363 -14402 20397 -14368
rect 20464 -14402 20498 -14368
rect 20363 -14492 20397 -14458
rect 20464 -14492 20498 -14458
rect 20363 -14582 20397 -14548
rect 20464 -14582 20498 -14548
rect 20363 -14672 20397 -14638
rect 20464 -14672 20498 -14638
rect 20363 -14762 20397 -14728
rect 20464 -14762 20498 -14728
rect 20363 -14852 20397 -14818
rect 20464 -14852 20498 -14818
rect 20363 -14942 20397 -14908
rect 20464 -14942 20498 -14908
rect 20363 -15032 20397 -14998
rect 20464 -15032 20498 -14998
rect 21651 -14042 21685 -14008
rect 21752 -14042 21786 -14008
rect 21651 -14132 21685 -14098
rect 21752 -14132 21786 -14098
rect 21651 -14222 21685 -14188
rect 21752 -14222 21786 -14188
rect 21651 -14312 21685 -14278
rect 21752 -14312 21786 -14278
rect 21651 -14402 21685 -14368
rect 21752 -14402 21786 -14368
rect 21651 -14492 21685 -14458
rect 21752 -14492 21786 -14458
rect 21651 -14582 21685 -14548
rect 21752 -14582 21786 -14548
rect 21651 -14672 21685 -14638
rect 21752 -14672 21786 -14638
rect 21651 -14762 21685 -14728
rect 21752 -14762 21786 -14728
rect 21651 -14852 21685 -14818
rect 21752 -14852 21786 -14818
rect 21651 -14942 21685 -14908
rect 21752 -14942 21786 -14908
rect 21651 -15032 21685 -14998
rect 21752 -15032 21786 -14998
rect 22939 -14042 22973 -14008
rect 23040 -14042 23074 -14008
rect 22939 -14132 22973 -14098
rect 23040 -14132 23074 -14098
rect 22939 -14222 22973 -14188
rect 23040 -14222 23074 -14188
rect 22939 -14312 22973 -14278
rect 23040 -14312 23074 -14278
rect 22939 -14402 22973 -14368
rect 23040 -14402 23074 -14368
rect 22939 -14492 22973 -14458
rect 23040 -14492 23074 -14458
rect 22939 -14582 22973 -14548
rect 23040 -14582 23074 -14548
rect 22939 -14672 22973 -14638
rect 23040 -14672 23074 -14638
rect 22939 -14762 22973 -14728
rect 23040 -14762 23074 -14728
rect 22939 -14852 22973 -14818
rect 23040 -14852 23074 -14818
rect 22939 -14942 22973 -14908
rect 23040 -14942 23074 -14908
rect 22939 -15032 22973 -14998
rect 23040 -15032 23074 -14998
rect 24227 -14042 24261 -14008
rect 24328 -14042 24362 -14008
rect 24227 -14132 24261 -14098
rect 24328 -14132 24362 -14098
rect 24227 -14222 24261 -14188
rect 24328 -14222 24362 -14188
rect 24227 -14312 24261 -14278
rect 24328 -14312 24362 -14278
rect 24227 -14402 24261 -14368
rect 24328 -14402 24362 -14368
rect 24227 -14492 24261 -14458
rect 24328 -14492 24362 -14458
rect 24227 -14582 24261 -14548
rect 24328 -14582 24362 -14548
rect 24227 -14672 24261 -14638
rect 24328 -14672 24362 -14638
rect 24227 -14762 24261 -14728
rect 24328 -14762 24362 -14728
rect 24227 -14852 24261 -14818
rect 24328 -14852 24362 -14818
rect 24227 -14942 24261 -14908
rect 24328 -14942 24362 -14908
rect 24227 -15032 24261 -14998
rect 24328 -15032 24362 -14998
rect 25515 -14042 25549 -14008
rect 25616 -14042 25650 -14008
rect 25515 -14132 25549 -14098
rect 25616 -14132 25650 -14098
rect 25515 -14222 25549 -14188
rect 25616 -14222 25650 -14188
rect 25515 -14312 25549 -14278
rect 25616 -14312 25650 -14278
rect 25515 -14402 25549 -14368
rect 25616 -14402 25650 -14368
rect 25515 -14492 25549 -14458
rect 25616 -14492 25650 -14458
rect 25515 -14582 25549 -14548
rect 25616 -14582 25650 -14548
rect 25515 -14672 25549 -14638
rect 25616 -14672 25650 -14638
rect 25515 -14762 25549 -14728
rect 25616 -14762 25650 -14728
rect 25515 -14852 25549 -14818
rect 25616 -14852 25650 -14818
rect 25515 -14942 25549 -14908
rect 25616 -14942 25650 -14908
rect 25515 -15032 25549 -14998
rect 25616 -15032 25650 -14998
rect 26803 -14042 26837 -14008
rect 26803 -14132 26837 -14098
rect 26803 -14222 26837 -14188
rect 26803 -14312 26837 -14278
rect 26803 -14402 26837 -14368
rect 26803 -14492 26837 -14458
rect 26803 -14582 26837 -14548
rect 26803 -14672 26837 -14638
rect 26803 -14762 26837 -14728
rect 26803 -14852 26837 -14818
rect 26803 -14942 26837 -14908
rect 26803 -15032 26837 -14998
rect 16684 -15133 16718 -15099
rect 16774 -15133 16808 -15099
rect 16864 -15133 16898 -15099
rect 16954 -15133 16988 -15099
rect 17044 -15133 17078 -15099
rect 17134 -15133 17168 -15099
rect 17224 -15133 17258 -15099
rect 17314 -15133 17348 -15099
rect 17404 -15133 17438 -15099
rect 17494 -15133 17528 -15099
rect 17584 -15133 17618 -15099
rect 17674 -15133 17708 -15099
rect 17764 -15133 17798 -15099
rect 17972 -15133 18006 -15099
rect 18062 -15133 18096 -15099
rect 18152 -15133 18186 -15099
rect 18242 -15133 18276 -15099
rect 18332 -15133 18366 -15099
rect 18422 -15133 18456 -15099
rect 18512 -15133 18546 -15099
rect 18602 -15133 18636 -15099
rect 18692 -15133 18726 -15099
rect 18782 -15133 18816 -15099
rect 18872 -15133 18906 -15099
rect 18962 -15133 18996 -15099
rect 19052 -15133 19086 -15099
rect 19260 -15133 19294 -15099
rect 19350 -15133 19384 -15099
rect 19440 -15133 19474 -15099
rect 19530 -15133 19564 -15099
rect 19620 -15133 19654 -15099
rect 19710 -15133 19744 -15099
rect 19800 -15133 19834 -15099
rect 19890 -15133 19924 -15099
rect 19980 -15133 20014 -15099
rect 20070 -15133 20104 -15099
rect 20160 -15133 20194 -15099
rect 20250 -15133 20284 -15099
rect 20340 -15133 20374 -15099
rect 20548 -15133 20582 -15099
rect 20638 -15133 20672 -15099
rect 20728 -15133 20762 -15099
rect 20818 -15133 20852 -15099
rect 20908 -15133 20942 -15099
rect 20998 -15133 21032 -15099
rect 21088 -15133 21122 -15099
rect 21178 -15133 21212 -15099
rect 21268 -15133 21302 -15099
rect 21358 -15133 21392 -15099
rect 21448 -15133 21482 -15099
rect 21538 -15133 21572 -15099
rect 21628 -15133 21662 -15099
rect 21836 -15133 21870 -15099
rect 21926 -15133 21960 -15099
rect 22016 -15133 22050 -15099
rect 22106 -15133 22140 -15099
rect 22196 -15133 22230 -15099
rect 22286 -15133 22320 -15099
rect 22376 -15133 22410 -15099
rect 22466 -15133 22500 -15099
rect 22556 -15133 22590 -15099
rect 22646 -15133 22680 -15099
rect 22736 -15133 22770 -15099
rect 22826 -15133 22860 -15099
rect 22916 -15133 22950 -15099
rect 23124 -15133 23158 -15099
rect 23214 -15133 23248 -15099
rect 23304 -15133 23338 -15099
rect 23394 -15133 23428 -15099
rect 23484 -15133 23518 -15099
rect 23574 -15133 23608 -15099
rect 23664 -15133 23698 -15099
rect 23754 -15133 23788 -15099
rect 23844 -15133 23878 -15099
rect 23934 -15133 23968 -15099
rect 24024 -15133 24058 -15099
rect 24114 -15133 24148 -15099
rect 24204 -15133 24238 -15099
rect 24412 -15133 24446 -15099
rect 24502 -15133 24536 -15099
rect 24592 -15133 24626 -15099
rect 24682 -15133 24716 -15099
rect 24772 -15133 24806 -15099
rect 24862 -15133 24896 -15099
rect 24952 -15133 24986 -15099
rect 25042 -15133 25076 -15099
rect 25132 -15133 25166 -15099
rect 25222 -15133 25256 -15099
rect 25312 -15133 25346 -15099
rect 25402 -15133 25436 -15099
rect 25492 -15133 25526 -15099
rect 25700 -15133 25734 -15099
rect 25790 -15133 25824 -15099
rect 25880 -15133 25914 -15099
rect 25970 -15133 26004 -15099
rect 26060 -15133 26094 -15099
rect 26150 -15133 26184 -15099
rect 26240 -15133 26274 -15099
rect 26330 -15133 26364 -15099
rect 26420 -15133 26454 -15099
rect 26510 -15133 26544 -15099
rect 26600 -15133 26634 -15099
rect 26690 -15133 26724 -15099
rect 26780 -15133 26814 -15099
rect 16684 -15234 16718 -15200
rect 16774 -15234 16808 -15200
rect 16864 -15234 16898 -15200
rect 16954 -15234 16988 -15200
rect 17044 -15234 17078 -15200
rect 17134 -15234 17168 -15200
rect 17224 -15234 17258 -15200
rect 17314 -15234 17348 -15200
rect 17404 -15234 17438 -15200
rect 17494 -15234 17528 -15200
rect 17584 -15234 17618 -15200
rect 17674 -15234 17708 -15200
rect 17764 -15234 17798 -15200
rect 17972 -15234 18006 -15200
rect 18062 -15234 18096 -15200
rect 18152 -15234 18186 -15200
rect 18242 -15234 18276 -15200
rect 18332 -15234 18366 -15200
rect 18422 -15234 18456 -15200
rect 18512 -15234 18546 -15200
rect 18602 -15234 18636 -15200
rect 18692 -15234 18726 -15200
rect 18782 -15234 18816 -15200
rect 18872 -15234 18906 -15200
rect 18962 -15234 18996 -15200
rect 19052 -15234 19086 -15200
rect 19260 -15234 19294 -15200
rect 19350 -15234 19384 -15200
rect 19440 -15234 19474 -15200
rect 19530 -15234 19564 -15200
rect 19620 -15234 19654 -15200
rect 19710 -15234 19744 -15200
rect 19800 -15234 19834 -15200
rect 19890 -15234 19924 -15200
rect 19980 -15234 20014 -15200
rect 20070 -15234 20104 -15200
rect 20160 -15234 20194 -15200
rect 20250 -15234 20284 -15200
rect 20340 -15234 20374 -15200
rect 20548 -15234 20582 -15200
rect 20638 -15234 20672 -15200
rect 20728 -15234 20762 -15200
rect 20818 -15234 20852 -15200
rect 20908 -15234 20942 -15200
rect 20998 -15234 21032 -15200
rect 21088 -15234 21122 -15200
rect 21178 -15234 21212 -15200
rect 21268 -15234 21302 -15200
rect 21358 -15234 21392 -15200
rect 21448 -15234 21482 -15200
rect 21538 -15234 21572 -15200
rect 21628 -15234 21662 -15200
rect 21836 -15234 21870 -15200
rect 21926 -15234 21960 -15200
rect 22016 -15234 22050 -15200
rect 22106 -15234 22140 -15200
rect 22196 -15234 22230 -15200
rect 22286 -15234 22320 -15200
rect 22376 -15234 22410 -15200
rect 22466 -15234 22500 -15200
rect 22556 -15234 22590 -15200
rect 22646 -15234 22680 -15200
rect 22736 -15234 22770 -15200
rect 22826 -15234 22860 -15200
rect 22916 -15234 22950 -15200
rect 23124 -15234 23158 -15200
rect 23214 -15234 23248 -15200
rect 23304 -15234 23338 -15200
rect 23394 -15234 23428 -15200
rect 23484 -15234 23518 -15200
rect 23574 -15234 23608 -15200
rect 23664 -15234 23698 -15200
rect 23754 -15234 23788 -15200
rect 23844 -15234 23878 -15200
rect 23934 -15234 23968 -15200
rect 24024 -15234 24058 -15200
rect 24114 -15234 24148 -15200
rect 24204 -15234 24238 -15200
rect 24412 -15234 24446 -15200
rect 24502 -15234 24536 -15200
rect 24592 -15234 24626 -15200
rect 24682 -15234 24716 -15200
rect 24772 -15234 24806 -15200
rect 24862 -15234 24896 -15200
rect 24952 -15234 24986 -15200
rect 25042 -15234 25076 -15200
rect 25132 -15234 25166 -15200
rect 25222 -15234 25256 -15200
rect 25312 -15234 25346 -15200
rect 25402 -15234 25436 -15200
rect 25492 -15234 25526 -15200
rect 25700 -15234 25734 -15200
rect 25790 -15234 25824 -15200
rect 25880 -15234 25914 -15200
rect 25970 -15234 26004 -15200
rect 26060 -15234 26094 -15200
rect 26150 -15234 26184 -15200
rect 26240 -15234 26274 -15200
rect 26330 -15234 26364 -15200
rect 26420 -15234 26454 -15200
rect 26510 -15234 26544 -15200
rect 26600 -15234 26634 -15200
rect 26690 -15234 26724 -15200
rect 26780 -15234 26814 -15200
rect 16600 -15330 16634 -15296
rect 16600 -15420 16634 -15386
rect 16600 -15510 16634 -15476
rect 16600 -15600 16634 -15566
rect 16600 -15690 16634 -15656
rect 16600 -15780 16634 -15746
rect 16600 -15870 16634 -15836
rect 16600 -15960 16634 -15926
rect 16600 -16050 16634 -16016
rect 16600 -16140 16634 -16106
rect 16600 -16230 16634 -16196
rect 16600 -16320 16634 -16286
rect 17787 -15330 17821 -15296
rect 17888 -15330 17922 -15296
rect 17787 -15420 17821 -15386
rect 17888 -15420 17922 -15386
rect 17787 -15510 17821 -15476
rect 17888 -15510 17922 -15476
rect 17787 -15600 17821 -15566
rect 17888 -15600 17922 -15566
rect 17787 -15690 17821 -15656
rect 17888 -15690 17922 -15656
rect 17787 -15780 17821 -15746
rect 17888 -15780 17922 -15746
rect 17787 -15870 17821 -15836
rect 17888 -15870 17922 -15836
rect 17787 -15960 17821 -15926
rect 17888 -15960 17922 -15926
rect 17787 -16050 17821 -16016
rect 17888 -16050 17922 -16016
rect 17787 -16140 17821 -16106
rect 17888 -16140 17922 -16106
rect 17787 -16230 17821 -16196
rect 17888 -16230 17922 -16196
rect 17787 -16320 17821 -16286
rect 17888 -16320 17922 -16286
rect 19075 -15330 19109 -15296
rect 19176 -15330 19210 -15296
rect 19075 -15420 19109 -15386
rect 19176 -15420 19210 -15386
rect 19075 -15510 19109 -15476
rect 19176 -15510 19210 -15476
rect 19075 -15600 19109 -15566
rect 19176 -15600 19210 -15566
rect 19075 -15690 19109 -15656
rect 19176 -15690 19210 -15656
rect 19075 -15780 19109 -15746
rect 19176 -15780 19210 -15746
rect 19075 -15870 19109 -15836
rect 19176 -15870 19210 -15836
rect 19075 -15960 19109 -15926
rect 19176 -15960 19210 -15926
rect 19075 -16050 19109 -16016
rect 19176 -16050 19210 -16016
rect 19075 -16140 19109 -16106
rect 19176 -16140 19210 -16106
rect 19075 -16230 19109 -16196
rect 19176 -16230 19210 -16196
rect 19075 -16320 19109 -16286
rect 19176 -16320 19210 -16286
rect 20363 -15330 20397 -15296
rect 20464 -15330 20498 -15296
rect 20363 -15420 20397 -15386
rect 20464 -15420 20498 -15386
rect 20363 -15510 20397 -15476
rect 20464 -15510 20498 -15476
rect 20363 -15600 20397 -15566
rect 20464 -15600 20498 -15566
rect 20363 -15690 20397 -15656
rect 20464 -15690 20498 -15656
rect 20363 -15780 20397 -15746
rect 20464 -15780 20498 -15746
rect 20363 -15870 20397 -15836
rect 20464 -15870 20498 -15836
rect 20363 -15960 20397 -15926
rect 20464 -15960 20498 -15926
rect 20363 -16050 20397 -16016
rect 20464 -16050 20498 -16016
rect 20363 -16140 20397 -16106
rect 20464 -16140 20498 -16106
rect 20363 -16230 20397 -16196
rect 20464 -16230 20498 -16196
rect 20363 -16320 20397 -16286
rect 20464 -16320 20498 -16286
rect 21651 -15330 21685 -15296
rect 21752 -15330 21786 -15296
rect 21651 -15420 21685 -15386
rect 21752 -15420 21786 -15386
rect 21651 -15510 21685 -15476
rect 21752 -15510 21786 -15476
rect 21651 -15600 21685 -15566
rect 21752 -15600 21786 -15566
rect 21651 -15690 21685 -15656
rect 21752 -15690 21786 -15656
rect 21651 -15780 21685 -15746
rect 21752 -15780 21786 -15746
rect 21651 -15870 21685 -15836
rect 21752 -15870 21786 -15836
rect 21651 -15960 21685 -15926
rect 21752 -15960 21786 -15926
rect 21651 -16050 21685 -16016
rect 21752 -16050 21786 -16016
rect 21651 -16140 21685 -16106
rect 21752 -16140 21786 -16106
rect 21651 -16230 21685 -16196
rect 21752 -16230 21786 -16196
rect 21651 -16320 21685 -16286
rect 21752 -16320 21786 -16286
rect 22939 -15330 22973 -15296
rect 23040 -15330 23074 -15296
rect 22939 -15420 22973 -15386
rect 23040 -15420 23074 -15386
rect 22939 -15510 22973 -15476
rect 23040 -15510 23074 -15476
rect 22939 -15600 22973 -15566
rect 23040 -15600 23074 -15566
rect 22939 -15690 22973 -15656
rect 23040 -15690 23074 -15656
rect 22939 -15780 22973 -15746
rect 23040 -15780 23074 -15746
rect 22939 -15870 22973 -15836
rect 23040 -15870 23074 -15836
rect 22939 -15960 22973 -15926
rect 23040 -15960 23074 -15926
rect 22939 -16050 22973 -16016
rect 23040 -16050 23074 -16016
rect 22939 -16140 22973 -16106
rect 23040 -16140 23074 -16106
rect 22939 -16230 22973 -16196
rect 23040 -16230 23074 -16196
rect 22939 -16320 22973 -16286
rect 23040 -16320 23074 -16286
rect 24227 -15330 24261 -15296
rect 24328 -15330 24362 -15296
rect 24227 -15420 24261 -15386
rect 24328 -15420 24362 -15386
rect 24227 -15510 24261 -15476
rect 24328 -15510 24362 -15476
rect 24227 -15600 24261 -15566
rect 24328 -15600 24362 -15566
rect 24227 -15690 24261 -15656
rect 24328 -15690 24362 -15656
rect 24227 -15780 24261 -15746
rect 24328 -15780 24362 -15746
rect 24227 -15870 24261 -15836
rect 24328 -15870 24362 -15836
rect 24227 -15960 24261 -15926
rect 24328 -15960 24362 -15926
rect 24227 -16050 24261 -16016
rect 24328 -16050 24362 -16016
rect 24227 -16140 24261 -16106
rect 24328 -16140 24362 -16106
rect 24227 -16230 24261 -16196
rect 24328 -16230 24362 -16196
rect 24227 -16320 24261 -16286
rect 24328 -16320 24362 -16286
rect 25515 -15330 25549 -15296
rect 25616 -15330 25650 -15296
rect 25515 -15420 25549 -15386
rect 25616 -15420 25650 -15386
rect 25515 -15510 25549 -15476
rect 25616 -15510 25650 -15476
rect 25515 -15600 25549 -15566
rect 25616 -15600 25650 -15566
rect 25515 -15690 25549 -15656
rect 25616 -15690 25650 -15656
rect 25515 -15780 25549 -15746
rect 25616 -15780 25650 -15746
rect 25515 -15870 25549 -15836
rect 25616 -15870 25650 -15836
rect 25515 -15960 25549 -15926
rect 25616 -15960 25650 -15926
rect 25515 -16050 25549 -16016
rect 25616 -16050 25650 -16016
rect 25515 -16140 25549 -16106
rect 25616 -16140 25650 -16106
rect 25515 -16230 25549 -16196
rect 25616 -16230 25650 -16196
rect 25515 -16320 25549 -16286
rect 25616 -16320 25650 -16286
rect 26803 -15330 26837 -15296
rect 26803 -15420 26837 -15386
rect 26803 -15510 26837 -15476
rect 26803 -15600 26837 -15566
rect 26803 -15690 26837 -15656
rect 26803 -15780 26837 -15746
rect 26803 -15870 26837 -15836
rect 26803 -15960 26837 -15926
rect 26803 -16050 26837 -16016
rect 26803 -16140 26837 -16106
rect 26803 -16230 26837 -16196
rect 26803 -16320 26837 -16286
rect 16684 -16421 16718 -16387
rect 16774 -16421 16808 -16387
rect 16864 -16421 16898 -16387
rect 16954 -16421 16988 -16387
rect 17044 -16421 17078 -16387
rect 17134 -16421 17168 -16387
rect 17224 -16421 17258 -16387
rect 17314 -16421 17348 -16387
rect 17404 -16421 17438 -16387
rect 17494 -16421 17528 -16387
rect 17584 -16421 17618 -16387
rect 17674 -16421 17708 -16387
rect 17764 -16421 17798 -16387
rect 17972 -16421 18006 -16387
rect 18062 -16421 18096 -16387
rect 18152 -16421 18186 -16387
rect 18242 -16421 18276 -16387
rect 18332 -16421 18366 -16387
rect 18422 -16421 18456 -16387
rect 18512 -16421 18546 -16387
rect 18602 -16421 18636 -16387
rect 18692 -16421 18726 -16387
rect 18782 -16421 18816 -16387
rect 18872 -16421 18906 -16387
rect 18962 -16421 18996 -16387
rect 19052 -16421 19086 -16387
rect 19260 -16421 19294 -16387
rect 19350 -16421 19384 -16387
rect 19440 -16421 19474 -16387
rect 19530 -16421 19564 -16387
rect 19620 -16421 19654 -16387
rect 19710 -16421 19744 -16387
rect 19800 -16421 19834 -16387
rect 19890 -16421 19924 -16387
rect 19980 -16421 20014 -16387
rect 20070 -16421 20104 -16387
rect 20160 -16421 20194 -16387
rect 20250 -16421 20284 -16387
rect 20340 -16421 20374 -16387
rect 20548 -16421 20582 -16387
rect 20638 -16421 20672 -16387
rect 20728 -16421 20762 -16387
rect 20818 -16421 20852 -16387
rect 20908 -16421 20942 -16387
rect 20998 -16421 21032 -16387
rect 21088 -16421 21122 -16387
rect 21178 -16421 21212 -16387
rect 21268 -16421 21302 -16387
rect 21358 -16421 21392 -16387
rect 21448 -16421 21482 -16387
rect 21538 -16421 21572 -16387
rect 21628 -16421 21662 -16387
rect 21836 -16421 21870 -16387
rect 21926 -16421 21960 -16387
rect 22016 -16421 22050 -16387
rect 22106 -16421 22140 -16387
rect 22196 -16421 22230 -16387
rect 22286 -16421 22320 -16387
rect 22376 -16421 22410 -16387
rect 22466 -16421 22500 -16387
rect 22556 -16421 22590 -16387
rect 22646 -16421 22680 -16387
rect 22736 -16421 22770 -16387
rect 22826 -16421 22860 -16387
rect 22916 -16421 22950 -16387
rect 23124 -16421 23158 -16387
rect 23214 -16421 23248 -16387
rect 23304 -16421 23338 -16387
rect 23394 -16421 23428 -16387
rect 23484 -16421 23518 -16387
rect 23574 -16421 23608 -16387
rect 23664 -16421 23698 -16387
rect 23754 -16421 23788 -16387
rect 23844 -16421 23878 -16387
rect 23934 -16421 23968 -16387
rect 24024 -16421 24058 -16387
rect 24114 -16421 24148 -16387
rect 24204 -16421 24238 -16387
rect 24412 -16421 24446 -16387
rect 24502 -16421 24536 -16387
rect 24592 -16421 24626 -16387
rect 24682 -16421 24716 -16387
rect 24772 -16421 24806 -16387
rect 24862 -16421 24896 -16387
rect 24952 -16421 24986 -16387
rect 25042 -16421 25076 -16387
rect 25132 -16421 25166 -16387
rect 25222 -16421 25256 -16387
rect 25312 -16421 25346 -16387
rect 25402 -16421 25436 -16387
rect 25492 -16421 25526 -16387
rect 25700 -16421 25734 -16387
rect 25790 -16421 25824 -16387
rect 25880 -16421 25914 -16387
rect 25970 -16421 26004 -16387
rect 26060 -16421 26094 -16387
rect 26150 -16421 26184 -16387
rect 26240 -16421 26274 -16387
rect 26330 -16421 26364 -16387
rect 26420 -16421 26454 -16387
rect 26510 -16421 26544 -16387
rect 26600 -16421 26634 -16387
rect 26690 -16421 26724 -16387
rect 26780 -16421 26814 -16387
rect 7302 -17050 13606 -16480
rect 16684 -16522 16718 -16488
rect 16774 -16522 16808 -16488
rect 16864 -16522 16898 -16488
rect 16954 -16522 16988 -16488
rect 17044 -16522 17078 -16488
rect 17134 -16522 17168 -16488
rect 17224 -16522 17258 -16488
rect 17314 -16522 17348 -16488
rect 17404 -16522 17438 -16488
rect 17494 -16522 17528 -16488
rect 17584 -16522 17618 -16488
rect 17674 -16522 17708 -16488
rect 17764 -16522 17798 -16488
rect 17972 -16522 18006 -16488
rect 18062 -16522 18096 -16488
rect 18152 -16522 18186 -16488
rect 18242 -16522 18276 -16488
rect 18332 -16522 18366 -16488
rect 18422 -16522 18456 -16488
rect 18512 -16522 18546 -16488
rect 18602 -16522 18636 -16488
rect 18692 -16522 18726 -16488
rect 18782 -16522 18816 -16488
rect 18872 -16522 18906 -16488
rect 18962 -16522 18996 -16488
rect 19052 -16522 19086 -16488
rect 19260 -16522 19294 -16488
rect 19350 -16522 19384 -16488
rect 19440 -16522 19474 -16488
rect 19530 -16522 19564 -16488
rect 19620 -16522 19654 -16488
rect 19710 -16522 19744 -16488
rect 19800 -16522 19834 -16488
rect 19890 -16522 19924 -16488
rect 19980 -16522 20014 -16488
rect 20070 -16522 20104 -16488
rect 20160 -16522 20194 -16488
rect 20250 -16522 20284 -16488
rect 20340 -16522 20374 -16488
rect 20548 -16522 20582 -16488
rect 20638 -16522 20672 -16488
rect 20728 -16522 20762 -16488
rect 20818 -16522 20852 -16488
rect 20908 -16522 20942 -16488
rect 20998 -16522 21032 -16488
rect 21088 -16522 21122 -16488
rect 21178 -16522 21212 -16488
rect 21268 -16522 21302 -16488
rect 21358 -16522 21392 -16488
rect 21448 -16522 21482 -16488
rect 21538 -16522 21572 -16488
rect 21628 -16522 21662 -16488
rect 21836 -16522 21870 -16488
rect 21926 -16522 21960 -16488
rect 22016 -16522 22050 -16488
rect 22106 -16522 22140 -16488
rect 22196 -16522 22230 -16488
rect 22286 -16522 22320 -16488
rect 22376 -16522 22410 -16488
rect 22466 -16522 22500 -16488
rect 22556 -16522 22590 -16488
rect 22646 -16522 22680 -16488
rect 22736 -16522 22770 -16488
rect 22826 -16522 22860 -16488
rect 22916 -16522 22950 -16488
rect 23124 -16522 23158 -16488
rect 23214 -16522 23248 -16488
rect 23304 -16522 23338 -16488
rect 23394 -16522 23428 -16488
rect 23484 -16522 23518 -16488
rect 23574 -16522 23608 -16488
rect 23664 -16522 23698 -16488
rect 23754 -16522 23788 -16488
rect 23844 -16522 23878 -16488
rect 23934 -16522 23968 -16488
rect 24024 -16522 24058 -16488
rect 24114 -16522 24148 -16488
rect 24204 -16522 24238 -16488
rect 24412 -16522 24446 -16488
rect 24502 -16522 24536 -16488
rect 24592 -16522 24626 -16488
rect 24682 -16522 24716 -16488
rect 24772 -16522 24806 -16488
rect 24862 -16522 24896 -16488
rect 24952 -16522 24986 -16488
rect 25042 -16522 25076 -16488
rect 25132 -16522 25166 -16488
rect 25222 -16522 25256 -16488
rect 25312 -16522 25346 -16488
rect 25402 -16522 25436 -16488
rect 25492 -16522 25526 -16488
rect 25700 -16522 25734 -16488
rect 25790 -16522 25824 -16488
rect 25880 -16522 25914 -16488
rect 25970 -16522 26004 -16488
rect 26060 -16522 26094 -16488
rect 26150 -16522 26184 -16488
rect 26240 -16522 26274 -16488
rect 26330 -16522 26364 -16488
rect 26420 -16522 26454 -16488
rect 26510 -16522 26544 -16488
rect 26600 -16522 26634 -16488
rect 26690 -16522 26724 -16488
rect 26780 -16522 26814 -16488
rect 16600 -16618 16634 -16584
rect 16600 -16708 16634 -16674
rect 16600 -16798 16634 -16764
rect 16600 -16888 16634 -16854
rect 16600 -16978 16634 -16944
rect 16600 -17068 16634 -17034
rect 16600 -17158 16634 -17124
rect 16600 -17248 16634 -17214
rect 16600 -17338 16634 -17304
rect 16600 -17428 16634 -17394
rect 16600 -17518 16634 -17484
rect 16600 -17608 16634 -17574
rect 17787 -16618 17821 -16584
rect 17888 -16618 17922 -16584
rect 17787 -16708 17821 -16674
rect 17888 -16708 17922 -16674
rect 17787 -16798 17821 -16764
rect 17888 -16798 17922 -16764
rect 17787 -16888 17821 -16854
rect 17888 -16888 17922 -16854
rect 17787 -16978 17821 -16944
rect 17888 -16978 17922 -16944
rect 17787 -17068 17821 -17034
rect 17888 -17068 17922 -17034
rect 17787 -17158 17821 -17124
rect 17888 -17158 17922 -17124
rect 17787 -17248 17821 -17214
rect 17888 -17248 17922 -17214
rect 17787 -17338 17821 -17304
rect 17888 -17338 17922 -17304
rect 17787 -17428 17821 -17394
rect 17888 -17428 17922 -17394
rect 17787 -17518 17821 -17484
rect 17888 -17518 17922 -17484
rect 17787 -17608 17821 -17574
rect 17888 -17608 17922 -17574
rect 19075 -16618 19109 -16584
rect 19176 -16618 19210 -16584
rect 19075 -16708 19109 -16674
rect 19176 -16708 19210 -16674
rect 19075 -16798 19109 -16764
rect 19176 -16798 19210 -16764
rect 19075 -16888 19109 -16854
rect 19176 -16888 19210 -16854
rect 19075 -16978 19109 -16944
rect 19176 -16978 19210 -16944
rect 19075 -17068 19109 -17034
rect 19176 -17068 19210 -17034
rect 19075 -17158 19109 -17124
rect 19176 -17158 19210 -17124
rect 19075 -17248 19109 -17214
rect 19176 -17248 19210 -17214
rect 19075 -17338 19109 -17304
rect 19176 -17338 19210 -17304
rect 19075 -17428 19109 -17394
rect 19176 -17428 19210 -17394
rect 19075 -17518 19109 -17484
rect 19176 -17518 19210 -17484
rect 19075 -17608 19109 -17574
rect 19176 -17608 19210 -17574
rect 20363 -16618 20397 -16584
rect 20464 -16618 20498 -16584
rect 20363 -16708 20397 -16674
rect 20464 -16708 20498 -16674
rect 20363 -16798 20397 -16764
rect 20464 -16798 20498 -16764
rect 20363 -16888 20397 -16854
rect 20464 -16888 20498 -16854
rect 20363 -16978 20397 -16944
rect 20464 -16978 20498 -16944
rect 20363 -17068 20397 -17034
rect 20464 -17068 20498 -17034
rect 20363 -17158 20397 -17124
rect 20464 -17158 20498 -17124
rect 20363 -17248 20397 -17214
rect 20464 -17248 20498 -17214
rect 20363 -17338 20397 -17304
rect 20464 -17338 20498 -17304
rect 20363 -17428 20397 -17394
rect 20464 -17428 20498 -17394
rect 20363 -17518 20397 -17484
rect 20464 -17518 20498 -17484
rect 20363 -17608 20397 -17574
rect 20464 -17608 20498 -17574
rect 21651 -16618 21685 -16584
rect 21752 -16618 21786 -16584
rect 21651 -16708 21685 -16674
rect 21752 -16708 21786 -16674
rect 21651 -16798 21685 -16764
rect 21752 -16798 21786 -16764
rect 21651 -16888 21685 -16854
rect 21752 -16888 21786 -16854
rect 21651 -16978 21685 -16944
rect 21752 -16978 21786 -16944
rect 21651 -17068 21685 -17034
rect 21752 -17068 21786 -17034
rect 21651 -17158 21685 -17124
rect 21752 -17158 21786 -17124
rect 21651 -17248 21685 -17214
rect 21752 -17248 21786 -17214
rect 21651 -17338 21685 -17304
rect 21752 -17338 21786 -17304
rect 21651 -17428 21685 -17394
rect 21752 -17428 21786 -17394
rect 21651 -17518 21685 -17484
rect 21752 -17518 21786 -17484
rect 21651 -17608 21685 -17574
rect 21752 -17608 21786 -17574
rect 22939 -16618 22973 -16584
rect 23040 -16618 23074 -16584
rect 22939 -16708 22973 -16674
rect 23040 -16708 23074 -16674
rect 22939 -16798 22973 -16764
rect 23040 -16798 23074 -16764
rect 22939 -16888 22973 -16854
rect 23040 -16888 23074 -16854
rect 22939 -16978 22973 -16944
rect 23040 -16978 23074 -16944
rect 22939 -17068 22973 -17034
rect 23040 -17068 23074 -17034
rect 22939 -17158 22973 -17124
rect 23040 -17158 23074 -17124
rect 22939 -17248 22973 -17214
rect 23040 -17248 23074 -17214
rect 22939 -17338 22973 -17304
rect 23040 -17338 23074 -17304
rect 22939 -17428 22973 -17394
rect 23040 -17428 23074 -17394
rect 22939 -17518 22973 -17484
rect 23040 -17518 23074 -17484
rect 22939 -17608 22973 -17574
rect 23040 -17608 23074 -17574
rect 24227 -16618 24261 -16584
rect 24328 -16618 24362 -16584
rect 24227 -16708 24261 -16674
rect 24328 -16708 24362 -16674
rect 24227 -16798 24261 -16764
rect 24328 -16798 24362 -16764
rect 24227 -16888 24261 -16854
rect 24328 -16888 24362 -16854
rect 24227 -16978 24261 -16944
rect 24328 -16978 24362 -16944
rect 24227 -17068 24261 -17034
rect 24328 -17068 24362 -17034
rect 24227 -17158 24261 -17124
rect 24328 -17158 24362 -17124
rect 24227 -17248 24261 -17214
rect 24328 -17248 24362 -17214
rect 24227 -17338 24261 -17304
rect 24328 -17338 24362 -17304
rect 24227 -17428 24261 -17394
rect 24328 -17428 24362 -17394
rect 24227 -17518 24261 -17484
rect 24328 -17518 24362 -17484
rect 24227 -17608 24261 -17574
rect 24328 -17608 24362 -17574
rect 25515 -16618 25549 -16584
rect 25616 -16618 25650 -16584
rect 25515 -16708 25549 -16674
rect 25616 -16708 25650 -16674
rect 25515 -16798 25549 -16764
rect 25616 -16798 25650 -16764
rect 25515 -16888 25549 -16854
rect 25616 -16888 25650 -16854
rect 25515 -16978 25549 -16944
rect 25616 -16978 25650 -16944
rect 25515 -17068 25549 -17034
rect 25616 -17068 25650 -17034
rect 25515 -17158 25549 -17124
rect 25616 -17158 25650 -17124
rect 25515 -17248 25549 -17214
rect 25616 -17248 25650 -17214
rect 25515 -17338 25549 -17304
rect 25616 -17338 25650 -17304
rect 25515 -17428 25549 -17394
rect 25616 -17428 25650 -17394
rect 25515 -17518 25549 -17484
rect 25616 -17518 25650 -17484
rect 25515 -17608 25549 -17574
rect 25616 -17608 25650 -17574
rect 26803 -16618 26837 -16584
rect 26803 -16708 26837 -16674
rect 26803 -16798 26837 -16764
rect 26803 -16888 26837 -16854
rect 26803 -16978 26837 -16944
rect 26803 -17068 26837 -17034
rect 26803 -17158 26837 -17124
rect 26803 -17248 26837 -17214
rect 26803 -17338 26837 -17304
rect 26803 -17428 26837 -17394
rect 26803 -17518 26837 -17484
rect 26803 -17608 26837 -17574
rect 16684 -17709 16718 -17675
rect 16774 -17709 16808 -17675
rect 16864 -17709 16898 -17675
rect 16954 -17709 16988 -17675
rect 17044 -17709 17078 -17675
rect 17134 -17709 17168 -17675
rect 17224 -17709 17258 -17675
rect 17314 -17709 17348 -17675
rect 17404 -17709 17438 -17675
rect 17494 -17709 17528 -17675
rect 17584 -17709 17618 -17675
rect 17674 -17709 17708 -17675
rect 17764 -17709 17798 -17675
rect 17972 -17709 18006 -17675
rect 18062 -17709 18096 -17675
rect 18152 -17709 18186 -17675
rect 18242 -17709 18276 -17675
rect 18332 -17709 18366 -17675
rect 18422 -17709 18456 -17675
rect 18512 -17709 18546 -17675
rect 18602 -17709 18636 -17675
rect 18692 -17709 18726 -17675
rect 18782 -17709 18816 -17675
rect 18872 -17709 18906 -17675
rect 18962 -17709 18996 -17675
rect 19052 -17709 19086 -17675
rect 19260 -17709 19294 -17675
rect 19350 -17709 19384 -17675
rect 19440 -17709 19474 -17675
rect 19530 -17709 19564 -17675
rect 19620 -17709 19654 -17675
rect 19710 -17709 19744 -17675
rect 19800 -17709 19834 -17675
rect 19890 -17709 19924 -17675
rect 19980 -17709 20014 -17675
rect 20070 -17709 20104 -17675
rect 20160 -17709 20194 -17675
rect 20250 -17709 20284 -17675
rect 20340 -17709 20374 -17675
rect 20548 -17709 20582 -17675
rect 20638 -17709 20672 -17675
rect 20728 -17709 20762 -17675
rect 20818 -17709 20852 -17675
rect 20908 -17709 20942 -17675
rect 20998 -17709 21032 -17675
rect 21088 -17709 21122 -17675
rect 21178 -17709 21212 -17675
rect 21268 -17709 21302 -17675
rect 21358 -17709 21392 -17675
rect 21448 -17709 21482 -17675
rect 21538 -17709 21572 -17675
rect 21628 -17709 21662 -17675
rect 21836 -17709 21870 -17675
rect 21926 -17709 21960 -17675
rect 22016 -17709 22050 -17675
rect 22106 -17709 22140 -17675
rect 22196 -17709 22230 -17675
rect 22286 -17709 22320 -17675
rect 22376 -17709 22410 -17675
rect 22466 -17709 22500 -17675
rect 22556 -17709 22590 -17675
rect 22646 -17709 22680 -17675
rect 22736 -17709 22770 -17675
rect 22826 -17709 22860 -17675
rect 22916 -17709 22950 -17675
rect 23124 -17709 23158 -17675
rect 23214 -17709 23248 -17675
rect 23304 -17709 23338 -17675
rect 23394 -17709 23428 -17675
rect 23484 -17709 23518 -17675
rect 23574 -17709 23608 -17675
rect 23664 -17709 23698 -17675
rect 23754 -17709 23788 -17675
rect 23844 -17709 23878 -17675
rect 23934 -17709 23968 -17675
rect 24024 -17709 24058 -17675
rect 24114 -17709 24148 -17675
rect 24204 -17709 24238 -17675
rect 24412 -17709 24446 -17675
rect 24502 -17709 24536 -17675
rect 24592 -17709 24626 -17675
rect 24682 -17709 24716 -17675
rect 24772 -17709 24806 -17675
rect 24862 -17709 24896 -17675
rect 24952 -17709 24986 -17675
rect 25042 -17709 25076 -17675
rect 25132 -17709 25166 -17675
rect 25222 -17709 25256 -17675
rect 25312 -17709 25346 -17675
rect 25402 -17709 25436 -17675
rect 25492 -17709 25526 -17675
rect 25700 -17709 25734 -17675
rect 25790 -17709 25824 -17675
rect 25880 -17709 25914 -17675
rect 25970 -17709 26004 -17675
rect 26060 -17709 26094 -17675
rect 26150 -17709 26184 -17675
rect 26240 -17709 26274 -17675
rect 26330 -17709 26364 -17675
rect 26420 -17709 26454 -17675
rect 26510 -17709 26544 -17675
rect 26600 -17709 26634 -17675
rect 26690 -17709 26724 -17675
rect 26780 -17709 26814 -17675
rect 7302 -31738 13606 -31168
rect 7302 -36698 13606 -36128
rect 7302 -39942 13606 -39372
<< nsubdiffcont >>
rect 16863 -11518 16897 -11484
rect 16953 -11518 16987 -11484
rect 17043 -11518 17077 -11484
rect 17133 -11518 17167 -11484
rect 17223 -11518 17257 -11484
rect 17313 -11518 17347 -11484
rect 17403 -11518 17437 -11484
rect 17493 -11518 17527 -11484
rect 17583 -11518 17617 -11484
rect 16750 -11596 16784 -11562
rect 16750 -11686 16784 -11652
rect 16750 -11776 16784 -11742
rect 16750 -11866 16784 -11832
rect 16750 -11956 16784 -11922
rect 16750 -12046 16784 -12012
rect 16750 -12136 16784 -12102
rect 16750 -12226 16784 -12192
rect 16750 -12316 16784 -12282
rect 17640 -11630 17674 -11596
rect 17640 -11720 17674 -11686
rect 17640 -11810 17674 -11776
rect 17640 -11900 17674 -11866
rect 17640 -11990 17674 -11956
rect 17640 -12080 17674 -12046
rect 17640 -12170 17674 -12136
rect 17640 -12260 17674 -12226
rect 17640 -12350 17674 -12316
rect 16844 -12408 16878 -12374
rect 16934 -12408 16968 -12374
rect 17024 -12408 17058 -12374
rect 17114 -12408 17148 -12374
rect 17204 -12408 17238 -12374
rect 17294 -12408 17328 -12374
rect 17384 -12408 17418 -12374
rect 17474 -12408 17508 -12374
rect 17564 -12408 17598 -12374
rect 18151 -11518 18185 -11484
rect 18241 -11518 18275 -11484
rect 18331 -11518 18365 -11484
rect 18421 -11518 18455 -11484
rect 18511 -11518 18545 -11484
rect 18601 -11518 18635 -11484
rect 18691 -11518 18725 -11484
rect 18781 -11518 18815 -11484
rect 18871 -11518 18905 -11484
rect 18038 -11596 18072 -11562
rect 18038 -11686 18072 -11652
rect 18038 -11776 18072 -11742
rect 18038 -11866 18072 -11832
rect 18038 -11956 18072 -11922
rect 18038 -12046 18072 -12012
rect 18038 -12136 18072 -12102
rect 18038 -12226 18072 -12192
rect 18038 -12316 18072 -12282
rect 18928 -11630 18962 -11596
rect 18928 -11720 18962 -11686
rect 18928 -11810 18962 -11776
rect 18928 -11900 18962 -11866
rect 18928 -11990 18962 -11956
rect 18928 -12080 18962 -12046
rect 18928 -12170 18962 -12136
rect 18928 -12260 18962 -12226
rect 18928 -12350 18962 -12316
rect 18132 -12408 18166 -12374
rect 18222 -12408 18256 -12374
rect 18312 -12408 18346 -12374
rect 18402 -12408 18436 -12374
rect 18492 -12408 18526 -12374
rect 18582 -12408 18616 -12374
rect 18672 -12408 18706 -12374
rect 18762 -12408 18796 -12374
rect 18852 -12408 18886 -12374
rect 19439 -11518 19473 -11484
rect 19529 -11518 19563 -11484
rect 19619 -11518 19653 -11484
rect 19709 -11518 19743 -11484
rect 19799 -11518 19833 -11484
rect 19889 -11518 19923 -11484
rect 19979 -11518 20013 -11484
rect 20069 -11518 20103 -11484
rect 20159 -11518 20193 -11484
rect 19326 -11596 19360 -11562
rect 19326 -11686 19360 -11652
rect 19326 -11776 19360 -11742
rect 19326 -11866 19360 -11832
rect 19326 -11956 19360 -11922
rect 19326 -12046 19360 -12012
rect 19326 -12136 19360 -12102
rect 19326 -12226 19360 -12192
rect 19326 -12316 19360 -12282
rect 20216 -11630 20250 -11596
rect 20216 -11720 20250 -11686
rect 20216 -11810 20250 -11776
rect 20216 -11900 20250 -11866
rect 20216 -11990 20250 -11956
rect 20216 -12080 20250 -12046
rect 20216 -12170 20250 -12136
rect 20216 -12260 20250 -12226
rect 20216 -12350 20250 -12316
rect 19420 -12408 19454 -12374
rect 19510 -12408 19544 -12374
rect 19600 -12408 19634 -12374
rect 19690 -12408 19724 -12374
rect 19780 -12408 19814 -12374
rect 19870 -12408 19904 -12374
rect 19960 -12408 19994 -12374
rect 20050 -12408 20084 -12374
rect 20140 -12408 20174 -12374
rect 20727 -11518 20761 -11484
rect 20817 -11518 20851 -11484
rect 20907 -11518 20941 -11484
rect 20997 -11518 21031 -11484
rect 21087 -11518 21121 -11484
rect 21177 -11518 21211 -11484
rect 21267 -11518 21301 -11484
rect 21357 -11518 21391 -11484
rect 21447 -11518 21481 -11484
rect 20614 -11596 20648 -11562
rect 20614 -11686 20648 -11652
rect 20614 -11776 20648 -11742
rect 20614 -11866 20648 -11832
rect 20614 -11956 20648 -11922
rect 20614 -12046 20648 -12012
rect 20614 -12136 20648 -12102
rect 20614 -12226 20648 -12192
rect 20614 -12316 20648 -12282
rect 21504 -11630 21538 -11596
rect 21504 -11720 21538 -11686
rect 21504 -11810 21538 -11776
rect 21504 -11900 21538 -11866
rect 21504 -11990 21538 -11956
rect 21504 -12080 21538 -12046
rect 21504 -12170 21538 -12136
rect 21504 -12260 21538 -12226
rect 21504 -12350 21538 -12316
rect 20708 -12408 20742 -12374
rect 20798 -12408 20832 -12374
rect 20888 -12408 20922 -12374
rect 20978 -12408 21012 -12374
rect 21068 -12408 21102 -12374
rect 21158 -12408 21192 -12374
rect 21248 -12408 21282 -12374
rect 21338 -12408 21372 -12374
rect 21428 -12408 21462 -12374
rect 22015 -11518 22049 -11484
rect 22105 -11518 22139 -11484
rect 22195 -11518 22229 -11484
rect 22285 -11518 22319 -11484
rect 22375 -11518 22409 -11484
rect 22465 -11518 22499 -11484
rect 22555 -11518 22589 -11484
rect 22645 -11518 22679 -11484
rect 22735 -11518 22769 -11484
rect 21902 -11596 21936 -11562
rect 21902 -11686 21936 -11652
rect 21902 -11776 21936 -11742
rect 21902 -11866 21936 -11832
rect 21902 -11956 21936 -11922
rect 21902 -12046 21936 -12012
rect 21902 -12136 21936 -12102
rect 21902 -12226 21936 -12192
rect 21902 -12316 21936 -12282
rect 22792 -11630 22826 -11596
rect 22792 -11720 22826 -11686
rect 22792 -11810 22826 -11776
rect 22792 -11900 22826 -11866
rect 22792 -11990 22826 -11956
rect 22792 -12080 22826 -12046
rect 22792 -12170 22826 -12136
rect 22792 -12260 22826 -12226
rect 22792 -12350 22826 -12316
rect 21996 -12408 22030 -12374
rect 22086 -12408 22120 -12374
rect 22176 -12408 22210 -12374
rect 22266 -12408 22300 -12374
rect 22356 -12408 22390 -12374
rect 22446 -12408 22480 -12374
rect 22536 -12408 22570 -12374
rect 22626 -12408 22660 -12374
rect 22716 -12408 22750 -12374
rect 23303 -11518 23337 -11484
rect 23393 -11518 23427 -11484
rect 23483 -11518 23517 -11484
rect 23573 -11518 23607 -11484
rect 23663 -11518 23697 -11484
rect 23753 -11518 23787 -11484
rect 23843 -11518 23877 -11484
rect 23933 -11518 23967 -11484
rect 24023 -11518 24057 -11484
rect 23190 -11596 23224 -11562
rect 23190 -11686 23224 -11652
rect 23190 -11776 23224 -11742
rect 23190 -11866 23224 -11832
rect 23190 -11956 23224 -11922
rect 23190 -12046 23224 -12012
rect 23190 -12136 23224 -12102
rect 23190 -12226 23224 -12192
rect 23190 -12316 23224 -12282
rect 24080 -11630 24114 -11596
rect 24080 -11720 24114 -11686
rect 24080 -11810 24114 -11776
rect 24080 -11900 24114 -11866
rect 24080 -11990 24114 -11956
rect 24080 -12080 24114 -12046
rect 24080 -12170 24114 -12136
rect 24080 -12260 24114 -12226
rect 24080 -12350 24114 -12316
rect 23284 -12408 23318 -12374
rect 23374 -12408 23408 -12374
rect 23464 -12408 23498 -12374
rect 23554 -12408 23588 -12374
rect 23644 -12408 23678 -12374
rect 23734 -12408 23768 -12374
rect 23824 -12408 23858 -12374
rect 23914 -12408 23948 -12374
rect 24004 -12408 24038 -12374
rect 24591 -11518 24625 -11484
rect 24681 -11518 24715 -11484
rect 24771 -11518 24805 -11484
rect 24861 -11518 24895 -11484
rect 24951 -11518 24985 -11484
rect 25041 -11518 25075 -11484
rect 25131 -11518 25165 -11484
rect 25221 -11518 25255 -11484
rect 25311 -11518 25345 -11484
rect 24478 -11596 24512 -11562
rect 24478 -11686 24512 -11652
rect 24478 -11776 24512 -11742
rect 24478 -11866 24512 -11832
rect 24478 -11956 24512 -11922
rect 24478 -12046 24512 -12012
rect 24478 -12136 24512 -12102
rect 24478 -12226 24512 -12192
rect 24478 -12316 24512 -12282
rect 25368 -11630 25402 -11596
rect 25368 -11720 25402 -11686
rect 25368 -11810 25402 -11776
rect 25368 -11900 25402 -11866
rect 25368 -11990 25402 -11956
rect 25368 -12080 25402 -12046
rect 25368 -12170 25402 -12136
rect 25368 -12260 25402 -12226
rect 25368 -12350 25402 -12316
rect 24572 -12408 24606 -12374
rect 24662 -12408 24696 -12374
rect 24752 -12408 24786 -12374
rect 24842 -12408 24876 -12374
rect 24932 -12408 24966 -12374
rect 25022 -12408 25056 -12374
rect 25112 -12408 25146 -12374
rect 25202 -12408 25236 -12374
rect 25292 -12408 25326 -12374
rect 25879 -11518 25913 -11484
rect 25969 -11518 26003 -11484
rect 26059 -11518 26093 -11484
rect 26149 -11518 26183 -11484
rect 26239 -11518 26273 -11484
rect 26329 -11518 26363 -11484
rect 26419 -11518 26453 -11484
rect 26509 -11518 26543 -11484
rect 26599 -11518 26633 -11484
rect 25766 -11596 25800 -11562
rect 25766 -11686 25800 -11652
rect 25766 -11776 25800 -11742
rect 25766 -11866 25800 -11832
rect 25766 -11956 25800 -11922
rect 25766 -12046 25800 -12012
rect 25766 -12136 25800 -12102
rect 25766 -12226 25800 -12192
rect 25766 -12316 25800 -12282
rect 26656 -11630 26690 -11596
rect 26656 -11720 26690 -11686
rect 26656 -11810 26690 -11776
rect 26656 -11900 26690 -11866
rect 26656 -11990 26690 -11956
rect 26656 -12080 26690 -12046
rect 26656 -12170 26690 -12136
rect 26656 -12260 26690 -12226
rect 26656 -12350 26690 -12316
rect 25860 -12408 25894 -12374
rect 25950 -12408 25984 -12374
rect 26040 -12408 26074 -12374
rect 26130 -12408 26164 -12374
rect 26220 -12408 26254 -12374
rect 26310 -12408 26344 -12374
rect 26400 -12408 26434 -12374
rect 26490 -12408 26524 -12374
rect 26580 -12408 26614 -12374
rect 16863 -12806 16897 -12772
rect 16953 -12806 16987 -12772
rect 17043 -12806 17077 -12772
rect 17133 -12806 17167 -12772
rect 17223 -12806 17257 -12772
rect 17313 -12806 17347 -12772
rect 17403 -12806 17437 -12772
rect 17493 -12806 17527 -12772
rect 17583 -12806 17617 -12772
rect 16750 -12884 16784 -12850
rect 16750 -12974 16784 -12940
rect 16750 -13064 16784 -13030
rect 16750 -13154 16784 -13120
rect 16750 -13244 16784 -13210
rect 16750 -13334 16784 -13300
rect 16750 -13424 16784 -13390
rect 16750 -13514 16784 -13480
rect 16750 -13604 16784 -13570
rect 17640 -12918 17674 -12884
rect 17640 -13008 17674 -12974
rect 17640 -13098 17674 -13064
rect 17640 -13188 17674 -13154
rect 17640 -13278 17674 -13244
rect 17640 -13368 17674 -13334
rect 17640 -13458 17674 -13424
rect 17640 -13548 17674 -13514
rect 17640 -13638 17674 -13604
rect 16844 -13696 16878 -13662
rect 16934 -13696 16968 -13662
rect 17024 -13696 17058 -13662
rect 17114 -13696 17148 -13662
rect 17204 -13696 17238 -13662
rect 17294 -13696 17328 -13662
rect 17384 -13696 17418 -13662
rect 17474 -13696 17508 -13662
rect 17564 -13696 17598 -13662
rect 18151 -12806 18185 -12772
rect 18241 -12806 18275 -12772
rect 18331 -12806 18365 -12772
rect 18421 -12806 18455 -12772
rect 18511 -12806 18545 -12772
rect 18601 -12806 18635 -12772
rect 18691 -12806 18725 -12772
rect 18781 -12806 18815 -12772
rect 18871 -12806 18905 -12772
rect 18038 -12884 18072 -12850
rect 18038 -12974 18072 -12940
rect 18038 -13064 18072 -13030
rect 18038 -13154 18072 -13120
rect 18038 -13244 18072 -13210
rect 18038 -13334 18072 -13300
rect 18038 -13424 18072 -13390
rect 18038 -13514 18072 -13480
rect 18038 -13604 18072 -13570
rect 18928 -12918 18962 -12884
rect 18928 -13008 18962 -12974
rect 18928 -13098 18962 -13064
rect 18928 -13188 18962 -13154
rect 18928 -13278 18962 -13244
rect 18928 -13368 18962 -13334
rect 18928 -13458 18962 -13424
rect 18928 -13548 18962 -13514
rect 18928 -13638 18962 -13604
rect 18132 -13696 18166 -13662
rect 18222 -13696 18256 -13662
rect 18312 -13696 18346 -13662
rect 18402 -13696 18436 -13662
rect 18492 -13696 18526 -13662
rect 18582 -13696 18616 -13662
rect 18672 -13696 18706 -13662
rect 18762 -13696 18796 -13662
rect 18852 -13696 18886 -13662
rect 19439 -12806 19473 -12772
rect 19529 -12806 19563 -12772
rect 19619 -12806 19653 -12772
rect 19709 -12806 19743 -12772
rect 19799 -12806 19833 -12772
rect 19889 -12806 19923 -12772
rect 19979 -12806 20013 -12772
rect 20069 -12806 20103 -12772
rect 20159 -12806 20193 -12772
rect 19326 -12884 19360 -12850
rect 19326 -12974 19360 -12940
rect 19326 -13064 19360 -13030
rect 19326 -13154 19360 -13120
rect 19326 -13244 19360 -13210
rect 19326 -13334 19360 -13300
rect 19326 -13424 19360 -13390
rect 19326 -13514 19360 -13480
rect 19326 -13604 19360 -13570
rect 20216 -12918 20250 -12884
rect 20216 -13008 20250 -12974
rect 20216 -13098 20250 -13064
rect 20216 -13188 20250 -13154
rect 20216 -13278 20250 -13244
rect 20216 -13368 20250 -13334
rect 20216 -13458 20250 -13424
rect 20216 -13548 20250 -13514
rect 20216 -13638 20250 -13604
rect 19420 -13696 19454 -13662
rect 19510 -13696 19544 -13662
rect 19600 -13696 19634 -13662
rect 19690 -13696 19724 -13662
rect 19780 -13696 19814 -13662
rect 19870 -13696 19904 -13662
rect 19960 -13696 19994 -13662
rect 20050 -13696 20084 -13662
rect 20140 -13696 20174 -13662
rect 20727 -12806 20761 -12772
rect 20817 -12806 20851 -12772
rect 20907 -12806 20941 -12772
rect 20997 -12806 21031 -12772
rect 21087 -12806 21121 -12772
rect 21177 -12806 21211 -12772
rect 21267 -12806 21301 -12772
rect 21357 -12806 21391 -12772
rect 21447 -12806 21481 -12772
rect 20614 -12884 20648 -12850
rect 20614 -12974 20648 -12940
rect 20614 -13064 20648 -13030
rect 20614 -13154 20648 -13120
rect 20614 -13244 20648 -13210
rect 20614 -13334 20648 -13300
rect 20614 -13424 20648 -13390
rect 20614 -13514 20648 -13480
rect 20614 -13604 20648 -13570
rect 21504 -12918 21538 -12884
rect 21504 -13008 21538 -12974
rect 21504 -13098 21538 -13064
rect 21504 -13188 21538 -13154
rect 21504 -13278 21538 -13244
rect 21504 -13368 21538 -13334
rect 21504 -13458 21538 -13424
rect 21504 -13548 21538 -13514
rect 21504 -13638 21538 -13604
rect 20708 -13696 20742 -13662
rect 20798 -13696 20832 -13662
rect 20888 -13696 20922 -13662
rect 20978 -13696 21012 -13662
rect 21068 -13696 21102 -13662
rect 21158 -13696 21192 -13662
rect 21248 -13696 21282 -13662
rect 21338 -13696 21372 -13662
rect 21428 -13696 21462 -13662
rect 22015 -12806 22049 -12772
rect 22105 -12806 22139 -12772
rect 22195 -12806 22229 -12772
rect 22285 -12806 22319 -12772
rect 22375 -12806 22409 -12772
rect 22465 -12806 22499 -12772
rect 22555 -12806 22589 -12772
rect 22645 -12806 22679 -12772
rect 22735 -12806 22769 -12772
rect 21902 -12884 21936 -12850
rect 21902 -12974 21936 -12940
rect 21902 -13064 21936 -13030
rect 21902 -13154 21936 -13120
rect 21902 -13244 21936 -13210
rect 21902 -13334 21936 -13300
rect 21902 -13424 21936 -13390
rect 21902 -13514 21936 -13480
rect 21902 -13604 21936 -13570
rect 22792 -12918 22826 -12884
rect 22792 -13008 22826 -12974
rect 22792 -13098 22826 -13064
rect 22792 -13188 22826 -13154
rect 22792 -13278 22826 -13244
rect 22792 -13368 22826 -13334
rect 22792 -13458 22826 -13424
rect 22792 -13548 22826 -13514
rect 22792 -13638 22826 -13604
rect 21996 -13696 22030 -13662
rect 22086 -13696 22120 -13662
rect 22176 -13696 22210 -13662
rect 22266 -13696 22300 -13662
rect 22356 -13696 22390 -13662
rect 22446 -13696 22480 -13662
rect 22536 -13696 22570 -13662
rect 22626 -13696 22660 -13662
rect 22716 -13696 22750 -13662
rect 23303 -12806 23337 -12772
rect 23393 -12806 23427 -12772
rect 23483 -12806 23517 -12772
rect 23573 -12806 23607 -12772
rect 23663 -12806 23697 -12772
rect 23753 -12806 23787 -12772
rect 23843 -12806 23877 -12772
rect 23933 -12806 23967 -12772
rect 24023 -12806 24057 -12772
rect 23190 -12884 23224 -12850
rect 23190 -12974 23224 -12940
rect 23190 -13064 23224 -13030
rect 23190 -13154 23224 -13120
rect 23190 -13244 23224 -13210
rect 23190 -13334 23224 -13300
rect 23190 -13424 23224 -13390
rect 23190 -13514 23224 -13480
rect 23190 -13604 23224 -13570
rect 24080 -12918 24114 -12884
rect 24080 -13008 24114 -12974
rect 24080 -13098 24114 -13064
rect 24080 -13188 24114 -13154
rect 24080 -13278 24114 -13244
rect 24080 -13368 24114 -13334
rect 24080 -13458 24114 -13424
rect 24080 -13548 24114 -13514
rect 24080 -13638 24114 -13604
rect 23284 -13696 23318 -13662
rect 23374 -13696 23408 -13662
rect 23464 -13696 23498 -13662
rect 23554 -13696 23588 -13662
rect 23644 -13696 23678 -13662
rect 23734 -13696 23768 -13662
rect 23824 -13696 23858 -13662
rect 23914 -13696 23948 -13662
rect 24004 -13696 24038 -13662
rect 24591 -12806 24625 -12772
rect 24681 -12806 24715 -12772
rect 24771 -12806 24805 -12772
rect 24861 -12806 24895 -12772
rect 24951 -12806 24985 -12772
rect 25041 -12806 25075 -12772
rect 25131 -12806 25165 -12772
rect 25221 -12806 25255 -12772
rect 25311 -12806 25345 -12772
rect 24478 -12884 24512 -12850
rect 24478 -12974 24512 -12940
rect 24478 -13064 24512 -13030
rect 24478 -13154 24512 -13120
rect 24478 -13244 24512 -13210
rect 24478 -13334 24512 -13300
rect 24478 -13424 24512 -13390
rect 24478 -13514 24512 -13480
rect 24478 -13604 24512 -13570
rect 25368 -12918 25402 -12884
rect 25368 -13008 25402 -12974
rect 25368 -13098 25402 -13064
rect 25368 -13188 25402 -13154
rect 25368 -13278 25402 -13244
rect 25368 -13368 25402 -13334
rect 25368 -13458 25402 -13424
rect 25368 -13548 25402 -13514
rect 25368 -13638 25402 -13604
rect 24572 -13696 24606 -13662
rect 24662 -13696 24696 -13662
rect 24752 -13696 24786 -13662
rect 24842 -13696 24876 -13662
rect 24932 -13696 24966 -13662
rect 25022 -13696 25056 -13662
rect 25112 -13696 25146 -13662
rect 25202 -13696 25236 -13662
rect 25292 -13696 25326 -13662
rect 25879 -12806 25913 -12772
rect 25969 -12806 26003 -12772
rect 26059 -12806 26093 -12772
rect 26149 -12806 26183 -12772
rect 26239 -12806 26273 -12772
rect 26329 -12806 26363 -12772
rect 26419 -12806 26453 -12772
rect 26509 -12806 26543 -12772
rect 26599 -12806 26633 -12772
rect 25766 -12884 25800 -12850
rect 25766 -12974 25800 -12940
rect 25766 -13064 25800 -13030
rect 25766 -13154 25800 -13120
rect 25766 -13244 25800 -13210
rect 25766 -13334 25800 -13300
rect 25766 -13424 25800 -13390
rect 25766 -13514 25800 -13480
rect 25766 -13604 25800 -13570
rect 26656 -12918 26690 -12884
rect 26656 -13008 26690 -12974
rect 26656 -13098 26690 -13064
rect 26656 -13188 26690 -13154
rect 26656 -13278 26690 -13244
rect 26656 -13368 26690 -13334
rect 26656 -13458 26690 -13424
rect 26656 -13548 26690 -13514
rect 26656 -13638 26690 -13604
rect 25860 -13696 25894 -13662
rect 25950 -13696 25984 -13662
rect 26040 -13696 26074 -13662
rect 26130 -13696 26164 -13662
rect 26220 -13696 26254 -13662
rect 26310 -13696 26344 -13662
rect 26400 -13696 26434 -13662
rect 26490 -13696 26524 -13662
rect 26580 -13696 26614 -13662
rect 16863 -14094 16897 -14060
rect 16953 -14094 16987 -14060
rect 17043 -14094 17077 -14060
rect 17133 -14094 17167 -14060
rect 17223 -14094 17257 -14060
rect 17313 -14094 17347 -14060
rect 17403 -14094 17437 -14060
rect 17493 -14094 17527 -14060
rect 17583 -14094 17617 -14060
rect 16750 -14172 16784 -14138
rect 16750 -14262 16784 -14228
rect 16750 -14352 16784 -14318
rect 16750 -14442 16784 -14408
rect 16750 -14532 16784 -14498
rect 16750 -14622 16784 -14588
rect 16750 -14712 16784 -14678
rect 16750 -14802 16784 -14768
rect 16750 -14892 16784 -14858
rect 17640 -14206 17674 -14172
rect 17640 -14296 17674 -14262
rect 17640 -14386 17674 -14352
rect 17640 -14476 17674 -14442
rect 17640 -14566 17674 -14532
rect 17640 -14656 17674 -14622
rect 17640 -14746 17674 -14712
rect 17640 -14836 17674 -14802
rect 17640 -14926 17674 -14892
rect 16844 -14984 16878 -14950
rect 16934 -14984 16968 -14950
rect 17024 -14984 17058 -14950
rect 17114 -14984 17148 -14950
rect 17204 -14984 17238 -14950
rect 17294 -14984 17328 -14950
rect 17384 -14984 17418 -14950
rect 17474 -14984 17508 -14950
rect 17564 -14984 17598 -14950
rect 18151 -14094 18185 -14060
rect 18241 -14094 18275 -14060
rect 18331 -14094 18365 -14060
rect 18421 -14094 18455 -14060
rect 18511 -14094 18545 -14060
rect 18601 -14094 18635 -14060
rect 18691 -14094 18725 -14060
rect 18781 -14094 18815 -14060
rect 18871 -14094 18905 -14060
rect 18038 -14172 18072 -14138
rect 18038 -14262 18072 -14228
rect 18038 -14352 18072 -14318
rect 18038 -14442 18072 -14408
rect 18038 -14532 18072 -14498
rect 18038 -14622 18072 -14588
rect 18038 -14712 18072 -14678
rect 18038 -14802 18072 -14768
rect 18038 -14892 18072 -14858
rect 18928 -14206 18962 -14172
rect 18928 -14296 18962 -14262
rect 18928 -14386 18962 -14352
rect 18928 -14476 18962 -14442
rect 18928 -14566 18962 -14532
rect 18928 -14656 18962 -14622
rect 18928 -14746 18962 -14712
rect 18928 -14836 18962 -14802
rect 18928 -14926 18962 -14892
rect 18132 -14984 18166 -14950
rect 18222 -14984 18256 -14950
rect 18312 -14984 18346 -14950
rect 18402 -14984 18436 -14950
rect 18492 -14984 18526 -14950
rect 18582 -14984 18616 -14950
rect 18672 -14984 18706 -14950
rect 18762 -14984 18796 -14950
rect 18852 -14984 18886 -14950
rect 19439 -14094 19473 -14060
rect 19529 -14094 19563 -14060
rect 19619 -14094 19653 -14060
rect 19709 -14094 19743 -14060
rect 19799 -14094 19833 -14060
rect 19889 -14094 19923 -14060
rect 19979 -14094 20013 -14060
rect 20069 -14094 20103 -14060
rect 20159 -14094 20193 -14060
rect 19326 -14172 19360 -14138
rect 19326 -14262 19360 -14228
rect 19326 -14352 19360 -14318
rect 19326 -14442 19360 -14408
rect 19326 -14532 19360 -14498
rect 19326 -14622 19360 -14588
rect 19326 -14712 19360 -14678
rect 19326 -14802 19360 -14768
rect 19326 -14892 19360 -14858
rect 20216 -14206 20250 -14172
rect 20216 -14296 20250 -14262
rect 20216 -14386 20250 -14352
rect 20216 -14476 20250 -14442
rect 20216 -14566 20250 -14532
rect 20216 -14656 20250 -14622
rect 20216 -14746 20250 -14712
rect 20216 -14836 20250 -14802
rect 20216 -14926 20250 -14892
rect 19420 -14984 19454 -14950
rect 19510 -14984 19544 -14950
rect 19600 -14984 19634 -14950
rect 19690 -14984 19724 -14950
rect 19780 -14984 19814 -14950
rect 19870 -14984 19904 -14950
rect 19960 -14984 19994 -14950
rect 20050 -14984 20084 -14950
rect 20140 -14984 20174 -14950
rect 20727 -14094 20761 -14060
rect 20817 -14094 20851 -14060
rect 20907 -14094 20941 -14060
rect 20997 -14094 21031 -14060
rect 21087 -14094 21121 -14060
rect 21177 -14094 21211 -14060
rect 21267 -14094 21301 -14060
rect 21357 -14094 21391 -14060
rect 21447 -14094 21481 -14060
rect 20614 -14172 20648 -14138
rect 20614 -14262 20648 -14228
rect 20614 -14352 20648 -14318
rect 20614 -14442 20648 -14408
rect 20614 -14532 20648 -14498
rect 20614 -14622 20648 -14588
rect 20614 -14712 20648 -14678
rect 20614 -14802 20648 -14768
rect 20614 -14892 20648 -14858
rect 21504 -14206 21538 -14172
rect 21504 -14296 21538 -14262
rect 21504 -14386 21538 -14352
rect 21504 -14476 21538 -14442
rect 21504 -14566 21538 -14532
rect 21504 -14656 21538 -14622
rect 21504 -14746 21538 -14712
rect 21504 -14836 21538 -14802
rect 21504 -14926 21538 -14892
rect 20708 -14984 20742 -14950
rect 20798 -14984 20832 -14950
rect 20888 -14984 20922 -14950
rect 20978 -14984 21012 -14950
rect 21068 -14984 21102 -14950
rect 21158 -14984 21192 -14950
rect 21248 -14984 21282 -14950
rect 21338 -14984 21372 -14950
rect 21428 -14984 21462 -14950
rect 22015 -14094 22049 -14060
rect 22105 -14094 22139 -14060
rect 22195 -14094 22229 -14060
rect 22285 -14094 22319 -14060
rect 22375 -14094 22409 -14060
rect 22465 -14094 22499 -14060
rect 22555 -14094 22589 -14060
rect 22645 -14094 22679 -14060
rect 22735 -14094 22769 -14060
rect 21902 -14172 21936 -14138
rect 21902 -14262 21936 -14228
rect 21902 -14352 21936 -14318
rect 21902 -14442 21936 -14408
rect 21902 -14532 21936 -14498
rect 21902 -14622 21936 -14588
rect 21902 -14712 21936 -14678
rect 21902 -14802 21936 -14768
rect 21902 -14892 21936 -14858
rect 22792 -14206 22826 -14172
rect 22792 -14296 22826 -14262
rect 22792 -14386 22826 -14352
rect 22792 -14476 22826 -14442
rect 22792 -14566 22826 -14532
rect 22792 -14656 22826 -14622
rect 22792 -14746 22826 -14712
rect 22792 -14836 22826 -14802
rect 22792 -14926 22826 -14892
rect 21996 -14984 22030 -14950
rect 22086 -14984 22120 -14950
rect 22176 -14984 22210 -14950
rect 22266 -14984 22300 -14950
rect 22356 -14984 22390 -14950
rect 22446 -14984 22480 -14950
rect 22536 -14984 22570 -14950
rect 22626 -14984 22660 -14950
rect 22716 -14984 22750 -14950
rect 23303 -14094 23337 -14060
rect 23393 -14094 23427 -14060
rect 23483 -14094 23517 -14060
rect 23573 -14094 23607 -14060
rect 23663 -14094 23697 -14060
rect 23753 -14094 23787 -14060
rect 23843 -14094 23877 -14060
rect 23933 -14094 23967 -14060
rect 24023 -14094 24057 -14060
rect 23190 -14172 23224 -14138
rect 23190 -14262 23224 -14228
rect 23190 -14352 23224 -14318
rect 23190 -14442 23224 -14408
rect 23190 -14532 23224 -14498
rect 23190 -14622 23224 -14588
rect 23190 -14712 23224 -14678
rect 23190 -14802 23224 -14768
rect 23190 -14892 23224 -14858
rect 24080 -14206 24114 -14172
rect 24080 -14296 24114 -14262
rect 24080 -14386 24114 -14352
rect 24080 -14476 24114 -14442
rect 24080 -14566 24114 -14532
rect 24080 -14656 24114 -14622
rect 24080 -14746 24114 -14712
rect 24080 -14836 24114 -14802
rect 24080 -14926 24114 -14892
rect 23284 -14984 23318 -14950
rect 23374 -14984 23408 -14950
rect 23464 -14984 23498 -14950
rect 23554 -14984 23588 -14950
rect 23644 -14984 23678 -14950
rect 23734 -14984 23768 -14950
rect 23824 -14984 23858 -14950
rect 23914 -14984 23948 -14950
rect 24004 -14984 24038 -14950
rect 24591 -14094 24625 -14060
rect 24681 -14094 24715 -14060
rect 24771 -14094 24805 -14060
rect 24861 -14094 24895 -14060
rect 24951 -14094 24985 -14060
rect 25041 -14094 25075 -14060
rect 25131 -14094 25165 -14060
rect 25221 -14094 25255 -14060
rect 25311 -14094 25345 -14060
rect 24478 -14172 24512 -14138
rect 24478 -14262 24512 -14228
rect 24478 -14352 24512 -14318
rect 24478 -14442 24512 -14408
rect 24478 -14532 24512 -14498
rect 24478 -14622 24512 -14588
rect 24478 -14712 24512 -14678
rect 24478 -14802 24512 -14768
rect 24478 -14892 24512 -14858
rect 25368 -14206 25402 -14172
rect 25368 -14296 25402 -14262
rect 25368 -14386 25402 -14352
rect 25368 -14476 25402 -14442
rect 25368 -14566 25402 -14532
rect 25368 -14656 25402 -14622
rect 25368 -14746 25402 -14712
rect 25368 -14836 25402 -14802
rect 25368 -14926 25402 -14892
rect 24572 -14984 24606 -14950
rect 24662 -14984 24696 -14950
rect 24752 -14984 24786 -14950
rect 24842 -14984 24876 -14950
rect 24932 -14984 24966 -14950
rect 25022 -14984 25056 -14950
rect 25112 -14984 25146 -14950
rect 25202 -14984 25236 -14950
rect 25292 -14984 25326 -14950
rect 25879 -14094 25913 -14060
rect 25969 -14094 26003 -14060
rect 26059 -14094 26093 -14060
rect 26149 -14094 26183 -14060
rect 26239 -14094 26273 -14060
rect 26329 -14094 26363 -14060
rect 26419 -14094 26453 -14060
rect 26509 -14094 26543 -14060
rect 26599 -14094 26633 -14060
rect 25766 -14172 25800 -14138
rect 25766 -14262 25800 -14228
rect 25766 -14352 25800 -14318
rect 25766 -14442 25800 -14408
rect 25766 -14532 25800 -14498
rect 25766 -14622 25800 -14588
rect 25766 -14712 25800 -14678
rect 25766 -14802 25800 -14768
rect 25766 -14892 25800 -14858
rect 26656 -14206 26690 -14172
rect 26656 -14296 26690 -14262
rect 26656 -14386 26690 -14352
rect 26656 -14476 26690 -14442
rect 26656 -14566 26690 -14532
rect 26656 -14656 26690 -14622
rect 26656 -14746 26690 -14712
rect 26656 -14836 26690 -14802
rect 26656 -14926 26690 -14892
rect 25860 -14984 25894 -14950
rect 25950 -14984 25984 -14950
rect 26040 -14984 26074 -14950
rect 26130 -14984 26164 -14950
rect 26220 -14984 26254 -14950
rect 26310 -14984 26344 -14950
rect 26400 -14984 26434 -14950
rect 26490 -14984 26524 -14950
rect 26580 -14984 26614 -14950
rect 16863 -15382 16897 -15348
rect 16953 -15382 16987 -15348
rect 17043 -15382 17077 -15348
rect 17133 -15382 17167 -15348
rect 17223 -15382 17257 -15348
rect 17313 -15382 17347 -15348
rect 17403 -15382 17437 -15348
rect 17493 -15382 17527 -15348
rect 17583 -15382 17617 -15348
rect 16750 -15460 16784 -15426
rect 16750 -15550 16784 -15516
rect 16750 -15640 16784 -15606
rect 16750 -15730 16784 -15696
rect 16750 -15820 16784 -15786
rect 16750 -15910 16784 -15876
rect 16750 -16000 16784 -15966
rect 16750 -16090 16784 -16056
rect 16750 -16180 16784 -16146
rect 17640 -15494 17674 -15460
rect 17640 -15584 17674 -15550
rect 17640 -15674 17674 -15640
rect 17640 -15764 17674 -15730
rect 17640 -15854 17674 -15820
rect 17640 -15944 17674 -15910
rect 17640 -16034 17674 -16000
rect 17640 -16124 17674 -16090
rect 17640 -16214 17674 -16180
rect 16844 -16272 16878 -16238
rect 16934 -16272 16968 -16238
rect 17024 -16272 17058 -16238
rect 17114 -16272 17148 -16238
rect 17204 -16272 17238 -16238
rect 17294 -16272 17328 -16238
rect 17384 -16272 17418 -16238
rect 17474 -16272 17508 -16238
rect 17564 -16272 17598 -16238
rect 18151 -15382 18185 -15348
rect 18241 -15382 18275 -15348
rect 18331 -15382 18365 -15348
rect 18421 -15382 18455 -15348
rect 18511 -15382 18545 -15348
rect 18601 -15382 18635 -15348
rect 18691 -15382 18725 -15348
rect 18781 -15382 18815 -15348
rect 18871 -15382 18905 -15348
rect 18038 -15460 18072 -15426
rect 18038 -15550 18072 -15516
rect 18038 -15640 18072 -15606
rect 18038 -15730 18072 -15696
rect 18038 -15820 18072 -15786
rect 18038 -15910 18072 -15876
rect 18038 -16000 18072 -15966
rect 18038 -16090 18072 -16056
rect 18038 -16180 18072 -16146
rect 18928 -15494 18962 -15460
rect 18928 -15584 18962 -15550
rect 18928 -15674 18962 -15640
rect 18928 -15764 18962 -15730
rect 18928 -15854 18962 -15820
rect 18928 -15944 18962 -15910
rect 18928 -16034 18962 -16000
rect 18928 -16124 18962 -16090
rect 18928 -16214 18962 -16180
rect 18132 -16272 18166 -16238
rect 18222 -16272 18256 -16238
rect 18312 -16272 18346 -16238
rect 18402 -16272 18436 -16238
rect 18492 -16272 18526 -16238
rect 18582 -16272 18616 -16238
rect 18672 -16272 18706 -16238
rect 18762 -16272 18796 -16238
rect 18852 -16272 18886 -16238
rect 19439 -15382 19473 -15348
rect 19529 -15382 19563 -15348
rect 19619 -15382 19653 -15348
rect 19709 -15382 19743 -15348
rect 19799 -15382 19833 -15348
rect 19889 -15382 19923 -15348
rect 19979 -15382 20013 -15348
rect 20069 -15382 20103 -15348
rect 20159 -15382 20193 -15348
rect 19326 -15460 19360 -15426
rect 19326 -15550 19360 -15516
rect 19326 -15640 19360 -15606
rect 19326 -15730 19360 -15696
rect 19326 -15820 19360 -15786
rect 19326 -15910 19360 -15876
rect 19326 -16000 19360 -15966
rect 19326 -16090 19360 -16056
rect 19326 -16180 19360 -16146
rect 20216 -15494 20250 -15460
rect 20216 -15584 20250 -15550
rect 20216 -15674 20250 -15640
rect 20216 -15764 20250 -15730
rect 20216 -15854 20250 -15820
rect 20216 -15944 20250 -15910
rect 20216 -16034 20250 -16000
rect 20216 -16124 20250 -16090
rect 20216 -16214 20250 -16180
rect 19420 -16272 19454 -16238
rect 19510 -16272 19544 -16238
rect 19600 -16272 19634 -16238
rect 19690 -16272 19724 -16238
rect 19780 -16272 19814 -16238
rect 19870 -16272 19904 -16238
rect 19960 -16272 19994 -16238
rect 20050 -16272 20084 -16238
rect 20140 -16272 20174 -16238
rect 20727 -15382 20761 -15348
rect 20817 -15382 20851 -15348
rect 20907 -15382 20941 -15348
rect 20997 -15382 21031 -15348
rect 21087 -15382 21121 -15348
rect 21177 -15382 21211 -15348
rect 21267 -15382 21301 -15348
rect 21357 -15382 21391 -15348
rect 21447 -15382 21481 -15348
rect 20614 -15460 20648 -15426
rect 20614 -15550 20648 -15516
rect 20614 -15640 20648 -15606
rect 20614 -15730 20648 -15696
rect 20614 -15820 20648 -15786
rect 20614 -15910 20648 -15876
rect 20614 -16000 20648 -15966
rect 20614 -16090 20648 -16056
rect 20614 -16180 20648 -16146
rect 21504 -15494 21538 -15460
rect 21504 -15584 21538 -15550
rect 21504 -15674 21538 -15640
rect 21504 -15764 21538 -15730
rect 21504 -15854 21538 -15820
rect 21504 -15944 21538 -15910
rect 21504 -16034 21538 -16000
rect 21504 -16124 21538 -16090
rect 21504 -16214 21538 -16180
rect 20708 -16272 20742 -16238
rect 20798 -16272 20832 -16238
rect 20888 -16272 20922 -16238
rect 20978 -16272 21012 -16238
rect 21068 -16272 21102 -16238
rect 21158 -16272 21192 -16238
rect 21248 -16272 21282 -16238
rect 21338 -16272 21372 -16238
rect 21428 -16272 21462 -16238
rect 22015 -15382 22049 -15348
rect 22105 -15382 22139 -15348
rect 22195 -15382 22229 -15348
rect 22285 -15382 22319 -15348
rect 22375 -15382 22409 -15348
rect 22465 -15382 22499 -15348
rect 22555 -15382 22589 -15348
rect 22645 -15382 22679 -15348
rect 22735 -15382 22769 -15348
rect 21902 -15460 21936 -15426
rect 21902 -15550 21936 -15516
rect 21902 -15640 21936 -15606
rect 21902 -15730 21936 -15696
rect 21902 -15820 21936 -15786
rect 21902 -15910 21936 -15876
rect 21902 -16000 21936 -15966
rect 21902 -16090 21936 -16056
rect 21902 -16180 21936 -16146
rect 22792 -15494 22826 -15460
rect 22792 -15584 22826 -15550
rect 22792 -15674 22826 -15640
rect 22792 -15764 22826 -15730
rect 22792 -15854 22826 -15820
rect 22792 -15944 22826 -15910
rect 22792 -16034 22826 -16000
rect 22792 -16124 22826 -16090
rect 22792 -16214 22826 -16180
rect 21996 -16272 22030 -16238
rect 22086 -16272 22120 -16238
rect 22176 -16272 22210 -16238
rect 22266 -16272 22300 -16238
rect 22356 -16272 22390 -16238
rect 22446 -16272 22480 -16238
rect 22536 -16272 22570 -16238
rect 22626 -16272 22660 -16238
rect 22716 -16272 22750 -16238
rect 23303 -15382 23337 -15348
rect 23393 -15382 23427 -15348
rect 23483 -15382 23517 -15348
rect 23573 -15382 23607 -15348
rect 23663 -15382 23697 -15348
rect 23753 -15382 23787 -15348
rect 23843 -15382 23877 -15348
rect 23933 -15382 23967 -15348
rect 24023 -15382 24057 -15348
rect 23190 -15460 23224 -15426
rect 23190 -15550 23224 -15516
rect 23190 -15640 23224 -15606
rect 23190 -15730 23224 -15696
rect 23190 -15820 23224 -15786
rect 23190 -15910 23224 -15876
rect 23190 -16000 23224 -15966
rect 23190 -16090 23224 -16056
rect 23190 -16180 23224 -16146
rect 24080 -15494 24114 -15460
rect 24080 -15584 24114 -15550
rect 24080 -15674 24114 -15640
rect 24080 -15764 24114 -15730
rect 24080 -15854 24114 -15820
rect 24080 -15944 24114 -15910
rect 24080 -16034 24114 -16000
rect 24080 -16124 24114 -16090
rect 24080 -16214 24114 -16180
rect 23284 -16272 23318 -16238
rect 23374 -16272 23408 -16238
rect 23464 -16272 23498 -16238
rect 23554 -16272 23588 -16238
rect 23644 -16272 23678 -16238
rect 23734 -16272 23768 -16238
rect 23824 -16272 23858 -16238
rect 23914 -16272 23948 -16238
rect 24004 -16272 24038 -16238
rect 24591 -15382 24625 -15348
rect 24681 -15382 24715 -15348
rect 24771 -15382 24805 -15348
rect 24861 -15382 24895 -15348
rect 24951 -15382 24985 -15348
rect 25041 -15382 25075 -15348
rect 25131 -15382 25165 -15348
rect 25221 -15382 25255 -15348
rect 25311 -15382 25345 -15348
rect 24478 -15460 24512 -15426
rect 24478 -15550 24512 -15516
rect 24478 -15640 24512 -15606
rect 24478 -15730 24512 -15696
rect 24478 -15820 24512 -15786
rect 24478 -15910 24512 -15876
rect 24478 -16000 24512 -15966
rect 24478 -16090 24512 -16056
rect 24478 -16180 24512 -16146
rect 25368 -15494 25402 -15460
rect 25368 -15584 25402 -15550
rect 25368 -15674 25402 -15640
rect 25368 -15764 25402 -15730
rect 25368 -15854 25402 -15820
rect 25368 -15944 25402 -15910
rect 25368 -16034 25402 -16000
rect 25368 -16124 25402 -16090
rect 25368 -16214 25402 -16180
rect 24572 -16272 24606 -16238
rect 24662 -16272 24696 -16238
rect 24752 -16272 24786 -16238
rect 24842 -16272 24876 -16238
rect 24932 -16272 24966 -16238
rect 25022 -16272 25056 -16238
rect 25112 -16272 25146 -16238
rect 25202 -16272 25236 -16238
rect 25292 -16272 25326 -16238
rect 25879 -15382 25913 -15348
rect 25969 -15382 26003 -15348
rect 26059 -15382 26093 -15348
rect 26149 -15382 26183 -15348
rect 26239 -15382 26273 -15348
rect 26329 -15382 26363 -15348
rect 26419 -15382 26453 -15348
rect 26509 -15382 26543 -15348
rect 26599 -15382 26633 -15348
rect 25766 -15460 25800 -15426
rect 25766 -15550 25800 -15516
rect 25766 -15640 25800 -15606
rect 25766 -15730 25800 -15696
rect 25766 -15820 25800 -15786
rect 25766 -15910 25800 -15876
rect 25766 -16000 25800 -15966
rect 25766 -16090 25800 -16056
rect 25766 -16180 25800 -16146
rect 26656 -15494 26690 -15460
rect 26656 -15584 26690 -15550
rect 26656 -15674 26690 -15640
rect 26656 -15764 26690 -15730
rect 26656 -15854 26690 -15820
rect 26656 -15944 26690 -15910
rect 26656 -16034 26690 -16000
rect 26656 -16124 26690 -16090
rect 26656 -16214 26690 -16180
rect 25860 -16272 25894 -16238
rect 25950 -16272 25984 -16238
rect 26040 -16272 26074 -16238
rect 26130 -16272 26164 -16238
rect 26220 -16272 26254 -16238
rect 26310 -16272 26344 -16238
rect 26400 -16272 26434 -16238
rect 26490 -16272 26524 -16238
rect 26580 -16272 26614 -16238
rect 16863 -16670 16897 -16636
rect 16953 -16670 16987 -16636
rect 17043 -16670 17077 -16636
rect 17133 -16670 17167 -16636
rect 17223 -16670 17257 -16636
rect 17313 -16670 17347 -16636
rect 17403 -16670 17437 -16636
rect 17493 -16670 17527 -16636
rect 17583 -16670 17617 -16636
rect 16750 -16748 16784 -16714
rect 16750 -16838 16784 -16804
rect 16750 -16928 16784 -16894
rect 16750 -17018 16784 -16984
rect 16750 -17108 16784 -17074
rect 16750 -17198 16784 -17164
rect 16750 -17288 16784 -17254
rect 16750 -17378 16784 -17344
rect 16750 -17468 16784 -17434
rect 17640 -16782 17674 -16748
rect 17640 -16872 17674 -16838
rect 17640 -16962 17674 -16928
rect 17640 -17052 17674 -17018
rect 17640 -17142 17674 -17108
rect 17640 -17232 17674 -17198
rect 17640 -17322 17674 -17288
rect 17640 -17412 17674 -17378
rect 17640 -17502 17674 -17468
rect 16844 -17560 16878 -17526
rect 16934 -17560 16968 -17526
rect 17024 -17560 17058 -17526
rect 17114 -17560 17148 -17526
rect 17204 -17560 17238 -17526
rect 17294 -17560 17328 -17526
rect 17384 -17560 17418 -17526
rect 17474 -17560 17508 -17526
rect 17564 -17560 17598 -17526
rect 18151 -16670 18185 -16636
rect 18241 -16670 18275 -16636
rect 18331 -16670 18365 -16636
rect 18421 -16670 18455 -16636
rect 18511 -16670 18545 -16636
rect 18601 -16670 18635 -16636
rect 18691 -16670 18725 -16636
rect 18781 -16670 18815 -16636
rect 18871 -16670 18905 -16636
rect 18038 -16748 18072 -16714
rect 18038 -16838 18072 -16804
rect 18038 -16928 18072 -16894
rect 18038 -17018 18072 -16984
rect 18038 -17108 18072 -17074
rect 18038 -17198 18072 -17164
rect 18038 -17288 18072 -17254
rect 18038 -17378 18072 -17344
rect 18038 -17468 18072 -17434
rect 18928 -16782 18962 -16748
rect 18928 -16872 18962 -16838
rect 18928 -16962 18962 -16928
rect 18928 -17052 18962 -17018
rect 18928 -17142 18962 -17108
rect 18928 -17232 18962 -17198
rect 18928 -17322 18962 -17288
rect 18928 -17412 18962 -17378
rect 18928 -17502 18962 -17468
rect 18132 -17560 18166 -17526
rect 18222 -17560 18256 -17526
rect 18312 -17560 18346 -17526
rect 18402 -17560 18436 -17526
rect 18492 -17560 18526 -17526
rect 18582 -17560 18616 -17526
rect 18672 -17560 18706 -17526
rect 18762 -17560 18796 -17526
rect 18852 -17560 18886 -17526
rect 19439 -16670 19473 -16636
rect 19529 -16670 19563 -16636
rect 19619 -16670 19653 -16636
rect 19709 -16670 19743 -16636
rect 19799 -16670 19833 -16636
rect 19889 -16670 19923 -16636
rect 19979 -16670 20013 -16636
rect 20069 -16670 20103 -16636
rect 20159 -16670 20193 -16636
rect 19326 -16748 19360 -16714
rect 19326 -16838 19360 -16804
rect 19326 -16928 19360 -16894
rect 19326 -17018 19360 -16984
rect 19326 -17108 19360 -17074
rect 19326 -17198 19360 -17164
rect 19326 -17288 19360 -17254
rect 19326 -17378 19360 -17344
rect 19326 -17468 19360 -17434
rect 20216 -16782 20250 -16748
rect 20216 -16872 20250 -16838
rect 20216 -16962 20250 -16928
rect 20216 -17052 20250 -17018
rect 20216 -17142 20250 -17108
rect 20216 -17232 20250 -17198
rect 20216 -17322 20250 -17288
rect 20216 -17412 20250 -17378
rect 20216 -17502 20250 -17468
rect 19420 -17560 19454 -17526
rect 19510 -17560 19544 -17526
rect 19600 -17560 19634 -17526
rect 19690 -17560 19724 -17526
rect 19780 -17560 19814 -17526
rect 19870 -17560 19904 -17526
rect 19960 -17560 19994 -17526
rect 20050 -17560 20084 -17526
rect 20140 -17560 20174 -17526
rect 20727 -16670 20761 -16636
rect 20817 -16670 20851 -16636
rect 20907 -16670 20941 -16636
rect 20997 -16670 21031 -16636
rect 21087 -16670 21121 -16636
rect 21177 -16670 21211 -16636
rect 21267 -16670 21301 -16636
rect 21357 -16670 21391 -16636
rect 21447 -16670 21481 -16636
rect 20614 -16748 20648 -16714
rect 20614 -16838 20648 -16804
rect 20614 -16928 20648 -16894
rect 20614 -17018 20648 -16984
rect 20614 -17108 20648 -17074
rect 20614 -17198 20648 -17164
rect 20614 -17288 20648 -17254
rect 20614 -17378 20648 -17344
rect 20614 -17468 20648 -17434
rect 21504 -16782 21538 -16748
rect 21504 -16872 21538 -16838
rect 21504 -16962 21538 -16928
rect 21504 -17052 21538 -17018
rect 21504 -17142 21538 -17108
rect 21504 -17232 21538 -17198
rect 21504 -17322 21538 -17288
rect 21504 -17412 21538 -17378
rect 21504 -17502 21538 -17468
rect 20708 -17560 20742 -17526
rect 20798 -17560 20832 -17526
rect 20888 -17560 20922 -17526
rect 20978 -17560 21012 -17526
rect 21068 -17560 21102 -17526
rect 21158 -17560 21192 -17526
rect 21248 -17560 21282 -17526
rect 21338 -17560 21372 -17526
rect 21428 -17560 21462 -17526
rect 22015 -16670 22049 -16636
rect 22105 -16670 22139 -16636
rect 22195 -16670 22229 -16636
rect 22285 -16670 22319 -16636
rect 22375 -16670 22409 -16636
rect 22465 -16670 22499 -16636
rect 22555 -16670 22589 -16636
rect 22645 -16670 22679 -16636
rect 22735 -16670 22769 -16636
rect 21902 -16748 21936 -16714
rect 21902 -16838 21936 -16804
rect 21902 -16928 21936 -16894
rect 21902 -17018 21936 -16984
rect 21902 -17108 21936 -17074
rect 21902 -17198 21936 -17164
rect 21902 -17288 21936 -17254
rect 21902 -17378 21936 -17344
rect 21902 -17468 21936 -17434
rect 22792 -16782 22826 -16748
rect 22792 -16872 22826 -16838
rect 22792 -16962 22826 -16928
rect 22792 -17052 22826 -17018
rect 22792 -17142 22826 -17108
rect 22792 -17232 22826 -17198
rect 22792 -17322 22826 -17288
rect 22792 -17412 22826 -17378
rect 22792 -17502 22826 -17468
rect 21996 -17560 22030 -17526
rect 22086 -17560 22120 -17526
rect 22176 -17560 22210 -17526
rect 22266 -17560 22300 -17526
rect 22356 -17560 22390 -17526
rect 22446 -17560 22480 -17526
rect 22536 -17560 22570 -17526
rect 22626 -17560 22660 -17526
rect 22716 -17560 22750 -17526
rect 23303 -16670 23337 -16636
rect 23393 -16670 23427 -16636
rect 23483 -16670 23517 -16636
rect 23573 -16670 23607 -16636
rect 23663 -16670 23697 -16636
rect 23753 -16670 23787 -16636
rect 23843 -16670 23877 -16636
rect 23933 -16670 23967 -16636
rect 24023 -16670 24057 -16636
rect 23190 -16748 23224 -16714
rect 23190 -16838 23224 -16804
rect 23190 -16928 23224 -16894
rect 23190 -17018 23224 -16984
rect 23190 -17108 23224 -17074
rect 23190 -17198 23224 -17164
rect 23190 -17288 23224 -17254
rect 23190 -17378 23224 -17344
rect 23190 -17468 23224 -17434
rect 24080 -16782 24114 -16748
rect 24080 -16872 24114 -16838
rect 24080 -16962 24114 -16928
rect 24080 -17052 24114 -17018
rect 24080 -17142 24114 -17108
rect 24080 -17232 24114 -17198
rect 24080 -17322 24114 -17288
rect 24080 -17412 24114 -17378
rect 24080 -17502 24114 -17468
rect 23284 -17560 23318 -17526
rect 23374 -17560 23408 -17526
rect 23464 -17560 23498 -17526
rect 23554 -17560 23588 -17526
rect 23644 -17560 23678 -17526
rect 23734 -17560 23768 -17526
rect 23824 -17560 23858 -17526
rect 23914 -17560 23948 -17526
rect 24004 -17560 24038 -17526
rect 24591 -16670 24625 -16636
rect 24681 -16670 24715 -16636
rect 24771 -16670 24805 -16636
rect 24861 -16670 24895 -16636
rect 24951 -16670 24985 -16636
rect 25041 -16670 25075 -16636
rect 25131 -16670 25165 -16636
rect 25221 -16670 25255 -16636
rect 25311 -16670 25345 -16636
rect 24478 -16748 24512 -16714
rect 24478 -16838 24512 -16804
rect 24478 -16928 24512 -16894
rect 24478 -17018 24512 -16984
rect 24478 -17108 24512 -17074
rect 24478 -17198 24512 -17164
rect 24478 -17288 24512 -17254
rect 24478 -17378 24512 -17344
rect 24478 -17468 24512 -17434
rect 25368 -16782 25402 -16748
rect 25368 -16872 25402 -16838
rect 25368 -16962 25402 -16928
rect 25368 -17052 25402 -17018
rect 25368 -17142 25402 -17108
rect 25368 -17232 25402 -17198
rect 25368 -17322 25402 -17288
rect 25368 -17412 25402 -17378
rect 25368 -17502 25402 -17468
rect 24572 -17560 24606 -17526
rect 24662 -17560 24696 -17526
rect 24752 -17560 24786 -17526
rect 24842 -17560 24876 -17526
rect 24932 -17560 24966 -17526
rect 25022 -17560 25056 -17526
rect 25112 -17560 25146 -17526
rect 25202 -17560 25236 -17526
rect 25292 -17560 25326 -17526
rect 25879 -16670 25913 -16636
rect 25969 -16670 26003 -16636
rect 26059 -16670 26093 -16636
rect 26149 -16670 26183 -16636
rect 26239 -16670 26273 -16636
rect 26329 -16670 26363 -16636
rect 26419 -16670 26453 -16636
rect 26509 -16670 26543 -16636
rect 26599 -16670 26633 -16636
rect 25766 -16748 25800 -16714
rect 25766 -16838 25800 -16804
rect 25766 -16928 25800 -16894
rect 25766 -17018 25800 -16984
rect 25766 -17108 25800 -17074
rect 25766 -17198 25800 -17164
rect 25766 -17288 25800 -17254
rect 25766 -17378 25800 -17344
rect 25766 -17468 25800 -17434
rect 26656 -16782 26690 -16748
rect 26656 -16872 26690 -16838
rect 26656 -16962 26690 -16928
rect 26656 -17052 26690 -17018
rect 26656 -17142 26690 -17108
rect 26656 -17232 26690 -17198
rect 26656 -17322 26690 -17288
rect 26656 -17412 26690 -17378
rect 26656 -17502 26690 -17468
rect 25860 -17560 25894 -17526
rect 25950 -17560 25984 -17526
rect 26040 -17560 26074 -17526
rect 26130 -17560 26164 -17526
rect 26220 -17560 26254 -17526
rect 26310 -17560 26344 -17526
rect 26400 -17560 26434 -17526
rect 26490 -17560 26524 -17526
rect 26580 -17560 26614 -17526
<< xpolycontact >>
rect 6870 -17850 7302 -17280
rect 13606 -17850 14038 -17280
rect 6870 -18668 7302 -18098
rect 13606 -18668 14038 -18098
rect 6870 -19486 7302 -18916
rect 13606 -19486 14038 -18916
rect 6870 -20304 7302 -19734
rect 13606 -20304 14038 -19734
rect 6870 -21122 7302 -20552
rect 13606 -21122 14038 -20552
rect 6870 -21940 7302 -21370
rect 13606 -21940 14038 -21370
rect 6870 -22758 7302 -22188
rect 13606 -22758 14038 -22188
rect 6870 -23576 7302 -23006
rect 13606 -23576 14038 -23006
rect 6870 -24394 7302 -23824
rect 13606 -24394 14038 -23824
rect 6870 -25212 7302 -24642
rect 13606 -25212 14038 -24642
rect 6870 -26030 7302 -25460
rect 13606 -26030 14038 -25460
rect 6870 -26848 7302 -26278
rect 13606 -26848 14038 -26278
rect 6870 -27666 7302 -27096
rect 13606 -27666 14038 -27096
rect 6870 -28484 7302 -27914
rect 13606 -28484 14038 -27914
rect 6870 -29302 7302 -28732
rect 13606 -29302 14038 -28732
rect 6870 -30120 7302 -29550
rect 13606 -30120 14038 -29550
rect 6870 -30938 7302 -30368
rect 13606 -30938 14038 -30368
rect 6808 -33392 7240 -32822
rect 11540 -33392 11972 -32822
rect 6808 -34210 7240 -33640
rect 11540 -34210 11972 -33640
rect 6808 -35028 7240 -34458
rect 11540 -35028 11972 -34458
rect 6808 -35846 7240 -35276
rect 11540 -35846 11972 -35276
rect 8194 -37482 8626 -36912
rect 11950 -37482 12382 -36912
rect 8194 -38300 8626 -37730
rect 11950 -38300 12382 -37730
rect 8194 -39118 8626 -38548
rect 11950 -39118 12382 -38548
<< xpolyres >>
rect 7302 -17850 13606 -17280
rect 7302 -18668 13606 -18098
rect 7302 -19486 13606 -18916
rect 7302 -20304 13606 -19734
rect 7302 -21122 13606 -20552
rect 7302 -21940 13606 -21370
rect 7302 -22758 13606 -22188
rect 7302 -23576 13606 -23006
rect 7302 -24394 13606 -23824
rect 7302 -25212 13606 -24642
rect 7302 -26030 13606 -25460
rect 7302 -26848 13606 -26278
rect 7302 -27666 13606 -27096
rect 7302 -28484 13606 -27914
rect 7302 -29302 13606 -28732
rect 7302 -30120 13606 -29550
rect 7302 -30938 13606 -30368
rect 7240 -33392 11540 -32822
rect 7240 -34210 11540 -33640
rect 7240 -35028 11540 -34458
rect 7240 -35846 11540 -35276
rect 8626 -37482 11950 -36912
rect 8626 -38300 11950 -37730
rect 8626 -39118 11950 -38548
<< locali >>
rect 16568 -11336 26884 -11302
rect 16568 -11370 16684 -11336
rect 16718 -11370 16774 -11336
rect 16808 -11370 16864 -11336
rect 16898 -11370 16954 -11336
rect 16988 -11370 17044 -11336
rect 17078 -11370 17134 -11336
rect 17168 -11370 17224 -11336
rect 17258 -11370 17314 -11336
rect 17348 -11370 17404 -11336
rect 17438 -11370 17494 -11336
rect 17528 -11370 17584 -11336
rect 17618 -11370 17674 -11336
rect 17708 -11370 17764 -11336
rect 17798 -11370 17972 -11336
rect 18006 -11370 18062 -11336
rect 18096 -11370 18152 -11336
rect 18186 -11370 18242 -11336
rect 18276 -11370 18332 -11336
rect 18366 -11370 18422 -11336
rect 18456 -11370 18512 -11336
rect 18546 -11370 18602 -11336
rect 18636 -11370 18692 -11336
rect 18726 -11370 18782 -11336
rect 18816 -11370 18872 -11336
rect 18906 -11370 18962 -11336
rect 18996 -11370 19052 -11336
rect 19086 -11370 19260 -11336
rect 19294 -11370 19350 -11336
rect 19384 -11370 19440 -11336
rect 19474 -11370 19530 -11336
rect 19564 -11370 19620 -11336
rect 19654 -11370 19710 -11336
rect 19744 -11370 19800 -11336
rect 19834 -11370 19890 -11336
rect 19924 -11370 19980 -11336
rect 20014 -11370 20070 -11336
rect 20104 -11370 20160 -11336
rect 20194 -11370 20250 -11336
rect 20284 -11370 20340 -11336
rect 20374 -11370 20548 -11336
rect 20582 -11370 20638 -11336
rect 20672 -11370 20728 -11336
rect 20762 -11370 20818 -11336
rect 20852 -11370 20908 -11336
rect 20942 -11370 20998 -11336
rect 21032 -11370 21088 -11336
rect 21122 -11370 21178 -11336
rect 21212 -11370 21268 -11336
rect 21302 -11370 21358 -11336
rect 21392 -11370 21448 -11336
rect 21482 -11370 21538 -11336
rect 21572 -11370 21628 -11336
rect 21662 -11370 21836 -11336
rect 21870 -11370 21926 -11336
rect 21960 -11370 22016 -11336
rect 22050 -11370 22106 -11336
rect 22140 -11370 22196 -11336
rect 22230 -11370 22286 -11336
rect 22320 -11370 22376 -11336
rect 22410 -11370 22466 -11336
rect 22500 -11370 22556 -11336
rect 22590 -11370 22646 -11336
rect 22680 -11370 22736 -11336
rect 22770 -11370 22826 -11336
rect 22860 -11370 22916 -11336
rect 22950 -11370 23124 -11336
rect 23158 -11370 23214 -11336
rect 23248 -11370 23304 -11336
rect 23338 -11370 23394 -11336
rect 23428 -11370 23484 -11336
rect 23518 -11370 23574 -11336
rect 23608 -11370 23664 -11336
rect 23698 -11370 23754 -11336
rect 23788 -11370 23844 -11336
rect 23878 -11370 23934 -11336
rect 23968 -11370 24024 -11336
rect 24058 -11370 24114 -11336
rect 24148 -11370 24204 -11336
rect 24238 -11370 24412 -11336
rect 24446 -11370 24502 -11336
rect 24536 -11370 24592 -11336
rect 24626 -11370 24682 -11336
rect 24716 -11370 24772 -11336
rect 24806 -11370 24862 -11336
rect 24896 -11370 24952 -11336
rect 24986 -11370 25042 -11336
rect 25076 -11370 25132 -11336
rect 25166 -11370 25222 -11336
rect 25256 -11370 25312 -11336
rect 25346 -11370 25402 -11336
rect 25436 -11370 25492 -11336
rect 25526 -11370 25700 -11336
rect 25734 -11370 25790 -11336
rect 25824 -11370 25880 -11336
rect 25914 -11370 25970 -11336
rect 26004 -11370 26060 -11336
rect 26094 -11370 26150 -11336
rect 26184 -11370 26240 -11336
rect 26274 -11370 26330 -11336
rect 26364 -11370 26420 -11336
rect 26454 -11370 26510 -11336
rect 26544 -11370 26600 -11336
rect 26634 -11370 26690 -11336
rect 26724 -11370 26780 -11336
rect 26814 -11370 26884 -11336
rect 16568 -11432 26884 -11370
rect 16568 -11466 16600 -11432
rect 16634 -11466 17787 -11432
rect 17821 -11466 17888 -11432
rect 17922 -11466 19075 -11432
rect 19109 -11466 19176 -11432
rect 19210 -11466 20363 -11432
rect 20397 -11466 20464 -11432
rect 20498 -11466 21651 -11432
rect 21685 -11466 21752 -11432
rect 21786 -11466 22939 -11432
rect 22973 -11466 23040 -11432
rect 23074 -11466 24227 -11432
rect 24261 -11466 24328 -11432
rect 24362 -11466 25515 -11432
rect 25549 -11466 25616 -11432
rect 25650 -11466 26803 -11432
rect 26837 -11466 26884 -11432
rect 16568 -11484 26884 -11466
rect 16568 -11502 16863 -11484
rect 16568 -11522 16667 -11502
rect 16568 -11556 16600 -11522
rect 16634 -11556 16667 -11522
rect 16568 -11612 16667 -11556
rect 16568 -11646 16600 -11612
rect 16634 -11646 16667 -11612
rect 16568 -11702 16667 -11646
rect 16568 -11736 16600 -11702
rect 16634 -11736 16667 -11702
rect 16568 -11792 16667 -11736
rect 16568 -11826 16600 -11792
rect 16634 -11826 16667 -11792
rect 16568 -11882 16667 -11826
rect 16568 -11916 16600 -11882
rect 16634 -11916 16667 -11882
rect 16568 -11972 16667 -11916
rect 16568 -12006 16600 -11972
rect 16634 -12006 16667 -11972
rect 16568 -12062 16667 -12006
rect 16568 -12096 16600 -12062
rect 16634 -12096 16667 -12062
rect 16568 -12152 16667 -12096
rect 16568 -12186 16600 -12152
rect 16634 -12186 16667 -12152
rect 16568 -12242 16667 -12186
rect 16568 -12276 16600 -12242
rect 16634 -12276 16667 -12242
rect 16568 -12332 16667 -12276
rect 16568 -12366 16600 -12332
rect 16634 -12366 16667 -12332
rect 16568 -12402 16667 -12366
rect 16731 -11518 16863 -11502
rect 16897 -11518 16953 -11484
rect 16987 -11518 17043 -11484
rect 17077 -11518 17133 -11484
rect 17167 -11518 17223 -11484
rect 17257 -11518 17313 -11484
rect 17347 -11518 17403 -11484
rect 17437 -11518 17493 -11484
rect 17527 -11518 17583 -11484
rect 17617 -11502 18151 -11484
rect 17617 -11518 17693 -11502
rect 16731 -11537 17693 -11518
rect 16731 -11562 16803 -11537
rect 16731 -11596 16750 -11562
rect 16784 -11596 16803 -11562
rect 16731 -11652 16803 -11596
rect 17621 -11596 17693 -11537
rect 16731 -11686 16750 -11652
rect 16784 -11686 16803 -11652
rect 16731 -11742 16803 -11686
rect 16731 -11776 16750 -11742
rect 16784 -11776 16803 -11742
rect 16731 -11832 16803 -11776
rect 16731 -11866 16750 -11832
rect 16784 -11866 16803 -11832
rect 16731 -11922 16803 -11866
rect 16731 -11956 16750 -11922
rect 16784 -11956 16803 -11922
rect 16731 -12012 16803 -11956
rect 16731 -12046 16750 -12012
rect 16784 -12046 16803 -12012
rect 16731 -12102 16803 -12046
rect 16731 -12136 16750 -12102
rect 16784 -12136 16803 -12102
rect 16731 -12192 16803 -12136
rect 16731 -12226 16750 -12192
rect 16784 -12226 16803 -12192
rect 16731 -12282 16803 -12226
rect 16731 -12316 16750 -12282
rect 16784 -12316 16803 -12282
rect 16865 -11660 17559 -11599
rect 16865 -11694 16926 -11660
rect 16960 -11672 17016 -11660
rect 17050 -11672 17106 -11660
rect 17140 -11672 17196 -11660
rect 16972 -11694 17016 -11672
rect 17072 -11694 17106 -11672
rect 17172 -11694 17196 -11672
rect 17230 -11672 17286 -11660
rect 17230 -11694 17238 -11672
rect 16865 -11706 16938 -11694
rect 16972 -11706 17038 -11694
rect 17072 -11706 17138 -11694
rect 17172 -11706 17238 -11694
rect 17272 -11694 17286 -11672
rect 17320 -11672 17376 -11660
rect 17320 -11694 17338 -11672
rect 17272 -11706 17338 -11694
rect 17372 -11694 17376 -11672
rect 17410 -11672 17466 -11660
rect 17410 -11694 17438 -11672
rect 17500 -11694 17559 -11660
rect 17372 -11706 17438 -11694
rect 17472 -11706 17559 -11694
rect 16865 -11750 17559 -11706
rect 16865 -11784 16926 -11750
rect 16960 -11772 17016 -11750
rect 17050 -11772 17106 -11750
rect 17140 -11772 17196 -11750
rect 16972 -11784 17016 -11772
rect 17072 -11784 17106 -11772
rect 17172 -11784 17196 -11772
rect 17230 -11772 17286 -11750
rect 17230 -11784 17238 -11772
rect 16865 -11806 16938 -11784
rect 16972 -11806 17038 -11784
rect 17072 -11806 17138 -11784
rect 17172 -11806 17238 -11784
rect 17272 -11784 17286 -11772
rect 17320 -11772 17376 -11750
rect 17320 -11784 17338 -11772
rect 17272 -11806 17338 -11784
rect 17372 -11784 17376 -11772
rect 17410 -11772 17466 -11750
rect 17410 -11784 17438 -11772
rect 17500 -11784 17559 -11750
rect 17372 -11806 17438 -11784
rect 17472 -11806 17559 -11784
rect 16865 -11840 17559 -11806
rect 16865 -11874 16926 -11840
rect 16960 -11872 17016 -11840
rect 17050 -11872 17106 -11840
rect 17140 -11872 17196 -11840
rect 16972 -11874 17016 -11872
rect 17072 -11874 17106 -11872
rect 17172 -11874 17196 -11872
rect 17230 -11872 17286 -11840
rect 17230 -11874 17238 -11872
rect 16865 -11906 16938 -11874
rect 16972 -11906 17038 -11874
rect 17072 -11906 17138 -11874
rect 17172 -11906 17238 -11874
rect 17272 -11874 17286 -11872
rect 17320 -11872 17376 -11840
rect 17320 -11874 17338 -11872
rect 17272 -11906 17338 -11874
rect 17372 -11874 17376 -11872
rect 17410 -11872 17466 -11840
rect 17410 -11874 17438 -11872
rect 17500 -11874 17559 -11840
rect 17372 -11906 17438 -11874
rect 17472 -11906 17559 -11874
rect 16865 -11930 17559 -11906
rect 16865 -11964 16926 -11930
rect 16960 -11964 17016 -11930
rect 17050 -11964 17106 -11930
rect 17140 -11964 17196 -11930
rect 17230 -11964 17286 -11930
rect 17320 -11964 17376 -11930
rect 17410 -11964 17466 -11930
rect 17500 -11964 17559 -11930
rect 16865 -11972 17559 -11964
rect 16865 -12006 16938 -11972
rect 16972 -12006 17038 -11972
rect 17072 -12006 17138 -11972
rect 17172 -12006 17238 -11972
rect 17272 -12006 17338 -11972
rect 17372 -12006 17438 -11972
rect 17472 -12006 17559 -11972
rect 16865 -12020 17559 -12006
rect 16865 -12054 16926 -12020
rect 16960 -12054 17016 -12020
rect 17050 -12054 17106 -12020
rect 17140 -12054 17196 -12020
rect 17230 -12054 17286 -12020
rect 17320 -12054 17376 -12020
rect 17410 -12054 17466 -12020
rect 17500 -12054 17559 -12020
rect 16865 -12072 17559 -12054
rect 16865 -12106 16938 -12072
rect 16972 -12106 17038 -12072
rect 17072 -12106 17138 -12072
rect 17172 -12106 17238 -12072
rect 17272 -12106 17338 -12072
rect 17372 -12106 17438 -12072
rect 17472 -12106 17559 -12072
rect 16865 -12110 17559 -12106
rect 16865 -12144 16926 -12110
rect 16960 -12144 17016 -12110
rect 17050 -12144 17106 -12110
rect 17140 -12144 17196 -12110
rect 17230 -12144 17286 -12110
rect 17320 -12144 17376 -12110
rect 17410 -12144 17466 -12110
rect 17500 -12144 17559 -12110
rect 16865 -12172 17559 -12144
rect 16865 -12200 16938 -12172
rect 16972 -12200 17038 -12172
rect 17072 -12200 17138 -12172
rect 17172 -12200 17238 -12172
rect 16865 -12234 16926 -12200
rect 16972 -12206 17016 -12200
rect 17072 -12206 17106 -12200
rect 17172 -12206 17196 -12200
rect 16960 -12234 17016 -12206
rect 17050 -12234 17106 -12206
rect 17140 -12234 17196 -12206
rect 17230 -12206 17238 -12200
rect 17272 -12200 17338 -12172
rect 17272 -12206 17286 -12200
rect 17230 -12234 17286 -12206
rect 17320 -12206 17338 -12200
rect 17372 -12200 17438 -12172
rect 17472 -12200 17559 -12172
rect 17372 -12206 17376 -12200
rect 17320 -12234 17376 -12206
rect 17410 -12206 17438 -12200
rect 17410 -12234 17466 -12206
rect 17500 -12234 17559 -12200
rect 16865 -12293 17559 -12234
rect 17621 -11630 17640 -11596
rect 17674 -11630 17693 -11596
rect 17621 -11686 17693 -11630
rect 17621 -11720 17640 -11686
rect 17674 -11720 17693 -11686
rect 17621 -11776 17693 -11720
rect 17621 -11810 17640 -11776
rect 17674 -11810 17693 -11776
rect 17621 -11866 17693 -11810
rect 17621 -11900 17640 -11866
rect 17674 -11900 17693 -11866
rect 17621 -11956 17693 -11900
rect 17621 -11990 17640 -11956
rect 17674 -11990 17693 -11956
rect 17621 -12046 17693 -11990
rect 17621 -12080 17640 -12046
rect 17674 -12080 17693 -12046
rect 17621 -12136 17693 -12080
rect 17621 -12170 17640 -12136
rect 17674 -12170 17693 -12136
rect 17621 -12226 17693 -12170
rect 17621 -12260 17640 -12226
rect 17674 -12260 17693 -12226
rect 16731 -12355 16803 -12316
rect 17621 -12316 17693 -12260
rect 17621 -12350 17640 -12316
rect 17674 -12350 17693 -12316
rect 17621 -12355 17693 -12350
rect 16731 -12374 17693 -12355
rect 16731 -12402 16844 -12374
rect 16568 -12408 16844 -12402
rect 16878 -12408 16934 -12374
rect 16968 -12408 17024 -12374
rect 17058 -12408 17114 -12374
rect 17148 -12408 17204 -12374
rect 17238 -12408 17294 -12374
rect 17328 -12408 17384 -12374
rect 17418 -12408 17474 -12374
rect 17508 -12408 17564 -12374
rect 17598 -12402 17693 -12374
rect 17757 -11522 17955 -11502
rect 17757 -11556 17787 -11522
rect 17821 -11556 17888 -11522
rect 17922 -11556 17955 -11522
rect 17757 -11612 17955 -11556
rect 17757 -11646 17787 -11612
rect 17821 -11646 17888 -11612
rect 17922 -11646 17955 -11612
rect 17757 -11702 17955 -11646
rect 17757 -11736 17787 -11702
rect 17821 -11736 17888 -11702
rect 17922 -11736 17955 -11702
rect 17757 -11792 17955 -11736
rect 17757 -11826 17787 -11792
rect 17821 -11826 17888 -11792
rect 17922 -11826 17955 -11792
rect 17757 -11882 17955 -11826
rect 17757 -11916 17787 -11882
rect 17821 -11916 17888 -11882
rect 17922 -11916 17955 -11882
rect 17757 -11972 17955 -11916
rect 17757 -12006 17787 -11972
rect 17821 -12006 17888 -11972
rect 17922 -12006 17955 -11972
rect 17757 -12062 17955 -12006
rect 17757 -12096 17787 -12062
rect 17821 -12096 17888 -12062
rect 17922 -12096 17955 -12062
rect 17757 -12152 17955 -12096
rect 17757 -12186 17787 -12152
rect 17821 -12186 17888 -12152
rect 17922 -12186 17955 -12152
rect 17757 -12242 17955 -12186
rect 17757 -12276 17787 -12242
rect 17821 -12276 17888 -12242
rect 17922 -12276 17955 -12242
rect 17757 -12332 17955 -12276
rect 17757 -12366 17787 -12332
rect 17821 -12366 17888 -12332
rect 17922 -12366 17955 -12332
rect 17757 -12402 17955 -12366
rect 18019 -11518 18151 -11502
rect 18185 -11518 18241 -11484
rect 18275 -11518 18331 -11484
rect 18365 -11518 18421 -11484
rect 18455 -11518 18511 -11484
rect 18545 -11518 18601 -11484
rect 18635 -11518 18691 -11484
rect 18725 -11518 18781 -11484
rect 18815 -11518 18871 -11484
rect 18905 -11502 19439 -11484
rect 18905 -11518 18981 -11502
rect 18019 -11537 18981 -11518
rect 18019 -11562 18091 -11537
rect 18019 -11596 18038 -11562
rect 18072 -11596 18091 -11562
rect 18019 -11652 18091 -11596
rect 18909 -11596 18981 -11537
rect 18019 -11686 18038 -11652
rect 18072 -11686 18091 -11652
rect 18019 -11742 18091 -11686
rect 18019 -11776 18038 -11742
rect 18072 -11776 18091 -11742
rect 18019 -11832 18091 -11776
rect 18019 -11866 18038 -11832
rect 18072 -11866 18091 -11832
rect 18019 -11922 18091 -11866
rect 18019 -11956 18038 -11922
rect 18072 -11956 18091 -11922
rect 18019 -12012 18091 -11956
rect 18019 -12046 18038 -12012
rect 18072 -12046 18091 -12012
rect 18019 -12102 18091 -12046
rect 18019 -12136 18038 -12102
rect 18072 -12136 18091 -12102
rect 18019 -12192 18091 -12136
rect 18019 -12226 18038 -12192
rect 18072 -12226 18091 -12192
rect 18019 -12282 18091 -12226
rect 18019 -12316 18038 -12282
rect 18072 -12316 18091 -12282
rect 18153 -11660 18847 -11599
rect 18153 -11694 18214 -11660
rect 18248 -11672 18304 -11660
rect 18338 -11672 18394 -11660
rect 18428 -11672 18484 -11660
rect 18260 -11694 18304 -11672
rect 18360 -11694 18394 -11672
rect 18460 -11694 18484 -11672
rect 18518 -11672 18574 -11660
rect 18518 -11694 18526 -11672
rect 18153 -11706 18226 -11694
rect 18260 -11706 18326 -11694
rect 18360 -11706 18426 -11694
rect 18460 -11706 18526 -11694
rect 18560 -11694 18574 -11672
rect 18608 -11672 18664 -11660
rect 18608 -11694 18626 -11672
rect 18560 -11706 18626 -11694
rect 18660 -11694 18664 -11672
rect 18698 -11672 18754 -11660
rect 18698 -11694 18726 -11672
rect 18788 -11694 18847 -11660
rect 18660 -11706 18726 -11694
rect 18760 -11706 18847 -11694
rect 18153 -11750 18847 -11706
rect 18153 -11784 18214 -11750
rect 18248 -11772 18304 -11750
rect 18338 -11772 18394 -11750
rect 18428 -11772 18484 -11750
rect 18260 -11784 18304 -11772
rect 18360 -11784 18394 -11772
rect 18460 -11784 18484 -11772
rect 18518 -11772 18574 -11750
rect 18518 -11784 18526 -11772
rect 18153 -11806 18226 -11784
rect 18260 -11806 18326 -11784
rect 18360 -11806 18426 -11784
rect 18460 -11806 18526 -11784
rect 18560 -11784 18574 -11772
rect 18608 -11772 18664 -11750
rect 18608 -11784 18626 -11772
rect 18560 -11806 18626 -11784
rect 18660 -11784 18664 -11772
rect 18698 -11772 18754 -11750
rect 18698 -11784 18726 -11772
rect 18788 -11784 18847 -11750
rect 18660 -11806 18726 -11784
rect 18760 -11806 18847 -11784
rect 18153 -11840 18847 -11806
rect 18153 -11874 18214 -11840
rect 18248 -11872 18304 -11840
rect 18338 -11872 18394 -11840
rect 18428 -11872 18484 -11840
rect 18260 -11874 18304 -11872
rect 18360 -11874 18394 -11872
rect 18460 -11874 18484 -11872
rect 18518 -11872 18574 -11840
rect 18518 -11874 18526 -11872
rect 18153 -11906 18226 -11874
rect 18260 -11906 18326 -11874
rect 18360 -11906 18426 -11874
rect 18460 -11906 18526 -11874
rect 18560 -11874 18574 -11872
rect 18608 -11872 18664 -11840
rect 18608 -11874 18626 -11872
rect 18560 -11906 18626 -11874
rect 18660 -11874 18664 -11872
rect 18698 -11872 18754 -11840
rect 18698 -11874 18726 -11872
rect 18788 -11874 18847 -11840
rect 18660 -11906 18726 -11874
rect 18760 -11906 18847 -11874
rect 18153 -11930 18847 -11906
rect 18153 -11964 18214 -11930
rect 18248 -11964 18304 -11930
rect 18338 -11964 18394 -11930
rect 18428 -11964 18484 -11930
rect 18518 -11964 18574 -11930
rect 18608 -11964 18664 -11930
rect 18698 -11964 18754 -11930
rect 18788 -11964 18847 -11930
rect 18153 -11972 18847 -11964
rect 18153 -12006 18226 -11972
rect 18260 -12006 18326 -11972
rect 18360 -12006 18426 -11972
rect 18460 -12006 18526 -11972
rect 18560 -12006 18626 -11972
rect 18660 -12006 18726 -11972
rect 18760 -12006 18847 -11972
rect 18153 -12020 18847 -12006
rect 18153 -12054 18214 -12020
rect 18248 -12054 18304 -12020
rect 18338 -12054 18394 -12020
rect 18428 -12054 18484 -12020
rect 18518 -12054 18574 -12020
rect 18608 -12054 18664 -12020
rect 18698 -12054 18754 -12020
rect 18788 -12054 18847 -12020
rect 18153 -12072 18847 -12054
rect 18153 -12106 18226 -12072
rect 18260 -12106 18326 -12072
rect 18360 -12106 18426 -12072
rect 18460 -12106 18526 -12072
rect 18560 -12106 18626 -12072
rect 18660 -12106 18726 -12072
rect 18760 -12106 18847 -12072
rect 18153 -12110 18847 -12106
rect 18153 -12144 18214 -12110
rect 18248 -12144 18304 -12110
rect 18338 -12144 18394 -12110
rect 18428 -12144 18484 -12110
rect 18518 -12144 18574 -12110
rect 18608 -12144 18664 -12110
rect 18698 -12144 18754 -12110
rect 18788 -12144 18847 -12110
rect 18153 -12172 18847 -12144
rect 18153 -12200 18226 -12172
rect 18260 -12200 18326 -12172
rect 18360 -12200 18426 -12172
rect 18460 -12200 18526 -12172
rect 18153 -12234 18214 -12200
rect 18260 -12206 18304 -12200
rect 18360 -12206 18394 -12200
rect 18460 -12206 18484 -12200
rect 18248 -12234 18304 -12206
rect 18338 -12234 18394 -12206
rect 18428 -12234 18484 -12206
rect 18518 -12206 18526 -12200
rect 18560 -12200 18626 -12172
rect 18560 -12206 18574 -12200
rect 18518 -12234 18574 -12206
rect 18608 -12206 18626 -12200
rect 18660 -12200 18726 -12172
rect 18760 -12200 18847 -12172
rect 18660 -12206 18664 -12200
rect 18608 -12234 18664 -12206
rect 18698 -12206 18726 -12200
rect 18698 -12234 18754 -12206
rect 18788 -12234 18847 -12200
rect 18153 -12293 18847 -12234
rect 18909 -11630 18928 -11596
rect 18962 -11630 18981 -11596
rect 18909 -11686 18981 -11630
rect 18909 -11720 18928 -11686
rect 18962 -11720 18981 -11686
rect 18909 -11776 18981 -11720
rect 18909 -11810 18928 -11776
rect 18962 -11810 18981 -11776
rect 18909 -11866 18981 -11810
rect 18909 -11900 18928 -11866
rect 18962 -11900 18981 -11866
rect 18909 -11956 18981 -11900
rect 18909 -11990 18928 -11956
rect 18962 -11990 18981 -11956
rect 18909 -12046 18981 -11990
rect 18909 -12080 18928 -12046
rect 18962 -12080 18981 -12046
rect 18909 -12136 18981 -12080
rect 18909 -12170 18928 -12136
rect 18962 -12170 18981 -12136
rect 18909 -12226 18981 -12170
rect 18909 -12260 18928 -12226
rect 18962 -12260 18981 -12226
rect 18019 -12355 18091 -12316
rect 18909 -12316 18981 -12260
rect 18909 -12350 18928 -12316
rect 18962 -12350 18981 -12316
rect 18909 -12355 18981 -12350
rect 18019 -12374 18981 -12355
rect 18019 -12402 18132 -12374
rect 17598 -12408 18132 -12402
rect 18166 -12408 18222 -12374
rect 18256 -12408 18312 -12374
rect 18346 -12408 18402 -12374
rect 18436 -12408 18492 -12374
rect 18526 -12408 18582 -12374
rect 18616 -12408 18672 -12374
rect 18706 -12408 18762 -12374
rect 18796 -12408 18852 -12374
rect 18886 -12402 18981 -12374
rect 19045 -11522 19243 -11502
rect 19045 -11556 19075 -11522
rect 19109 -11556 19176 -11522
rect 19210 -11556 19243 -11522
rect 19045 -11612 19243 -11556
rect 19045 -11646 19075 -11612
rect 19109 -11646 19176 -11612
rect 19210 -11646 19243 -11612
rect 19045 -11702 19243 -11646
rect 19045 -11736 19075 -11702
rect 19109 -11736 19176 -11702
rect 19210 -11736 19243 -11702
rect 19045 -11792 19243 -11736
rect 19045 -11826 19075 -11792
rect 19109 -11826 19176 -11792
rect 19210 -11826 19243 -11792
rect 19045 -11882 19243 -11826
rect 19045 -11916 19075 -11882
rect 19109 -11916 19176 -11882
rect 19210 -11916 19243 -11882
rect 19045 -11972 19243 -11916
rect 19045 -12006 19075 -11972
rect 19109 -12006 19176 -11972
rect 19210 -12006 19243 -11972
rect 19045 -12062 19243 -12006
rect 19045 -12096 19075 -12062
rect 19109 -12096 19176 -12062
rect 19210 -12096 19243 -12062
rect 19045 -12152 19243 -12096
rect 19045 -12186 19075 -12152
rect 19109 -12186 19176 -12152
rect 19210 -12186 19243 -12152
rect 19045 -12242 19243 -12186
rect 19045 -12276 19075 -12242
rect 19109 -12276 19176 -12242
rect 19210 -12276 19243 -12242
rect 19045 -12332 19243 -12276
rect 19045 -12366 19075 -12332
rect 19109 -12366 19176 -12332
rect 19210 -12366 19243 -12332
rect 19045 -12402 19243 -12366
rect 19307 -11518 19439 -11502
rect 19473 -11518 19529 -11484
rect 19563 -11518 19619 -11484
rect 19653 -11518 19709 -11484
rect 19743 -11518 19799 -11484
rect 19833 -11518 19889 -11484
rect 19923 -11518 19979 -11484
rect 20013 -11518 20069 -11484
rect 20103 -11518 20159 -11484
rect 20193 -11502 20727 -11484
rect 20193 -11518 20269 -11502
rect 19307 -11537 20269 -11518
rect 19307 -11562 19379 -11537
rect 19307 -11596 19326 -11562
rect 19360 -11596 19379 -11562
rect 19307 -11652 19379 -11596
rect 20197 -11596 20269 -11537
rect 19307 -11686 19326 -11652
rect 19360 -11686 19379 -11652
rect 19307 -11742 19379 -11686
rect 19307 -11776 19326 -11742
rect 19360 -11776 19379 -11742
rect 19307 -11832 19379 -11776
rect 19307 -11866 19326 -11832
rect 19360 -11866 19379 -11832
rect 19307 -11922 19379 -11866
rect 19307 -11956 19326 -11922
rect 19360 -11956 19379 -11922
rect 19307 -12012 19379 -11956
rect 19307 -12046 19326 -12012
rect 19360 -12046 19379 -12012
rect 19307 -12102 19379 -12046
rect 19307 -12136 19326 -12102
rect 19360 -12136 19379 -12102
rect 19307 -12192 19379 -12136
rect 19307 -12226 19326 -12192
rect 19360 -12226 19379 -12192
rect 19307 -12282 19379 -12226
rect 19307 -12316 19326 -12282
rect 19360 -12316 19379 -12282
rect 19441 -11660 20135 -11599
rect 19441 -11694 19502 -11660
rect 19536 -11672 19592 -11660
rect 19626 -11672 19682 -11660
rect 19716 -11672 19772 -11660
rect 19548 -11694 19592 -11672
rect 19648 -11694 19682 -11672
rect 19748 -11694 19772 -11672
rect 19806 -11672 19862 -11660
rect 19806 -11694 19814 -11672
rect 19441 -11706 19514 -11694
rect 19548 -11706 19614 -11694
rect 19648 -11706 19714 -11694
rect 19748 -11706 19814 -11694
rect 19848 -11694 19862 -11672
rect 19896 -11672 19952 -11660
rect 19896 -11694 19914 -11672
rect 19848 -11706 19914 -11694
rect 19948 -11694 19952 -11672
rect 19986 -11672 20042 -11660
rect 19986 -11694 20014 -11672
rect 20076 -11694 20135 -11660
rect 19948 -11706 20014 -11694
rect 20048 -11706 20135 -11694
rect 19441 -11750 20135 -11706
rect 19441 -11784 19502 -11750
rect 19536 -11772 19592 -11750
rect 19626 -11772 19682 -11750
rect 19716 -11772 19772 -11750
rect 19548 -11784 19592 -11772
rect 19648 -11784 19682 -11772
rect 19748 -11784 19772 -11772
rect 19806 -11772 19862 -11750
rect 19806 -11784 19814 -11772
rect 19441 -11806 19514 -11784
rect 19548 -11806 19614 -11784
rect 19648 -11806 19714 -11784
rect 19748 -11806 19814 -11784
rect 19848 -11784 19862 -11772
rect 19896 -11772 19952 -11750
rect 19896 -11784 19914 -11772
rect 19848 -11806 19914 -11784
rect 19948 -11784 19952 -11772
rect 19986 -11772 20042 -11750
rect 19986 -11784 20014 -11772
rect 20076 -11784 20135 -11750
rect 19948 -11806 20014 -11784
rect 20048 -11806 20135 -11784
rect 19441 -11840 20135 -11806
rect 19441 -11874 19502 -11840
rect 19536 -11872 19592 -11840
rect 19626 -11872 19682 -11840
rect 19716 -11872 19772 -11840
rect 19548 -11874 19592 -11872
rect 19648 -11874 19682 -11872
rect 19748 -11874 19772 -11872
rect 19806 -11872 19862 -11840
rect 19806 -11874 19814 -11872
rect 19441 -11906 19514 -11874
rect 19548 -11906 19614 -11874
rect 19648 -11906 19714 -11874
rect 19748 -11906 19814 -11874
rect 19848 -11874 19862 -11872
rect 19896 -11872 19952 -11840
rect 19896 -11874 19914 -11872
rect 19848 -11906 19914 -11874
rect 19948 -11874 19952 -11872
rect 19986 -11872 20042 -11840
rect 19986 -11874 20014 -11872
rect 20076 -11874 20135 -11840
rect 19948 -11906 20014 -11874
rect 20048 -11906 20135 -11874
rect 19441 -11930 20135 -11906
rect 19441 -11964 19502 -11930
rect 19536 -11964 19592 -11930
rect 19626 -11964 19682 -11930
rect 19716 -11964 19772 -11930
rect 19806 -11964 19862 -11930
rect 19896 -11964 19952 -11930
rect 19986 -11964 20042 -11930
rect 20076 -11964 20135 -11930
rect 19441 -11972 20135 -11964
rect 19441 -12006 19514 -11972
rect 19548 -12006 19614 -11972
rect 19648 -12006 19714 -11972
rect 19748 -12006 19814 -11972
rect 19848 -12006 19914 -11972
rect 19948 -12006 20014 -11972
rect 20048 -12006 20135 -11972
rect 19441 -12020 20135 -12006
rect 19441 -12054 19502 -12020
rect 19536 -12054 19592 -12020
rect 19626 -12054 19682 -12020
rect 19716 -12054 19772 -12020
rect 19806 -12054 19862 -12020
rect 19896 -12054 19952 -12020
rect 19986 -12054 20042 -12020
rect 20076 -12054 20135 -12020
rect 19441 -12072 20135 -12054
rect 19441 -12106 19514 -12072
rect 19548 -12106 19614 -12072
rect 19648 -12106 19714 -12072
rect 19748 -12106 19814 -12072
rect 19848 -12106 19914 -12072
rect 19948 -12106 20014 -12072
rect 20048 -12106 20135 -12072
rect 19441 -12110 20135 -12106
rect 19441 -12144 19502 -12110
rect 19536 -12144 19592 -12110
rect 19626 -12144 19682 -12110
rect 19716 -12144 19772 -12110
rect 19806 -12144 19862 -12110
rect 19896 -12144 19952 -12110
rect 19986 -12144 20042 -12110
rect 20076 -12144 20135 -12110
rect 19441 -12172 20135 -12144
rect 19441 -12200 19514 -12172
rect 19548 -12200 19614 -12172
rect 19648 -12200 19714 -12172
rect 19748 -12200 19814 -12172
rect 19441 -12234 19502 -12200
rect 19548 -12206 19592 -12200
rect 19648 -12206 19682 -12200
rect 19748 -12206 19772 -12200
rect 19536 -12234 19592 -12206
rect 19626 -12234 19682 -12206
rect 19716 -12234 19772 -12206
rect 19806 -12206 19814 -12200
rect 19848 -12200 19914 -12172
rect 19848 -12206 19862 -12200
rect 19806 -12234 19862 -12206
rect 19896 -12206 19914 -12200
rect 19948 -12200 20014 -12172
rect 20048 -12200 20135 -12172
rect 19948 -12206 19952 -12200
rect 19896 -12234 19952 -12206
rect 19986 -12206 20014 -12200
rect 19986 -12234 20042 -12206
rect 20076 -12234 20135 -12200
rect 19441 -12293 20135 -12234
rect 20197 -11630 20216 -11596
rect 20250 -11630 20269 -11596
rect 20197 -11686 20269 -11630
rect 20197 -11720 20216 -11686
rect 20250 -11720 20269 -11686
rect 20197 -11776 20269 -11720
rect 20197 -11810 20216 -11776
rect 20250 -11810 20269 -11776
rect 20197 -11866 20269 -11810
rect 20197 -11900 20216 -11866
rect 20250 -11900 20269 -11866
rect 20197 -11956 20269 -11900
rect 20197 -11990 20216 -11956
rect 20250 -11990 20269 -11956
rect 20197 -12046 20269 -11990
rect 20197 -12080 20216 -12046
rect 20250 -12080 20269 -12046
rect 20197 -12136 20269 -12080
rect 20197 -12170 20216 -12136
rect 20250 -12170 20269 -12136
rect 20197 -12226 20269 -12170
rect 20197 -12260 20216 -12226
rect 20250 -12260 20269 -12226
rect 19307 -12355 19379 -12316
rect 20197 -12316 20269 -12260
rect 20197 -12350 20216 -12316
rect 20250 -12350 20269 -12316
rect 20197 -12355 20269 -12350
rect 19307 -12374 20269 -12355
rect 19307 -12402 19420 -12374
rect 18886 -12408 19420 -12402
rect 19454 -12408 19510 -12374
rect 19544 -12408 19600 -12374
rect 19634 -12408 19690 -12374
rect 19724 -12408 19780 -12374
rect 19814 -12408 19870 -12374
rect 19904 -12408 19960 -12374
rect 19994 -12408 20050 -12374
rect 20084 -12408 20140 -12374
rect 20174 -12402 20269 -12374
rect 20333 -11522 20531 -11502
rect 20333 -11556 20363 -11522
rect 20397 -11556 20464 -11522
rect 20498 -11556 20531 -11522
rect 20333 -11612 20531 -11556
rect 20333 -11646 20363 -11612
rect 20397 -11646 20464 -11612
rect 20498 -11646 20531 -11612
rect 20333 -11702 20531 -11646
rect 20333 -11736 20363 -11702
rect 20397 -11736 20464 -11702
rect 20498 -11736 20531 -11702
rect 20333 -11792 20531 -11736
rect 20333 -11826 20363 -11792
rect 20397 -11826 20464 -11792
rect 20498 -11826 20531 -11792
rect 20333 -11882 20531 -11826
rect 20333 -11916 20363 -11882
rect 20397 -11916 20464 -11882
rect 20498 -11916 20531 -11882
rect 20333 -11972 20531 -11916
rect 20333 -12006 20363 -11972
rect 20397 -12006 20464 -11972
rect 20498 -12006 20531 -11972
rect 20333 -12062 20531 -12006
rect 20333 -12096 20363 -12062
rect 20397 -12096 20464 -12062
rect 20498 -12096 20531 -12062
rect 20333 -12152 20531 -12096
rect 20333 -12186 20363 -12152
rect 20397 -12186 20464 -12152
rect 20498 -12186 20531 -12152
rect 20333 -12242 20531 -12186
rect 20333 -12276 20363 -12242
rect 20397 -12276 20464 -12242
rect 20498 -12276 20531 -12242
rect 20333 -12332 20531 -12276
rect 20333 -12366 20363 -12332
rect 20397 -12366 20464 -12332
rect 20498 -12366 20531 -12332
rect 20333 -12402 20531 -12366
rect 20595 -11518 20727 -11502
rect 20761 -11518 20817 -11484
rect 20851 -11518 20907 -11484
rect 20941 -11518 20997 -11484
rect 21031 -11518 21087 -11484
rect 21121 -11518 21177 -11484
rect 21211 -11518 21267 -11484
rect 21301 -11518 21357 -11484
rect 21391 -11518 21447 -11484
rect 21481 -11502 22015 -11484
rect 21481 -11518 21557 -11502
rect 20595 -11537 21557 -11518
rect 20595 -11562 20667 -11537
rect 20595 -11596 20614 -11562
rect 20648 -11596 20667 -11562
rect 20595 -11652 20667 -11596
rect 21485 -11596 21557 -11537
rect 20595 -11686 20614 -11652
rect 20648 -11686 20667 -11652
rect 20595 -11742 20667 -11686
rect 20595 -11776 20614 -11742
rect 20648 -11776 20667 -11742
rect 20595 -11832 20667 -11776
rect 20595 -11866 20614 -11832
rect 20648 -11866 20667 -11832
rect 20595 -11922 20667 -11866
rect 20595 -11956 20614 -11922
rect 20648 -11956 20667 -11922
rect 20595 -12012 20667 -11956
rect 20595 -12046 20614 -12012
rect 20648 -12046 20667 -12012
rect 20595 -12102 20667 -12046
rect 20595 -12136 20614 -12102
rect 20648 -12136 20667 -12102
rect 20595 -12192 20667 -12136
rect 20595 -12226 20614 -12192
rect 20648 -12226 20667 -12192
rect 20595 -12282 20667 -12226
rect 20595 -12316 20614 -12282
rect 20648 -12316 20667 -12282
rect 20729 -11660 21423 -11599
rect 20729 -11694 20790 -11660
rect 20824 -11672 20880 -11660
rect 20914 -11672 20970 -11660
rect 21004 -11672 21060 -11660
rect 20836 -11694 20880 -11672
rect 20936 -11694 20970 -11672
rect 21036 -11694 21060 -11672
rect 21094 -11672 21150 -11660
rect 21094 -11694 21102 -11672
rect 20729 -11706 20802 -11694
rect 20836 -11706 20902 -11694
rect 20936 -11706 21002 -11694
rect 21036 -11706 21102 -11694
rect 21136 -11694 21150 -11672
rect 21184 -11672 21240 -11660
rect 21184 -11694 21202 -11672
rect 21136 -11706 21202 -11694
rect 21236 -11694 21240 -11672
rect 21274 -11672 21330 -11660
rect 21274 -11694 21302 -11672
rect 21364 -11694 21423 -11660
rect 21236 -11706 21302 -11694
rect 21336 -11706 21423 -11694
rect 20729 -11750 21423 -11706
rect 20729 -11784 20790 -11750
rect 20824 -11772 20880 -11750
rect 20914 -11772 20970 -11750
rect 21004 -11772 21060 -11750
rect 20836 -11784 20880 -11772
rect 20936 -11784 20970 -11772
rect 21036 -11784 21060 -11772
rect 21094 -11772 21150 -11750
rect 21094 -11784 21102 -11772
rect 20729 -11806 20802 -11784
rect 20836 -11806 20902 -11784
rect 20936 -11806 21002 -11784
rect 21036 -11806 21102 -11784
rect 21136 -11784 21150 -11772
rect 21184 -11772 21240 -11750
rect 21184 -11784 21202 -11772
rect 21136 -11806 21202 -11784
rect 21236 -11784 21240 -11772
rect 21274 -11772 21330 -11750
rect 21274 -11784 21302 -11772
rect 21364 -11784 21423 -11750
rect 21236 -11806 21302 -11784
rect 21336 -11806 21423 -11784
rect 20729 -11840 21423 -11806
rect 20729 -11874 20790 -11840
rect 20824 -11872 20880 -11840
rect 20914 -11872 20970 -11840
rect 21004 -11872 21060 -11840
rect 20836 -11874 20880 -11872
rect 20936 -11874 20970 -11872
rect 21036 -11874 21060 -11872
rect 21094 -11872 21150 -11840
rect 21094 -11874 21102 -11872
rect 20729 -11906 20802 -11874
rect 20836 -11906 20902 -11874
rect 20936 -11906 21002 -11874
rect 21036 -11906 21102 -11874
rect 21136 -11874 21150 -11872
rect 21184 -11872 21240 -11840
rect 21184 -11874 21202 -11872
rect 21136 -11906 21202 -11874
rect 21236 -11874 21240 -11872
rect 21274 -11872 21330 -11840
rect 21274 -11874 21302 -11872
rect 21364 -11874 21423 -11840
rect 21236 -11906 21302 -11874
rect 21336 -11906 21423 -11874
rect 20729 -11930 21423 -11906
rect 20729 -11964 20790 -11930
rect 20824 -11964 20880 -11930
rect 20914 -11964 20970 -11930
rect 21004 -11964 21060 -11930
rect 21094 -11964 21150 -11930
rect 21184 -11964 21240 -11930
rect 21274 -11964 21330 -11930
rect 21364 -11964 21423 -11930
rect 20729 -11972 21423 -11964
rect 20729 -12006 20802 -11972
rect 20836 -12006 20902 -11972
rect 20936 -12006 21002 -11972
rect 21036 -12006 21102 -11972
rect 21136 -12006 21202 -11972
rect 21236 -12006 21302 -11972
rect 21336 -12006 21423 -11972
rect 20729 -12020 21423 -12006
rect 20729 -12054 20790 -12020
rect 20824 -12054 20880 -12020
rect 20914 -12054 20970 -12020
rect 21004 -12054 21060 -12020
rect 21094 -12054 21150 -12020
rect 21184 -12054 21240 -12020
rect 21274 -12054 21330 -12020
rect 21364 -12054 21423 -12020
rect 20729 -12072 21423 -12054
rect 20729 -12106 20802 -12072
rect 20836 -12106 20902 -12072
rect 20936 -12106 21002 -12072
rect 21036 -12106 21102 -12072
rect 21136 -12106 21202 -12072
rect 21236 -12106 21302 -12072
rect 21336 -12106 21423 -12072
rect 20729 -12110 21423 -12106
rect 20729 -12144 20790 -12110
rect 20824 -12144 20880 -12110
rect 20914 -12144 20970 -12110
rect 21004 -12144 21060 -12110
rect 21094 -12144 21150 -12110
rect 21184 -12144 21240 -12110
rect 21274 -12144 21330 -12110
rect 21364 -12144 21423 -12110
rect 20729 -12172 21423 -12144
rect 20729 -12200 20802 -12172
rect 20836 -12200 20902 -12172
rect 20936 -12200 21002 -12172
rect 21036 -12200 21102 -12172
rect 20729 -12234 20790 -12200
rect 20836 -12206 20880 -12200
rect 20936 -12206 20970 -12200
rect 21036 -12206 21060 -12200
rect 20824 -12234 20880 -12206
rect 20914 -12234 20970 -12206
rect 21004 -12234 21060 -12206
rect 21094 -12206 21102 -12200
rect 21136 -12200 21202 -12172
rect 21136 -12206 21150 -12200
rect 21094 -12234 21150 -12206
rect 21184 -12206 21202 -12200
rect 21236 -12200 21302 -12172
rect 21336 -12200 21423 -12172
rect 21236 -12206 21240 -12200
rect 21184 -12234 21240 -12206
rect 21274 -12206 21302 -12200
rect 21274 -12234 21330 -12206
rect 21364 -12234 21423 -12200
rect 20729 -12293 21423 -12234
rect 21485 -11630 21504 -11596
rect 21538 -11630 21557 -11596
rect 21485 -11686 21557 -11630
rect 21485 -11720 21504 -11686
rect 21538 -11720 21557 -11686
rect 21485 -11776 21557 -11720
rect 21485 -11810 21504 -11776
rect 21538 -11810 21557 -11776
rect 21485 -11866 21557 -11810
rect 21485 -11900 21504 -11866
rect 21538 -11900 21557 -11866
rect 21485 -11956 21557 -11900
rect 21485 -11990 21504 -11956
rect 21538 -11990 21557 -11956
rect 21485 -12046 21557 -11990
rect 21485 -12080 21504 -12046
rect 21538 -12080 21557 -12046
rect 21485 -12136 21557 -12080
rect 21485 -12170 21504 -12136
rect 21538 -12170 21557 -12136
rect 21485 -12226 21557 -12170
rect 21485 -12260 21504 -12226
rect 21538 -12260 21557 -12226
rect 20595 -12355 20667 -12316
rect 21485 -12316 21557 -12260
rect 21485 -12350 21504 -12316
rect 21538 -12350 21557 -12316
rect 21485 -12355 21557 -12350
rect 20595 -12374 21557 -12355
rect 20595 -12402 20708 -12374
rect 20174 -12408 20708 -12402
rect 20742 -12408 20798 -12374
rect 20832 -12408 20888 -12374
rect 20922 -12408 20978 -12374
rect 21012 -12408 21068 -12374
rect 21102 -12408 21158 -12374
rect 21192 -12408 21248 -12374
rect 21282 -12408 21338 -12374
rect 21372 -12408 21428 -12374
rect 21462 -12402 21557 -12374
rect 21621 -11522 21819 -11502
rect 21621 -11556 21651 -11522
rect 21685 -11556 21752 -11522
rect 21786 -11556 21819 -11522
rect 21621 -11612 21819 -11556
rect 21621 -11646 21651 -11612
rect 21685 -11646 21752 -11612
rect 21786 -11646 21819 -11612
rect 21621 -11702 21819 -11646
rect 21621 -11736 21651 -11702
rect 21685 -11736 21752 -11702
rect 21786 -11736 21819 -11702
rect 21621 -11792 21819 -11736
rect 21621 -11826 21651 -11792
rect 21685 -11826 21752 -11792
rect 21786 -11826 21819 -11792
rect 21621 -11882 21819 -11826
rect 21621 -11916 21651 -11882
rect 21685 -11916 21752 -11882
rect 21786 -11916 21819 -11882
rect 21621 -11972 21819 -11916
rect 21621 -12006 21651 -11972
rect 21685 -12006 21752 -11972
rect 21786 -12006 21819 -11972
rect 21621 -12062 21819 -12006
rect 21621 -12096 21651 -12062
rect 21685 -12096 21752 -12062
rect 21786 -12096 21819 -12062
rect 21621 -12152 21819 -12096
rect 21621 -12186 21651 -12152
rect 21685 -12186 21752 -12152
rect 21786 -12186 21819 -12152
rect 21621 -12242 21819 -12186
rect 21621 -12276 21651 -12242
rect 21685 -12276 21752 -12242
rect 21786 -12276 21819 -12242
rect 21621 -12332 21819 -12276
rect 21621 -12366 21651 -12332
rect 21685 -12366 21752 -12332
rect 21786 -12366 21819 -12332
rect 21621 -12402 21819 -12366
rect 21883 -11518 22015 -11502
rect 22049 -11518 22105 -11484
rect 22139 -11518 22195 -11484
rect 22229 -11518 22285 -11484
rect 22319 -11518 22375 -11484
rect 22409 -11518 22465 -11484
rect 22499 -11518 22555 -11484
rect 22589 -11518 22645 -11484
rect 22679 -11518 22735 -11484
rect 22769 -11502 23303 -11484
rect 22769 -11518 22845 -11502
rect 21883 -11537 22845 -11518
rect 21883 -11562 21955 -11537
rect 21883 -11596 21902 -11562
rect 21936 -11596 21955 -11562
rect 21883 -11652 21955 -11596
rect 22773 -11596 22845 -11537
rect 21883 -11686 21902 -11652
rect 21936 -11686 21955 -11652
rect 21883 -11742 21955 -11686
rect 21883 -11776 21902 -11742
rect 21936 -11776 21955 -11742
rect 21883 -11832 21955 -11776
rect 21883 -11866 21902 -11832
rect 21936 -11866 21955 -11832
rect 21883 -11922 21955 -11866
rect 21883 -11956 21902 -11922
rect 21936 -11956 21955 -11922
rect 21883 -12012 21955 -11956
rect 21883 -12046 21902 -12012
rect 21936 -12046 21955 -12012
rect 21883 -12102 21955 -12046
rect 21883 -12136 21902 -12102
rect 21936 -12136 21955 -12102
rect 21883 -12192 21955 -12136
rect 21883 -12226 21902 -12192
rect 21936 -12226 21955 -12192
rect 21883 -12282 21955 -12226
rect 21883 -12316 21902 -12282
rect 21936 -12316 21955 -12282
rect 22017 -11660 22711 -11599
rect 22017 -11694 22078 -11660
rect 22112 -11672 22168 -11660
rect 22202 -11672 22258 -11660
rect 22292 -11672 22348 -11660
rect 22124 -11694 22168 -11672
rect 22224 -11694 22258 -11672
rect 22324 -11694 22348 -11672
rect 22382 -11672 22438 -11660
rect 22382 -11694 22390 -11672
rect 22017 -11706 22090 -11694
rect 22124 -11706 22190 -11694
rect 22224 -11706 22290 -11694
rect 22324 -11706 22390 -11694
rect 22424 -11694 22438 -11672
rect 22472 -11672 22528 -11660
rect 22472 -11694 22490 -11672
rect 22424 -11706 22490 -11694
rect 22524 -11694 22528 -11672
rect 22562 -11672 22618 -11660
rect 22562 -11694 22590 -11672
rect 22652 -11694 22711 -11660
rect 22524 -11706 22590 -11694
rect 22624 -11706 22711 -11694
rect 22017 -11750 22711 -11706
rect 22017 -11784 22078 -11750
rect 22112 -11772 22168 -11750
rect 22202 -11772 22258 -11750
rect 22292 -11772 22348 -11750
rect 22124 -11784 22168 -11772
rect 22224 -11784 22258 -11772
rect 22324 -11784 22348 -11772
rect 22382 -11772 22438 -11750
rect 22382 -11784 22390 -11772
rect 22017 -11806 22090 -11784
rect 22124 -11806 22190 -11784
rect 22224 -11806 22290 -11784
rect 22324 -11806 22390 -11784
rect 22424 -11784 22438 -11772
rect 22472 -11772 22528 -11750
rect 22472 -11784 22490 -11772
rect 22424 -11806 22490 -11784
rect 22524 -11784 22528 -11772
rect 22562 -11772 22618 -11750
rect 22562 -11784 22590 -11772
rect 22652 -11784 22711 -11750
rect 22524 -11806 22590 -11784
rect 22624 -11806 22711 -11784
rect 22017 -11840 22711 -11806
rect 22017 -11874 22078 -11840
rect 22112 -11872 22168 -11840
rect 22202 -11872 22258 -11840
rect 22292 -11872 22348 -11840
rect 22124 -11874 22168 -11872
rect 22224 -11874 22258 -11872
rect 22324 -11874 22348 -11872
rect 22382 -11872 22438 -11840
rect 22382 -11874 22390 -11872
rect 22017 -11906 22090 -11874
rect 22124 -11906 22190 -11874
rect 22224 -11906 22290 -11874
rect 22324 -11906 22390 -11874
rect 22424 -11874 22438 -11872
rect 22472 -11872 22528 -11840
rect 22472 -11874 22490 -11872
rect 22424 -11906 22490 -11874
rect 22524 -11874 22528 -11872
rect 22562 -11872 22618 -11840
rect 22562 -11874 22590 -11872
rect 22652 -11874 22711 -11840
rect 22524 -11906 22590 -11874
rect 22624 -11906 22711 -11874
rect 22017 -11930 22711 -11906
rect 22017 -11964 22078 -11930
rect 22112 -11964 22168 -11930
rect 22202 -11964 22258 -11930
rect 22292 -11964 22348 -11930
rect 22382 -11964 22438 -11930
rect 22472 -11964 22528 -11930
rect 22562 -11964 22618 -11930
rect 22652 -11964 22711 -11930
rect 22017 -11972 22711 -11964
rect 22017 -12006 22090 -11972
rect 22124 -12006 22190 -11972
rect 22224 -12006 22290 -11972
rect 22324 -12006 22390 -11972
rect 22424 -12006 22490 -11972
rect 22524 -12006 22590 -11972
rect 22624 -12006 22711 -11972
rect 22017 -12020 22711 -12006
rect 22017 -12054 22078 -12020
rect 22112 -12054 22168 -12020
rect 22202 -12054 22258 -12020
rect 22292 -12054 22348 -12020
rect 22382 -12054 22438 -12020
rect 22472 -12054 22528 -12020
rect 22562 -12054 22618 -12020
rect 22652 -12054 22711 -12020
rect 22017 -12072 22711 -12054
rect 22017 -12106 22090 -12072
rect 22124 -12106 22190 -12072
rect 22224 -12106 22290 -12072
rect 22324 -12106 22390 -12072
rect 22424 -12106 22490 -12072
rect 22524 -12106 22590 -12072
rect 22624 -12106 22711 -12072
rect 22017 -12110 22711 -12106
rect 22017 -12144 22078 -12110
rect 22112 -12144 22168 -12110
rect 22202 -12144 22258 -12110
rect 22292 -12144 22348 -12110
rect 22382 -12144 22438 -12110
rect 22472 -12144 22528 -12110
rect 22562 -12144 22618 -12110
rect 22652 -12144 22711 -12110
rect 22017 -12172 22711 -12144
rect 22017 -12200 22090 -12172
rect 22124 -12200 22190 -12172
rect 22224 -12200 22290 -12172
rect 22324 -12200 22390 -12172
rect 22017 -12234 22078 -12200
rect 22124 -12206 22168 -12200
rect 22224 -12206 22258 -12200
rect 22324 -12206 22348 -12200
rect 22112 -12234 22168 -12206
rect 22202 -12234 22258 -12206
rect 22292 -12234 22348 -12206
rect 22382 -12206 22390 -12200
rect 22424 -12200 22490 -12172
rect 22424 -12206 22438 -12200
rect 22382 -12234 22438 -12206
rect 22472 -12206 22490 -12200
rect 22524 -12200 22590 -12172
rect 22624 -12200 22711 -12172
rect 22524 -12206 22528 -12200
rect 22472 -12234 22528 -12206
rect 22562 -12206 22590 -12200
rect 22562 -12234 22618 -12206
rect 22652 -12234 22711 -12200
rect 22017 -12293 22711 -12234
rect 22773 -11630 22792 -11596
rect 22826 -11630 22845 -11596
rect 22773 -11686 22845 -11630
rect 22773 -11720 22792 -11686
rect 22826 -11720 22845 -11686
rect 22773 -11776 22845 -11720
rect 22773 -11810 22792 -11776
rect 22826 -11810 22845 -11776
rect 22773 -11866 22845 -11810
rect 22773 -11900 22792 -11866
rect 22826 -11900 22845 -11866
rect 22773 -11956 22845 -11900
rect 22773 -11990 22792 -11956
rect 22826 -11990 22845 -11956
rect 22773 -12046 22845 -11990
rect 22773 -12080 22792 -12046
rect 22826 -12080 22845 -12046
rect 22773 -12136 22845 -12080
rect 22773 -12170 22792 -12136
rect 22826 -12170 22845 -12136
rect 22773 -12226 22845 -12170
rect 22773 -12260 22792 -12226
rect 22826 -12260 22845 -12226
rect 21883 -12355 21955 -12316
rect 22773 -12316 22845 -12260
rect 22773 -12350 22792 -12316
rect 22826 -12350 22845 -12316
rect 22773 -12355 22845 -12350
rect 21883 -12374 22845 -12355
rect 21883 -12402 21996 -12374
rect 21462 -12408 21996 -12402
rect 22030 -12408 22086 -12374
rect 22120 -12408 22176 -12374
rect 22210 -12408 22266 -12374
rect 22300 -12408 22356 -12374
rect 22390 -12408 22446 -12374
rect 22480 -12408 22536 -12374
rect 22570 -12408 22626 -12374
rect 22660 -12408 22716 -12374
rect 22750 -12402 22845 -12374
rect 22909 -11522 23107 -11502
rect 22909 -11556 22939 -11522
rect 22973 -11556 23040 -11522
rect 23074 -11556 23107 -11522
rect 22909 -11612 23107 -11556
rect 22909 -11646 22939 -11612
rect 22973 -11646 23040 -11612
rect 23074 -11646 23107 -11612
rect 22909 -11702 23107 -11646
rect 22909 -11736 22939 -11702
rect 22973 -11736 23040 -11702
rect 23074 -11736 23107 -11702
rect 22909 -11792 23107 -11736
rect 22909 -11826 22939 -11792
rect 22973 -11826 23040 -11792
rect 23074 -11826 23107 -11792
rect 22909 -11882 23107 -11826
rect 22909 -11916 22939 -11882
rect 22973 -11916 23040 -11882
rect 23074 -11916 23107 -11882
rect 22909 -11972 23107 -11916
rect 22909 -12006 22939 -11972
rect 22973 -12006 23040 -11972
rect 23074 -12006 23107 -11972
rect 22909 -12062 23107 -12006
rect 22909 -12096 22939 -12062
rect 22973 -12096 23040 -12062
rect 23074 -12096 23107 -12062
rect 22909 -12152 23107 -12096
rect 22909 -12186 22939 -12152
rect 22973 -12186 23040 -12152
rect 23074 -12186 23107 -12152
rect 22909 -12242 23107 -12186
rect 22909 -12276 22939 -12242
rect 22973 -12276 23040 -12242
rect 23074 -12276 23107 -12242
rect 22909 -12332 23107 -12276
rect 22909 -12366 22939 -12332
rect 22973 -12366 23040 -12332
rect 23074 -12366 23107 -12332
rect 22909 -12402 23107 -12366
rect 23171 -11518 23303 -11502
rect 23337 -11518 23393 -11484
rect 23427 -11518 23483 -11484
rect 23517 -11518 23573 -11484
rect 23607 -11518 23663 -11484
rect 23697 -11518 23753 -11484
rect 23787 -11518 23843 -11484
rect 23877 -11518 23933 -11484
rect 23967 -11518 24023 -11484
rect 24057 -11502 24591 -11484
rect 24057 -11518 24133 -11502
rect 23171 -11537 24133 -11518
rect 23171 -11562 23243 -11537
rect 23171 -11596 23190 -11562
rect 23224 -11596 23243 -11562
rect 23171 -11652 23243 -11596
rect 24061 -11596 24133 -11537
rect 23171 -11686 23190 -11652
rect 23224 -11686 23243 -11652
rect 23171 -11742 23243 -11686
rect 23171 -11776 23190 -11742
rect 23224 -11776 23243 -11742
rect 23171 -11832 23243 -11776
rect 23171 -11866 23190 -11832
rect 23224 -11866 23243 -11832
rect 23171 -11922 23243 -11866
rect 23171 -11956 23190 -11922
rect 23224 -11956 23243 -11922
rect 23171 -12012 23243 -11956
rect 23171 -12046 23190 -12012
rect 23224 -12046 23243 -12012
rect 23171 -12102 23243 -12046
rect 23171 -12136 23190 -12102
rect 23224 -12136 23243 -12102
rect 23171 -12192 23243 -12136
rect 23171 -12226 23190 -12192
rect 23224 -12226 23243 -12192
rect 23171 -12282 23243 -12226
rect 23171 -12316 23190 -12282
rect 23224 -12316 23243 -12282
rect 23305 -11660 23999 -11599
rect 23305 -11694 23366 -11660
rect 23400 -11672 23456 -11660
rect 23490 -11672 23546 -11660
rect 23580 -11672 23636 -11660
rect 23412 -11694 23456 -11672
rect 23512 -11694 23546 -11672
rect 23612 -11694 23636 -11672
rect 23670 -11672 23726 -11660
rect 23670 -11694 23678 -11672
rect 23305 -11706 23378 -11694
rect 23412 -11706 23478 -11694
rect 23512 -11706 23578 -11694
rect 23612 -11706 23678 -11694
rect 23712 -11694 23726 -11672
rect 23760 -11672 23816 -11660
rect 23760 -11694 23778 -11672
rect 23712 -11706 23778 -11694
rect 23812 -11694 23816 -11672
rect 23850 -11672 23906 -11660
rect 23850 -11694 23878 -11672
rect 23940 -11694 23999 -11660
rect 23812 -11706 23878 -11694
rect 23912 -11706 23999 -11694
rect 23305 -11750 23999 -11706
rect 23305 -11784 23366 -11750
rect 23400 -11772 23456 -11750
rect 23490 -11772 23546 -11750
rect 23580 -11772 23636 -11750
rect 23412 -11784 23456 -11772
rect 23512 -11784 23546 -11772
rect 23612 -11784 23636 -11772
rect 23670 -11772 23726 -11750
rect 23670 -11784 23678 -11772
rect 23305 -11806 23378 -11784
rect 23412 -11806 23478 -11784
rect 23512 -11806 23578 -11784
rect 23612 -11806 23678 -11784
rect 23712 -11784 23726 -11772
rect 23760 -11772 23816 -11750
rect 23760 -11784 23778 -11772
rect 23712 -11806 23778 -11784
rect 23812 -11784 23816 -11772
rect 23850 -11772 23906 -11750
rect 23850 -11784 23878 -11772
rect 23940 -11784 23999 -11750
rect 23812 -11806 23878 -11784
rect 23912 -11806 23999 -11784
rect 23305 -11840 23999 -11806
rect 23305 -11874 23366 -11840
rect 23400 -11872 23456 -11840
rect 23490 -11872 23546 -11840
rect 23580 -11872 23636 -11840
rect 23412 -11874 23456 -11872
rect 23512 -11874 23546 -11872
rect 23612 -11874 23636 -11872
rect 23670 -11872 23726 -11840
rect 23670 -11874 23678 -11872
rect 23305 -11906 23378 -11874
rect 23412 -11906 23478 -11874
rect 23512 -11906 23578 -11874
rect 23612 -11906 23678 -11874
rect 23712 -11874 23726 -11872
rect 23760 -11872 23816 -11840
rect 23760 -11874 23778 -11872
rect 23712 -11906 23778 -11874
rect 23812 -11874 23816 -11872
rect 23850 -11872 23906 -11840
rect 23850 -11874 23878 -11872
rect 23940 -11874 23999 -11840
rect 23812 -11906 23878 -11874
rect 23912 -11906 23999 -11874
rect 23305 -11930 23999 -11906
rect 23305 -11964 23366 -11930
rect 23400 -11964 23456 -11930
rect 23490 -11964 23546 -11930
rect 23580 -11964 23636 -11930
rect 23670 -11964 23726 -11930
rect 23760 -11964 23816 -11930
rect 23850 -11964 23906 -11930
rect 23940 -11964 23999 -11930
rect 23305 -11972 23999 -11964
rect 23305 -12006 23378 -11972
rect 23412 -12006 23478 -11972
rect 23512 -12006 23578 -11972
rect 23612 -12006 23678 -11972
rect 23712 -12006 23778 -11972
rect 23812 -12006 23878 -11972
rect 23912 -12006 23999 -11972
rect 23305 -12020 23999 -12006
rect 23305 -12054 23366 -12020
rect 23400 -12054 23456 -12020
rect 23490 -12054 23546 -12020
rect 23580 -12054 23636 -12020
rect 23670 -12054 23726 -12020
rect 23760 -12054 23816 -12020
rect 23850 -12054 23906 -12020
rect 23940 -12054 23999 -12020
rect 23305 -12072 23999 -12054
rect 23305 -12106 23378 -12072
rect 23412 -12106 23478 -12072
rect 23512 -12106 23578 -12072
rect 23612 -12106 23678 -12072
rect 23712 -12106 23778 -12072
rect 23812 -12106 23878 -12072
rect 23912 -12106 23999 -12072
rect 23305 -12110 23999 -12106
rect 23305 -12144 23366 -12110
rect 23400 -12144 23456 -12110
rect 23490 -12144 23546 -12110
rect 23580 -12144 23636 -12110
rect 23670 -12144 23726 -12110
rect 23760 -12144 23816 -12110
rect 23850 -12144 23906 -12110
rect 23940 -12144 23999 -12110
rect 23305 -12172 23999 -12144
rect 23305 -12200 23378 -12172
rect 23412 -12200 23478 -12172
rect 23512 -12200 23578 -12172
rect 23612 -12200 23678 -12172
rect 23305 -12234 23366 -12200
rect 23412 -12206 23456 -12200
rect 23512 -12206 23546 -12200
rect 23612 -12206 23636 -12200
rect 23400 -12234 23456 -12206
rect 23490 -12234 23546 -12206
rect 23580 -12234 23636 -12206
rect 23670 -12206 23678 -12200
rect 23712 -12200 23778 -12172
rect 23712 -12206 23726 -12200
rect 23670 -12234 23726 -12206
rect 23760 -12206 23778 -12200
rect 23812 -12200 23878 -12172
rect 23912 -12200 23999 -12172
rect 23812 -12206 23816 -12200
rect 23760 -12234 23816 -12206
rect 23850 -12206 23878 -12200
rect 23850 -12234 23906 -12206
rect 23940 -12234 23999 -12200
rect 23305 -12293 23999 -12234
rect 24061 -11630 24080 -11596
rect 24114 -11630 24133 -11596
rect 24061 -11686 24133 -11630
rect 24061 -11720 24080 -11686
rect 24114 -11720 24133 -11686
rect 24061 -11776 24133 -11720
rect 24061 -11810 24080 -11776
rect 24114 -11810 24133 -11776
rect 24061 -11866 24133 -11810
rect 24061 -11900 24080 -11866
rect 24114 -11900 24133 -11866
rect 24061 -11956 24133 -11900
rect 24061 -11990 24080 -11956
rect 24114 -11990 24133 -11956
rect 24061 -12046 24133 -11990
rect 24061 -12080 24080 -12046
rect 24114 -12080 24133 -12046
rect 24061 -12136 24133 -12080
rect 24061 -12170 24080 -12136
rect 24114 -12170 24133 -12136
rect 24061 -12226 24133 -12170
rect 24061 -12260 24080 -12226
rect 24114 -12260 24133 -12226
rect 23171 -12355 23243 -12316
rect 24061 -12316 24133 -12260
rect 24061 -12350 24080 -12316
rect 24114 -12350 24133 -12316
rect 24061 -12355 24133 -12350
rect 23171 -12374 24133 -12355
rect 23171 -12402 23284 -12374
rect 22750 -12408 23284 -12402
rect 23318 -12408 23374 -12374
rect 23408 -12408 23464 -12374
rect 23498 -12408 23554 -12374
rect 23588 -12408 23644 -12374
rect 23678 -12408 23734 -12374
rect 23768 -12408 23824 -12374
rect 23858 -12408 23914 -12374
rect 23948 -12408 24004 -12374
rect 24038 -12402 24133 -12374
rect 24197 -11522 24395 -11502
rect 24197 -11556 24227 -11522
rect 24261 -11556 24328 -11522
rect 24362 -11556 24395 -11522
rect 24197 -11612 24395 -11556
rect 24197 -11646 24227 -11612
rect 24261 -11646 24328 -11612
rect 24362 -11646 24395 -11612
rect 24197 -11702 24395 -11646
rect 24197 -11736 24227 -11702
rect 24261 -11736 24328 -11702
rect 24362 -11736 24395 -11702
rect 24197 -11792 24395 -11736
rect 24197 -11826 24227 -11792
rect 24261 -11826 24328 -11792
rect 24362 -11826 24395 -11792
rect 24197 -11882 24395 -11826
rect 24197 -11916 24227 -11882
rect 24261 -11916 24328 -11882
rect 24362 -11916 24395 -11882
rect 24197 -11972 24395 -11916
rect 24197 -12006 24227 -11972
rect 24261 -12006 24328 -11972
rect 24362 -12006 24395 -11972
rect 24197 -12062 24395 -12006
rect 24197 -12096 24227 -12062
rect 24261 -12096 24328 -12062
rect 24362 -12096 24395 -12062
rect 24197 -12152 24395 -12096
rect 24197 -12186 24227 -12152
rect 24261 -12186 24328 -12152
rect 24362 -12186 24395 -12152
rect 24197 -12242 24395 -12186
rect 24197 -12276 24227 -12242
rect 24261 -12276 24328 -12242
rect 24362 -12276 24395 -12242
rect 24197 -12332 24395 -12276
rect 24197 -12366 24227 -12332
rect 24261 -12366 24328 -12332
rect 24362 -12366 24395 -12332
rect 24197 -12402 24395 -12366
rect 24459 -11518 24591 -11502
rect 24625 -11518 24681 -11484
rect 24715 -11518 24771 -11484
rect 24805 -11518 24861 -11484
rect 24895 -11518 24951 -11484
rect 24985 -11518 25041 -11484
rect 25075 -11518 25131 -11484
rect 25165 -11518 25221 -11484
rect 25255 -11518 25311 -11484
rect 25345 -11502 25879 -11484
rect 25345 -11518 25421 -11502
rect 24459 -11537 25421 -11518
rect 24459 -11562 24531 -11537
rect 24459 -11596 24478 -11562
rect 24512 -11596 24531 -11562
rect 24459 -11652 24531 -11596
rect 25349 -11596 25421 -11537
rect 24459 -11686 24478 -11652
rect 24512 -11686 24531 -11652
rect 24459 -11742 24531 -11686
rect 24459 -11776 24478 -11742
rect 24512 -11776 24531 -11742
rect 24459 -11832 24531 -11776
rect 24459 -11866 24478 -11832
rect 24512 -11866 24531 -11832
rect 24459 -11922 24531 -11866
rect 24459 -11956 24478 -11922
rect 24512 -11956 24531 -11922
rect 24459 -12012 24531 -11956
rect 24459 -12046 24478 -12012
rect 24512 -12046 24531 -12012
rect 24459 -12102 24531 -12046
rect 24459 -12136 24478 -12102
rect 24512 -12136 24531 -12102
rect 24459 -12192 24531 -12136
rect 24459 -12226 24478 -12192
rect 24512 -12226 24531 -12192
rect 24459 -12282 24531 -12226
rect 24459 -12316 24478 -12282
rect 24512 -12316 24531 -12282
rect 24593 -11660 25287 -11599
rect 24593 -11694 24654 -11660
rect 24688 -11672 24744 -11660
rect 24778 -11672 24834 -11660
rect 24868 -11672 24924 -11660
rect 24700 -11694 24744 -11672
rect 24800 -11694 24834 -11672
rect 24900 -11694 24924 -11672
rect 24958 -11672 25014 -11660
rect 24958 -11694 24966 -11672
rect 24593 -11706 24666 -11694
rect 24700 -11706 24766 -11694
rect 24800 -11706 24866 -11694
rect 24900 -11706 24966 -11694
rect 25000 -11694 25014 -11672
rect 25048 -11672 25104 -11660
rect 25048 -11694 25066 -11672
rect 25000 -11706 25066 -11694
rect 25100 -11694 25104 -11672
rect 25138 -11672 25194 -11660
rect 25138 -11694 25166 -11672
rect 25228 -11694 25287 -11660
rect 25100 -11706 25166 -11694
rect 25200 -11706 25287 -11694
rect 24593 -11750 25287 -11706
rect 24593 -11784 24654 -11750
rect 24688 -11772 24744 -11750
rect 24778 -11772 24834 -11750
rect 24868 -11772 24924 -11750
rect 24700 -11784 24744 -11772
rect 24800 -11784 24834 -11772
rect 24900 -11784 24924 -11772
rect 24958 -11772 25014 -11750
rect 24958 -11784 24966 -11772
rect 24593 -11806 24666 -11784
rect 24700 -11806 24766 -11784
rect 24800 -11806 24866 -11784
rect 24900 -11806 24966 -11784
rect 25000 -11784 25014 -11772
rect 25048 -11772 25104 -11750
rect 25048 -11784 25066 -11772
rect 25000 -11806 25066 -11784
rect 25100 -11784 25104 -11772
rect 25138 -11772 25194 -11750
rect 25138 -11784 25166 -11772
rect 25228 -11784 25287 -11750
rect 25100 -11806 25166 -11784
rect 25200 -11806 25287 -11784
rect 24593 -11840 25287 -11806
rect 24593 -11874 24654 -11840
rect 24688 -11872 24744 -11840
rect 24778 -11872 24834 -11840
rect 24868 -11872 24924 -11840
rect 24700 -11874 24744 -11872
rect 24800 -11874 24834 -11872
rect 24900 -11874 24924 -11872
rect 24958 -11872 25014 -11840
rect 24958 -11874 24966 -11872
rect 24593 -11906 24666 -11874
rect 24700 -11906 24766 -11874
rect 24800 -11906 24866 -11874
rect 24900 -11906 24966 -11874
rect 25000 -11874 25014 -11872
rect 25048 -11872 25104 -11840
rect 25048 -11874 25066 -11872
rect 25000 -11906 25066 -11874
rect 25100 -11874 25104 -11872
rect 25138 -11872 25194 -11840
rect 25138 -11874 25166 -11872
rect 25228 -11874 25287 -11840
rect 25100 -11906 25166 -11874
rect 25200 -11906 25287 -11874
rect 24593 -11930 25287 -11906
rect 24593 -11964 24654 -11930
rect 24688 -11964 24744 -11930
rect 24778 -11964 24834 -11930
rect 24868 -11964 24924 -11930
rect 24958 -11964 25014 -11930
rect 25048 -11964 25104 -11930
rect 25138 -11964 25194 -11930
rect 25228 -11964 25287 -11930
rect 24593 -11972 25287 -11964
rect 24593 -12006 24666 -11972
rect 24700 -12006 24766 -11972
rect 24800 -12006 24866 -11972
rect 24900 -12006 24966 -11972
rect 25000 -12006 25066 -11972
rect 25100 -12006 25166 -11972
rect 25200 -12006 25287 -11972
rect 24593 -12020 25287 -12006
rect 24593 -12054 24654 -12020
rect 24688 -12054 24744 -12020
rect 24778 -12054 24834 -12020
rect 24868 -12054 24924 -12020
rect 24958 -12054 25014 -12020
rect 25048 -12054 25104 -12020
rect 25138 -12054 25194 -12020
rect 25228 -12054 25287 -12020
rect 24593 -12072 25287 -12054
rect 24593 -12106 24666 -12072
rect 24700 -12106 24766 -12072
rect 24800 -12106 24866 -12072
rect 24900 -12106 24966 -12072
rect 25000 -12106 25066 -12072
rect 25100 -12106 25166 -12072
rect 25200 -12106 25287 -12072
rect 24593 -12110 25287 -12106
rect 24593 -12144 24654 -12110
rect 24688 -12144 24744 -12110
rect 24778 -12144 24834 -12110
rect 24868 -12144 24924 -12110
rect 24958 -12144 25014 -12110
rect 25048 -12144 25104 -12110
rect 25138 -12144 25194 -12110
rect 25228 -12144 25287 -12110
rect 24593 -12172 25287 -12144
rect 24593 -12200 24666 -12172
rect 24700 -12200 24766 -12172
rect 24800 -12200 24866 -12172
rect 24900 -12200 24966 -12172
rect 24593 -12234 24654 -12200
rect 24700 -12206 24744 -12200
rect 24800 -12206 24834 -12200
rect 24900 -12206 24924 -12200
rect 24688 -12234 24744 -12206
rect 24778 -12234 24834 -12206
rect 24868 -12234 24924 -12206
rect 24958 -12206 24966 -12200
rect 25000 -12200 25066 -12172
rect 25000 -12206 25014 -12200
rect 24958 -12234 25014 -12206
rect 25048 -12206 25066 -12200
rect 25100 -12200 25166 -12172
rect 25200 -12200 25287 -12172
rect 25100 -12206 25104 -12200
rect 25048 -12234 25104 -12206
rect 25138 -12206 25166 -12200
rect 25138 -12234 25194 -12206
rect 25228 -12234 25287 -12200
rect 24593 -12293 25287 -12234
rect 25349 -11630 25368 -11596
rect 25402 -11630 25421 -11596
rect 25349 -11686 25421 -11630
rect 25349 -11720 25368 -11686
rect 25402 -11720 25421 -11686
rect 25349 -11776 25421 -11720
rect 25349 -11810 25368 -11776
rect 25402 -11810 25421 -11776
rect 25349 -11866 25421 -11810
rect 25349 -11900 25368 -11866
rect 25402 -11900 25421 -11866
rect 25349 -11956 25421 -11900
rect 25349 -11990 25368 -11956
rect 25402 -11990 25421 -11956
rect 25349 -12046 25421 -11990
rect 25349 -12080 25368 -12046
rect 25402 -12080 25421 -12046
rect 25349 -12136 25421 -12080
rect 25349 -12170 25368 -12136
rect 25402 -12170 25421 -12136
rect 25349 -12226 25421 -12170
rect 25349 -12260 25368 -12226
rect 25402 -12260 25421 -12226
rect 24459 -12355 24531 -12316
rect 25349 -12316 25421 -12260
rect 25349 -12350 25368 -12316
rect 25402 -12350 25421 -12316
rect 25349 -12355 25421 -12350
rect 24459 -12374 25421 -12355
rect 24459 -12402 24572 -12374
rect 24038 -12408 24572 -12402
rect 24606 -12408 24662 -12374
rect 24696 -12408 24752 -12374
rect 24786 -12408 24842 -12374
rect 24876 -12408 24932 -12374
rect 24966 -12408 25022 -12374
rect 25056 -12408 25112 -12374
rect 25146 -12408 25202 -12374
rect 25236 -12408 25292 -12374
rect 25326 -12402 25421 -12374
rect 25485 -11522 25683 -11502
rect 25485 -11556 25515 -11522
rect 25549 -11556 25616 -11522
rect 25650 -11556 25683 -11522
rect 25485 -11612 25683 -11556
rect 25485 -11646 25515 -11612
rect 25549 -11646 25616 -11612
rect 25650 -11646 25683 -11612
rect 25485 -11702 25683 -11646
rect 25485 -11736 25515 -11702
rect 25549 -11736 25616 -11702
rect 25650 -11736 25683 -11702
rect 25485 -11792 25683 -11736
rect 25485 -11826 25515 -11792
rect 25549 -11826 25616 -11792
rect 25650 -11826 25683 -11792
rect 25485 -11882 25683 -11826
rect 25485 -11916 25515 -11882
rect 25549 -11916 25616 -11882
rect 25650 -11916 25683 -11882
rect 25485 -11972 25683 -11916
rect 25485 -12006 25515 -11972
rect 25549 -12006 25616 -11972
rect 25650 -12006 25683 -11972
rect 25485 -12062 25683 -12006
rect 25485 -12096 25515 -12062
rect 25549 -12096 25616 -12062
rect 25650 -12096 25683 -12062
rect 25485 -12152 25683 -12096
rect 25485 -12186 25515 -12152
rect 25549 -12186 25616 -12152
rect 25650 -12186 25683 -12152
rect 25485 -12242 25683 -12186
rect 25485 -12276 25515 -12242
rect 25549 -12276 25616 -12242
rect 25650 -12276 25683 -12242
rect 25485 -12332 25683 -12276
rect 25485 -12366 25515 -12332
rect 25549 -12366 25616 -12332
rect 25650 -12366 25683 -12332
rect 25485 -12402 25683 -12366
rect 25747 -11518 25879 -11502
rect 25913 -11518 25969 -11484
rect 26003 -11518 26059 -11484
rect 26093 -11518 26149 -11484
rect 26183 -11518 26239 -11484
rect 26273 -11518 26329 -11484
rect 26363 -11518 26419 -11484
rect 26453 -11518 26509 -11484
rect 26543 -11518 26599 -11484
rect 26633 -11502 26884 -11484
rect 26633 -11518 26709 -11502
rect 25747 -11537 26709 -11518
rect 25747 -11562 25819 -11537
rect 25747 -11596 25766 -11562
rect 25800 -11596 25819 -11562
rect 25747 -11652 25819 -11596
rect 26637 -11596 26709 -11537
rect 25747 -11686 25766 -11652
rect 25800 -11686 25819 -11652
rect 25747 -11742 25819 -11686
rect 25747 -11776 25766 -11742
rect 25800 -11776 25819 -11742
rect 25747 -11832 25819 -11776
rect 25747 -11866 25766 -11832
rect 25800 -11866 25819 -11832
rect 25747 -11922 25819 -11866
rect 25747 -11956 25766 -11922
rect 25800 -11956 25819 -11922
rect 25747 -12012 25819 -11956
rect 25747 -12046 25766 -12012
rect 25800 -12046 25819 -12012
rect 25747 -12102 25819 -12046
rect 25747 -12136 25766 -12102
rect 25800 -12136 25819 -12102
rect 25747 -12192 25819 -12136
rect 25747 -12226 25766 -12192
rect 25800 -12226 25819 -12192
rect 25747 -12282 25819 -12226
rect 25747 -12316 25766 -12282
rect 25800 -12316 25819 -12282
rect 25881 -11660 26575 -11599
rect 25881 -11694 25942 -11660
rect 25976 -11672 26032 -11660
rect 26066 -11672 26122 -11660
rect 26156 -11672 26212 -11660
rect 25988 -11694 26032 -11672
rect 26088 -11694 26122 -11672
rect 26188 -11694 26212 -11672
rect 26246 -11672 26302 -11660
rect 26246 -11694 26254 -11672
rect 25881 -11706 25954 -11694
rect 25988 -11706 26054 -11694
rect 26088 -11706 26154 -11694
rect 26188 -11706 26254 -11694
rect 26288 -11694 26302 -11672
rect 26336 -11672 26392 -11660
rect 26336 -11694 26354 -11672
rect 26288 -11706 26354 -11694
rect 26388 -11694 26392 -11672
rect 26426 -11672 26482 -11660
rect 26426 -11694 26454 -11672
rect 26516 -11694 26575 -11660
rect 26388 -11706 26454 -11694
rect 26488 -11706 26575 -11694
rect 25881 -11750 26575 -11706
rect 25881 -11784 25942 -11750
rect 25976 -11772 26032 -11750
rect 26066 -11772 26122 -11750
rect 26156 -11772 26212 -11750
rect 25988 -11784 26032 -11772
rect 26088 -11784 26122 -11772
rect 26188 -11784 26212 -11772
rect 26246 -11772 26302 -11750
rect 26246 -11784 26254 -11772
rect 25881 -11806 25954 -11784
rect 25988 -11806 26054 -11784
rect 26088 -11806 26154 -11784
rect 26188 -11806 26254 -11784
rect 26288 -11784 26302 -11772
rect 26336 -11772 26392 -11750
rect 26336 -11784 26354 -11772
rect 26288 -11806 26354 -11784
rect 26388 -11784 26392 -11772
rect 26426 -11772 26482 -11750
rect 26426 -11784 26454 -11772
rect 26516 -11784 26575 -11750
rect 26388 -11806 26454 -11784
rect 26488 -11806 26575 -11784
rect 25881 -11840 26575 -11806
rect 25881 -11874 25942 -11840
rect 25976 -11872 26032 -11840
rect 26066 -11872 26122 -11840
rect 26156 -11872 26212 -11840
rect 25988 -11874 26032 -11872
rect 26088 -11874 26122 -11872
rect 26188 -11874 26212 -11872
rect 26246 -11872 26302 -11840
rect 26246 -11874 26254 -11872
rect 25881 -11906 25954 -11874
rect 25988 -11906 26054 -11874
rect 26088 -11906 26154 -11874
rect 26188 -11906 26254 -11874
rect 26288 -11874 26302 -11872
rect 26336 -11872 26392 -11840
rect 26336 -11874 26354 -11872
rect 26288 -11906 26354 -11874
rect 26388 -11874 26392 -11872
rect 26426 -11872 26482 -11840
rect 26426 -11874 26454 -11872
rect 26516 -11874 26575 -11840
rect 26388 -11906 26454 -11874
rect 26488 -11906 26575 -11874
rect 25881 -11930 26575 -11906
rect 25881 -11964 25942 -11930
rect 25976 -11964 26032 -11930
rect 26066 -11964 26122 -11930
rect 26156 -11964 26212 -11930
rect 26246 -11964 26302 -11930
rect 26336 -11964 26392 -11930
rect 26426 -11964 26482 -11930
rect 26516 -11964 26575 -11930
rect 25881 -11972 26575 -11964
rect 25881 -12006 25954 -11972
rect 25988 -12006 26054 -11972
rect 26088 -12006 26154 -11972
rect 26188 -12006 26254 -11972
rect 26288 -12006 26354 -11972
rect 26388 -12006 26454 -11972
rect 26488 -12006 26575 -11972
rect 25881 -12020 26575 -12006
rect 25881 -12054 25942 -12020
rect 25976 -12054 26032 -12020
rect 26066 -12054 26122 -12020
rect 26156 -12054 26212 -12020
rect 26246 -12054 26302 -12020
rect 26336 -12054 26392 -12020
rect 26426 -12054 26482 -12020
rect 26516 -12054 26575 -12020
rect 25881 -12072 26575 -12054
rect 25881 -12106 25954 -12072
rect 25988 -12106 26054 -12072
rect 26088 -12106 26154 -12072
rect 26188 -12106 26254 -12072
rect 26288 -12106 26354 -12072
rect 26388 -12106 26454 -12072
rect 26488 -12106 26575 -12072
rect 25881 -12110 26575 -12106
rect 25881 -12144 25942 -12110
rect 25976 -12144 26032 -12110
rect 26066 -12144 26122 -12110
rect 26156 -12144 26212 -12110
rect 26246 -12144 26302 -12110
rect 26336 -12144 26392 -12110
rect 26426 -12144 26482 -12110
rect 26516 -12144 26575 -12110
rect 25881 -12172 26575 -12144
rect 25881 -12200 25954 -12172
rect 25988 -12200 26054 -12172
rect 26088 -12200 26154 -12172
rect 26188 -12200 26254 -12172
rect 25881 -12234 25942 -12200
rect 25988 -12206 26032 -12200
rect 26088 -12206 26122 -12200
rect 26188 -12206 26212 -12200
rect 25976 -12234 26032 -12206
rect 26066 -12234 26122 -12206
rect 26156 -12234 26212 -12206
rect 26246 -12206 26254 -12200
rect 26288 -12200 26354 -12172
rect 26288 -12206 26302 -12200
rect 26246 -12234 26302 -12206
rect 26336 -12206 26354 -12200
rect 26388 -12200 26454 -12172
rect 26488 -12200 26575 -12172
rect 26388 -12206 26392 -12200
rect 26336 -12234 26392 -12206
rect 26426 -12206 26454 -12200
rect 26426 -12234 26482 -12206
rect 26516 -12234 26575 -12200
rect 25881 -12293 26575 -12234
rect 26637 -11630 26656 -11596
rect 26690 -11630 26709 -11596
rect 26637 -11686 26709 -11630
rect 26637 -11720 26656 -11686
rect 26690 -11720 26709 -11686
rect 26637 -11776 26709 -11720
rect 26637 -11810 26656 -11776
rect 26690 -11810 26709 -11776
rect 26637 -11866 26709 -11810
rect 26637 -11900 26656 -11866
rect 26690 -11900 26709 -11866
rect 26637 -11956 26709 -11900
rect 26637 -11990 26656 -11956
rect 26690 -11990 26709 -11956
rect 26637 -12046 26709 -11990
rect 26637 -12080 26656 -12046
rect 26690 -12080 26709 -12046
rect 26637 -12136 26709 -12080
rect 26637 -12170 26656 -12136
rect 26690 -12170 26709 -12136
rect 26637 -12226 26709 -12170
rect 26637 -12260 26656 -12226
rect 26690 -12260 26709 -12226
rect 25747 -12355 25819 -12316
rect 26637 -12316 26709 -12260
rect 26637 -12350 26656 -12316
rect 26690 -12350 26709 -12316
rect 26637 -12355 26709 -12350
rect 25747 -12374 26709 -12355
rect 25747 -12402 25860 -12374
rect 25326 -12408 25860 -12402
rect 25894 -12408 25950 -12374
rect 25984 -12408 26040 -12374
rect 26074 -12408 26130 -12374
rect 26164 -12408 26220 -12374
rect 26254 -12408 26310 -12374
rect 26344 -12408 26400 -12374
rect 26434 -12408 26490 -12374
rect 26524 -12408 26580 -12374
rect 26614 -12402 26709 -12374
rect 26773 -11522 26872 -11502
rect 26773 -11556 26803 -11522
rect 26837 -11556 26872 -11522
rect 26773 -11612 26872 -11556
rect 26773 -11646 26803 -11612
rect 26837 -11646 26872 -11612
rect 26773 -11702 26872 -11646
rect 26773 -11736 26803 -11702
rect 26837 -11736 26872 -11702
rect 26773 -11792 26872 -11736
rect 26773 -11826 26803 -11792
rect 26837 -11826 26872 -11792
rect 26773 -11882 26872 -11826
rect 26773 -11916 26803 -11882
rect 26837 -11916 26872 -11882
rect 26773 -11972 26872 -11916
rect 26773 -12006 26803 -11972
rect 26837 -12006 26872 -11972
rect 26773 -12062 26872 -12006
rect 26773 -12096 26803 -12062
rect 26837 -12096 26872 -12062
rect 26773 -12152 26872 -12096
rect 26773 -12186 26803 -12152
rect 26837 -12186 26872 -12152
rect 26773 -12242 26872 -12186
rect 26773 -12276 26803 -12242
rect 26837 -12276 26872 -12242
rect 26773 -12332 26872 -12276
rect 26773 -12366 26803 -12332
rect 26837 -12366 26872 -12332
rect 26773 -12402 26872 -12366
rect 26614 -12408 26872 -12402
rect 16568 -12422 26872 -12408
rect 16568 -12456 16600 -12422
rect 16634 -12456 17787 -12422
rect 17821 -12456 17888 -12422
rect 17922 -12456 19075 -12422
rect 19109 -12456 19176 -12422
rect 19210 -12456 20363 -12422
rect 20397 -12456 20464 -12422
rect 20498 -12456 21651 -12422
rect 21685 -12456 21752 -12422
rect 21786 -12456 22939 -12422
rect 22973 -12456 23040 -12422
rect 23074 -12456 24227 -12422
rect 24261 -12456 24328 -12422
rect 24362 -12456 25515 -12422
rect 25549 -12456 25616 -12422
rect 25650 -12456 26803 -12422
rect 26837 -12456 26872 -12422
rect 16568 -12523 26872 -12456
rect 16568 -12557 16684 -12523
rect 16718 -12557 16774 -12523
rect 16808 -12557 16864 -12523
rect 16898 -12557 16954 -12523
rect 16988 -12557 17044 -12523
rect 17078 -12557 17134 -12523
rect 17168 -12557 17224 -12523
rect 17258 -12557 17314 -12523
rect 17348 -12557 17404 -12523
rect 17438 -12557 17494 -12523
rect 17528 -12557 17584 -12523
rect 17618 -12557 17674 -12523
rect 17708 -12557 17764 -12523
rect 17798 -12557 17972 -12523
rect 18006 -12557 18062 -12523
rect 18096 -12557 18152 -12523
rect 18186 -12557 18242 -12523
rect 18276 -12557 18332 -12523
rect 18366 -12557 18422 -12523
rect 18456 -12557 18512 -12523
rect 18546 -12557 18602 -12523
rect 18636 -12557 18692 -12523
rect 18726 -12557 18782 -12523
rect 18816 -12557 18872 -12523
rect 18906 -12557 18962 -12523
rect 18996 -12557 19052 -12523
rect 19086 -12557 19260 -12523
rect 19294 -12557 19350 -12523
rect 19384 -12557 19440 -12523
rect 19474 -12557 19530 -12523
rect 19564 -12557 19620 -12523
rect 19654 -12557 19710 -12523
rect 19744 -12557 19800 -12523
rect 19834 -12557 19890 -12523
rect 19924 -12557 19980 -12523
rect 20014 -12557 20070 -12523
rect 20104 -12557 20160 -12523
rect 20194 -12557 20250 -12523
rect 20284 -12557 20340 -12523
rect 20374 -12557 20548 -12523
rect 20582 -12557 20638 -12523
rect 20672 -12557 20728 -12523
rect 20762 -12557 20818 -12523
rect 20852 -12557 20908 -12523
rect 20942 -12557 20998 -12523
rect 21032 -12557 21088 -12523
rect 21122 -12557 21178 -12523
rect 21212 -12557 21268 -12523
rect 21302 -12557 21358 -12523
rect 21392 -12557 21448 -12523
rect 21482 -12557 21538 -12523
rect 21572 -12557 21628 -12523
rect 21662 -12557 21836 -12523
rect 21870 -12557 21926 -12523
rect 21960 -12557 22016 -12523
rect 22050 -12557 22106 -12523
rect 22140 -12557 22196 -12523
rect 22230 -12557 22286 -12523
rect 22320 -12557 22376 -12523
rect 22410 -12557 22466 -12523
rect 22500 -12557 22556 -12523
rect 22590 -12557 22646 -12523
rect 22680 -12557 22736 -12523
rect 22770 -12557 22826 -12523
rect 22860 -12557 22916 -12523
rect 22950 -12557 23124 -12523
rect 23158 -12557 23214 -12523
rect 23248 -12557 23304 -12523
rect 23338 -12557 23394 -12523
rect 23428 -12557 23484 -12523
rect 23518 -12557 23574 -12523
rect 23608 -12557 23664 -12523
rect 23698 -12557 23754 -12523
rect 23788 -12557 23844 -12523
rect 23878 -12557 23934 -12523
rect 23968 -12557 24024 -12523
rect 24058 -12557 24114 -12523
rect 24148 -12557 24204 -12523
rect 24238 -12557 24412 -12523
rect 24446 -12557 24502 -12523
rect 24536 -12557 24592 -12523
rect 24626 -12557 24682 -12523
rect 24716 -12557 24772 -12523
rect 24806 -12557 24862 -12523
rect 24896 -12557 24952 -12523
rect 24986 -12557 25042 -12523
rect 25076 -12557 25132 -12523
rect 25166 -12557 25222 -12523
rect 25256 -12557 25312 -12523
rect 25346 -12557 25402 -12523
rect 25436 -12557 25492 -12523
rect 25526 -12557 25700 -12523
rect 25734 -12557 25790 -12523
rect 25824 -12557 25880 -12523
rect 25914 -12557 25970 -12523
rect 26004 -12557 26060 -12523
rect 26094 -12557 26150 -12523
rect 26184 -12557 26240 -12523
rect 26274 -12557 26330 -12523
rect 26364 -12557 26420 -12523
rect 26454 -12557 26510 -12523
rect 26544 -12557 26600 -12523
rect 26634 -12557 26690 -12523
rect 26724 -12557 26780 -12523
rect 26814 -12557 26872 -12523
rect 16568 -12624 26872 -12557
rect 16568 -12658 16684 -12624
rect 16718 -12658 16774 -12624
rect 16808 -12658 16864 -12624
rect 16898 -12658 16954 -12624
rect 16988 -12658 17044 -12624
rect 17078 -12658 17134 -12624
rect 17168 -12658 17224 -12624
rect 17258 -12658 17314 -12624
rect 17348 -12658 17404 -12624
rect 17438 -12658 17494 -12624
rect 17528 -12658 17584 -12624
rect 17618 -12658 17674 -12624
rect 17708 -12658 17764 -12624
rect 17798 -12658 17972 -12624
rect 18006 -12658 18062 -12624
rect 18096 -12658 18152 -12624
rect 18186 -12658 18242 -12624
rect 18276 -12658 18332 -12624
rect 18366 -12658 18422 -12624
rect 18456 -12658 18512 -12624
rect 18546 -12658 18602 -12624
rect 18636 -12658 18692 -12624
rect 18726 -12658 18782 -12624
rect 18816 -12658 18872 -12624
rect 18906 -12658 18962 -12624
rect 18996 -12658 19052 -12624
rect 19086 -12658 19260 -12624
rect 19294 -12658 19350 -12624
rect 19384 -12658 19440 -12624
rect 19474 -12658 19530 -12624
rect 19564 -12658 19620 -12624
rect 19654 -12658 19710 -12624
rect 19744 -12658 19800 -12624
rect 19834 -12658 19890 -12624
rect 19924 -12658 19980 -12624
rect 20014 -12658 20070 -12624
rect 20104 -12658 20160 -12624
rect 20194 -12658 20250 -12624
rect 20284 -12658 20340 -12624
rect 20374 -12658 20548 -12624
rect 20582 -12658 20638 -12624
rect 20672 -12658 20728 -12624
rect 20762 -12658 20818 -12624
rect 20852 -12658 20908 -12624
rect 20942 -12658 20998 -12624
rect 21032 -12658 21088 -12624
rect 21122 -12658 21178 -12624
rect 21212 -12658 21268 -12624
rect 21302 -12658 21358 -12624
rect 21392 -12658 21448 -12624
rect 21482 -12658 21538 -12624
rect 21572 -12658 21628 -12624
rect 21662 -12658 21836 -12624
rect 21870 -12658 21926 -12624
rect 21960 -12658 22016 -12624
rect 22050 -12658 22106 -12624
rect 22140 -12658 22196 -12624
rect 22230 -12658 22286 -12624
rect 22320 -12658 22376 -12624
rect 22410 -12658 22466 -12624
rect 22500 -12658 22556 -12624
rect 22590 -12658 22646 -12624
rect 22680 -12658 22736 -12624
rect 22770 -12658 22826 -12624
rect 22860 -12658 22916 -12624
rect 22950 -12658 23124 -12624
rect 23158 -12658 23214 -12624
rect 23248 -12658 23304 -12624
rect 23338 -12658 23394 -12624
rect 23428 -12658 23484 -12624
rect 23518 -12658 23574 -12624
rect 23608 -12658 23664 -12624
rect 23698 -12658 23754 -12624
rect 23788 -12658 23844 -12624
rect 23878 -12658 23934 -12624
rect 23968 -12658 24024 -12624
rect 24058 -12658 24114 -12624
rect 24148 -12658 24204 -12624
rect 24238 -12658 24412 -12624
rect 24446 -12658 24502 -12624
rect 24536 -12658 24592 -12624
rect 24626 -12658 24682 -12624
rect 24716 -12658 24772 -12624
rect 24806 -12658 24862 -12624
rect 24896 -12658 24952 -12624
rect 24986 -12658 25042 -12624
rect 25076 -12658 25132 -12624
rect 25166 -12658 25222 -12624
rect 25256 -12658 25312 -12624
rect 25346 -12658 25402 -12624
rect 25436 -12658 25492 -12624
rect 25526 -12658 25700 -12624
rect 25734 -12658 25790 -12624
rect 25824 -12658 25880 -12624
rect 25914 -12658 25970 -12624
rect 26004 -12658 26060 -12624
rect 26094 -12658 26150 -12624
rect 26184 -12658 26240 -12624
rect 26274 -12658 26330 -12624
rect 26364 -12658 26420 -12624
rect 26454 -12658 26510 -12624
rect 26544 -12658 26600 -12624
rect 26634 -12658 26690 -12624
rect 26724 -12658 26780 -12624
rect 26814 -12658 26872 -12624
rect 16568 -12720 26872 -12658
rect 16568 -12754 16600 -12720
rect 16634 -12754 17787 -12720
rect 17821 -12754 17888 -12720
rect 17922 -12754 19075 -12720
rect 19109 -12754 19176 -12720
rect 19210 -12754 20363 -12720
rect 20397 -12754 20464 -12720
rect 20498 -12754 21651 -12720
rect 21685 -12754 21752 -12720
rect 21786 -12754 22939 -12720
rect 22973 -12754 23040 -12720
rect 23074 -12754 24227 -12720
rect 24261 -12754 24328 -12720
rect 24362 -12754 25515 -12720
rect 25549 -12754 25616 -12720
rect 25650 -12754 26803 -12720
rect 26837 -12754 26872 -12720
rect 16568 -12772 26872 -12754
rect 16568 -12802 16863 -12772
rect 16568 -12810 16667 -12802
rect 16568 -12844 16600 -12810
rect 16634 -12844 16667 -12810
rect 16568 -12900 16667 -12844
rect 16568 -12934 16600 -12900
rect 16634 -12934 16667 -12900
rect 16568 -12990 16667 -12934
rect 16568 -13024 16600 -12990
rect 16634 -13024 16667 -12990
rect 16568 -13080 16667 -13024
rect 16568 -13114 16600 -13080
rect 16634 -13114 16667 -13080
rect 16568 -13170 16667 -13114
rect 16568 -13204 16600 -13170
rect 16634 -13204 16667 -13170
rect 16568 -13260 16667 -13204
rect 16568 -13294 16600 -13260
rect 16634 -13294 16667 -13260
rect 16568 -13350 16667 -13294
rect 16568 -13384 16600 -13350
rect 16634 -13384 16667 -13350
rect 16568 -13440 16667 -13384
rect 16568 -13474 16600 -13440
rect 16634 -13474 16667 -13440
rect 16568 -13530 16667 -13474
rect 16568 -13564 16600 -13530
rect 16634 -13564 16667 -13530
rect 16568 -13620 16667 -13564
rect 16568 -13654 16600 -13620
rect 16634 -13654 16667 -13620
rect 16568 -13702 16667 -13654
rect 16731 -12806 16863 -12802
rect 16897 -12806 16953 -12772
rect 16987 -12806 17043 -12772
rect 17077 -12806 17133 -12772
rect 17167 -12806 17223 -12772
rect 17257 -12806 17313 -12772
rect 17347 -12806 17403 -12772
rect 17437 -12806 17493 -12772
rect 17527 -12806 17583 -12772
rect 17617 -12802 18151 -12772
rect 17617 -12806 17693 -12802
rect 16731 -12825 17693 -12806
rect 16731 -12850 16803 -12825
rect 16731 -12884 16750 -12850
rect 16784 -12884 16803 -12850
rect 16731 -12940 16803 -12884
rect 17621 -12884 17693 -12825
rect 16731 -12974 16750 -12940
rect 16784 -12974 16803 -12940
rect 16731 -13030 16803 -12974
rect 16731 -13064 16750 -13030
rect 16784 -13064 16803 -13030
rect 16731 -13120 16803 -13064
rect 16731 -13154 16750 -13120
rect 16784 -13154 16803 -13120
rect 16731 -13210 16803 -13154
rect 16731 -13244 16750 -13210
rect 16784 -13244 16803 -13210
rect 16731 -13300 16803 -13244
rect 16731 -13334 16750 -13300
rect 16784 -13334 16803 -13300
rect 16731 -13390 16803 -13334
rect 16731 -13424 16750 -13390
rect 16784 -13424 16803 -13390
rect 16731 -13480 16803 -13424
rect 16731 -13514 16750 -13480
rect 16784 -13514 16803 -13480
rect 16731 -13570 16803 -13514
rect 16731 -13604 16750 -13570
rect 16784 -13604 16803 -13570
rect 16865 -12948 17559 -12887
rect 16865 -12982 16926 -12948
rect 16960 -12960 17016 -12948
rect 17050 -12960 17106 -12948
rect 17140 -12960 17196 -12948
rect 16972 -12982 17016 -12960
rect 17072 -12982 17106 -12960
rect 17172 -12982 17196 -12960
rect 17230 -12960 17286 -12948
rect 17230 -12982 17238 -12960
rect 16865 -12994 16938 -12982
rect 16972 -12994 17038 -12982
rect 17072 -12994 17138 -12982
rect 17172 -12994 17238 -12982
rect 17272 -12982 17286 -12960
rect 17320 -12960 17376 -12948
rect 17320 -12982 17338 -12960
rect 17272 -12994 17338 -12982
rect 17372 -12982 17376 -12960
rect 17410 -12960 17466 -12948
rect 17410 -12982 17438 -12960
rect 17500 -12982 17559 -12948
rect 17372 -12994 17438 -12982
rect 17472 -12994 17559 -12982
rect 16865 -13038 17559 -12994
rect 16865 -13072 16926 -13038
rect 16960 -13060 17016 -13038
rect 17050 -13060 17106 -13038
rect 17140 -13060 17196 -13038
rect 16972 -13072 17016 -13060
rect 17072 -13072 17106 -13060
rect 17172 -13072 17196 -13060
rect 17230 -13060 17286 -13038
rect 17230 -13072 17238 -13060
rect 16865 -13094 16938 -13072
rect 16972 -13094 17038 -13072
rect 17072 -13094 17138 -13072
rect 17172 -13094 17238 -13072
rect 17272 -13072 17286 -13060
rect 17320 -13060 17376 -13038
rect 17320 -13072 17338 -13060
rect 17272 -13094 17338 -13072
rect 17372 -13072 17376 -13060
rect 17410 -13060 17466 -13038
rect 17410 -13072 17438 -13060
rect 17500 -13072 17559 -13038
rect 17372 -13094 17438 -13072
rect 17472 -13094 17559 -13072
rect 16865 -13128 17559 -13094
rect 16865 -13162 16926 -13128
rect 16960 -13160 17016 -13128
rect 17050 -13160 17106 -13128
rect 17140 -13160 17196 -13128
rect 16972 -13162 17016 -13160
rect 17072 -13162 17106 -13160
rect 17172 -13162 17196 -13160
rect 17230 -13160 17286 -13128
rect 17230 -13162 17238 -13160
rect 16865 -13194 16938 -13162
rect 16972 -13194 17038 -13162
rect 17072 -13194 17138 -13162
rect 17172 -13194 17238 -13162
rect 17272 -13162 17286 -13160
rect 17320 -13160 17376 -13128
rect 17320 -13162 17338 -13160
rect 17272 -13194 17338 -13162
rect 17372 -13162 17376 -13160
rect 17410 -13160 17466 -13128
rect 17410 -13162 17438 -13160
rect 17500 -13162 17559 -13128
rect 17372 -13194 17438 -13162
rect 17472 -13194 17559 -13162
rect 16865 -13218 17559 -13194
rect 16865 -13252 16926 -13218
rect 16960 -13252 17016 -13218
rect 17050 -13252 17106 -13218
rect 17140 -13252 17196 -13218
rect 17230 -13252 17286 -13218
rect 17320 -13252 17376 -13218
rect 17410 -13252 17466 -13218
rect 17500 -13252 17559 -13218
rect 16865 -13260 17559 -13252
rect 16865 -13294 16938 -13260
rect 16972 -13294 17038 -13260
rect 17072 -13294 17138 -13260
rect 17172 -13294 17238 -13260
rect 17272 -13294 17338 -13260
rect 17372 -13294 17438 -13260
rect 17472 -13294 17559 -13260
rect 16865 -13308 17559 -13294
rect 16865 -13342 16926 -13308
rect 16960 -13342 17016 -13308
rect 17050 -13342 17106 -13308
rect 17140 -13342 17196 -13308
rect 17230 -13342 17286 -13308
rect 17320 -13342 17376 -13308
rect 17410 -13342 17466 -13308
rect 17500 -13342 17559 -13308
rect 16865 -13360 17559 -13342
rect 16865 -13394 16938 -13360
rect 16972 -13394 17038 -13360
rect 17072 -13394 17138 -13360
rect 17172 -13394 17238 -13360
rect 17272 -13394 17338 -13360
rect 17372 -13394 17438 -13360
rect 17472 -13394 17559 -13360
rect 16865 -13398 17559 -13394
rect 16865 -13432 16926 -13398
rect 16960 -13432 17016 -13398
rect 17050 -13432 17106 -13398
rect 17140 -13432 17196 -13398
rect 17230 -13432 17286 -13398
rect 17320 -13432 17376 -13398
rect 17410 -13432 17466 -13398
rect 17500 -13432 17559 -13398
rect 16865 -13460 17559 -13432
rect 16865 -13488 16938 -13460
rect 16972 -13488 17038 -13460
rect 17072 -13488 17138 -13460
rect 17172 -13488 17238 -13460
rect 16865 -13522 16926 -13488
rect 16972 -13494 17016 -13488
rect 17072 -13494 17106 -13488
rect 17172 -13494 17196 -13488
rect 16960 -13522 17016 -13494
rect 17050 -13522 17106 -13494
rect 17140 -13522 17196 -13494
rect 17230 -13494 17238 -13488
rect 17272 -13488 17338 -13460
rect 17272 -13494 17286 -13488
rect 17230 -13522 17286 -13494
rect 17320 -13494 17338 -13488
rect 17372 -13488 17438 -13460
rect 17472 -13488 17559 -13460
rect 17372 -13494 17376 -13488
rect 17320 -13522 17376 -13494
rect 17410 -13494 17438 -13488
rect 17410 -13522 17466 -13494
rect 17500 -13522 17559 -13488
rect 16865 -13581 17559 -13522
rect 17621 -12918 17640 -12884
rect 17674 -12918 17693 -12884
rect 17621 -12974 17693 -12918
rect 17621 -13008 17640 -12974
rect 17674 -13008 17693 -12974
rect 17621 -13064 17693 -13008
rect 17621 -13098 17640 -13064
rect 17674 -13098 17693 -13064
rect 17621 -13154 17693 -13098
rect 17621 -13188 17640 -13154
rect 17674 -13188 17693 -13154
rect 17621 -13244 17693 -13188
rect 17621 -13278 17640 -13244
rect 17674 -13278 17693 -13244
rect 17621 -13334 17693 -13278
rect 17621 -13368 17640 -13334
rect 17674 -13368 17693 -13334
rect 17621 -13424 17693 -13368
rect 17621 -13458 17640 -13424
rect 17674 -13458 17693 -13424
rect 17621 -13514 17693 -13458
rect 17621 -13548 17640 -13514
rect 17674 -13548 17693 -13514
rect 16731 -13643 16803 -13604
rect 17621 -13604 17693 -13548
rect 17621 -13638 17640 -13604
rect 17674 -13638 17693 -13604
rect 17621 -13643 17693 -13638
rect 16731 -13662 17693 -13643
rect 16731 -13696 16844 -13662
rect 16878 -13696 16934 -13662
rect 16968 -13696 17024 -13662
rect 17058 -13696 17114 -13662
rect 17148 -13696 17204 -13662
rect 17238 -13696 17294 -13662
rect 17328 -13696 17384 -13662
rect 17418 -13696 17474 -13662
rect 17508 -13696 17564 -13662
rect 17598 -13696 17693 -13662
rect 16731 -13702 17693 -13696
rect 17757 -12810 17955 -12802
rect 17757 -12844 17787 -12810
rect 17821 -12844 17888 -12810
rect 17922 -12844 17955 -12810
rect 17757 -12900 17955 -12844
rect 17757 -12934 17787 -12900
rect 17821 -12934 17888 -12900
rect 17922 -12934 17955 -12900
rect 17757 -12990 17955 -12934
rect 17757 -13024 17787 -12990
rect 17821 -13024 17888 -12990
rect 17922 -13024 17955 -12990
rect 17757 -13080 17955 -13024
rect 17757 -13114 17787 -13080
rect 17821 -13114 17888 -13080
rect 17922 -13114 17955 -13080
rect 17757 -13170 17955 -13114
rect 17757 -13204 17787 -13170
rect 17821 -13204 17888 -13170
rect 17922 -13204 17955 -13170
rect 17757 -13260 17955 -13204
rect 17757 -13294 17787 -13260
rect 17821 -13294 17888 -13260
rect 17922 -13294 17955 -13260
rect 17757 -13350 17955 -13294
rect 17757 -13384 17787 -13350
rect 17821 -13384 17888 -13350
rect 17922 -13384 17955 -13350
rect 17757 -13440 17955 -13384
rect 17757 -13474 17787 -13440
rect 17821 -13474 17888 -13440
rect 17922 -13474 17955 -13440
rect 17757 -13530 17955 -13474
rect 17757 -13564 17787 -13530
rect 17821 -13564 17888 -13530
rect 17922 -13564 17955 -13530
rect 17757 -13620 17955 -13564
rect 17757 -13654 17787 -13620
rect 17821 -13654 17888 -13620
rect 17922 -13654 17955 -13620
rect 17757 -13702 17955 -13654
rect 18019 -12806 18151 -12802
rect 18185 -12806 18241 -12772
rect 18275 -12806 18331 -12772
rect 18365 -12806 18421 -12772
rect 18455 -12806 18511 -12772
rect 18545 -12806 18601 -12772
rect 18635 -12806 18691 -12772
rect 18725 -12806 18781 -12772
rect 18815 -12806 18871 -12772
rect 18905 -12802 19439 -12772
rect 18905 -12806 18981 -12802
rect 18019 -12825 18981 -12806
rect 18019 -12850 18091 -12825
rect 18019 -12884 18038 -12850
rect 18072 -12884 18091 -12850
rect 18019 -12940 18091 -12884
rect 18909 -12884 18981 -12825
rect 18019 -12974 18038 -12940
rect 18072 -12974 18091 -12940
rect 18019 -13030 18091 -12974
rect 18019 -13064 18038 -13030
rect 18072 -13064 18091 -13030
rect 18019 -13120 18091 -13064
rect 18019 -13154 18038 -13120
rect 18072 -13154 18091 -13120
rect 18019 -13210 18091 -13154
rect 18019 -13244 18038 -13210
rect 18072 -13244 18091 -13210
rect 18019 -13300 18091 -13244
rect 18019 -13334 18038 -13300
rect 18072 -13334 18091 -13300
rect 18019 -13390 18091 -13334
rect 18019 -13424 18038 -13390
rect 18072 -13424 18091 -13390
rect 18019 -13480 18091 -13424
rect 18019 -13514 18038 -13480
rect 18072 -13514 18091 -13480
rect 18019 -13570 18091 -13514
rect 18019 -13604 18038 -13570
rect 18072 -13604 18091 -13570
rect 18153 -12948 18847 -12887
rect 18153 -12982 18214 -12948
rect 18248 -12960 18304 -12948
rect 18338 -12960 18394 -12948
rect 18428 -12960 18484 -12948
rect 18260 -12982 18304 -12960
rect 18360 -12982 18394 -12960
rect 18460 -12982 18484 -12960
rect 18518 -12960 18574 -12948
rect 18518 -12982 18526 -12960
rect 18153 -12994 18226 -12982
rect 18260 -12994 18326 -12982
rect 18360 -12994 18426 -12982
rect 18460 -12994 18526 -12982
rect 18560 -12982 18574 -12960
rect 18608 -12960 18664 -12948
rect 18608 -12982 18626 -12960
rect 18560 -12994 18626 -12982
rect 18660 -12982 18664 -12960
rect 18698 -12960 18754 -12948
rect 18698 -12982 18726 -12960
rect 18788 -12982 18847 -12948
rect 18660 -12994 18726 -12982
rect 18760 -12994 18847 -12982
rect 18153 -13038 18847 -12994
rect 18153 -13072 18214 -13038
rect 18248 -13060 18304 -13038
rect 18338 -13060 18394 -13038
rect 18428 -13060 18484 -13038
rect 18260 -13072 18304 -13060
rect 18360 -13072 18394 -13060
rect 18460 -13072 18484 -13060
rect 18518 -13060 18574 -13038
rect 18518 -13072 18526 -13060
rect 18153 -13094 18226 -13072
rect 18260 -13094 18326 -13072
rect 18360 -13094 18426 -13072
rect 18460 -13094 18526 -13072
rect 18560 -13072 18574 -13060
rect 18608 -13060 18664 -13038
rect 18608 -13072 18626 -13060
rect 18560 -13094 18626 -13072
rect 18660 -13072 18664 -13060
rect 18698 -13060 18754 -13038
rect 18698 -13072 18726 -13060
rect 18788 -13072 18847 -13038
rect 18660 -13094 18726 -13072
rect 18760 -13094 18847 -13072
rect 18153 -13128 18847 -13094
rect 18153 -13162 18214 -13128
rect 18248 -13160 18304 -13128
rect 18338 -13160 18394 -13128
rect 18428 -13160 18484 -13128
rect 18260 -13162 18304 -13160
rect 18360 -13162 18394 -13160
rect 18460 -13162 18484 -13160
rect 18518 -13160 18574 -13128
rect 18518 -13162 18526 -13160
rect 18153 -13194 18226 -13162
rect 18260 -13194 18326 -13162
rect 18360 -13194 18426 -13162
rect 18460 -13194 18526 -13162
rect 18560 -13162 18574 -13160
rect 18608 -13160 18664 -13128
rect 18608 -13162 18626 -13160
rect 18560 -13194 18626 -13162
rect 18660 -13162 18664 -13160
rect 18698 -13160 18754 -13128
rect 18698 -13162 18726 -13160
rect 18788 -13162 18847 -13128
rect 18660 -13194 18726 -13162
rect 18760 -13194 18847 -13162
rect 18153 -13218 18847 -13194
rect 18153 -13252 18214 -13218
rect 18248 -13252 18304 -13218
rect 18338 -13252 18394 -13218
rect 18428 -13252 18484 -13218
rect 18518 -13252 18574 -13218
rect 18608 -13252 18664 -13218
rect 18698 -13252 18754 -13218
rect 18788 -13252 18847 -13218
rect 18153 -13260 18847 -13252
rect 18153 -13294 18226 -13260
rect 18260 -13294 18326 -13260
rect 18360 -13294 18426 -13260
rect 18460 -13294 18526 -13260
rect 18560 -13294 18626 -13260
rect 18660 -13294 18726 -13260
rect 18760 -13294 18847 -13260
rect 18153 -13308 18847 -13294
rect 18153 -13342 18214 -13308
rect 18248 -13342 18304 -13308
rect 18338 -13342 18394 -13308
rect 18428 -13342 18484 -13308
rect 18518 -13342 18574 -13308
rect 18608 -13342 18664 -13308
rect 18698 -13342 18754 -13308
rect 18788 -13342 18847 -13308
rect 18153 -13360 18847 -13342
rect 18153 -13394 18226 -13360
rect 18260 -13394 18326 -13360
rect 18360 -13394 18426 -13360
rect 18460 -13394 18526 -13360
rect 18560 -13394 18626 -13360
rect 18660 -13394 18726 -13360
rect 18760 -13394 18847 -13360
rect 18153 -13398 18847 -13394
rect 18153 -13432 18214 -13398
rect 18248 -13432 18304 -13398
rect 18338 -13432 18394 -13398
rect 18428 -13432 18484 -13398
rect 18518 -13432 18574 -13398
rect 18608 -13432 18664 -13398
rect 18698 -13432 18754 -13398
rect 18788 -13432 18847 -13398
rect 18153 -13460 18847 -13432
rect 18153 -13488 18226 -13460
rect 18260 -13488 18326 -13460
rect 18360 -13488 18426 -13460
rect 18460 -13488 18526 -13460
rect 18153 -13522 18214 -13488
rect 18260 -13494 18304 -13488
rect 18360 -13494 18394 -13488
rect 18460 -13494 18484 -13488
rect 18248 -13522 18304 -13494
rect 18338 -13522 18394 -13494
rect 18428 -13522 18484 -13494
rect 18518 -13494 18526 -13488
rect 18560 -13488 18626 -13460
rect 18560 -13494 18574 -13488
rect 18518 -13522 18574 -13494
rect 18608 -13494 18626 -13488
rect 18660 -13488 18726 -13460
rect 18760 -13488 18847 -13460
rect 18660 -13494 18664 -13488
rect 18608 -13522 18664 -13494
rect 18698 -13494 18726 -13488
rect 18698 -13522 18754 -13494
rect 18788 -13522 18847 -13488
rect 18153 -13581 18847 -13522
rect 18909 -12918 18928 -12884
rect 18962 -12918 18981 -12884
rect 18909 -12974 18981 -12918
rect 18909 -13008 18928 -12974
rect 18962 -13008 18981 -12974
rect 18909 -13064 18981 -13008
rect 18909 -13098 18928 -13064
rect 18962 -13098 18981 -13064
rect 18909 -13154 18981 -13098
rect 18909 -13188 18928 -13154
rect 18962 -13188 18981 -13154
rect 18909 -13244 18981 -13188
rect 18909 -13278 18928 -13244
rect 18962 -13278 18981 -13244
rect 18909 -13334 18981 -13278
rect 18909 -13368 18928 -13334
rect 18962 -13368 18981 -13334
rect 18909 -13424 18981 -13368
rect 18909 -13458 18928 -13424
rect 18962 -13458 18981 -13424
rect 18909 -13514 18981 -13458
rect 18909 -13548 18928 -13514
rect 18962 -13548 18981 -13514
rect 18019 -13643 18091 -13604
rect 18909 -13604 18981 -13548
rect 18909 -13638 18928 -13604
rect 18962 -13638 18981 -13604
rect 18909 -13643 18981 -13638
rect 18019 -13662 18981 -13643
rect 18019 -13696 18132 -13662
rect 18166 -13696 18222 -13662
rect 18256 -13696 18312 -13662
rect 18346 -13696 18402 -13662
rect 18436 -13696 18492 -13662
rect 18526 -13696 18582 -13662
rect 18616 -13696 18672 -13662
rect 18706 -13696 18762 -13662
rect 18796 -13696 18852 -13662
rect 18886 -13696 18981 -13662
rect 18019 -13702 18981 -13696
rect 19045 -12810 19243 -12802
rect 19045 -12844 19075 -12810
rect 19109 -12844 19176 -12810
rect 19210 -12844 19243 -12810
rect 19045 -12900 19243 -12844
rect 19045 -12934 19075 -12900
rect 19109 -12934 19176 -12900
rect 19210 -12934 19243 -12900
rect 19045 -12990 19243 -12934
rect 19045 -13024 19075 -12990
rect 19109 -13024 19176 -12990
rect 19210 -13024 19243 -12990
rect 19045 -13080 19243 -13024
rect 19045 -13114 19075 -13080
rect 19109 -13114 19176 -13080
rect 19210 -13114 19243 -13080
rect 19045 -13170 19243 -13114
rect 19045 -13204 19075 -13170
rect 19109 -13204 19176 -13170
rect 19210 -13204 19243 -13170
rect 19045 -13260 19243 -13204
rect 19045 -13294 19075 -13260
rect 19109 -13294 19176 -13260
rect 19210 -13294 19243 -13260
rect 19045 -13350 19243 -13294
rect 19045 -13384 19075 -13350
rect 19109 -13384 19176 -13350
rect 19210 -13384 19243 -13350
rect 19045 -13440 19243 -13384
rect 19045 -13474 19075 -13440
rect 19109 -13474 19176 -13440
rect 19210 -13474 19243 -13440
rect 19045 -13530 19243 -13474
rect 19045 -13564 19075 -13530
rect 19109 -13564 19176 -13530
rect 19210 -13564 19243 -13530
rect 19045 -13620 19243 -13564
rect 19045 -13654 19075 -13620
rect 19109 -13654 19176 -13620
rect 19210 -13654 19243 -13620
rect 19045 -13702 19243 -13654
rect 19307 -12806 19439 -12802
rect 19473 -12806 19529 -12772
rect 19563 -12806 19619 -12772
rect 19653 -12806 19709 -12772
rect 19743 -12806 19799 -12772
rect 19833 -12806 19889 -12772
rect 19923 -12806 19979 -12772
rect 20013 -12806 20069 -12772
rect 20103 -12806 20159 -12772
rect 20193 -12802 20727 -12772
rect 20193 -12806 20269 -12802
rect 19307 -12825 20269 -12806
rect 19307 -12850 19379 -12825
rect 19307 -12884 19326 -12850
rect 19360 -12884 19379 -12850
rect 19307 -12940 19379 -12884
rect 20197 -12884 20269 -12825
rect 19307 -12974 19326 -12940
rect 19360 -12974 19379 -12940
rect 19307 -13030 19379 -12974
rect 19307 -13064 19326 -13030
rect 19360 -13064 19379 -13030
rect 19307 -13120 19379 -13064
rect 19307 -13154 19326 -13120
rect 19360 -13154 19379 -13120
rect 19307 -13210 19379 -13154
rect 19307 -13244 19326 -13210
rect 19360 -13244 19379 -13210
rect 19307 -13300 19379 -13244
rect 19307 -13334 19326 -13300
rect 19360 -13334 19379 -13300
rect 19307 -13390 19379 -13334
rect 19307 -13424 19326 -13390
rect 19360 -13424 19379 -13390
rect 19307 -13480 19379 -13424
rect 19307 -13514 19326 -13480
rect 19360 -13514 19379 -13480
rect 19307 -13570 19379 -13514
rect 19307 -13604 19326 -13570
rect 19360 -13604 19379 -13570
rect 19441 -12948 20135 -12887
rect 19441 -12982 19502 -12948
rect 19536 -12960 19592 -12948
rect 19626 -12960 19682 -12948
rect 19716 -12960 19772 -12948
rect 19548 -12982 19592 -12960
rect 19648 -12982 19682 -12960
rect 19748 -12982 19772 -12960
rect 19806 -12960 19862 -12948
rect 19806 -12982 19814 -12960
rect 19441 -12994 19514 -12982
rect 19548 -12994 19614 -12982
rect 19648 -12994 19714 -12982
rect 19748 -12994 19814 -12982
rect 19848 -12982 19862 -12960
rect 19896 -12960 19952 -12948
rect 19896 -12982 19914 -12960
rect 19848 -12994 19914 -12982
rect 19948 -12982 19952 -12960
rect 19986 -12960 20042 -12948
rect 19986 -12982 20014 -12960
rect 20076 -12982 20135 -12948
rect 19948 -12994 20014 -12982
rect 20048 -12994 20135 -12982
rect 19441 -13038 20135 -12994
rect 19441 -13072 19502 -13038
rect 19536 -13060 19592 -13038
rect 19626 -13060 19682 -13038
rect 19716 -13060 19772 -13038
rect 19548 -13072 19592 -13060
rect 19648 -13072 19682 -13060
rect 19748 -13072 19772 -13060
rect 19806 -13060 19862 -13038
rect 19806 -13072 19814 -13060
rect 19441 -13094 19514 -13072
rect 19548 -13094 19614 -13072
rect 19648 -13094 19714 -13072
rect 19748 -13094 19814 -13072
rect 19848 -13072 19862 -13060
rect 19896 -13060 19952 -13038
rect 19896 -13072 19914 -13060
rect 19848 -13094 19914 -13072
rect 19948 -13072 19952 -13060
rect 19986 -13060 20042 -13038
rect 19986 -13072 20014 -13060
rect 20076 -13072 20135 -13038
rect 19948 -13094 20014 -13072
rect 20048 -13094 20135 -13072
rect 19441 -13128 20135 -13094
rect 19441 -13162 19502 -13128
rect 19536 -13160 19592 -13128
rect 19626 -13160 19682 -13128
rect 19716 -13160 19772 -13128
rect 19548 -13162 19592 -13160
rect 19648 -13162 19682 -13160
rect 19748 -13162 19772 -13160
rect 19806 -13160 19862 -13128
rect 19806 -13162 19814 -13160
rect 19441 -13194 19514 -13162
rect 19548 -13194 19614 -13162
rect 19648 -13194 19714 -13162
rect 19748 -13194 19814 -13162
rect 19848 -13162 19862 -13160
rect 19896 -13160 19952 -13128
rect 19896 -13162 19914 -13160
rect 19848 -13194 19914 -13162
rect 19948 -13162 19952 -13160
rect 19986 -13160 20042 -13128
rect 19986 -13162 20014 -13160
rect 20076 -13162 20135 -13128
rect 19948 -13194 20014 -13162
rect 20048 -13194 20135 -13162
rect 19441 -13218 20135 -13194
rect 19441 -13252 19502 -13218
rect 19536 -13252 19592 -13218
rect 19626 -13252 19682 -13218
rect 19716 -13252 19772 -13218
rect 19806 -13252 19862 -13218
rect 19896 -13252 19952 -13218
rect 19986 -13252 20042 -13218
rect 20076 -13252 20135 -13218
rect 19441 -13260 20135 -13252
rect 19441 -13294 19514 -13260
rect 19548 -13294 19614 -13260
rect 19648 -13294 19714 -13260
rect 19748 -13294 19814 -13260
rect 19848 -13294 19914 -13260
rect 19948 -13294 20014 -13260
rect 20048 -13294 20135 -13260
rect 19441 -13308 20135 -13294
rect 19441 -13342 19502 -13308
rect 19536 -13342 19592 -13308
rect 19626 -13342 19682 -13308
rect 19716 -13342 19772 -13308
rect 19806 -13342 19862 -13308
rect 19896 -13342 19952 -13308
rect 19986 -13342 20042 -13308
rect 20076 -13342 20135 -13308
rect 19441 -13360 20135 -13342
rect 19441 -13394 19514 -13360
rect 19548 -13394 19614 -13360
rect 19648 -13394 19714 -13360
rect 19748 -13394 19814 -13360
rect 19848 -13394 19914 -13360
rect 19948 -13394 20014 -13360
rect 20048 -13394 20135 -13360
rect 19441 -13398 20135 -13394
rect 19441 -13432 19502 -13398
rect 19536 -13432 19592 -13398
rect 19626 -13432 19682 -13398
rect 19716 -13432 19772 -13398
rect 19806 -13432 19862 -13398
rect 19896 -13432 19952 -13398
rect 19986 -13432 20042 -13398
rect 20076 -13432 20135 -13398
rect 19441 -13460 20135 -13432
rect 19441 -13488 19514 -13460
rect 19548 -13488 19614 -13460
rect 19648 -13488 19714 -13460
rect 19748 -13488 19814 -13460
rect 19441 -13522 19502 -13488
rect 19548 -13494 19592 -13488
rect 19648 -13494 19682 -13488
rect 19748 -13494 19772 -13488
rect 19536 -13522 19592 -13494
rect 19626 -13522 19682 -13494
rect 19716 -13522 19772 -13494
rect 19806 -13494 19814 -13488
rect 19848 -13488 19914 -13460
rect 19848 -13494 19862 -13488
rect 19806 -13522 19862 -13494
rect 19896 -13494 19914 -13488
rect 19948 -13488 20014 -13460
rect 20048 -13488 20135 -13460
rect 19948 -13494 19952 -13488
rect 19896 -13522 19952 -13494
rect 19986 -13494 20014 -13488
rect 19986 -13522 20042 -13494
rect 20076 -13522 20135 -13488
rect 19441 -13581 20135 -13522
rect 20197 -12918 20216 -12884
rect 20250 -12918 20269 -12884
rect 20197 -12974 20269 -12918
rect 20197 -13008 20216 -12974
rect 20250 -13008 20269 -12974
rect 20197 -13064 20269 -13008
rect 20197 -13098 20216 -13064
rect 20250 -13098 20269 -13064
rect 20197 -13154 20269 -13098
rect 20197 -13188 20216 -13154
rect 20250 -13188 20269 -13154
rect 20197 -13244 20269 -13188
rect 20197 -13278 20216 -13244
rect 20250 -13278 20269 -13244
rect 20197 -13334 20269 -13278
rect 20197 -13368 20216 -13334
rect 20250 -13368 20269 -13334
rect 20197 -13424 20269 -13368
rect 20197 -13458 20216 -13424
rect 20250 -13458 20269 -13424
rect 20197 -13514 20269 -13458
rect 20197 -13548 20216 -13514
rect 20250 -13548 20269 -13514
rect 19307 -13643 19379 -13604
rect 20197 -13604 20269 -13548
rect 20197 -13638 20216 -13604
rect 20250 -13638 20269 -13604
rect 20197 -13643 20269 -13638
rect 19307 -13662 20269 -13643
rect 19307 -13696 19420 -13662
rect 19454 -13696 19510 -13662
rect 19544 -13696 19600 -13662
rect 19634 -13696 19690 -13662
rect 19724 -13696 19780 -13662
rect 19814 -13696 19870 -13662
rect 19904 -13696 19960 -13662
rect 19994 -13696 20050 -13662
rect 20084 -13696 20140 -13662
rect 20174 -13696 20269 -13662
rect 19307 -13702 20269 -13696
rect 20333 -12810 20531 -12802
rect 20333 -12844 20363 -12810
rect 20397 -12844 20464 -12810
rect 20498 -12844 20531 -12810
rect 20333 -12900 20531 -12844
rect 20333 -12934 20363 -12900
rect 20397 -12934 20464 -12900
rect 20498 -12934 20531 -12900
rect 20333 -12990 20531 -12934
rect 20333 -13024 20363 -12990
rect 20397 -13024 20464 -12990
rect 20498 -13024 20531 -12990
rect 20333 -13080 20531 -13024
rect 20333 -13114 20363 -13080
rect 20397 -13114 20464 -13080
rect 20498 -13114 20531 -13080
rect 20333 -13170 20531 -13114
rect 20333 -13204 20363 -13170
rect 20397 -13204 20464 -13170
rect 20498 -13204 20531 -13170
rect 20333 -13260 20531 -13204
rect 20333 -13294 20363 -13260
rect 20397 -13294 20464 -13260
rect 20498 -13294 20531 -13260
rect 20333 -13350 20531 -13294
rect 20333 -13384 20363 -13350
rect 20397 -13384 20464 -13350
rect 20498 -13384 20531 -13350
rect 20333 -13440 20531 -13384
rect 20333 -13474 20363 -13440
rect 20397 -13474 20464 -13440
rect 20498 -13474 20531 -13440
rect 20333 -13530 20531 -13474
rect 20333 -13564 20363 -13530
rect 20397 -13564 20464 -13530
rect 20498 -13564 20531 -13530
rect 20333 -13620 20531 -13564
rect 20333 -13654 20363 -13620
rect 20397 -13654 20464 -13620
rect 20498 -13654 20531 -13620
rect 20333 -13702 20531 -13654
rect 20595 -12806 20727 -12802
rect 20761 -12806 20817 -12772
rect 20851 -12806 20907 -12772
rect 20941 -12806 20997 -12772
rect 21031 -12806 21087 -12772
rect 21121 -12806 21177 -12772
rect 21211 -12806 21267 -12772
rect 21301 -12806 21357 -12772
rect 21391 -12806 21447 -12772
rect 21481 -12802 22015 -12772
rect 21481 -12806 21557 -12802
rect 20595 -12825 21557 -12806
rect 20595 -12850 20667 -12825
rect 20595 -12884 20614 -12850
rect 20648 -12884 20667 -12850
rect 20595 -12940 20667 -12884
rect 21485 -12884 21557 -12825
rect 20595 -12974 20614 -12940
rect 20648 -12974 20667 -12940
rect 20595 -13030 20667 -12974
rect 20595 -13064 20614 -13030
rect 20648 -13064 20667 -13030
rect 20595 -13120 20667 -13064
rect 20595 -13154 20614 -13120
rect 20648 -13154 20667 -13120
rect 20595 -13210 20667 -13154
rect 20595 -13244 20614 -13210
rect 20648 -13244 20667 -13210
rect 20595 -13300 20667 -13244
rect 20595 -13334 20614 -13300
rect 20648 -13334 20667 -13300
rect 20595 -13390 20667 -13334
rect 20595 -13424 20614 -13390
rect 20648 -13424 20667 -13390
rect 20595 -13480 20667 -13424
rect 20595 -13514 20614 -13480
rect 20648 -13514 20667 -13480
rect 20595 -13570 20667 -13514
rect 20595 -13604 20614 -13570
rect 20648 -13604 20667 -13570
rect 20729 -12948 21423 -12887
rect 20729 -12982 20790 -12948
rect 20824 -12960 20880 -12948
rect 20914 -12960 20970 -12948
rect 21004 -12960 21060 -12948
rect 20836 -12982 20880 -12960
rect 20936 -12982 20970 -12960
rect 21036 -12982 21060 -12960
rect 21094 -12960 21150 -12948
rect 21094 -12982 21102 -12960
rect 20729 -12994 20802 -12982
rect 20836 -12994 20902 -12982
rect 20936 -12994 21002 -12982
rect 21036 -12994 21102 -12982
rect 21136 -12982 21150 -12960
rect 21184 -12960 21240 -12948
rect 21184 -12982 21202 -12960
rect 21136 -12994 21202 -12982
rect 21236 -12982 21240 -12960
rect 21274 -12960 21330 -12948
rect 21274 -12982 21302 -12960
rect 21364 -12982 21423 -12948
rect 21236 -12994 21302 -12982
rect 21336 -12994 21423 -12982
rect 20729 -13038 21423 -12994
rect 20729 -13072 20790 -13038
rect 20824 -13060 20880 -13038
rect 20914 -13060 20970 -13038
rect 21004 -13060 21060 -13038
rect 20836 -13072 20880 -13060
rect 20936 -13072 20970 -13060
rect 21036 -13072 21060 -13060
rect 21094 -13060 21150 -13038
rect 21094 -13072 21102 -13060
rect 20729 -13094 20802 -13072
rect 20836 -13094 20902 -13072
rect 20936 -13094 21002 -13072
rect 21036 -13094 21102 -13072
rect 21136 -13072 21150 -13060
rect 21184 -13060 21240 -13038
rect 21184 -13072 21202 -13060
rect 21136 -13094 21202 -13072
rect 21236 -13072 21240 -13060
rect 21274 -13060 21330 -13038
rect 21274 -13072 21302 -13060
rect 21364 -13072 21423 -13038
rect 21236 -13094 21302 -13072
rect 21336 -13094 21423 -13072
rect 20729 -13128 21423 -13094
rect 20729 -13162 20790 -13128
rect 20824 -13160 20880 -13128
rect 20914 -13160 20970 -13128
rect 21004 -13160 21060 -13128
rect 20836 -13162 20880 -13160
rect 20936 -13162 20970 -13160
rect 21036 -13162 21060 -13160
rect 21094 -13160 21150 -13128
rect 21094 -13162 21102 -13160
rect 20729 -13194 20802 -13162
rect 20836 -13194 20902 -13162
rect 20936 -13194 21002 -13162
rect 21036 -13194 21102 -13162
rect 21136 -13162 21150 -13160
rect 21184 -13160 21240 -13128
rect 21184 -13162 21202 -13160
rect 21136 -13194 21202 -13162
rect 21236 -13162 21240 -13160
rect 21274 -13160 21330 -13128
rect 21274 -13162 21302 -13160
rect 21364 -13162 21423 -13128
rect 21236 -13194 21302 -13162
rect 21336 -13194 21423 -13162
rect 20729 -13218 21423 -13194
rect 20729 -13252 20790 -13218
rect 20824 -13252 20880 -13218
rect 20914 -13252 20970 -13218
rect 21004 -13252 21060 -13218
rect 21094 -13252 21150 -13218
rect 21184 -13252 21240 -13218
rect 21274 -13252 21330 -13218
rect 21364 -13252 21423 -13218
rect 20729 -13260 21423 -13252
rect 20729 -13294 20802 -13260
rect 20836 -13294 20902 -13260
rect 20936 -13294 21002 -13260
rect 21036 -13294 21102 -13260
rect 21136 -13294 21202 -13260
rect 21236 -13294 21302 -13260
rect 21336 -13294 21423 -13260
rect 20729 -13308 21423 -13294
rect 20729 -13342 20790 -13308
rect 20824 -13342 20880 -13308
rect 20914 -13342 20970 -13308
rect 21004 -13342 21060 -13308
rect 21094 -13342 21150 -13308
rect 21184 -13342 21240 -13308
rect 21274 -13342 21330 -13308
rect 21364 -13342 21423 -13308
rect 20729 -13360 21423 -13342
rect 20729 -13394 20802 -13360
rect 20836 -13394 20902 -13360
rect 20936 -13394 21002 -13360
rect 21036 -13394 21102 -13360
rect 21136 -13394 21202 -13360
rect 21236 -13394 21302 -13360
rect 21336 -13394 21423 -13360
rect 20729 -13398 21423 -13394
rect 20729 -13432 20790 -13398
rect 20824 -13432 20880 -13398
rect 20914 -13432 20970 -13398
rect 21004 -13432 21060 -13398
rect 21094 -13432 21150 -13398
rect 21184 -13432 21240 -13398
rect 21274 -13432 21330 -13398
rect 21364 -13432 21423 -13398
rect 20729 -13460 21423 -13432
rect 20729 -13488 20802 -13460
rect 20836 -13488 20902 -13460
rect 20936 -13488 21002 -13460
rect 21036 -13488 21102 -13460
rect 20729 -13522 20790 -13488
rect 20836 -13494 20880 -13488
rect 20936 -13494 20970 -13488
rect 21036 -13494 21060 -13488
rect 20824 -13522 20880 -13494
rect 20914 -13522 20970 -13494
rect 21004 -13522 21060 -13494
rect 21094 -13494 21102 -13488
rect 21136 -13488 21202 -13460
rect 21136 -13494 21150 -13488
rect 21094 -13522 21150 -13494
rect 21184 -13494 21202 -13488
rect 21236 -13488 21302 -13460
rect 21336 -13488 21423 -13460
rect 21236 -13494 21240 -13488
rect 21184 -13522 21240 -13494
rect 21274 -13494 21302 -13488
rect 21274 -13522 21330 -13494
rect 21364 -13522 21423 -13488
rect 20729 -13581 21423 -13522
rect 21485 -12918 21504 -12884
rect 21538 -12918 21557 -12884
rect 21485 -12974 21557 -12918
rect 21485 -13008 21504 -12974
rect 21538 -13008 21557 -12974
rect 21485 -13064 21557 -13008
rect 21485 -13098 21504 -13064
rect 21538 -13098 21557 -13064
rect 21485 -13154 21557 -13098
rect 21485 -13188 21504 -13154
rect 21538 -13188 21557 -13154
rect 21485 -13244 21557 -13188
rect 21485 -13278 21504 -13244
rect 21538 -13278 21557 -13244
rect 21485 -13334 21557 -13278
rect 21485 -13368 21504 -13334
rect 21538 -13368 21557 -13334
rect 21485 -13424 21557 -13368
rect 21485 -13458 21504 -13424
rect 21538 -13458 21557 -13424
rect 21485 -13514 21557 -13458
rect 21485 -13548 21504 -13514
rect 21538 -13548 21557 -13514
rect 20595 -13643 20667 -13604
rect 21485 -13604 21557 -13548
rect 21485 -13638 21504 -13604
rect 21538 -13638 21557 -13604
rect 21485 -13643 21557 -13638
rect 20595 -13662 21557 -13643
rect 20595 -13696 20708 -13662
rect 20742 -13696 20798 -13662
rect 20832 -13696 20888 -13662
rect 20922 -13696 20978 -13662
rect 21012 -13696 21068 -13662
rect 21102 -13696 21158 -13662
rect 21192 -13696 21248 -13662
rect 21282 -13696 21338 -13662
rect 21372 -13696 21428 -13662
rect 21462 -13696 21557 -13662
rect 20595 -13702 21557 -13696
rect 21621 -12810 21819 -12802
rect 21621 -12844 21651 -12810
rect 21685 -12844 21752 -12810
rect 21786 -12844 21819 -12810
rect 21621 -12900 21819 -12844
rect 21621 -12934 21651 -12900
rect 21685 -12934 21752 -12900
rect 21786 -12934 21819 -12900
rect 21621 -12990 21819 -12934
rect 21621 -13024 21651 -12990
rect 21685 -13024 21752 -12990
rect 21786 -13024 21819 -12990
rect 21621 -13080 21819 -13024
rect 21621 -13114 21651 -13080
rect 21685 -13114 21752 -13080
rect 21786 -13114 21819 -13080
rect 21621 -13170 21819 -13114
rect 21621 -13204 21651 -13170
rect 21685 -13204 21752 -13170
rect 21786 -13204 21819 -13170
rect 21621 -13260 21819 -13204
rect 21621 -13294 21651 -13260
rect 21685 -13294 21752 -13260
rect 21786 -13294 21819 -13260
rect 21621 -13350 21819 -13294
rect 21621 -13384 21651 -13350
rect 21685 -13384 21752 -13350
rect 21786 -13384 21819 -13350
rect 21621 -13440 21819 -13384
rect 21621 -13474 21651 -13440
rect 21685 -13474 21752 -13440
rect 21786 -13474 21819 -13440
rect 21621 -13530 21819 -13474
rect 21621 -13564 21651 -13530
rect 21685 -13564 21752 -13530
rect 21786 -13564 21819 -13530
rect 21621 -13620 21819 -13564
rect 21621 -13654 21651 -13620
rect 21685 -13654 21752 -13620
rect 21786 -13654 21819 -13620
rect 21621 -13702 21819 -13654
rect 21883 -12806 22015 -12802
rect 22049 -12806 22105 -12772
rect 22139 -12806 22195 -12772
rect 22229 -12806 22285 -12772
rect 22319 -12806 22375 -12772
rect 22409 -12806 22465 -12772
rect 22499 -12806 22555 -12772
rect 22589 -12806 22645 -12772
rect 22679 -12806 22735 -12772
rect 22769 -12802 23303 -12772
rect 22769 -12806 22845 -12802
rect 21883 -12825 22845 -12806
rect 21883 -12850 21955 -12825
rect 21883 -12884 21902 -12850
rect 21936 -12884 21955 -12850
rect 21883 -12940 21955 -12884
rect 22773 -12884 22845 -12825
rect 21883 -12974 21902 -12940
rect 21936 -12974 21955 -12940
rect 21883 -13030 21955 -12974
rect 21883 -13064 21902 -13030
rect 21936 -13064 21955 -13030
rect 21883 -13120 21955 -13064
rect 21883 -13154 21902 -13120
rect 21936 -13154 21955 -13120
rect 21883 -13210 21955 -13154
rect 21883 -13244 21902 -13210
rect 21936 -13244 21955 -13210
rect 21883 -13300 21955 -13244
rect 21883 -13334 21902 -13300
rect 21936 -13334 21955 -13300
rect 21883 -13390 21955 -13334
rect 21883 -13424 21902 -13390
rect 21936 -13424 21955 -13390
rect 21883 -13480 21955 -13424
rect 21883 -13514 21902 -13480
rect 21936 -13514 21955 -13480
rect 21883 -13570 21955 -13514
rect 21883 -13604 21902 -13570
rect 21936 -13604 21955 -13570
rect 22017 -12948 22711 -12887
rect 22017 -12982 22078 -12948
rect 22112 -12960 22168 -12948
rect 22202 -12960 22258 -12948
rect 22292 -12960 22348 -12948
rect 22124 -12982 22168 -12960
rect 22224 -12982 22258 -12960
rect 22324 -12982 22348 -12960
rect 22382 -12960 22438 -12948
rect 22382 -12982 22390 -12960
rect 22017 -12994 22090 -12982
rect 22124 -12994 22190 -12982
rect 22224 -12994 22290 -12982
rect 22324 -12994 22390 -12982
rect 22424 -12982 22438 -12960
rect 22472 -12960 22528 -12948
rect 22472 -12982 22490 -12960
rect 22424 -12994 22490 -12982
rect 22524 -12982 22528 -12960
rect 22562 -12960 22618 -12948
rect 22562 -12982 22590 -12960
rect 22652 -12982 22711 -12948
rect 22524 -12994 22590 -12982
rect 22624 -12994 22711 -12982
rect 22017 -13038 22711 -12994
rect 22017 -13072 22078 -13038
rect 22112 -13060 22168 -13038
rect 22202 -13060 22258 -13038
rect 22292 -13060 22348 -13038
rect 22124 -13072 22168 -13060
rect 22224 -13072 22258 -13060
rect 22324 -13072 22348 -13060
rect 22382 -13060 22438 -13038
rect 22382 -13072 22390 -13060
rect 22017 -13094 22090 -13072
rect 22124 -13094 22190 -13072
rect 22224 -13094 22290 -13072
rect 22324 -13094 22390 -13072
rect 22424 -13072 22438 -13060
rect 22472 -13060 22528 -13038
rect 22472 -13072 22490 -13060
rect 22424 -13094 22490 -13072
rect 22524 -13072 22528 -13060
rect 22562 -13060 22618 -13038
rect 22562 -13072 22590 -13060
rect 22652 -13072 22711 -13038
rect 22524 -13094 22590 -13072
rect 22624 -13094 22711 -13072
rect 22017 -13128 22711 -13094
rect 22017 -13162 22078 -13128
rect 22112 -13160 22168 -13128
rect 22202 -13160 22258 -13128
rect 22292 -13160 22348 -13128
rect 22124 -13162 22168 -13160
rect 22224 -13162 22258 -13160
rect 22324 -13162 22348 -13160
rect 22382 -13160 22438 -13128
rect 22382 -13162 22390 -13160
rect 22017 -13194 22090 -13162
rect 22124 -13194 22190 -13162
rect 22224 -13194 22290 -13162
rect 22324 -13194 22390 -13162
rect 22424 -13162 22438 -13160
rect 22472 -13160 22528 -13128
rect 22472 -13162 22490 -13160
rect 22424 -13194 22490 -13162
rect 22524 -13162 22528 -13160
rect 22562 -13160 22618 -13128
rect 22562 -13162 22590 -13160
rect 22652 -13162 22711 -13128
rect 22524 -13194 22590 -13162
rect 22624 -13194 22711 -13162
rect 22017 -13218 22711 -13194
rect 22017 -13252 22078 -13218
rect 22112 -13252 22168 -13218
rect 22202 -13252 22258 -13218
rect 22292 -13252 22348 -13218
rect 22382 -13252 22438 -13218
rect 22472 -13252 22528 -13218
rect 22562 -13252 22618 -13218
rect 22652 -13252 22711 -13218
rect 22017 -13260 22711 -13252
rect 22017 -13294 22090 -13260
rect 22124 -13294 22190 -13260
rect 22224 -13294 22290 -13260
rect 22324 -13294 22390 -13260
rect 22424 -13294 22490 -13260
rect 22524 -13294 22590 -13260
rect 22624 -13294 22711 -13260
rect 22017 -13308 22711 -13294
rect 22017 -13342 22078 -13308
rect 22112 -13342 22168 -13308
rect 22202 -13342 22258 -13308
rect 22292 -13342 22348 -13308
rect 22382 -13342 22438 -13308
rect 22472 -13342 22528 -13308
rect 22562 -13342 22618 -13308
rect 22652 -13342 22711 -13308
rect 22017 -13360 22711 -13342
rect 22017 -13394 22090 -13360
rect 22124 -13394 22190 -13360
rect 22224 -13394 22290 -13360
rect 22324 -13394 22390 -13360
rect 22424 -13394 22490 -13360
rect 22524 -13394 22590 -13360
rect 22624 -13394 22711 -13360
rect 22017 -13398 22711 -13394
rect 22017 -13432 22078 -13398
rect 22112 -13432 22168 -13398
rect 22202 -13432 22258 -13398
rect 22292 -13432 22348 -13398
rect 22382 -13432 22438 -13398
rect 22472 -13432 22528 -13398
rect 22562 -13432 22618 -13398
rect 22652 -13432 22711 -13398
rect 22017 -13460 22711 -13432
rect 22017 -13488 22090 -13460
rect 22124 -13488 22190 -13460
rect 22224 -13488 22290 -13460
rect 22324 -13488 22390 -13460
rect 22017 -13522 22078 -13488
rect 22124 -13494 22168 -13488
rect 22224 -13494 22258 -13488
rect 22324 -13494 22348 -13488
rect 22112 -13522 22168 -13494
rect 22202 -13522 22258 -13494
rect 22292 -13522 22348 -13494
rect 22382 -13494 22390 -13488
rect 22424 -13488 22490 -13460
rect 22424 -13494 22438 -13488
rect 22382 -13522 22438 -13494
rect 22472 -13494 22490 -13488
rect 22524 -13488 22590 -13460
rect 22624 -13488 22711 -13460
rect 22524 -13494 22528 -13488
rect 22472 -13522 22528 -13494
rect 22562 -13494 22590 -13488
rect 22562 -13522 22618 -13494
rect 22652 -13522 22711 -13488
rect 22017 -13581 22711 -13522
rect 22773 -12918 22792 -12884
rect 22826 -12918 22845 -12884
rect 22773 -12974 22845 -12918
rect 22773 -13008 22792 -12974
rect 22826 -13008 22845 -12974
rect 22773 -13064 22845 -13008
rect 22773 -13098 22792 -13064
rect 22826 -13098 22845 -13064
rect 22773 -13154 22845 -13098
rect 22773 -13188 22792 -13154
rect 22826 -13188 22845 -13154
rect 22773 -13244 22845 -13188
rect 22773 -13278 22792 -13244
rect 22826 -13278 22845 -13244
rect 22773 -13334 22845 -13278
rect 22773 -13368 22792 -13334
rect 22826 -13368 22845 -13334
rect 22773 -13424 22845 -13368
rect 22773 -13458 22792 -13424
rect 22826 -13458 22845 -13424
rect 22773 -13514 22845 -13458
rect 22773 -13548 22792 -13514
rect 22826 -13548 22845 -13514
rect 21883 -13643 21955 -13604
rect 22773 -13604 22845 -13548
rect 22773 -13638 22792 -13604
rect 22826 -13638 22845 -13604
rect 22773 -13643 22845 -13638
rect 21883 -13662 22845 -13643
rect 21883 -13696 21996 -13662
rect 22030 -13696 22086 -13662
rect 22120 -13696 22176 -13662
rect 22210 -13696 22266 -13662
rect 22300 -13696 22356 -13662
rect 22390 -13696 22446 -13662
rect 22480 -13696 22536 -13662
rect 22570 -13696 22626 -13662
rect 22660 -13696 22716 -13662
rect 22750 -13696 22845 -13662
rect 21883 -13702 22845 -13696
rect 22909 -12810 23107 -12802
rect 22909 -12844 22939 -12810
rect 22973 -12844 23040 -12810
rect 23074 -12844 23107 -12810
rect 22909 -12900 23107 -12844
rect 22909 -12934 22939 -12900
rect 22973 -12934 23040 -12900
rect 23074 -12934 23107 -12900
rect 22909 -12990 23107 -12934
rect 22909 -13024 22939 -12990
rect 22973 -13024 23040 -12990
rect 23074 -13024 23107 -12990
rect 22909 -13080 23107 -13024
rect 22909 -13114 22939 -13080
rect 22973 -13114 23040 -13080
rect 23074 -13114 23107 -13080
rect 22909 -13170 23107 -13114
rect 22909 -13204 22939 -13170
rect 22973 -13204 23040 -13170
rect 23074 -13204 23107 -13170
rect 22909 -13260 23107 -13204
rect 22909 -13294 22939 -13260
rect 22973 -13294 23040 -13260
rect 23074 -13294 23107 -13260
rect 22909 -13350 23107 -13294
rect 22909 -13384 22939 -13350
rect 22973 -13384 23040 -13350
rect 23074 -13384 23107 -13350
rect 22909 -13440 23107 -13384
rect 22909 -13474 22939 -13440
rect 22973 -13474 23040 -13440
rect 23074 -13474 23107 -13440
rect 22909 -13530 23107 -13474
rect 22909 -13564 22939 -13530
rect 22973 -13564 23040 -13530
rect 23074 -13564 23107 -13530
rect 22909 -13620 23107 -13564
rect 22909 -13654 22939 -13620
rect 22973 -13654 23040 -13620
rect 23074 -13654 23107 -13620
rect 22909 -13702 23107 -13654
rect 23171 -12806 23303 -12802
rect 23337 -12806 23393 -12772
rect 23427 -12806 23483 -12772
rect 23517 -12806 23573 -12772
rect 23607 -12806 23663 -12772
rect 23697 -12806 23753 -12772
rect 23787 -12806 23843 -12772
rect 23877 -12806 23933 -12772
rect 23967 -12806 24023 -12772
rect 24057 -12802 24591 -12772
rect 24057 -12806 24133 -12802
rect 23171 -12825 24133 -12806
rect 23171 -12850 23243 -12825
rect 23171 -12884 23190 -12850
rect 23224 -12884 23243 -12850
rect 23171 -12940 23243 -12884
rect 24061 -12884 24133 -12825
rect 23171 -12974 23190 -12940
rect 23224 -12974 23243 -12940
rect 23171 -13030 23243 -12974
rect 23171 -13064 23190 -13030
rect 23224 -13064 23243 -13030
rect 23171 -13120 23243 -13064
rect 23171 -13154 23190 -13120
rect 23224 -13154 23243 -13120
rect 23171 -13210 23243 -13154
rect 23171 -13244 23190 -13210
rect 23224 -13244 23243 -13210
rect 23171 -13300 23243 -13244
rect 23171 -13334 23190 -13300
rect 23224 -13334 23243 -13300
rect 23171 -13390 23243 -13334
rect 23171 -13424 23190 -13390
rect 23224 -13424 23243 -13390
rect 23171 -13480 23243 -13424
rect 23171 -13514 23190 -13480
rect 23224 -13514 23243 -13480
rect 23171 -13570 23243 -13514
rect 23171 -13604 23190 -13570
rect 23224 -13604 23243 -13570
rect 23305 -12948 23999 -12887
rect 23305 -12982 23366 -12948
rect 23400 -12960 23456 -12948
rect 23490 -12960 23546 -12948
rect 23580 -12960 23636 -12948
rect 23412 -12982 23456 -12960
rect 23512 -12982 23546 -12960
rect 23612 -12982 23636 -12960
rect 23670 -12960 23726 -12948
rect 23670 -12982 23678 -12960
rect 23305 -12994 23378 -12982
rect 23412 -12994 23478 -12982
rect 23512 -12994 23578 -12982
rect 23612 -12994 23678 -12982
rect 23712 -12982 23726 -12960
rect 23760 -12960 23816 -12948
rect 23760 -12982 23778 -12960
rect 23712 -12994 23778 -12982
rect 23812 -12982 23816 -12960
rect 23850 -12960 23906 -12948
rect 23850 -12982 23878 -12960
rect 23940 -12982 23999 -12948
rect 23812 -12994 23878 -12982
rect 23912 -12994 23999 -12982
rect 23305 -13038 23999 -12994
rect 23305 -13072 23366 -13038
rect 23400 -13060 23456 -13038
rect 23490 -13060 23546 -13038
rect 23580 -13060 23636 -13038
rect 23412 -13072 23456 -13060
rect 23512 -13072 23546 -13060
rect 23612 -13072 23636 -13060
rect 23670 -13060 23726 -13038
rect 23670 -13072 23678 -13060
rect 23305 -13094 23378 -13072
rect 23412 -13094 23478 -13072
rect 23512 -13094 23578 -13072
rect 23612 -13094 23678 -13072
rect 23712 -13072 23726 -13060
rect 23760 -13060 23816 -13038
rect 23760 -13072 23778 -13060
rect 23712 -13094 23778 -13072
rect 23812 -13072 23816 -13060
rect 23850 -13060 23906 -13038
rect 23850 -13072 23878 -13060
rect 23940 -13072 23999 -13038
rect 23812 -13094 23878 -13072
rect 23912 -13094 23999 -13072
rect 23305 -13128 23999 -13094
rect 23305 -13162 23366 -13128
rect 23400 -13160 23456 -13128
rect 23490 -13160 23546 -13128
rect 23580 -13160 23636 -13128
rect 23412 -13162 23456 -13160
rect 23512 -13162 23546 -13160
rect 23612 -13162 23636 -13160
rect 23670 -13160 23726 -13128
rect 23670 -13162 23678 -13160
rect 23305 -13194 23378 -13162
rect 23412 -13194 23478 -13162
rect 23512 -13194 23578 -13162
rect 23612 -13194 23678 -13162
rect 23712 -13162 23726 -13160
rect 23760 -13160 23816 -13128
rect 23760 -13162 23778 -13160
rect 23712 -13194 23778 -13162
rect 23812 -13162 23816 -13160
rect 23850 -13160 23906 -13128
rect 23850 -13162 23878 -13160
rect 23940 -13162 23999 -13128
rect 23812 -13194 23878 -13162
rect 23912 -13194 23999 -13162
rect 23305 -13218 23999 -13194
rect 23305 -13252 23366 -13218
rect 23400 -13252 23456 -13218
rect 23490 -13252 23546 -13218
rect 23580 -13252 23636 -13218
rect 23670 -13252 23726 -13218
rect 23760 -13252 23816 -13218
rect 23850 -13252 23906 -13218
rect 23940 -13252 23999 -13218
rect 23305 -13260 23999 -13252
rect 23305 -13294 23378 -13260
rect 23412 -13294 23478 -13260
rect 23512 -13294 23578 -13260
rect 23612 -13294 23678 -13260
rect 23712 -13294 23778 -13260
rect 23812 -13294 23878 -13260
rect 23912 -13294 23999 -13260
rect 23305 -13308 23999 -13294
rect 23305 -13342 23366 -13308
rect 23400 -13342 23456 -13308
rect 23490 -13342 23546 -13308
rect 23580 -13342 23636 -13308
rect 23670 -13342 23726 -13308
rect 23760 -13342 23816 -13308
rect 23850 -13342 23906 -13308
rect 23940 -13342 23999 -13308
rect 23305 -13360 23999 -13342
rect 23305 -13394 23378 -13360
rect 23412 -13394 23478 -13360
rect 23512 -13394 23578 -13360
rect 23612 -13394 23678 -13360
rect 23712 -13394 23778 -13360
rect 23812 -13394 23878 -13360
rect 23912 -13394 23999 -13360
rect 23305 -13398 23999 -13394
rect 23305 -13432 23366 -13398
rect 23400 -13432 23456 -13398
rect 23490 -13432 23546 -13398
rect 23580 -13432 23636 -13398
rect 23670 -13432 23726 -13398
rect 23760 -13432 23816 -13398
rect 23850 -13432 23906 -13398
rect 23940 -13432 23999 -13398
rect 23305 -13460 23999 -13432
rect 23305 -13488 23378 -13460
rect 23412 -13488 23478 -13460
rect 23512 -13488 23578 -13460
rect 23612 -13488 23678 -13460
rect 23305 -13522 23366 -13488
rect 23412 -13494 23456 -13488
rect 23512 -13494 23546 -13488
rect 23612 -13494 23636 -13488
rect 23400 -13522 23456 -13494
rect 23490 -13522 23546 -13494
rect 23580 -13522 23636 -13494
rect 23670 -13494 23678 -13488
rect 23712 -13488 23778 -13460
rect 23712 -13494 23726 -13488
rect 23670 -13522 23726 -13494
rect 23760 -13494 23778 -13488
rect 23812 -13488 23878 -13460
rect 23912 -13488 23999 -13460
rect 23812 -13494 23816 -13488
rect 23760 -13522 23816 -13494
rect 23850 -13494 23878 -13488
rect 23850 -13522 23906 -13494
rect 23940 -13522 23999 -13488
rect 23305 -13581 23999 -13522
rect 24061 -12918 24080 -12884
rect 24114 -12918 24133 -12884
rect 24061 -12974 24133 -12918
rect 24061 -13008 24080 -12974
rect 24114 -13008 24133 -12974
rect 24061 -13064 24133 -13008
rect 24061 -13098 24080 -13064
rect 24114 -13098 24133 -13064
rect 24061 -13154 24133 -13098
rect 24061 -13188 24080 -13154
rect 24114 -13188 24133 -13154
rect 24061 -13244 24133 -13188
rect 24061 -13278 24080 -13244
rect 24114 -13278 24133 -13244
rect 24061 -13334 24133 -13278
rect 24061 -13368 24080 -13334
rect 24114 -13368 24133 -13334
rect 24061 -13424 24133 -13368
rect 24061 -13458 24080 -13424
rect 24114 -13458 24133 -13424
rect 24061 -13514 24133 -13458
rect 24061 -13548 24080 -13514
rect 24114 -13548 24133 -13514
rect 23171 -13643 23243 -13604
rect 24061 -13604 24133 -13548
rect 24061 -13638 24080 -13604
rect 24114 -13638 24133 -13604
rect 24061 -13643 24133 -13638
rect 23171 -13662 24133 -13643
rect 23171 -13696 23284 -13662
rect 23318 -13696 23374 -13662
rect 23408 -13696 23464 -13662
rect 23498 -13696 23554 -13662
rect 23588 -13696 23644 -13662
rect 23678 -13696 23734 -13662
rect 23768 -13696 23824 -13662
rect 23858 -13696 23914 -13662
rect 23948 -13696 24004 -13662
rect 24038 -13696 24133 -13662
rect 23171 -13702 24133 -13696
rect 24197 -12810 24395 -12802
rect 24197 -12844 24227 -12810
rect 24261 -12844 24328 -12810
rect 24362 -12844 24395 -12810
rect 24197 -12900 24395 -12844
rect 24197 -12934 24227 -12900
rect 24261 -12934 24328 -12900
rect 24362 -12934 24395 -12900
rect 24197 -12990 24395 -12934
rect 24197 -13024 24227 -12990
rect 24261 -13024 24328 -12990
rect 24362 -13024 24395 -12990
rect 24197 -13080 24395 -13024
rect 24197 -13114 24227 -13080
rect 24261 -13114 24328 -13080
rect 24362 -13114 24395 -13080
rect 24197 -13170 24395 -13114
rect 24197 -13204 24227 -13170
rect 24261 -13204 24328 -13170
rect 24362 -13204 24395 -13170
rect 24197 -13260 24395 -13204
rect 24197 -13294 24227 -13260
rect 24261 -13294 24328 -13260
rect 24362 -13294 24395 -13260
rect 24197 -13350 24395 -13294
rect 24197 -13384 24227 -13350
rect 24261 -13384 24328 -13350
rect 24362 -13384 24395 -13350
rect 24197 -13440 24395 -13384
rect 24197 -13474 24227 -13440
rect 24261 -13474 24328 -13440
rect 24362 -13474 24395 -13440
rect 24197 -13530 24395 -13474
rect 24197 -13564 24227 -13530
rect 24261 -13564 24328 -13530
rect 24362 -13564 24395 -13530
rect 24197 -13620 24395 -13564
rect 24197 -13654 24227 -13620
rect 24261 -13654 24328 -13620
rect 24362 -13654 24395 -13620
rect 24197 -13702 24395 -13654
rect 24459 -12806 24591 -12802
rect 24625 -12806 24681 -12772
rect 24715 -12806 24771 -12772
rect 24805 -12806 24861 -12772
rect 24895 -12806 24951 -12772
rect 24985 -12806 25041 -12772
rect 25075 -12806 25131 -12772
rect 25165 -12806 25221 -12772
rect 25255 -12806 25311 -12772
rect 25345 -12802 25879 -12772
rect 25345 -12806 25421 -12802
rect 24459 -12825 25421 -12806
rect 24459 -12850 24531 -12825
rect 24459 -12884 24478 -12850
rect 24512 -12884 24531 -12850
rect 24459 -12940 24531 -12884
rect 25349 -12884 25421 -12825
rect 24459 -12974 24478 -12940
rect 24512 -12974 24531 -12940
rect 24459 -13030 24531 -12974
rect 24459 -13064 24478 -13030
rect 24512 -13064 24531 -13030
rect 24459 -13120 24531 -13064
rect 24459 -13154 24478 -13120
rect 24512 -13154 24531 -13120
rect 24459 -13210 24531 -13154
rect 24459 -13244 24478 -13210
rect 24512 -13244 24531 -13210
rect 24459 -13300 24531 -13244
rect 24459 -13334 24478 -13300
rect 24512 -13334 24531 -13300
rect 24459 -13390 24531 -13334
rect 24459 -13424 24478 -13390
rect 24512 -13424 24531 -13390
rect 24459 -13480 24531 -13424
rect 24459 -13514 24478 -13480
rect 24512 -13514 24531 -13480
rect 24459 -13570 24531 -13514
rect 24459 -13604 24478 -13570
rect 24512 -13604 24531 -13570
rect 24593 -12948 25287 -12887
rect 24593 -12982 24654 -12948
rect 24688 -12960 24744 -12948
rect 24778 -12960 24834 -12948
rect 24868 -12960 24924 -12948
rect 24700 -12982 24744 -12960
rect 24800 -12982 24834 -12960
rect 24900 -12982 24924 -12960
rect 24958 -12960 25014 -12948
rect 24958 -12982 24966 -12960
rect 24593 -12994 24666 -12982
rect 24700 -12994 24766 -12982
rect 24800 -12994 24866 -12982
rect 24900 -12994 24966 -12982
rect 25000 -12982 25014 -12960
rect 25048 -12960 25104 -12948
rect 25048 -12982 25066 -12960
rect 25000 -12994 25066 -12982
rect 25100 -12982 25104 -12960
rect 25138 -12960 25194 -12948
rect 25138 -12982 25166 -12960
rect 25228 -12982 25287 -12948
rect 25100 -12994 25166 -12982
rect 25200 -12994 25287 -12982
rect 24593 -13038 25287 -12994
rect 24593 -13072 24654 -13038
rect 24688 -13060 24744 -13038
rect 24778 -13060 24834 -13038
rect 24868 -13060 24924 -13038
rect 24700 -13072 24744 -13060
rect 24800 -13072 24834 -13060
rect 24900 -13072 24924 -13060
rect 24958 -13060 25014 -13038
rect 24958 -13072 24966 -13060
rect 24593 -13094 24666 -13072
rect 24700 -13094 24766 -13072
rect 24800 -13094 24866 -13072
rect 24900 -13094 24966 -13072
rect 25000 -13072 25014 -13060
rect 25048 -13060 25104 -13038
rect 25048 -13072 25066 -13060
rect 25000 -13094 25066 -13072
rect 25100 -13072 25104 -13060
rect 25138 -13060 25194 -13038
rect 25138 -13072 25166 -13060
rect 25228 -13072 25287 -13038
rect 25100 -13094 25166 -13072
rect 25200 -13094 25287 -13072
rect 24593 -13128 25287 -13094
rect 24593 -13162 24654 -13128
rect 24688 -13160 24744 -13128
rect 24778 -13160 24834 -13128
rect 24868 -13160 24924 -13128
rect 24700 -13162 24744 -13160
rect 24800 -13162 24834 -13160
rect 24900 -13162 24924 -13160
rect 24958 -13160 25014 -13128
rect 24958 -13162 24966 -13160
rect 24593 -13194 24666 -13162
rect 24700 -13194 24766 -13162
rect 24800 -13194 24866 -13162
rect 24900 -13194 24966 -13162
rect 25000 -13162 25014 -13160
rect 25048 -13160 25104 -13128
rect 25048 -13162 25066 -13160
rect 25000 -13194 25066 -13162
rect 25100 -13162 25104 -13160
rect 25138 -13160 25194 -13128
rect 25138 -13162 25166 -13160
rect 25228 -13162 25287 -13128
rect 25100 -13194 25166 -13162
rect 25200 -13194 25287 -13162
rect 24593 -13218 25287 -13194
rect 24593 -13252 24654 -13218
rect 24688 -13252 24744 -13218
rect 24778 -13252 24834 -13218
rect 24868 -13252 24924 -13218
rect 24958 -13252 25014 -13218
rect 25048 -13252 25104 -13218
rect 25138 -13252 25194 -13218
rect 25228 -13252 25287 -13218
rect 24593 -13260 25287 -13252
rect 24593 -13294 24666 -13260
rect 24700 -13294 24766 -13260
rect 24800 -13294 24866 -13260
rect 24900 -13294 24966 -13260
rect 25000 -13294 25066 -13260
rect 25100 -13294 25166 -13260
rect 25200 -13294 25287 -13260
rect 24593 -13308 25287 -13294
rect 24593 -13342 24654 -13308
rect 24688 -13342 24744 -13308
rect 24778 -13342 24834 -13308
rect 24868 -13342 24924 -13308
rect 24958 -13342 25014 -13308
rect 25048 -13342 25104 -13308
rect 25138 -13342 25194 -13308
rect 25228 -13342 25287 -13308
rect 24593 -13360 25287 -13342
rect 24593 -13394 24666 -13360
rect 24700 -13394 24766 -13360
rect 24800 -13394 24866 -13360
rect 24900 -13394 24966 -13360
rect 25000 -13394 25066 -13360
rect 25100 -13394 25166 -13360
rect 25200 -13394 25287 -13360
rect 24593 -13398 25287 -13394
rect 24593 -13432 24654 -13398
rect 24688 -13432 24744 -13398
rect 24778 -13432 24834 -13398
rect 24868 -13432 24924 -13398
rect 24958 -13432 25014 -13398
rect 25048 -13432 25104 -13398
rect 25138 -13432 25194 -13398
rect 25228 -13432 25287 -13398
rect 24593 -13460 25287 -13432
rect 24593 -13488 24666 -13460
rect 24700 -13488 24766 -13460
rect 24800 -13488 24866 -13460
rect 24900 -13488 24966 -13460
rect 24593 -13522 24654 -13488
rect 24700 -13494 24744 -13488
rect 24800 -13494 24834 -13488
rect 24900 -13494 24924 -13488
rect 24688 -13522 24744 -13494
rect 24778 -13522 24834 -13494
rect 24868 -13522 24924 -13494
rect 24958 -13494 24966 -13488
rect 25000 -13488 25066 -13460
rect 25000 -13494 25014 -13488
rect 24958 -13522 25014 -13494
rect 25048 -13494 25066 -13488
rect 25100 -13488 25166 -13460
rect 25200 -13488 25287 -13460
rect 25100 -13494 25104 -13488
rect 25048 -13522 25104 -13494
rect 25138 -13494 25166 -13488
rect 25138 -13522 25194 -13494
rect 25228 -13522 25287 -13488
rect 24593 -13581 25287 -13522
rect 25349 -12918 25368 -12884
rect 25402 -12918 25421 -12884
rect 25349 -12974 25421 -12918
rect 25349 -13008 25368 -12974
rect 25402 -13008 25421 -12974
rect 25349 -13064 25421 -13008
rect 25349 -13098 25368 -13064
rect 25402 -13098 25421 -13064
rect 25349 -13154 25421 -13098
rect 25349 -13188 25368 -13154
rect 25402 -13188 25421 -13154
rect 25349 -13244 25421 -13188
rect 25349 -13278 25368 -13244
rect 25402 -13278 25421 -13244
rect 25349 -13334 25421 -13278
rect 25349 -13368 25368 -13334
rect 25402 -13368 25421 -13334
rect 25349 -13424 25421 -13368
rect 25349 -13458 25368 -13424
rect 25402 -13458 25421 -13424
rect 25349 -13514 25421 -13458
rect 25349 -13548 25368 -13514
rect 25402 -13548 25421 -13514
rect 24459 -13643 24531 -13604
rect 25349 -13604 25421 -13548
rect 25349 -13638 25368 -13604
rect 25402 -13638 25421 -13604
rect 25349 -13643 25421 -13638
rect 24459 -13662 25421 -13643
rect 24459 -13696 24572 -13662
rect 24606 -13696 24662 -13662
rect 24696 -13696 24752 -13662
rect 24786 -13696 24842 -13662
rect 24876 -13696 24932 -13662
rect 24966 -13696 25022 -13662
rect 25056 -13696 25112 -13662
rect 25146 -13696 25202 -13662
rect 25236 -13696 25292 -13662
rect 25326 -13696 25421 -13662
rect 24459 -13702 25421 -13696
rect 25485 -12810 25683 -12802
rect 25485 -12844 25515 -12810
rect 25549 -12844 25616 -12810
rect 25650 -12844 25683 -12810
rect 25485 -12900 25683 -12844
rect 25485 -12934 25515 -12900
rect 25549 -12934 25616 -12900
rect 25650 -12934 25683 -12900
rect 25485 -12990 25683 -12934
rect 25485 -13024 25515 -12990
rect 25549 -13024 25616 -12990
rect 25650 -13024 25683 -12990
rect 25485 -13080 25683 -13024
rect 25485 -13114 25515 -13080
rect 25549 -13114 25616 -13080
rect 25650 -13114 25683 -13080
rect 25485 -13170 25683 -13114
rect 25485 -13204 25515 -13170
rect 25549 -13204 25616 -13170
rect 25650 -13204 25683 -13170
rect 25485 -13260 25683 -13204
rect 25485 -13294 25515 -13260
rect 25549 -13294 25616 -13260
rect 25650 -13294 25683 -13260
rect 25485 -13350 25683 -13294
rect 25485 -13384 25515 -13350
rect 25549 -13384 25616 -13350
rect 25650 -13384 25683 -13350
rect 25485 -13440 25683 -13384
rect 25485 -13474 25515 -13440
rect 25549 -13474 25616 -13440
rect 25650 -13474 25683 -13440
rect 25485 -13530 25683 -13474
rect 25485 -13564 25515 -13530
rect 25549 -13564 25616 -13530
rect 25650 -13564 25683 -13530
rect 25485 -13620 25683 -13564
rect 25485 -13654 25515 -13620
rect 25549 -13654 25616 -13620
rect 25650 -13654 25683 -13620
rect 25485 -13702 25683 -13654
rect 25747 -12806 25879 -12802
rect 25913 -12806 25969 -12772
rect 26003 -12806 26059 -12772
rect 26093 -12806 26149 -12772
rect 26183 -12806 26239 -12772
rect 26273 -12806 26329 -12772
rect 26363 -12806 26419 -12772
rect 26453 -12806 26509 -12772
rect 26543 -12806 26599 -12772
rect 26633 -12802 26872 -12772
rect 26633 -12806 26709 -12802
rect 25747 -12825 26709 -12806
rect 25747 -12850 25819 -12825
rect 25747 -12884 25766 -12850
rect 25800 -12884 25819 -12850
rect 25747 -12940 25819 -12884
rect 26637 -12884 26709 -12825
rect 25747 -12974 25766 -12940
rect 25800 -12974 25819 -12940
rect 25747 -13030 25819 -12974
rect 25747 -13064 25766 -13030
rect 25800 -13064 25819 -13030
rect 25747 -13120 25819 -13064
rect 25747 -13154 25766 -13120
rect 25800 -13154 25819 -13120
rect 25747 -13210 25819 -13154
rect 25747 -13244 25766 -13210
rect 25800 -13244 25819 -13210
rect 25747 -13300 25819 -13244
rect 25747 -13334 25766 -13300
rect 25800 -13334 25819 -13300
rect 25747 -13390 25819 -13334
rect 25747 -13424 25766 -13390
rect 25800 -13424 25819 -13390
rect 25747 -13480 25819 -13424
rect 25747 -13514 25766 -13480
rect 25800 -13514 25819 -13480
rect 25747 -13570 25819 -13514
rect 25747 -13604 25766 -13570
rect 25800 -13604 25819 -13570
rect 25881 -12948 26575 -12887
rect 25881 -12982 25942 -12948
rect 25976 -12960 26032 -12948
rect 26066 -12960 26122 -12948
rect 26156 -12960 26212 -12948
rect 25988 -12982 26032 -12960
rect 26088 -12982 26122 -12960
rect 26188 -12982 26212 -12960
rect 26246 -12960 26302 -12948
rect 26246 -12982 26254 -12960
rect 25881 -12994 25954 -12982
rect 25988 -12994 26054 -12982
rect 26088 -12994 26154 -12982
rect 26188 -12994 26254 -12982
rect 26288 -12982 26302 -12960
rect 26336 -12960 26392 -12948
rect 26336 -12982 26354 -12960
rect 26288 -12994 26354 -12982
rect 26388 -12982 26392 -12960
rect 26426 -12960 26482 -12948
rect 26426 -12982 26454 -12960
rect 26516 -12982 26575 -12948
rect 26388 -12994 26454 -12982
rect 26488 -12994 26575 -12982
rect 25881 -13038 26575 -12994
rect 25881 -13072 25942 -13038
rect 25976 -13060 26032 -13038
rect 26066 -13060 26122 -13038
rect 26156 -13060 26212 -13038
rect 25988 -13072 26032 -13060
rect 26088 -13072 26122 -13060
rect 26188 -13072 26212 -13060
rect 26246 -13060 26302 -13038
rect 26246 -13072 26254 -13060
rect 25881 -13094 25954 -13072
rect 25988 -13094 26054 -13072
rect 26088 -13094 26154 -13072
rect 26188 -13094 26254 -13072
rect 26288 -13072 26302 -13060
rect 26336 -13060 26392 -13038
rect 26336 -13072 26354 -13060
rect 26288 -13094 26354 -13072
rect 26388 -13072 26392 -13060
rect 26426 -13060 26482 -13038
rect 26426 -13072 26454 -13060
rect 26516 -13072 26575 -13038
rect 26388 -13094 26454 -13072
rect 26488 -13094 26575 -13072
rect 25881 -13128 26575 -13094
rect 25881 -13162 25942 -13128
rect 25976 -13160 26032 -13128
rect 26066 -13160 26122 -13128
rect 26156 -13160 26212 -13128
rect 25988 -13162 26032 -13160
rect 26088 -13162 26122 -13160
rect 26188 -13162 26212 -13160
rect 26246 -13160 26302 -13128
rect 26246 -13162 26254 -13160
rect 25881 -13194 25954 -13162
rect 25988 -13194 26054 -13162
rect 26088 -13194 26154 -13162
rect 26188 -13194 26254 -13162
rect 26288 -13162 26302 -13160
rect 26336 -13160 26392 -13128
rect 26336 -13162 26354 -13160
rect 26288 -13194 26354 -13162
rect 26388 -13162 26392 -13160
rect 26426 -13160 26482 -13128
rect 26426 -13162 26454 -13160
rect 26516 -13162 26575 -13128
rect 26388 -13194 26454 -13162
rect 26488 -13194 26575 -13162
rect 25881 -13218 26575 -13194
rect 25881 -13252 25942 -13218
rect 25976 -13252 26032 -13218
rect 26066 -13252 26122 -13218
rect 26156 -13252 26212 -13218
rect 26246 -13252 26302 -13218
rect 26336 -13252 26392 -13218
rect 26426 -13252 26482 -13218
rect 26516 -13252 26575 -13218
rect 25881 -13260 26575 -13252
rect 25881 -13294 25954 -13260
rect 25988 -13294 26054 -13260
rect 26088 -13294 26154 -13260
rect 26188 -13294 26254 -13260
rect 26288 -13294 26354 -13260
rect 26388 -13294 26454 -13260
rect 26488 -13294 26575 -13260
rect 25881 -13308 26575 -13294
rect 25881 -13342 25942 -13308
rect 25976 -13342 26032 -13308
rect 26066 -13342 26122 -13308
rect 26156 -13342 26212 -13308
rect 26246 -13342 26302 -13308
rect 26336 -13342 26392 -13308
rect 26426 -13342 26482 -13308
rect 26516 -13342 26575 -13308
rect 25881 -13360 26575 -13342
rect 25881 -13394 25954 -13360
rect 25988 -13394 26054 -13360
rect 26088 -13394 26154 -13360
rect 26188 -13394 26254 -13360
rect 26288 -13394 26354 -13360
rect 26388 -13394 26454 -13360
rect 26488 -13394 26575 -13360
rect 25881 -13398 26575 -13394
rect 25881 -13432 25942 -13398
rect 25976 -13432 26032 -13398
rect 26066 -13432 26122 -13398
rect 26156 -13432 26212 -13398
rect 26246 -13432 26302 -13398
rect 26336 -13432 26392 -13398
rect 26426 -13432 26482 -13398
rect 26516 -13432 26575 -13398
rect 25881 -13460 26575 -13432
rect 25881 -13488 25954 -13460
rect 25988 -13488 26054 -13460
rect 26088 -13488 26154 -13460
rect 26188 -13488 26254 -13460
rect 25881 -13522 25942 -13488
rect 25988 -13494 26032 -13488
rect 26088 -13494 26122 -13488
rect 26188 -13494 26212 -13488
rect 25976 -13522 26032 -13494
rect 26066 -13522 26122 -13494
rect 26156 -13522 26212 -13494
rect 26246 -13494 26254 -13488
rect 26288 -13488 26354 -13460
rect 26288 -13494 26302 -13488
rect 26246 -13522 26302 -13494
rect 26336 -13494 26354 -13488
rect 26388 -13488 26454 -13460
rect 26488 -13488 26575 -13460
rect 26388 -13494 26392 -13488
rect 26336 -13522 26392 -13494
rect 26426 -13494 26454 -13488
rect 26426 -13522 26482 -13494
rect 26516 -13522 26575 -13488
rect 25881 -13581 26575 -13522
rect 26637 -12918 26656 -12884
rect 26690 -12918 26709 -12884
rect 26637 -12974 26709 -12918
rect 26637 -13008 26656 -12974
rect 26690 -13008 26709 -12974
rect 26637 -13064 26709 -13008
rect 26637 -13098 26656 -13064
rect 26690 -13098 26709 -13064
rect 26637 -13154 26709 -13098
rect 26637 -13188 26656 -13154
rect 26690 -13188 26709 -13154
rect 26637 -13244 26709 -13188
rect 26637 -13278 26656 -13244
rect 26690 -13278 26709 -13244
rect 26637 -13334 26709 -13278
rect 26637 -13368 26656 -13334
rect 26690 -13368 26709 -13334
rect 26637 -13424 26709 -13368
rect 26637 -13458 26656 -13424
rect 26690 -13458 26709 -13424
rect 26637 -13514 26709 -13458
rect 26637 -13548 26656 -13514
rect 26690 -13548 26709 -13514
rect 25747 -13643 25819 -13604
rect 26637 -13604 26709 -13548
rect 26637 -13638 26656 -13604
rect 26690 -13638 26709 -13604
rect 26637 -13643 26709 -13638
rect 25747 -13662 26709 -13643
rect 25747 -13696 25860 -13662
rect 25894 -13696 25950 -13662
rect 25984 -13696 26040 -13662
rect 26074 -13696 26130 -13662
rect 26164 -13696 26220 -13662
rect 26254 -13696 26310 -13662
rect 26344 -13696 26400 -13662
rect 26434 -13696 26490 -13662
rect 26524 -13696 26580 -13662
rect 26614 -13696 26709 -13662
rect 25747 -13702 26709 -13696
rect 26773 -12810 26872 -12802
rect 26773 -12844 26803 -12810
rect 26837 -12844 26872 -12810
rect 26773 -12900 26872 -12844
rect 26773 -12934 26803 -12900
rect 26837 -12934 26872 -12900
rect 26773 -12990 26872 -12934
rect 26773 -13024 26803 -12990
rect 26837 -13024 26872 -12990
rect 26773 -13080 26872 -13024
rect 26773 -13114 26803 -13080
rect 26837 -13114 26872 -13080
rect 26773 -13170 26872 -13114
rect 26773 -13204 26803 -13170
rect 26837 -13204 26872 -13170
rect 26773 -13260 26872 -13204
rect 26773 -13294 26803 -13260
rect 26837 -13294 26872 -13260
rect 26773 -13350 26872 -13294
rect 26773 -13384 26803 -13350
rect 26837 -13384 26872 -13350
rect 26773 -13440 26872 -13384
rect 26773 -13474 26803 -13440
rect 26837 -13474 26872 -13440
rect 26773 -13530 26872 -13474
rect 26773 -13564 26803 -13530
rect 26837 -13564 26872 -13530
rect 26773 -13620 26872 -13564
rect 26773 -13654 26803 -13620
rect 26837 -13654 26872 -13620
rect 26773 -13702 26872 -13654
rect 16568 -13710 26872 -13702
rect 16568 -13744 16600 -13710
rect 16634 -13744 17787 -13710
rect 17821 -13744 17888 -13710
rect 17922 -13744 19075 -13710
rect 19109 -13744 19176 -13710
rect 19210 -13744 20363 -13710
rect 20397 -13744 20464 -13710
rect 20498 -13744 21651 -13710
rect 21685 -13744 21752 -13710
rect 21786 -13744 22939 -13710
rect 22973 -13744 23040 -13710
rect 23074 -13744 24227 -13710
rect 24261 -13744 24328 -13710
rect 24362 -13744 25515 -13710
rect 25549 -13744 25616 -13710
rect 25650 -13744 26803 -13710
rect 26837 -13744 26872 -13710
rect 16568 -13811 26872 -13744
rect 16568 -13845 16684 -13811
rect 16718 -13845 16774 -13811
rect 16808 -13845 16864 -13811
rect 16898 -13845 16954 -13811
rect 16988 -13845 17044 -13811
rect 17078 -13845 17134 -13811
rect 17168 -13845 17224 -13811
rect 17258 -13845 17314 -13811
rect 17348 -13845 17404 -13811
rect 17438 -13845 17494 -13811
rect 17528 -13845 17584 -13811
rect 17618 -13845 17674 -13811
rect 17708 -13845 17764 -13811
rect 17798 -13845 17972 -13811
rect 18006 -13845 18062 -13811
rect 18096 -13845 18152 -13811
rect 18186 -13845 18242 -13811
rect 18276 -13845 18332 -13811
rect 18366 -13845 18422 -13811
rect 18456 -13845 18512 -13811
rect 18546 -13845 18602 -13811
rect 18636 -13845 18692 -13811
rect 18726 -13845 18782 -13811
rect 18816 -13845 18872 -13811
rect 18906 -13845 18962 -13811
rect 18996 -13845 19052 -13811
rect 19086 -13845 19260 -13811
rect 19294 -13845 19350 -13811
rect 19384 -13845 19440 -13811
rect 19474 -13845 19530 -13811
rect 19564 -13845 19620 -13811
rect 19654 -13845 19710 -13811
rect 19744 -13845 19800 -13811
rect 19834 -13845 19890 -13811
rect 19924 -13845 19980 -13811
rect 20014 -13845 20070 -13811
rect 20104 -13845 20160 -13811
rect 20194 -13845 20250 -13811
rect 20284 -13845 20340 -13811
rect 20374 -13845 20548 -13811
rect 20582 -13845 20638 -13811
rect 20672 -13845 20728 -13811
rect 20762 -13845 20818 -13811
rect 20852 -13845 20908 -13811
rect 20942 -13845 20998 -13811
rect 21032 -13845 21088 -13811
rect 21122 -13845 21178 -13811
rect 21212 -13845 21268 -13811
rect 21302 -13845 21358 -13811
rect 21392 -13845 21448 -13811
rect 21482 -13845 21538 -13811
rect 21572 -13845 21628 -13811
rect 21662 -13845 21836 -13811
rect 21870 -13845 21926 -13811
rect 21960 -13845 22016 -13811
rect 22050 -13845 22106 -13811
rect 22140 -13845 22196 -13811
rect 22230 -13845 22286 -13811
rect 22320 -13845 22376 -13811
rect 22410 -13845 22466 -13811
rect 22500 -13845 22556 -13811
rect 22590 -13845 22646 -13811
rect 22680 -13845 22736 -13811
rect 22770 -13845 22826 -13811
rect 22860 -13845 22916 -13811
rect 22950 -13845 23124 -13811
rect 23158 -13845 23214 -13811
rect 23248 -13845 23304 -13811
rect 23338 -13845 23394 -13811
rect 23428 -13845 23484 -13811
rect 23518 -13845 23574 -13811
rect 23608 -13845 23664 -13811
rect 23698 -13845 23754 -13811
rect 23788 -13845 23844 -13811
rect 23878 -13845 23934 -13811
rect 23968 -13845 24024 -13811
rect 24058 -13845 24114 -13811
rect 24148 -13845 24204 -13811
rect 24238 -13845 24412 -13811
rect 24446 -13845 24502 -13811
rect 24536 -13845 24592 -13811
rect 24626 -13845 24682 -13811
rect 24716 -13845 24772 -13811
rect 24806 -13845 24862 -13811
rect 24896 -13845 24952 -13811
rect 24986 -13845 25042 -13811
rect 25076 -13845 25132 -13811
rect 25166 -13845 25222 -13811
rect 25256 -13845 25312 -13811
rect 25346 -13845 25402 -13811
rect 25436 -13845 25492 -13811
rect 25526 -13845 25700 -13811
rect 25734 -13845 25790 -13811
rect 25824 -13845 25880 -13811
rect 25914 -13845 25970 -13811
rect 26004 -13845 26060 -13811
rect 26094 -13845 26150 -13811
rect 26184 -13845 26240 -13811
rect 26274 -13845 26330 -13811
rect 26364 -13845 26420 -13811
rect 26454 -13845 26510 -13811
rect 26544 -13845 26600 -13811
rect 26634 -13845 26690 -13811
rect 26724 -13845 26780 -13811
rect 26814 -13845 26872 -13811
rect 16568 -13912 26872 -13845
rect 16568 -13946 16684 -13912
rect 16718 -13946 16774 -13912
rect 16808 -13946 16864 -13912
rect 16898 -13946 16954 -13912
rect 16988 -13946 17044 -13912
rect 17078 -13946 17134 -13912
rect 17168 -13946 17224 -13912
rect 17258 -13946 17314 -13912
rect 17348 -13946 17404 -13912
rect 17438 -13946 17494 -13912
rect 17528 -13946 17584 -13912
rect 17618 -13946 17674 -13912
rect 17708 -13946 17764 -13912
rect 17798 -13946 17972 -13912
rect 18006 -13946 18062 -13912
rect 18096 -13946 18152 -13912
rect 18186 -13946 18242 -13912
rect 18276 -13946 18332 -13912
rect 18366 -13946 18422 -13912
rect 18456 -13946 18512 -13912
rect 18546 -13946 18602 -13912
rect 18636 -13946 18692 -13912
rect 18726 -13946 18782 -13912
rect 18816 -13946 18872 -13912
rect 18906 -13946 18962 -13912
rect 18996 -13946 19052 -13912
rect 19086 -13946 19260 -13912
rect 19294 -13946 19350 -13912
rect 19384 -13946 19440 -13912
rect 19474 -13946 19530 -13912
rect 19564 -13946 19620 -13912
rect 19654 -13946 19710 -13912
rect 19744 -13946 19800 -13912
rect 19834 -13946 19890 -13912
rect 19924 -13946 19980 -13912
rect 20014 -13946 20070 -13912
rect 20104 -13946 20160 -13912
rect 20194 -13946 20250 -13912
rect 20284 -13946 20340 -13912
rect 20374 -13946 20548 -13912
rect 20582 -13946 20638 -13912
rect 20672 -13946 20728 -13912
rect 20762 -13946 20818 -13912
rect 20852 -13946 20908 -13912
rect 20942 -13946 20998 -13912
rect 21032 -13946 21088 -13912
rect 21122 -13946 21178 -13912
rect 21212 -13946 21268 -13912
rect 21302 -13946 21358 -13912
rect 21392 -13946 21448 -13912
rect 21482 -13946 21538 -13912
rect 21572 -13946 21628 -13912
rect 21662 -13946 21836 -13912
rect 21870 -13946 21926 -13912
rect 21960 -13946 22016 -13912
rect 22050 -13946 22106 -13912
rect 22140 -13946 22196 -13912
rect 22230 -13946 22286 -13912
rect 22320 -13946 22376 -13912
rect 22410 -13946 22466 -13912
rect 22500 -13946 22556 -13912
rect 22590 -13946 22646 -13912
rect 22680 -13946 22736 -13912
rect 22770 -13946 22826 -13912
rect 22860 -13946 22916 -13912
rect 22950 -13946 23124 -13912
rect 23158 -13946 23214 -13912
rect 23248 -13946 23304 -13912
rect 23338 -13946 23394 -13912
rect 23428 -13946 23484 -13912
rect 23518 -13946 23574 -13912
rect 23608 -13946 23664 -13912
rect 23698 -13946 23754 -13912
rect 23788 -13946 23844 -13912
rect 23878 -13946 23934 -13912
rect 23968 -13946 24024 -13912
rect 24058 -13946 24114 -13912
rect 24148 -13946 24204 -13912
rect 24238 -13946 24412 -13912
rect 24446 -13946 24502 -13912
rect 24536 -13946 24592 -13912
rect 24626 -13946 24682 -13912
rect 24716 -13946 24772 -13912
rect 24806 -13946 24862 -13912
rect 24896 -13946 24952 -13912
rect 24986 -13946 25042 -13912
rect 25076 -13946 25132 -13912
rect 25166 -13946 25222 -13912
rect 25256 -13946 25312 -13912
rect 25346 -13946 25402 -13912
rect 25436 -13946 25492 -13912
rect 25526 -13946 25700 -13912
rect 25734 -13946 25790 -13912
rect 25824 -13946 25880 -13912
rect 25914 -13946 25970 -13912
rect 26004 -13946 26060 -13912
rect 26094 -13946 26150 -13912
rect 26184 -13946 26240 -13912
rect 26274 -13946 26330 -13912
rect 26364 -13946 26420 -13912
rect 26454 -13946 26510 -13912
rect 26544 -13946 26600 -13912
rect 26634 -13946 26690 -13912
rect 26724 -13946 26780 -13912
rect 26814 -13946 26872 -13912
rect 16568 -14008 26872 -13946
rect 16568 -14042 16600 -14008
rect 16634 -14042 17787 -14008
rect 17821 -14042 17888 -14008
rect 17922 -14042 19075 -14008
rect 19109 -14042 19176 -14008
rect 19210 -14042 20363 -14008
rect 20397 -14042 20464 -14008
rect 20498 -14042 21651 -14008
rect 21685 -14042 21752 -14008
rect 21786 -14042 22939 -14008
rect 22973 -14042 23040 -14008
rect 23074 -14042 24227 -14008
rect 24261 -14042 24328 -14008
rect 24362 -14042 25515 -14008
rect 25549 -14042 25616 -14008
rect 25650 -14042 26803 -14008
rect 26837 -14042 26872 -14008
rect 16568 -14060 26872 -14042
rect 16568 -14094 16863 -14060
rect 16897 -14094 16953 -14060
rect 16987 -14094 17043 -14060
rect 17077 -14094 17133 -14060
rect 17167 -14094 17223 -14060
rect 17257 -14094 17313 -14060
rect 17347 -14094 17403 -14060
rect 17437 -14094 17493 -14060
rect 17527 -14094 17583 -14060
rect 17617 -14094 18151 -14060
rect 18185 -14094 18241 -14060
rect 18275 -14094 18331 -14060
rect 18365 -14094 18421 -14060
rect 18455 -14094 18511 -14060
rect 18545 -14094 18601 -14060
rect 18635 -14094 18691 -14060
rect 18725 -14094 18781 -14060
rect 18815 -14094 18871 -14060
rect 18905 -14094 19439 -14060
rect 19473 -14094 19529 -14060
rect 19563 -14094 19619 -14060
rect 19653 -14094 19709 -14060
rect 19743 -14094 19799 -14060
rect 19833 -14094 19889 -14060
rect 19923 -14094 19979 -14060
rect 20013 -14094 20069 -14060
rect 20103 -14094 20159 -14060
rect 20193 -14094 20727 -14060
rect 20761 -14094 20817 -14060
rect 20851 -14094 20907 -14060
rect 20941 -14094 20997 -14060
rect 21031 -14094 21087 -14060
rect 21121 -14094 21177 -14060
rect 21211 -14094 21267 -14060
rect 21301 -14094 21357 -14060
rect 21391 -14094 21447 -14060
rect 21481 -14094 22015 -14060
rect 22049 -14094 22105 -14060
rect 22139 -14094 22195 -14060
rect 22229 -14094 22285 -14060
rect 22319 -14094 22375 -14060
rect 22409 -14094 22465 -14060
rect 22499 -14094 22555 -14060
rect 22589 -14094 22645 -14060
rect 22679 -14094 22735 -14060
rect 22769 -14094 23303 -14060
rect 23337 -14094 23393 -14060
rect 23427 -14094 23483 -14060
rect 23517 -14094 23573 -14060
rect 23607 -14094 23663 -14060
rect 23697 -14094 23753 -14060
rect 23787 -14094 23843 -14060
rect 23877 -14094 23933 -14060
rect 23967 -14094 24023 -14060
rect 24057 -14094 24591 -14060
rect 24625 -14094 24681 -14060
rect 24715 -14094 24771 -14060
rect 24805 -14094 24861 -14060
rect 24895 -14094 24951 -14060
rect 24985 -14094 25041 -14060
rect 25075 -14094 25131 -14060
rect 25165 -14094 25221 -14060
rect 25255 -14094 25311 -14060
rect 25345 -14094 25879 -14060
rect 25913 -14094 25969 -14060
rect 26003 -14094 26059 -14060
rect 26093 -14094 26149 -14060
rect 26183 -14094 26239 -14060
rect 26273 -14094 26329 -14060
rect 26363 -14094 26419 -14060
rect 26453 -14094 26509 -14060
rect 26543 -14094 26599 -14060
rect 26633 -14094 26872 -14060
rect 16568 -14098 26872 -14094
rect 16568 -14132 16600 -14098
rect 16634 -14102 17787 -14098
rect 16634 -14132 16667 -14102
rect 16568 -14188 16667 -14132
rect 16568 -14222 16600 -14188
rect 16634 -14222 16667 -14188
rect 16568 -14278 16667 -14222
rect 16568 -14312 16600 -14278
rect 16634 -14312 16667 -14278
rect 16568 -14368 16667 -14312
rect 16568 -14402 16600 -14368
rect 16634 -14402 16667 -14368
rect 16568 -14458 16667 -14402
rect 16568 -14492 16600 -14458
rect 16634 -14492 16667 -14458
rect 16568 -14548 16667 -14492
rect 16568 -14582 16600 -14548
rect 16634 -14582 16667 -14548
rect 16568 -14638 16667 -14582
rect 16568 -14672 16600 -14638
rect 16634 -14672 16667 -14638
rect 16568 -14728 16667 -14672
rect 16568 -14762 16600 -14728
rect 16634 -14762 16667 -14728
rect 16568 -14818 16667 -14762
rect 16568 -14852 16600 -14818
rect 16634 -14852 16667 -14818
rect 16568 -14908 16667 -14852
rect 16568 -14942 16600 -14908
rect 16634 -14942 16667 -14908
rect 16568 -14998 16667 -14942
rect 16568 -15032 16600 -14998
rect 16634 -15002 16667 -14998
rect 16731 -14113 17693 -14102
rect 16731 -14138 16803 -14113
rect 16731 -14172 16750 -14138
rect 16784 -14172 16803 -14138
rect 16731 -14228 16803 -14172
rect 17621 -14172 17693 -14113
rect 16731 -14262 16750 -14228
rect 16784 -14262 16803 -14228
rect 16731 -14318 16803 -14262
rect 16731 -14352 16750 -14318
rect 16784 -14352 16803 -14318
rect 16731 -14408 16803 -14352
rect 16731 -14442 16750 -14408
rect 16784 -14442 16803 -14408
rect 16731 -14498 16803 -14442
rect 16731 -14532 16750 -14498
rect 16784 -14532 16803 -14498
rect 16731 -14588 16803 -14532
rect 16731 -14622 16750 -14588
rect 16784 -14622 16803 -14588
rect 16731 -14678 16803 -14622
rect 16731 -14712 16750 -14678
rect 16784 -14712 16803 -14678
rect 16731 -14768 16803 -14712
rect 16731 -14802 16750 -14768
rect 16784 -14802 16803 -14768
rect 16731 -14858 16803 -14802
rect 16731 -14892 16750 -14858
rect 16784 -14892 16803 -14858
rect 16865 -14236 17559 -14175
rect 16865 -14270 16926 -14236
rect 16960 -14248 17016 -14236
rect 17050 -14248 17106 -14236
rect 17140 -14248 17196 -14236
rect 16972 -14270 17016 -14248
rect 17072 -14270 17106 -14248
rect 17172 -14270 17196 -14248
rect 17230 -14248 17286 -14236
rect 17230 -14270 17238 -14248
rect 16865 -14282 16938 -14270
rect 16972 -14282 17038 -14270
rect 17072 -14282 17138 -14270
rect 17172 -14282 17238 -14270
rect 17272 -14270 17286 -14248
rect 17320 -14248 17376 -14236
rect 17320 -14270 17338 -14248
rect 17272 -14282 17338 -14270
rect 17372 -14270 17376 -14248
rect 17410 -14248 17466 -14236
rect 17410 -14270 17438 -14248
rect 17500 -14270 17559 -14236
rect 17372 -14282 17438 -14270
rect 17472 -14282 17559 -14270
rect 16865 -14326 17559 -14282
rect 16865 -14360 16926 -14326
rect 16960 -14348 17016 -14326
rect 17050 -14348 17106 -14326
rect 17140 -14348 17196 -14326
rect 16972 -14360 17016 -14348
rect 17072 -14360 17106 -14348
rect 17172 -14360 17196 -14348
rect 17230 -14348 17286 -14326
rect 17230 -14360 17238 -14348
rect 16865 -14382 16938 -14360
rect 16972 -14382 17038 -14360
rect 17072 -14382 17138 -14360
rect 17172 -14382 17238 -14360
rect 17272 -14360 17286 -14348
rect 17320 -14348 17376 -14326
rect 17320 -14360 17338 -14348
rect 17272 -14382 17338 -14360
rect 17372 -14360 17376 -14348
rect 17410 -14348 17466 -14326
rect 17410 -14360 17438 -14348
rect 17500 -14360 17559 -14326
rect 17372 -14382 17438 -14360
rect 17472 -14382 17559 -14360
rect 16865 -14416 17559 -14382
rect 16865 -14450 16926 -14416
rect 16960 -14448 17016 -14416
rect 17050 -14448 17106 -14416
rect 17140 -14448 17196 -14416
rect 16972 -14450 17016 -14448
rect 17072 -14450 17106 -14448
rect 17172 -14450 17196 -14448
rect 17230 -14448 17286 -14416
rect 17230 -14450 17238 -14448
rect 16865 -14482 16938 -14450
rect 16972 -14482 17038 -14450
rect 17072 -14482 17138 -14450
rect 17172 -14482 17238 -14450
rect 17272 -14450 17286 -14448
rect 17320 -14448 17376 -14416
rect 17320 -14450 17338 -14448
rect 17272 -14482 17338 -14450
rect 17372 -14450 17376 -14448
rect 17410 -14448 17466 -14416
rect 17410 -14450 17438 -14448
rect 17500 -14450 17559 -14416
rect 17372 -14482 17438 -14450
rect 17472 -14482 17559 -14450
rect 16865 -14506 17559 -14482
rect 16865 -14540 16926 -14506
rect 16960 -14540 17016 -14506
rect 17050 -14540 17106 -14506
rect 17140 -14540 17196 -14506
rect 17230 -14540 17286 -14506
rect 17320 -14540 17376 -14506
rect 17410 -14540 17466 -14506
rect 17500 -14540 17559 -14506
rect 16865 -14548 17559 -14540
rect 16865 -14582 16938 -14548
rect 16972 -14582 17038 -14548
rect 17072 -14582 17138 -14548
rect 17172 -14582 17238 -14548
rect 17272 -14582 17338 -14548
rect 17372 -14582 17438 -14548
rect 17472 -14582 17559 -14548
rect 16865 -14596 17559 -14582
rect 16865 -14630 16926 -14596
rect 16960 -14630 17016 -14596
rect 17050 -14630 17106 -14596
rect 17140 -14630 17196 -14596
rect 17230 -14630 17286 -14596
rect 17320 -14630 17376 -14596
rect 17410 -14630 17466 -14596
rect 17500 -14630 17559 -14596
rect 16865 -14648 17559 -14630
rect 16865 -14682 16938 -14648
rect 16972 -14682 17038 -14648
rect 17072 -14682 17138 -14648
rect 17172 -14682 17238 -14648
rect 17272 -14682 17338 -14648
rect 17372 -14682 17438 -14648
rect 17472 -14682 17559 -14648
rect 16865 -14686 17559 -14682
rect 16865 -14720 16926 -14686
rect 16960 -14720 17016 -14686
rect 17050 -14720 17106 -14686
rect 17140 -14720 17196 -14686
rect 17230 -14720 17286 -14686
rect 17320 -14720 17376 -14686
rect 17410 -14720 17466 -14686
rect 17500 -14720 17559 -14686
rect 16865 -14748 17559 -14720
rect 16865 -14776 16938 -14748
rect 16972 -14776 17038 -14748
rect 17072 -14776 17138 -14748
rect 17172 -14776 17238 -14748
rect 16865 -14810 16926 -14776
rect 16972 -14782 17016 -14776
rect 17072 -14782 17106 -14776
rect 17172 -14782 17196 -14776
rect 16960 -14810 17016 -14782
rect 17050 -14810 17106 -14782
rect 17140 -14810 17196 -14782
rect 17230 -14782 17238 -14776
rect 17272 -14776 17338 -14748
rect 17272 -14782 17286 -14776
rect 17230 -14810 17286 -14782
rect 17320 -14782 17338 -14776
rect 17372 -14776 17438 -14748
rect 17472 -14776 17559 -14748
rect 17372 -14782 17376 -14776
rect 17320 -14810 17376 -14782
rect 17410 -14782 17438 -14776
rect 17410 -14810 17466 -14782
rect 17500 -14810 17559 -14776
rect 16865 -14869 17559 -14810
rect 17621 -14206 17640 -14172
rect 17674 -14206 17693 -14172
rect 17621 -14262 17693 -14206
rect 17621 -14296 17640 -14262
rect 17674 -14296 17693 -14262
rect 17621 -14352 17693 -14296
rect 17621 -14386 17640 -14352
rect 17674 -14386 17693 -14352
rect 17621 -14442 17693 -14386
rect 17621 -14476 17640 -14442
rect 17674 -14476 17693 -14442
rect 17621 -14532 17693 -14476
rect 17621 -14566 17640 -14532
rect 17674 -14566 17693 -14532
rect 17621 -14622 17693 -14566
rect 17621 -14656 17640 -14622
rect 17674 -14656 17693 -14622
rect 17621 -14712 17693 -14656
rect 17621 -14746 17640 -14712
rect 17674 -14746 17693 -14712
rect 17621 -14802 17693 -14746
rect 17621 -14836 17640 -14802
rect 17674 -14836 17693 -14802
rect 16731 -14931 16803 -14892
rect 17621 -14892 17693 -14836
rect 17621 -14926 17640 -14892
rect 17674 -14926 17693 -14892
rect 17621 -14931 17693 -14926
rect 16731 -14950 17693 -14931
rect 16731 -14984 16844 -14950
rect 16878 -14984 16934 -14950
rect 16968 -14984 17024 -14950
rect 17058 -14984 17114 -14950
rect 17148 -14984 17204 -14950
rect 17238 -14984 17294 -14950
rect 17328 -14984 17384 -14950
rect 17418 -14984 17474 -14950
rect 17508 -14984 17564 -14950
rect 17598 -14984 17693 -14950
rect 16731 -15002 17693 -14984
rect 17757 -14132 17787 -14102
rect 17821 -14132 17888 -14098
rect 17922 -14102 19075 -14098
rect 17922 -14132 17955 -14102
rect 17757 -14188 17955 -14132
rect 17757 -14222 17787 -14188
rect 17821 -14222 17888 -14188
rect 17922 -14222 17955 -14188
rect 17757 -14278 17955 -14222
rect 17757 -14312 17787 -14278
rect 17821 -14312 17888 -14278
rect 17922 -14312 17955 -14278
rect 17757 -14368 17955 -14312
rect 17757 -14402 17787 -14368
rect 17821 -14402 17888 -14368
rect 17922 -14402 17955 -14368
rect 17757 -14458 17955 -14402
rect 17757 -14492 17787 -14458
rect 17821 -14492 17888 -14458
rect 17922 -14492 17955 -14458
rect 17757 -14548 17955 -14492
rect 17757 -14582 17787 -14548
rect 17821 -14582 17888 -14548
rect 17922 -14582 17955 -14548
rect 17757 -14638 17955 -14582
rect 17757 -14672 17787 -14638
rect 17821 -14672 17888 -14638
rect 17922 -14672 17955 -14638
rect 17757 -14728 17955 -14672
rect 17757 -14762 17787 -14728
rect 17821 -14762 17888 -14728
rect 17922 -14762 17955 -14728
rect 17757 -14818 17955 -14762
rect 17757 -14852 17787 -14818
rect 17821 -14852 17888 -14818
rect 17922 -14852 17955 -14818
rect 17757 -14908 17955 -14852
rect 17757 -14942 17787 -14908
rect 17821 -14942 17888 -14908
rect 17922 -14942 17955 -14908
rect 17757 -14998 17955 -14942
rect 17757 -15002 17787 -14998
rect 16634 -15032 17787 -15002
rect 17821 -15032 17888 -14998
rect 17922 -15002 17955 -14998
rect 18019 -14113 18981 -14102
rect 18019 -14138 18091 -14113
rect 18019 -14172 18038 -14138
rect 18072 -14172 18091 -14138
rect 18019 -14228 18091 -14172
rect 18909 -14172 18981 -14113
rect 18019 -14262 18038 -14228
rect 18072 -14262 18091 -14228
rect 18019 -14318 18091 -14262
rect 18019 -14352 18038 -14318
rect 18072 -14352 18091 -14318
rect 18019 -14408 18091 -14352
rect 18019 -14442 18038 -14408
rect 18072 -14442 18091 -14408
rect 18019 -14498 18091 -14442
rect 18019 -14532 18038 -14498
rect 18072 -14532 18091 -14498
rect 18019 -14588 18091 -14532
rect 18019 -14622 18038 -14588
rect 18072 -14622 18091 -14588
rect 18019 -14678 18091 -14622
rect 18019 -14712 18038 -14678
rect 18072 -14712 18091 -14678
rect 18019 -14768 18091 -14712
rect 18019 -14802 18038 -14768
rect 18072 -14802 18091 -14768
rect 18019 -14858 18091 -14802
rect 18019 -14892 18038 -14858
rect 18072 -14892 18091 -14858
rect 18153 -14236 18847 -14175
rect 18153 -14270 18214 -14236
rect 18248 -14248 18304 -14236
rect 18338 -14248 18394 -14236
rect 18428 -14248 18484 -14236
rect 18260 -14270 18304 -14248
rect 18360 -14270 18394 -14248
rect 18460 -14270 18484 -14248
rect 18518 -14248 18574 -14236
rect 18518 -14270 18526 -14248
rect 18153 -14282 18226 -14270
rect 18260 -14282 18326 -14270
rect 18360 -14282 18426 -14270
rect 18460 -14282 18526 -14270
rect 18560 -14270 18574 -14248
rect 18608 -14248 18664 -14236
rect 18608 -14270 18626 -14248
rect 18560 -14282 18626 -14270
rect 18660 -14270 18664 -14248
rect 18698 -14248 18754 -14236
rect 18698 -14270 18726 -14248
rect 18788 -14270 18847 -14236
rect 18660 -14282 18726 -14270
rect 18760 -14282 18847 -14270
rect 18153 -14326 18847 -14282
rect 18153 -14360 18214 -14326
rect 18248 -14348 18304 -14326
rect 18338 -14348 18394 -14326
rect 18428 -14348 18484 -14326
rect 18260 -14360 18304 -14348
rect 18360 -14360 18394 -14348
rect 18460 -14360 18484 -14348
rect 18518 -14348 18574 -14326
rect 18518 -14360 18526 -14348
rect 18153 -14382 18226 -14360
rect 18260 -14382 18326 -14360
rect 18360 -14382 18426 -14360
rect 18460 -14382 18526 -14360
rect 18560 -14360 18574 -14348
rect 18608 -14348 18664 -14326
rect 18608 -14360 18626 -14348
rect 18560 -14382 18626 -14360
rect 18660 -14360 18664 -14348
rect 18698 -14348 18754 -14326
rect 18698 -14360 18726 -14348
rect 18788 -14360 18847 -14326
rect 18660 -14382 18726 -14360
rect 18760 -14382 18847 -14360
rect 18153 -14416 18847 -14382
rect 18153 -14450 18214 -14416
rect 18248 -14448 18304 -14416
rect 18338 -14448 18394 -14416
rect 18428 -14448 18484 -14416
rect 18260 -14450 18304 -14448
rect 18360 -14450 18394 -14448
rect 18460 -14450 18484 -14448
rect 18518 -14448 18574 -14416
rect 18518 -14450 18526 -14448
rect 18153 -14482 18226 -14450
rect 18260 -14482 18326 -14450
rect 18360 -14482 18426 -14450
rect 18460 -14482 18526 -14450
rect 18560 -14450 18574 -14448
rect 18608 -14448 18664 -14416
rect 18608 -14450 18626 -14448
rect 18560 -14482 18626 -14450
rect 18660 -14450 18664 -14448
rect 18698 -14448 18754 -14416
rect 18698 -14450 18726 -14448
rect 18788 -14450 18847 -14416
rect 18660 -14482 18726 -14450
rect 18760 -14482 18847 -14450
rect 18153 -14506 18847 -14482
rect 18153 -14540 18214 -14506
rect 18248 -14540 18304 -14506
rect 18338 -14540 18394 -14506
rect 18428 -14540 18484 -14506
rect 18518 -14540 18574 -14506
rect 18608 -14540 18664 -14506
rect 18698 -14540 18754 -14506
rect 18788 -14540 18847 -14506
rect 18153 -14548 18847 -14540
rect 18153 -14582 18226 -14548
rect 18260 -14582 18326 -14548
rect 18360 -14582 18426 -14548
rect 18460 -14582 18526 -14548
rect 18560 -14582 18626 -14548
rect 18660 -14582 18726 -14548
rect 18760 -14582 18847 -14548
rect 18153 -14596 18847 -14582
rect 18153 -14630 18214 -14596
rect 18248 -14630 18304 -14596
rect 18338 -14630 18394 -14596
rect 18428 -14630 18484 -14596
rect 18518 -14630 18574 -14596
rect 18608 -14630 18664 -14596
rect 18698 -14630 18754 -14596
rect 18788 -14630 18847 -14596
rect 18153 -14648 18847 -14630
rect 18153 -14682 18226 -14648
rect 18260 -14682 18326 -14648
rect 18360 -14682 18426 -14648
rect 18460 -14682 18526 -14648
rect 18560 -14682 18626 -14648
rect 18660 -14682 18726 -14648
rect 18760 -14682 18847 -14648
rect 18153 -14686 18847 -14682
rect 18153 -14720 18214 -14686
rect 18248 -14720 18304 -14686
rect 18338 -14720 18394 -14686
rect 18428 -14720 18484 -14686
rect 18518 -14720 18574 -14686
rect 18608 -14720 18664 -14686
rect 18698 -14720 18754 -14686
rect 18788 -14720 18847 -14686
rect 18153 -14748 18847 -14720
rect 18153 -14776 18226 -14748
rect 18260 -14776 18326 -14748
rect 18360 -14776 18426 -14748
rect 18460 -14776 18526 -14748
rect 18153 -14810 18214 -14776
rect 18260 -14782 18304 -14776
rect 18360 -14782 18394 -14776
rect 18460 -14782 18484 -14776
rect 18248 -14810 18304 -14782
rect 18338 -14810 18394 -14782
rect 18428 -14810 18484 -14782
rect 18518 -14782 18526 -14776
rect 18560 -14776 18626 -14748
rect 18560 -14782 18574 -14776
rect 18518 -14810 18574 -14782
rect 18608 -14782 18626 -14776
rect 18660 -14776 18726 -14748
rect 18760 -14776 18847 -14748
rect 18660 -14782 18664 -14776
rect 18608 -14810 18664 -14782
rect 18698 -14782 18726 -14776
rect 18698 -14810 18754 -14782
rect 18788 -14810 18847 -14776
rect 18153 -14869 18847 -14810
rect 18909 -14206 18928 -14172
rect 18962 -14206 18981 -14172
rect 18909 -14262 18981 -14206
rect 18909 -14296 18928 -14262
rect 18962 -14296 18981 -14262
rect 18909 -14352 18981 -14296
rect 18909 -14386 18928 -14352
rect 18962 -14386 18981 -14352
rect 18909 -14442 18981 -14386
rect 18909 -14476 18928 -14442
rect 18962 -14476 18981 -14442
rect 18909 -14532 18981 -14476
rect 18909 -14566 18928 -14532
rect 18962 -14566 18981 -14532
rect 18909 -14622 18981 -14566
rect 18909 -14656 18928 -14622
rect 18962 -14656 18981 -14622
rect 18909 -14712 18981 -14656
rect 18909 -14746 18928 -14712
rect 18962 -14746 18981 -14712
rect 18909 -14802 18981 -14746
rect 18909 -14836 18928 -14802
rect 18962 -14836 18981 -14802
rect 18019 -14931 18091 -14892
rect 18909 -14892 18981 -14836
rect 18909 -14926 18928 -14892
rect 18962 -14926 18981 -14892
rect 18909 -14931 18981 -14926
rect 18019 -14950 18981 -14931
rect 18019 -14984 18132 -14950
rect 18166 -14984 18222 -14950
rect 18256 -14984 18312 -14950
rect 18346 -14984 18402 -14950
rect 18436 -14984 18492 -14950
rect 18526 -14984 18582 -14950
rect 18616 -14984 18672 -14950
rect 18706 -14984 18762 -14950
rect 18796 -14984 18852 -14950
rect 18886 -14984 18981 -14950
rect 18019 -15002 18981 -14984
rect 19045 -14132 19075 -14102
rect 19109 -14132 19176 -14098
rect 19210 -14102 20363 -14098
rect 19210 -14132 19243 -14102
rect 19045 -14188 19243 -14132
rect 19045 -14222 19075 -14188
rect 19109 -14222 19176 -14188
rect 19210 -14222 19243 -14188
rect 19045 -14278 19243 -14222
rect 19045 -14312 19075 -14278
rect 19109 -14312 19176 -14278
rect 19210 -14312 19243 -14278
rect 19045 -14368 19243 -14312
rect 19045 -14402 19075 -14368
rect 19109 -14402 19176 -14368
rect 19210 -14402 19243 -14368
rect 19045 -14458 19243 -14402
rect 19045 -14492 19075 -14458
rect 19109 -14492 19176 -14458
rect 19210 -14492 19243 -14458
rect 19045 -14548 19243 -14492
rect 19045 -14582 19075 -14548
rect 19109 -14582 19176 -14548
rect 19210 -14582 19243 -14548
rect 19045 -14638 19243 -14582
rect 19045 -14672 19075 -14638
rect 19109 -14672 19176 -14638
rect 19210 -14672 19243 -14638
rect 19045 -14728 19243 -14672
rect 19045 -14762 19075 -14728
rect 19109 -14762 19176 -14728
rect 19210 -14762 19243 -14728
rect 19045 -14818 19243 -14762
rect 19045 -14852 19075 -14818
rect 19109 -14852 19176 -14818
rect 19210 -14852 19243 -14818
rect 19045 -14908 19243 -14852
rect 19045 -14942 19075 -14908
rect 19109 -14942 19176 -14908
rect 19210 -14942 19243 -14908
rect 19045 -14998 19243 -14942
rect 19045 -15002 19075 -14998
rect 17922 -15032 19075 -15002
rect 19109 -15032 19176 -14998
rect 19210 -15002 19243 -14998
rect 19307 -14113 20269 -14102
rect 19307 -14138 19379 -14113
rect 19307 -14172 19326 -14138
rect 19360 -14172 19379 -14138
rect 19307 -14228 19379 -14172
rect 20197 -14172 20269 -14113
rect 19307 -14262 19326 -14228
rect 19360 -14262 19379 -14228
rect 19307 -14318 19379 -14262
rect 19307 -14352 19326 -14318
rect 19360 -14352 19379 -14318
rect 19307 -14408 19379 -14352
rect 19307 -14442 19326 -14408
rect 19360 -14442 19379 -14408
rect 19307 -14498 19379 -14442
rect 19307 -14532 19326 -14498
rect 19360 -14532 19379 -14498
rect 19307 -14588 19379 -14532
rect 19307 -14622 19326 -14588
rect 19360 -14622 19379 -14588
rect 19307 -14678 19379 -14622
rect 19307 -14712 19326 -14678
rect 19360 -14712 19379 -14678
rect 19307 -14768 19379 -14712
rect 19307 -14802 19326 -14768
rect 19360 -14802 19379 -14768
rect 19307 -14858 19379 -14802
rect 19307 -14892 19326 -14858
rect 19360 -14892 19379 -14858
rect 19441 -14236 20135 -14175
rect 19441 -14270 19502 -14236
rect 19536 -14248 19592 -14236
rect 19626 -14248 19682 -14236
rect 19716 -14248 19772 -14236
rect 19548 -14270 19592 -14248
rect 19648 -14270 19682 -14248
rect 19748 -14270 19772 -14248
rect 19806 -14248 19862 -14236
rect 19806 -14270 19814 -14248
rect 19441 -14282 19514 -14270
rect 19548 -14282 19614 -14270
rect 19648 -14282 19714 -14270
rect 19748 -14282 19814 -14270
rect 19848 -14270 19862 -14248
rect 19896 -14248 19952 -14236
rect 19896 -14270 19914 -14248
rect 19848 -14282 19914 -14270
rect 19948 -14270 19952 -14248
rect 19986 -14248 20042 -14236
rect 19986 -14270 20014 -14248
rect 20076 -14270 20135 -14236
rect 19948 -14282 20014 -14270
rect 20048 -14282 20135 -14270
rect 19441 -14326 20135 -14282
rect 19441 -14360 19502 -14326
rect 19536 -14348 19592 -14326
rect 19626 -14348 19682 -14326
rect 19716 -14348 19772 -14326
rect 19548 -14360 19592 -14348
rect 19648 -14360 19682 -14348
rect 19748 -14360 19772 -14348
rect 19806 -14348 19862 -14326
rect 19806 -14360 19814 -14348
rect 19441 -14382 19514 -14360
rect 19548 -14382 19614 -14360
rect 19648 -14382 19714 -14360
rect 19748 -14382 19814 -14360
rect 19848 -14360 19862 -14348
rect 19896 -14348 19952 -14326
rect 19896 -14360 19914 -14348
rect 19848 -14382 19914 -14360
rect 19948 -14360 19952 -14348
rect 19986 -14348 20042 -14326
rect 19986 -14360 20014 -14348
rect 20076 -14360 20135 -14326
rect 19948 -14382 20014 -14360
rect 20048 -14382 20135 -14360
rect 19441 -14416 20135 -14382
rect 19441 -14450 19502 -14416
rect 19536 -14448 19592 -14416
rect 19626 -14448 19682 -14416
rect 19716 -14448 19772 -14416
rect 19548 -14450 19592 -14448
rect 19648 -14450 19682 -14448
rect 19748 -14450 19772 -14448
rect 19806 -14448 19862 -14416
rect 19806 -14450 19814 -14448
rect 19441 -14482 19514 -14450
rect 19548 -14482 19614 -14450
rect 19648 -14482 19714 -14450
rect 19748 -14482 19814 -14450
rect 19848 -14450 19862 -14448
rect 19896 -14448 19952 -14416
rect 19896 -14450 19914 -14448
rect 19848 -14482 19914 -14450
rect 19948 -14450 19952 -14448
rect 19986 -14448 20042 -14416
rect 19986 -14450 20014 -14448
rect 20076 -14450 20135 -14416
rect 19948 -14482 20014 -14450
rect 20048 -14482 20135 -14450
rect 19441 -14506 20135 -14482
rect 19441 -14540 19502 -14506
rect 19536 -14540 19592 -14506
rect 19626 -14540 19682 -14506
rect 19716 -14540 19772 -14506
rect 19806 -14540 19862 -14506
rect 19896 -14540 19952 -14506
rect 19986 -14540 20042 -14506
rect 20076 -14540 20135 -14506
rect 19441 -14548 20135 -14540
rect 19441 -14582 19514 -14548
rect 19548 -14582 19614 -14548
rect 19648 -14582 19714 -14548
rect 19748 -14582 19814 -14548
rect 19848 -14582 19914 -14548
rect 19948 -14582 20014 -14548
rect 20048 -14582 20135 -14548
rect 19441 -14596 20135 -14582
rect 19441 -14630 19502 -14596
rect 19536 -14630 19592 -14596
rect 19626 -14630 19682 -14596
rect 19716 -14630 19772 -14596
rect 19806 -14630 19862 -14596
rect 19896 -14630 19952 -14596
rect 19986 -14630 20042 -14596
rect 20076 -14630 20135 -14596
rect 19441 -14648 20135 -14630
rect 19441 -14682 19514 -14648
rect 19548 -14682 19614 -14648
rect 19648 -14682 19714 -14648
rect 19748 -14682 19814 -14648
rect 19848 -14682 19914 -14648
rect 19948 -14682 20014 -14648
rect 20048 -14682 20135 -14648
rect 19441 -14686 20135 -14682
rect 19441 -14720 19502 -14686
rect 19536 -14720 19592 -14686
rect 19626 -14720 19682 -14686
rect 19716 -14720 19772 -14686
rect 19806 -14720 19862 -14686
rect 19896 -14720 19952 -14686
rect 19986 -14720 20042 -14686
rect 20076 -14720 20135 -14686
rect 19441 -14748 20135 -14720
rect 19441 -14776 19514 -14748
rect 19548 -14776 19614 -14748
rect 19648 -14776 19714 -14748
rect 19748 -14776 19814 -14748
rect 19441 -14810 19502 -14776
rect 19548 -14782 19592 -14776
rect 19648 -14782 19682 -14776
rect 19748 -14782 19772 -14776
rect 19536 -14810 19592 -14782
rect 19626 -14810 19682 -14782
rect 19716 -14810 19772 -14782
rect 19806 -14782 19814 -14776
rect 19848 -14776 19914 -14748
rect 19848 -14782 19862 -14776
rect 19806 -14810 19862 -14782
rect 19896 -14782 19914 -14776
rect 19948 -14776 20014 -14748
rect 20048 -14776 20135 -14748
rect 19948 -14782 19952 -14776
rect 19896 -14810 19952 -14782
rect 19986 -14782 20014 -14776
rect 19986 -14810 20042 -14782
rect 20076 -14810 20135 -14776
rect 19441 -14869 20135 -14810
rect 20197 -14206 20216 -14172
rect 20250 -14206 20269 -14172
rect 20197 -14262 20269 -14206
rect 20197 -14296 20216 -14262
rect 20250 -14296 20269 -14262
rect 20197 -14352 20269 -14296
rect 20197 -14386 20216 -14352
rect 20250 -14386 20269 -14352
rect 20197 -14442 20269 -14386
rect 20197 -14476 20216 -14442
rect 20250 -14476 20269 -14442
rect 20197 -14532 20269 -14476
rect 20197 -14566 20216 -14532
rect 20250 -14566 20269 -14532
rect 20197 -14622 20269 -14566
rect 20197 -14656 20216 -14622
rect 20250 -14656 20269 -14622
rect 20197 -14712 20269 -14656
rect 20197 -14746 20216 -14712
rect 20250 -14746 20269 -14712
rect 20197 -14802 20269 -14746
rect 20197 -14836 20216 -14802
rect 20250 -14836 20269 -14802
rect 19307 -14931 19379 -14892
rect 20197 -14892 20269 -14836
rect 20197 -14926 20216 -14892
rect 20250 -14926 20269 -14892
rect 20197 -14931 20269 -14926
rect 19307 -14950 20269 -14931
rect 19307 -14984 19420 -14950
rect 19454 -14984 19510 -14950
rect 19544 -14984 19600 -14950
rect 19634 -14984 19690 -14950
rect 19724 -14984 19780 -14950
rect 19814 -14984 19870 -14950
rect 19904 -14984 19960 -14950
rect 19994 -14984 20050 -14950
rect 20084 -14984 20140 -14950
rect 20174 -14984 20269 -14950
rect 19307 -15002 20269 -14984
rect 20333 -14132 20363 -14102
rect 20397 -14132 20464 -14098
rect 20498 -14102 21651 -14098
rect 20498 -14132 20531 -14102
rect 20333 -14188 20531 -14132
rect 20333 -14222 20363 -14188
rect 20397 -14222 20464 -14188
rect 20498 -14222 20531 -14188
rect 20333 -14278 20531 -14222
rect 20333 -14312 20363 -14278
rect 20397 -14312 20464 -14278
rect 20498 -14312 20531 -14278
rect 20333 -14368 20531 -14312
rect 20333 -14402 20363 -14368
rect 20397 -14402 20464 -14368
rect 20498 -14402 20531 -14368
rect 20333 -14458 20531 -14402
rect 20333 -14492 20363 -14458
rect 20397 -14492 20464 -14458
rect 20498 -14492 20531 -14458
rect 20333 -14548 20531 -14492
rect 20333 -14582 20363 -14548
rect 20397 -14582 20464 -14548
rect 20498 -14582 20531 -14548
rect 20333 -14638 20531 -14582
rect 20333 -14672 20363 -14638
rect 20397 -14672 20464 -14638
rect 20498 -14672 20531 -14638
rect 20333 -14728 20531 -14672
rect 20333 -14762 20363 -14728
rect 20397 -14762 20464 -14728
rect 20498 -14762 20531 -14728
rect 20333 -14818 20531 -14762
rect 20333 -14852 20363 -14818
rect 20397 -14852 20464 -14818
rect 20498 -14852 20531 -14818
rect 20333 -14908 20531 -14852
rect 20333 -14942 20363 -14908
rect 20397 -14942 20464 -14908
rect 20498 -14942 20531 -14908
rect 20333 -14998 20531 -14942
rect 20333 -15002 20363 -14998
rect 19210 -15032 20363 -15002
rect 20397 -15032 20464 -14998
rect 20498 -15002 20531 -14998
rect 20595 -14113 21557 -14102
rect 20595 -14138 20667 -14113
rect 20595 -14172 20614 -14138
rect 20648 -14172 20667 -14138
rect 20595 -14228 20667 -14172
rect 21485 -14172 21557 -14113
rect 20595 -14262 20614 -14228
rect 20648 -14262 20667 -14228
rect 20595 -14318 20667 -14262
rect 20595 -14352 20614 -14318
rect 20648 -14352 20667 -14318
rect 20595 -14408 20667 -14352
rect 20595 -14442 20614 -14408
rect 20648 -14442 20667 -14408
rect 20595 -14498 20667 -14442
rect 20595 -14532 20614 -14498
rect 20648 -14532 20667 -14498
rect 20595 -14588 20667 -14532
rect 20595 -14622 20614 -14588
rect 20648 -14622 20667 -14588
rect 20595 -14678 20667 -14622
rect 20595 -14712 20614 -14678
rect 20648 -14712 20667 -14678
rect 20595 -14768 20667 -14712
rect 20595 -14802 20614 -14768
rect 20648 -14802 20667 -14768
rect 20595 -14858 20667 -14802
rect 20595 -14892 20614 -14858
rect 20648 -14892 20667 -14858
rect 20729 -14236 21423 -14175
rect 20729 -14270 20790 -14236
rect 20824 -14248 20880 -14236
rect 20914 -14248 20970 -14236
rect 21004 -14248 21060 -14236
rect 20836 -14270 20880 -14248
rect 20936 -14270 20970 -14248
rect 21036 -14270 21060 -14248
rect 21094 -14248 21150 -14236
rect 21094 -14270 21102 -14248
rect 20729 -14282 20802 -14270
rect 20836 -14282 20902 -14270
rect 20936 -14282 21002 -14270
rect 21036 -14282 21102 -14270
rect 21136 -14270 21150 -14248
rect 21184 -14248 21240 -14236
rect 21184 -14270 21202 -14248
rect 21136 -14282 21202 -14270
rect 21236 -14270 21240 -14248
rect 21274 -14248 21330 -14236
rect 21274 -14270 21302 -14248
rect 21364 -14270 21423 -14236
rect 21236 -14282 21302 -14270
rect 21336 -14282 21423 -14270
rect 20729 -14326 21423 -14282
rect 20729 -14360 20790 -14326
rect 20824 -14348 20880 -14326
rect 20914 -14348 20970 -14326
rect 21004 -14348 21060 -14326
rect 20836 -14360 20880 -14348
rect 20936 -14360 20970 -14348
rect 21036 -14360 21060 -14348
rect 21094 -14348 21150 -14326
rect 21094 -14360 21102 -14348
rect 20729 -14382 20802 -14360
rect 20836 -14382 20902 -14360
rect 20936 -14382 21002 -14360
rect 21036 -14382 21102 -14360
rect 21136 -14360 21150 -14348
rect 21184 -14348 21240 -14326
rect 21184 -14360 21202 -14348
rect 21136 -14382 21202 -14360
rect 21236 -14360 21240 -14348
rect 21274 -14348 21330 -14326
rect 21274 -14360 21302 -14348
rect 21364 -14360 21423 -14326
rect 21236 -14382 21302 -14360
rect 21336 -14382 21423 -14360
rect 20729 -14416 21423 -14382
rect 20729 -14450 20790 -14416
rect 20824 -14448 20880 -14416
rect 20914 -14448 20970 -14416
rect 21004 -14448 21060 -14416
rect 20836 -14450 20880 -14448
rect 20936 -14450 20970 -14448
rect 21036 -14450 21060 -14448
rect 21094 -14448 21150 -14416
rect 21094 -14450 21102 -14448
rect 20729 -14482 20802 -14450
rect 20836 -14482 20902 -14450
rect 20936 -14482 21002 -14450
rect 21036 -14482 21102 -14450
rect 21136 -14450 21150 -14448
rect 21184 -14448 21240 -14416
rect 21184 -14450 21202 -14448
rect 21136 -14482 21202 -14450
rect 21236 -14450 21240 -14448
rect 21274 -14448 21330 -14416
rect 21274 -14450 21302 -14448
rect 21364 -14450 21423 -14416
rect 21236 -14482 21302 -14450
rect 21336 -14482 21423 -14450
rect 20729 -14506 21423 -14482
rect 20729 -14540 20790 -14506
rect 20824 -14540 20880 -14506
rect 20914 -14540 20970 -14506
rect 21004 -14540 21060 -14506
rect 21094 -14540 21150 -14506
rect 21184 -14540 21240 -14506
rect 21274 -14540 21330 -14506
rect 21364 -14540 21423 -14506
rect 20729 -14548 21423 -14540
rect 20729 -14582 20802 -14548
rect 20836 -14582 20902 -14548
rect 20936 -14582 21002 -14548
rect 21036 -14582 21102 -14548
rect 21136 -14582 21202 -14548
rect 21236 -14582 21302 -14548
rect 21336 -14582 21423 -14548
rect 20729 -14596 21423 -14582
rect 20729 -14630 20790 -14596
rect 20824 -14630 20880 -14596
rect 20914 -14630 20970 -14596
rect 21004 -14630 21060 -14596
rect 21094 -14630 21150 -14596
rect 21184 -14630 21240 -14596
rect 21274 -14630 21330 -14596
rect 21364 -14630 21423 -14596
rect 20729 -14648 21423 -14630
rect 20729 -14682 20802 -14648
rect 20836 -14682 20902 -14648
rect 20936 -14682 21002 -14648
rect 21036 -14682 21102 -14648
rect 21136 -14682 21202 -14648
rect 21236 -14682 21302 -14648
rect 21336 -14682 21423 -14648
rect 20729 -14686 21423 -14682
rect 20729 -14720 20790 -14686
rect 20824 -14720 20880 -14686
rect 20914 -14720 20970 -14686
rect 21004 -14720 21060 -14686
rect 21094 -14720 21150 -14686
rect 21184 -14720 21240 -14686
rect 21274 -14720 21330 -14686
rect 21364 -14720 21423 -14686
rect 20729 -14748 21423 -14720
rect 20729 -14776 20802 -14748
rect 20836 -14776 20902 -14748
rect 20936 -14776 21002 -14748
rect 21036 -14776 21102 -14748
rect 20729 -14810 20790 -14776
rect 20836 -14782 20880 -14776
rect 20936 -14782 20970 -14776
rect 21036 -14782 21060 -14776
rect 20824 -14810 20880 -14782
rect 20914 -14810 20970 -14782
rect 21004 -14810 21060 -14782
rect 21094 -14782 21102 -14776
rect 21136 -14776 21202 -14748
rect 21136 -14782 21150 -14776
rect 21094 -14810 21150 -14782
rect 21184 -14782 21202 -14776
rect 21236 -14776 21302 -14748
rect 21336 -14776 21423 -14748
rect 21236 -14782 21240 -14776
rect 21184 -14810 21240 -14782
rect 21274 -14782 21302 -14776
rect 21274 -14810 21330 -14782
rect 21364 -14810 21423 -14776
rect 20729 -14869 21423 -14810
rect 21485 -14206 21504 -14172
rect 21538 -14206 21557 -14172
rect 21485 -14262 21557 -14206
rect 21485 -14296 21504 -14262
rect 21538 -14296 21557 -14262
rect 21485 -14352 21557 -14296
rect 21485 -14386 21504 -14352
rect 21538 -14386 21557 -14352
rect 21485 -14442 21557 -14386
rect 21485 -14476 21504 -14442
rect 21538 -14476 21557 -14442
rect 21485 -14532 21557 -14476
rect 21485 -14566 21504 -14532
rect 21538 -14566 21557 -14532
rect 21485 -14622 21557 -14566
rect 21485 -14656 21504 -14622
rect 21538 -14656 21557 -14622
rect 21485 -14712 21557 -14656
rect 21485 -14746 21504 -14712
rect 21538 -14746 21557 -14712
rect 21485 -14802 21557 -14746
rect 21485 -14836 21504 -14802
rect 21538 -14836 21557 -14802
rect 20595 -14931 20667 -14892
rect 21485 -14892 21557 -14836
rect 21485 -14926 21504 -14892
rect 21538 -14926 21557 -14892
rect 21485 -14931 21557 -14926
rect 20595 -14950 21557 -14931
rect 20595 -14984 20708 -14950
rect 20742 -14984 20798 -14950
rect 20832 -14984 20888 -14950
rect 20922 -14984 20978 -14950
rect 21012 -14984 21068 -14950
rect 21102 -14984 21158 -14950
rect 21192 -14984 21248 -14950
rect 21282 -14984 21338 -14950
rect 21372 -14984 21428 -14950
rect 21462 -14984 21557 -14950
rect 20595 -15002 21557 -14984
rect 21621 -14132 21651 -14102
rect 21685 -14132 21752 -14098
rect 21786 -14102 22939 -14098
rect 21786 -14132 21819 -14102
rect 21621 -14188 21819 -14132
rect 21621 -14222 21651 -14188
rect 21685 -14222 21752 -14188
rect 21786 -14222 21819 -14188
rect 21621 -14278 21819 -14222
rect 21621 -14312 21651 -14278
rect 21685 -14312 21752 -14278
rect 21786 -14312 21819 -14278
rect 21621 -14368 21819 -14312
rect 21621 -14402 21651 -14368
rect 21685 -14402 21752 -14368
rect 21786 -14402 21819 -14368
rect 21621 -14458 21819 -14402
rect 21621 -14492 21651 -14458
rect 21685 -14492 21752 -14458
rect 21786 -14492 21819 -14458
rect 21621 -14548 21819 -14492
rect 21621 -14582 21651 -14548
rect 21685 -14582 21752 -14548
rect 21786 -14582 21819 -14548
rect 21621 -14638 21819 -14582
rect 21621 -14672 21651 -14638
rect 21685 -14672 21752 -14638
rect 21786 -14672 21819 -14638
rect 21621 -14728 21819 -14672
rect 21621 -14762 21651 -14728
rect 21685 -14762 21752 -14728
rect 21786 -14762 21819 -14728
rect 21621 -14818 21819 -14762
rect 21621 -14852 21651 -14818
rect 21685 -14852 21752 -14818
rect 21786 -14852 21819 -14818
rect 21621 -14908 21819 -14852
rect 21621 -14942 21651 -14908
rect 21685 -14942 21752 -14908
rect 21786 -14942 21819 -14908
rect 21621 -14998 21819 -14942
rect 21621 -15002 21651 -14998
rect 20498 -15032 21651 -15002
rect 21685 -15032 21752 -14998
rect 21786 -15002 21819 -14998
rect 21883 -14113 22845 -14102
rect 21883 -14138 21955 -14113
rect 21883 -14172 21902 -14138
rect 21936 -14172 21955 -14138
rect 21883 -14228 21955 -14172
rect 22773 -14172 22845 -14113
rect 21883 -14262 21902 -14228
rect 21936 -14262 21955 -14228
rect 21883 -14318 21955 -14262
rect 21883 -14352 21902 -14318
rect 21936 -14352 21955 -14318
rect 21883 -14408 21955 -14352
rect 21883 -14442 21902 -14408
rect 21936 -14442 21955 -14408
rect 21883 -14498 21955 -14442
rect 21883 -14532 21902 -14498
rect 21936 -14532 21955 -14498
rect 21883 -14588 21955 -14532
rect 21883 -14622 21902 -14588
rect 21936 -14622 21955 -14588
rect 21883 -14678 21955 -14622
rect 21883 -14712 21902 -14678
rect 21936 -14712 21955 -14678
rect 21883 -14768 21955 -14712
rect 21883 -14802 21902 -14768
rect 21936 -14802 21955 -14768
rect 21883 -14858 21955 -14802
rect 21883 -14892 21902 -14858
rect 21936 -14892 21955 -14858
rect 22017 -14236 22711 -14175
rect 22017 -14270 22078 -14236
rect 22112 -14248 22168 -14236
rect 22202 -14248 22258 -14236
rect 22292 -14248 22348 -14236
rect 22124 -14270 22168 -14248
rect 22224 -14270 22258 -14248
rect 22324 -14270 22348 -14248
rect 22382 -14248 22438 -14236
rect 22382 -14270 22390 -14248
rect 22017 -14282 22090 -14270
rect 22124 -14282 22190 -14270
rect 22224 -14282 22290 -14270
rect 22324 -14282 22390 -14270
rect 22424 -14270 22438 -14248
rect 22472 -14248 22528 -14236
rect 22472 -14270 22490 -14248
rect 22424 -14282 22490 -14270
rect 22524 -14270 22528 -14248
rect 22562 -14248 22618 -14236
rect 22562 -14270 22590 -14248
rect 22652 -14270 22711 -14236
rect 22524 -14282 22590 -14270
rect 22624 -14282 22711 -14270
rect 22017 -14326 22711 -14282
rect 22017 -14360 22078 -14326
rect 22112 -14348 22168 -14326
rect 22202 -14348 22258 -14326
rect 22292 -14348 22348 -14326
rect 22124 -14360 22168 -14348
rect 22224 -14360 22258 -14348
rect 22324 -14360 22348 -14348
rect 22382 -14348 22438 -14326
rect 22382 -14360 22390 -14348
rect 22017 -14382 22090 -14360
rect 22124 -14382 22190 -14360
rect 22224 -14382 22290 -14360
rect 22324 -14382 22390 -14360
rect 22424 -14360 22438 -14348
rect 22472 -14348 22528 -14326
rect 22472 -14360 22490 -14348
rect 22424 -14382 22490 -14360
rect 22524 -14360 22528 -14348
rect 22562 -14348 22618 -14326
rect 22562 -14360 22590 -14348
rect 22652 -14360 22711 -14326
rect 22524 -14382 22590 -14360
rect 22624 -14382 22711 -14360
rect 22017 -14416 22711 -14382
rect 22017 -14450 22078 -14416
rect 22112 -14448 22168 -14416
rect 22202 -14448 22258 -14416
rect 22292 -14448 22348 -14416
rect 22124 -14450 22168 -14448
rect 22224 -14450 22258 -14448
rect 22324 -14450 22348 -14448
rect 22382 -14448 22438 -14416
rect 22382 -14450 22390 -14448
rect 22017 -14482 22090 -14450
rect 22124 -14482 22190 -14450
rect 22224 -14482 22290 -14450
rect 22324 -14482 22390 -14450
rect 22424 -14450 22438 -14448
rect 22472 -14448 22528 -14416
rect 22472 -14450 22490 -14448
rect 22424 -14482 22490 -14450
rect 22524 -14450 22528 -14448
rect 22562 -14448 22618 -14416
rect 22562 -14450 22590 -14448
rect 22652 -14450 22711 -14416
rect 22524 -14482 22590 -14450
rect 22624 -14482 22711 -14450
rect 22017 -14506 22711 -14482
rect 22017 -14540 22078 -14506
rect 22112 -14540 22168 -14506
rect 22202 -14540 22258 -14506
rect 22292 -14540 22348 -14506
rect 22382 -14540 22438 -14506
rect 22472 -14540 22528 -14506
rect 22562 -14540 22618 -14506
rect 22652 -14540 22711 -14506
rect 22017 -14548 22711 -14540
rect 22017 -14582 22090 -14548
rect 22124 -14582 22190 -14548
rect 22224 -14582 22290 -14548
rect 22324 -14582 22390 -14548
rect 22424 -14582 22490 -14548
rect 22524 -14582 22590 -14548
rect 22624 -14582 22711 -14548
rect 22017 -14596 22711 -14582
rect 22017 -14630 22078 -14596
rect 22112 -14630 22168 -14596
rect 22202 -14630 22258 -14596
rect 22292 -14630 22348 -14596
rect 22382 -14630 22438 -14596
rect 22472 -14630 22528 -14596
rect 22562 -14630 22618 -14596
rect 22652 -14630 22711 -14596
rect 22017 -14648 22711 -14630
rect 22017 -14682 22090 -14648
rect 22124 -14682 22190 -14648
rect 22224 -14682 22290 -14648
rect 22324 -14682 22390 -14648
rect 22424 -14682 22490 -14648
rect 22524 -14682 22590 -14648
rect 22624 -14682 22711 -14648
rect 22017 -14686 22711 -14682
rect 22017 -14720 22078 -14686
rect 22112 -14720 22168 -14686
rect 22202 -14720 22258 -14686
rect 22292 -14720 22348 -14686
rect 22382 -14720 22438 -14686
rect 22472 -14720 22528 -14686
rect 22562 -14720 22618 -14686
rect 22652 -14720 22711 -14686
rect 22017 -14748 22711 -14720
rect 22017 -14776 22090 -14748
rect 22124 -14776 22190 -14748
rect 22224 -14776 22290 -14748
rect 22324 -14776 22390 -14748
rect 22017 -14810 22078 -14776
rect 22124 -14782 22168 -14776
rect 22224 -14782 22258 -14776
rect 22324 -14782 22348 -14776
rect 22112 -14810 22168 -14782
rect 22202 -14810 22258 -14782
rect 22292 -14810 22348 -14782
rect 22382 -14782 22390 -14776
rect 22424 -14776 22490 -14748
rect 22424 -14782 22438 -14776
rect 22382 -14810 22438 -14782
rect 22472 -14782 22490 -14776
rect 22524 -14776 22590 -14748
rect 22624 -14776 22711 -14748
rect 22524 -14782 22528 -14776
rect 22472 -14810 22528 -14782
rect 22562 -14782 22590 -14776
rect 22562 -14810 22618 -14782
rect 22652 -14810 22711 -14776
rect 22017 -14869 22711 -14810
rect 22773 -14206 22792 -14172
rect 22826 -14206 22845 -14172
rect 22773 -14262 22845 -14206
rect 22773 -14296 22792 -14262
rect 22826 -14296 22845 -14262
rect 22773 -14352 22845 -14296
rect 22773 -14386 22792 -14352
rect 22826 -14386 22845 -14352
rect 22773 -14442 22845 -14386
rect 22773 -14476 22792 -14442
rect 22826 -14476 22845 -14442
rect 22773 -14532 22845 -14476
rect 22773 -14566 22792 -14532
rect 22826 -14566 22845 -14532
rect 22773 -14622 22845 -14566
rect 22773 -14656 22792 -14622
rect 22826 -14656 22845 -14622
rect 22773 -14712 22845 -14656
rect 22773 -14746 22792 -14712
rect 22826 -14746 22845 -14712
rect 22773 -14802 22845 -14746
rect 22773 -14836 22792 -14802
rect 22826 -14836 22845 -14802
rect 21883 -14931 21955 -14892
rect 22773 -14892 22845 -14836
rect 22773 -14926 22792 -14892
rect 22826 -14926 22845 -14892
rect 22773 -14931 22845 -14926
rect 21883 -14950 22845 -14931
rect 21883 -14984 21996 -14950
rect 22030 -14984 22086 -14950
rect 22120 -14984 22176 -14950
rect 22210 -14984 22266 -14950
rect 22300 -14984 22356 -14950
rect 22390 -14984 22446 -14950
rect 22480 -14984 22536 -14950
rect 22570 -14984 22626 -14950
rect 22660 -14984 22716 -14950
rect 22750 -14984 22845 -14950
rect 21883 -15002 22845 -14984
rect 22909 -14132 22939 -14102
rect 22973 -14132 23040 -14098
rect 23074 -14102 24227 -14098
rect 23074 -14132 23107 -14102
rect 22909 -14188 23107 -14132
rect 22909 -14222 22939 -14188
rect 22973 -14222 23040 -14188
rect 23074 -14222 23107 -14188
rect 22909 -14278 23107 -14222
rect 22909 -14312 22939 -14278
rect 22973 -14312 23040 -14278
rect 23074 -14312 23107 -14278
rect 22909 -14368 23107 -14312
rect 22909 -14402 22939 -14368
rect 22973 -14402 23040 -14368
rect 23074 -14402 23107 -14368
rect 22909 -14458 23107 -14402
rect 22909 -14492 22939 -14458
rect 22973 -14492 23040 -14458
rect 23074 -14492 23107 -14458
rect 22909 -14548 23107 -14492
rect 22909 -14582 22939 -14548
rect 22973 -14582 23040 -14548
rect 23074 -14582 23107 -14548
rect 22909 -14638 23107 -14582
rect 22909 -14672 22939 -14638
rect 22973 -14672 23040 -14638
rect 23074 -14672 23107 -14638
rect 22909 -14728 23107 -14672
rect 22909 -14762 22939 -14728
rect 22973 -14762 23040 -14728
rect 23074 -14762 23107 -14728
rect 22909 -14818 23107 -14762
rect 22909 -14852 22939 -14818
rect 22973 -14852 23040 -14818
rect 23074 -14852 23107 -14818
rect 22909 -14908 23107 -14852
rect 22909 -14942 22939 -14908
rect 22973 -14942 23040 -14908
rect 23074 -14942 23107 -14908
rect 22909 -14998 23107 -14942
rect 22909 -15002 22939 -14998
rect 21786 -15032 22939 -15002
rect 22973 -15032 23040 -14998
rect 23074 -15002 23107 -14998
rect 23171 -14113 24133 -14102
rect 23171 -14138 23243 -14113
rect 23171 -14172 23190 -14138
rect 23224 -14172 23243 -14138
rect 23171 -14228 23243 -14172
rect 24061 -14172 24133 -14113
rect 23171 -14262 23190 -14228
rect 23224 -14262 23243 -14228
rect 23171 -14318 23243 -14262
rect 23171 -14352 23190 -14318
rect 23224 -14352 23243 -14318
rect 23171 -14408 23243 -14352
rect 23171 -14442 23190 -14408
rect 23224 -14442 23243 -14408
rect 23171 -14498 23243 -14442
rect 23171 -14532 23190 -14498
rect 23224 -14532 23243 -14498
rect 23171 -14588 23243 -14532
rect 23171 -14622 23190 -14588
rect 23224 -14622 23243 -14588
rect 23171 -14678 23243 -14622
rect 23171 -14712 23190 -14678
rect 23224 -14712 23243 -14678
rect 23171 -14768 23243 -14712
rect 23171 -14802 23190 -14768
rect 23224 -14802 23243 -14768
rect 23171 -14858 23243 -14802
rect 23171 -14892 23190 -14858
rect 23224 -14892 23243 -14858
rect 23305 -14236 23999 -14175
rect 23305 -14270 23366 -14236
rect 23400 -14248 23456 -14236
rect 23490 -14248 23546 -14236
rect 23580 -14248 23636 -14236
rect 23412 -14270 23456 -14248
rect 23512 -14270 23546 -14248
rect 23612 -14270 23636 -14248
rect 23670 -14248 23726 -14236
rect 23670 -14270 23678 -14248
rect 23305 -14282 23378 -14270
rect 23412 -14282 23478 -14270
rect 23512 -14282 23578 -14270
rect 23612 -14282 23678 -14270
rect 23712 -14270 23726 -14248
rect 23760 -14248 23816 -14236
rect 23760 -14270 23778 -14248
rect 23712 -14282 23778 -14270
rect 23812 -14270 23816 -14248
rect 23850 -14248 23906 -14236
rect 23850 -14270 23878 -14248
rect 23940 -14270 23999 -14236
rect 23812 -14282 23878 -14270
rect 23912 -14282 23999 -14270
rect 23305 -14326 23999 -14282
rect 23305 -14360 23366 -14326
rect 23400 -14348 23456 -14326
rect 23490 -14348 23546 -14326
rect 23580 -14348 23636 -14326
rect 23412 -14360 23456 -14348
rect 23512 -14360 23546 -14348
rect 23612 -14360 23636 -14348
rect 23670 -14348 23726 -14326
rect 23670 -14360 23678 -14348
rect 23305 -14382 23378 -14360
rect 23412 -14382 23478 -14360
rect 23512 -14382 23578 -14360
rect 23612 -14382 23678 -14360
rect 23712 -14360 23726 -14348
rect 23760 -14348 23816 -14326
rect 23760 -14360 23778 -14348
rect 23712 -14382 23778 -14360
rect 23812 -14360 23816 -14348
rect 23850 -14348 23906 -14326
rect 23850 -14360 23878 -14348
rect 23940 -14360 23999 -14326
rect 23812 -14382 23878 -14360
rect 23912 -14382 23999 -14360
rect 23305 -14416 23999 -14382
rect 23305 -14450 23366 -14416
rect 23400 -14448 23456 -14416
rect 23490 -14448 23546 -14416
rect 23580 -14448 23636 -14416
rect 23412 -14450 23456 -14448
rect 23512 -14450 23546 -14448
rect 23612 -14450 23636 -14448
rect 23670 -14448 23726 -14416
rect 23670 -14450 23678 -14448
rect 23305 -14482 23378 -14450
rect 23412 -14482 23478 -14450
rect 23512 -14482 23578 -14450
rect 23612 -14482 23678 -14450
rect 23712 -14450 23726 -14448
rect 23760 -14448 23816 -14416
rect 23760 -14450 23778 -14448
rect 23712 -14482 23778 -14450
rect 23812 -14450 23816 -14448
rect 23850 -14448 23906 -14416
rect 23850 -14450 23878 -14448
rect 23940 -14450 23999 -14416
rect 23812 -14482 23878 -14450
rect 23912 -14482 23999 -14450
rect 23305 -14506 23999 -14482
rect 23305 -14540 23366 -14506
rect 23400 -14540 23456 -14506
rect 23490 -14540 23546 -14506
rect 23580 -14540 23636 -14506
rect 23670 -14540 23726 -14506
rect 23760 -14540 23816 -14506
rect 23850 -14540 23906 -14506
rect 23940 -14540 23999 -14506
rect 23305 -14548 23999 -14540
rect 23305 -14582 23378 -14548
rect 23412 -14582 23478 -14548
rect 23512 -14582 23578 -14548
rect 23612 -14582 23678 -14548
rect 23712 -14582 23778 -14548
rect 23812 -14582 23878 -14548
rect 23912 -14582 23999 -14548
rect 23305 -14596 23999 -14582
rect 23305 -14630 23366 -14596
rect 23400 -14630 23456 -14596
rect 23490 -14630 23546 -14596
rect 23580 -14630 23636 -14596
rect 23670 -14630 23726 -14596
rect 23760 -14630 23816 -14596
rect 23850 -14630 23906 -14596
rect 23940 -14630 23999 -14596
rect 23305 -14648 23999 -14630
rect 23305 -14682 23378 -14648
rect 23412 -14682 23478 -14648
rect 23512 -14682 23578 -14648
rect 23612 -14682 23678 -14648
rect 23712 -14682 23778 -14648
rect 23812 -14682 23878 -14648
rect 23912 -14682 23999 -14648
rect 23305 -14686 23999 -14682
rect 23305 -14720 23366 -14686
rect 23400 -14720 23456 -14686
rect 23490 -14720 23546 -14686
rect 23580 -14720 23636 -14686
rect 23670 -14720 23726 -14686
rect 23760 -14720 23816 -14686
rect 23850 -14720 23906 -14686
rect 23940 -14720 23999 -14686
rect 23305 -14748 23999 -14720
rect 23305 -14776 23378 -14748
rect 23412 -14776 23478 -14748
rect 23512 -14776 23578 -14748
rect 23612 -14776 23678 -14748
rect 23305 -14810 23366 -14776
rect 23412 -14782 23456 -14776
rect 23512 -14782 23546 -14776
rect 23612 -14782 23636 -14776
rect 23400 -14810 23456 -14782
rect 23490 -14810 23546 -14782
rect 23580 -14810 23636 -14782
rect 23670 -14782 23678 -14776
rect 23712 -14776 23778 -14748
rect 23712 -14782 23726 -14776
rect 23670 -14810 23726 -14782
rect 23760 -14782 23778 -14776
rect 23812 -14776 23878 -14748
rect 23912 -14776 23999 -14748
rect 23812 -14782 23816 -14776
rect 23760 -14810 23816 -14782
rect 23850 -14782 23878 -14776
rect 23850 -14810 23906 -14782
rect 23940 -14810 23999 -14776
rect 23305 -14869 23999 -14810
rect 24061 -14206 24080 -14172
rect 24114 -14206 24133 -14172
rect 24061 -14262 24133 -14206
rect 24061 -14296 24080 -14262
rect 24114 -14296 24133 -14262
rect 24061 -14352 24133 -14296
rect 24061 -14386 24080 -14352
rect 24114 -14386 24133 -14352
rect 24061 -14442 24133 -14386
rect 24061 -14476 24080 -14442
rect 24114 -14476 24133 -14442
rect 24061 -14532 24133 -14476
rect 24061 -14566 24080 -14532
rect 24114 -14566 24133 -14532
rect 24061 -14622 24133 -14566
rect 24061 -14656 24080 -14622
rect 24114 -14656 24133 -14622
rect 24061 -14712 24133 -14656
rect 24061 -14746 24080 -14712
rect 24114 -14746 24133 -14712
rect 24061 -14802 24133 -14746
rect 24061 -14836 24080 -14802
rect 24114 -14836 24133 -14802
rect 23171 -14931 23243 -14892
rect 24061 -14892 24133 -14836
rect 24061 -14926 24080 -14892
rect 24114 -14926 24133 -14892
rect 24061 -14931 24133 -14926
rect 23171 -14950 24133 -14931
rect 23171 -14984 23284 -14950
rect 23318 -14984 23374 -14950
rect 23408 -14984 23464 -14950
rect 23498 -14984 23554 -14950
rect 23588 -14984 23644 -14950
rect 23678 -14984 23734 -14950
rect 23768 -14984 23824 -14950
rect 23858 -14984 23914 -14950
rect 23948 -14984 24004 -14950
rect 24038 -14984 24133 -14950
rect 23171 -15002 24133 -14984
rect 24197 -14132 24227 -14102
rect 24261 -14132 24328 -14098
rect 24362 -14102 25515 -14098
rect 24362 -14132 24395 -14102
rect 24197 -14188 24395 -14132
rect 24197 -14222 24227 -14188
rect 24261 -14222 24328 -14188
rect 24362 -14222 24395 -14188
rect 24197 -14278 24395 -14222
rect 24197 -14312 24227 -14278
rect 24261 -14312 24328 -14278
rect 24362 -14312 24395 -14278
rect 24197 -14368 24395 -14312
rect 24197 -14402 24227 -14368
rect 24261 -14402 24328 -14368
rect 24362 -14402 24395 -14368
rect 24197 -14458 24395 -14402
rect 24197 -14492 24227 -14458
rect 24261 -14492 24328 -14458
rect 24362 -14492 24395 -14458
rect 24197 -14548 24395 -14492
rect 24197 -14582 24227 -14548
rect 24261 -14582 24328 -14548
rect 24362 -14582 24395 -14548
rect 24197 -14638 24395 -14582
rect 24197 -14672 24227 -14638
rect 24261 -14672 24328 -14638
rect 24362 -14672 24395 -14638
rect 24197 -14728 24395 -14672
rect 24197 -14762 24227 -14728
rect 24261 -14762 24328 -14728
rect 24362 -14762 24395 -14728
rect 24197 -14818 24395 -14762
rect 24197 -14852 24227 -14818
rect 24261 -14852 24328 -14818
rect 24362 -14852 24395 -14818
rect 24197 -14908 24395 -14852
rect 24197 -14942 24227 -14908
rect 24261 -14942 24328 -14908
rect 24362 -14942 24395 -14908
rect 24197 -14998 24395 -14942
rect 24197 -15002 24227 -14998
rect 23074 -15032 24227 -15002
rect 24261 -15032 24328 -14998
rect 24362 -15002 24395 -14998
rect 24459 -14113 25421 -14102
rect 24459 -14138 24531 -14113
rect 24459 -14172 24478 -14138
rect 24512 -14172 24531 -14138
rect 24459 -14228 24531 -14172
rect 25349 -14172 25421 -14113
rect 24459 -14262 24478 -14228
rect 24512 -14262 24531 -14228
rect 24459 -14318 24531 -14262
rect 24459 -14352 24478 -14318
rect 24512 -14352 24531 -14318
rect 24459 -14408 24531 -14352
rect 24459 -14442 24478 -14408
rect 24512 -14442 24531 -14408
rect 24459 -14498 24531 -14442
rect 24459 -14532 24478 -14498
rect 24512 -14532 24531 -14498
rect 24459 -14588 24531 -14532
rect 24459 -14622 24478 -14588
rect 24512 -14622 24531 -14588
rect 24459 -14678 24531 -14622
rect 24459 -14712 24478 -14678
rect 24512 -14712 24531 -14678
rect 24459 -14768 24531 -14712
rect 24459 -14802 24478 -14768
rect 24512 -14802 24531 -14768
rect 24459 -14858 24531 -14802
rect 24459 -14892 24478 -14858
rect 24512 -14892 24531 -14858
rect 24593 -14236 25287 -14175
rect 24593 -14270 24654 -14236
rect 24688 -14248 24744 -14236
rect 24778 -14248 24834 -14236
rect 24868 -14248 24924 -14236
rect 24700 -14270 24744 -14248
rect 24800 -14270 24834 -14248
rect 24900 -14270 24924 -14248
rect 24958 -14248 25014 -14236
rect 24958 -14270 24966 -14248
rect 24593 -14282 24666 -14270
rect 24700 -14282 24766 -14270
rect 24800 -14282 24866 -14270
rect 24900 -14282 24966 -14270
rect 25000 -14270 25014 -14248
rect 25048 -14248 25104 -14236
rect 25048 -14270 25066 -14248
rect 25000 -14282 25066 -14270
rect 25100 -14270 25104 -14248
rect 25138 -14248 25194 -14236
rect 25138 -14270 25166 -14248
rect 25228 -14270 25287 -14236
rect 25100 -14282 25166 -14270
rect 25200 -14282 25287 -14270
rect 24593 -14326 25287 -14282
rect 24593 -14360 24654 -14326
rect 24688 -14348 24744 -14326
rect 24778 -14348 24834 -14326
rect 24868 -14348 24924 -14326
rect 24700 -14360 24744 -14348
rect 24800 -14360 24834 -14348
rect 24900 -14360 24924 -14348
rect 24958 -14348 25014 -14326
rect 24958 -14360 24966 -14348
rect 24593 -14382 24666 -14360
rect 24700 -14382 24766 -14360
rect 24800 -14382 24866 -14360
rect 24900 -14382 24966 -14360
rect 25000 -14360 25014 -14348
rect 25048 -14348 25104 -14326
rect 25048 -14360 25066 -14348
rect 25000 -14382 25066 -14360
rect 25100 -14360 25104 -14348
rect 25138 -14348 25194 -14326
rect 25138 -14360 25166 -14348
rect 25228 -14360 25287 -14326
rect 25100 -14382 25166 -14360
rect 25200 -14382 25287 -14360
rect 24593 -14416 25287 -14382
rect 24593 -14450 24654 -14416
rect 24688 -14448 24744 -14416
rect 24778 -14448 24834 -14416
rect 24868 -14448 24924 -14416
rect 24700 -14450 24744 -14448
rect 24800 -14450 24834 -14448
rect 24900 -14450 24924 -14448
rect 24958 -14448 25014 -14416
rect 24958 -14450 24966 -14448
rect 24593 -14482 24666 -14450
rect 24700 -14482 24766 -14450
rect 24800 -14482 24866 -14450
rect 24900 -14482 24966 -14450
rect 25000 -14450 25014 -14448
rect 25048 -14448 25104 -14416
rect 25048 -14450 25066 -14448
rect 25000 -14482 25066 -14450
rect 25100 -14450 25104 -14448
rect 25138 -14448 25194 -14416
rect 25138 -14450 25166 -14448
rect 25228 -14450 25287 -14416
rect 25100 -14482 25166 -14450
rect 25200 -14482 25287 -14450
rect 24593 -14506 25287 -14482
rect 24593 -14540 24654 -14506
rect 24688 -14540 24744 -14506
rect 24778 -14540 24834 -14506
rect 24868 -14540 24924 -14506
rect 24958 -14540 25014 -14506
rect 25048 -14540 25104 -14506
rect 25138 -14540 25194 -14506
rect 25228 -14540 25287 -14506
rect 24593 -14548 25287 -14540
rect 24593 -14582 24666 -14548
rect 24700 -14582 24766 -14548
rect 24800 -14582 24866 -14548
rect 24900 -14582 24966 -14548
rect 25000 -14582 25066 -14548
rect 25100 -14582 25166 -14548
rect 25200 -14582 25287 -14548
rect 24593 -14596 25287 -14582
rect 24593 -14630 24654 -14596
rect 24688 -14630 24744 -14596
rect 24778 -14630 24834 -14596
rect 24868 -14630 24924 -14596
rect 24958 -14630 25014 -14596
rect 25048 -14630 25104 -14596
rect 25138 -14630 25194 -14596
rect 25228 -14630 25287 -14596
rect 24593 -14648 25287 -14630
rect 24593 -14682 24666 -14648
rect 24700 -14682 24766 -14648
rect 24800 -14682 24866 -14648
rect 24900 -14682 24966 -14648
rect 25000 -14682 25066 -14648
rect 25100 -14682 25166 -14648
rect 25200 -14682 25287 -14648
rect 24593 -14686 25287 -14682
rect 24593 -14720 24654 -14686
rect 24688 -14720 24744 -14686
rect 24778 -14720 24834 -14686
rect 24868 -14720 24924 -14686
rect 24958 -14720 25014 -14686
rect 25048 -14720 25104 -14686
rect 25138 -14720 25194 -14686
rect 25228 -14720 25287 -14686
rect 24593 -14748 25287 -14720
rect 24593 -14776 24666 -14748
rect 24700 -14776 24766 -14748
rect 24800 -14776 24866 -14748
rect 24900 -14776 24966 -14748
rect 24593 -14810 24654 -14776
rect 24700 -14782 24744 -14776
rect 24800 -14782 24834 -14776
rect 24900 -14782 24924 -14776
rect 24688 -14810 24744 -14782
rect 24778 -14810 24834 -14782
rect 24868 -14810 24924 -14782
rect 24958 -14782 24966 -14776
rect 25000 -14776 25066 -14748
rect 25000 -14782 25014 -14776
rect 24958 -14810 25014 -14782
rect 25048 -14782 25066 -14776
rect 25100 -14776 25166 -14748
rect 25200 -14776 25287 -14748
rect 25100 -14782 25104 -14776
rect 25048 -14810 25104 -14782
rect 25138 -14782 25166 -14776
rect 25138 -14810 25194 -14782
rect 25228 -14810 25287 -14776
rect 24593 -14869 25287 -14810
rect 25349 -14206 25368 -14172
rect 25402 -14206 25421 -14172
rect 25349 -14262 25421 -14206
rect 25349 -14296 25368 -14262
rect 25402 -14296 25421 -14262
rect 25349 -14352 25421 -14296
rect 25349 -14386 25368 -14352
rect 25402 -14386 25421 -14352
rect 25349 -14442 25421 -14386
rect 25349 -14476 25368 -14442
rect 25402 -14476 25421 -14442
rect 25349 -14532 25421 -14476
rect 25349 -14566 25368 -14532
rect 25402 -14566 25421 -14532
rect 25349 -14622 25421 -14566
rect 25349 -14656 25368 -14622
rect 25402 -14656 25421 -14622
rect 25349 -14712 25421 -14656
rect 25349 -14746 25368 -14712
rect 25402 -14746 25421 -14712
rect 25349 -14802 25421 -14746
rect 25349 -14836 25368 -14802
rect 25402 -14836 25421 -14802
rect 24459 -14931 24531 -14892
rect 25349 -14892 25421 -14836
rect 25349 -14926 25368 -14892
rect 25402 -14926 25421 -14892
rect 25349 -14931 25421 -14926
rect 24459 -14950 25421 -14931
rect 24459 -14984 24572 -14950
rect 24606 -14984 24662 -14950
rect 24696 -14984 24752 -14950
rect 24786 -14984 24842 -14950
rect 24876 -14984 24932 -14950
rect 24966 -14984 25022 -14950
rect 25056 -14984 25112 -14950
rect 25146 -14984 25202 -14950
rect 25236 -14984 25292 -14950
rect 25326 -14984 25421 -14950
rect 24459 -15002 25421 -14984
rect 25485 -14132 25515 -14102
rect 25549 -14132 25616 -14098
rect 25650 -14102 26803 -14098
rect 25650 -14132 25683 -14102
rect 25485 -14188 25683 -14132
rect 25485 -14222 25515 -14188
rect 25549 -14222 25616 -14188
rect 25650 -14222 25683 -14188
rect 25485 -14278 25683 -14222
rect 25485 -14312 25515 -14278
rect 25549 -14312 25616 -14278
rect 25650 -14312 25683 -14278
rect 25485 -14368 25683 -14312
rect 25485 -14402 25515 -14368
rect 25549 -14402 25616 -14368
rect 25650 -14402 25683 -14368
rect 25485 -14458 25683 -14402
rect 25485 -14492 25515 -14458
rect 25549 -14492 25616 -14458
rect 25650 -14492 25683 -14458
rect 25485 -14548 25683 -14492
rect 25485 -14582 25515 -14548
rect 25549 -14582 25616 -14548
rect 25650 -14582 25683 -14548
rect 25485 -14638 25683 -14582
rect 25485 -14672 25515 -14638
rect 25549 -14672 25616 -14638
rect 25650 -14672 25683 -14638
rect 25485 -14728 25683 -14672
rect 25485 -14762 25515 -14728
rect 25549 -14762 25616 -14728
rect 25650 -14762 25683 -14728
rect 25485 -14818 25683 -14762
rect 25485 -14852 25515 -14818
rect 25549 -14852 25616 -14818
rect 25650 -14852 25683 -14818
rect 25485 -14908 25683 -14852
rect 25485 -14942 25515 -14908
rect 25549 -14942 25616 -14908
rect 25650 -14942 25683 -14908
rect 25485 -14998 25683 -14942
rect 25485 -15002 25515 -14998
rect 24362 -15032 25515 -15002
rect 25549 -15032 25616 -14998
rect 25650 -15002 25683 -14998
rect 25747 -14113 26709 -14102
rect 25747 -14138 25819 -14113
rect 25747 -14172 25766 -14138
rect 25800 -14172 25819 -14138
rect 25747 -14228 25819 -14172
rect 26637 -14172 26709 -14113
rect 25747 -14262 25766 -14228
rect 25800 -14262 25819 -14228
rect 25747 -14318 25819 -14262
rect 25747 -14352 25766 -14318
rect 25800 -14352 25819 -14318
rect 25747 -14408 25819 -14352
rect 25747 -14442 25766 -14408
rect 25800 -14442 25819 -14408
rect 25747 -14498 25819 -14442
rect 25747 -14532 25766 -14498
rect 25800 -14532 25819 -14498
rect 25747 -14588 25819 -14532
rect 25747 -14622 25766 -14588
rect 25800 -14622 25819 -14588
rect 25747 -14678 25819 -14622
rect 25747 -14712 25766 -14678
rect 25800 -14712 25819 -14678
rect 25747 -14768 25819 -14712
rect 25747 -14802 25766 -14768
rect 25800 -14802 25819 -14768
rect 25747 -14858 25819 -14802
rect 25747 -14892 25766 -14858
rect 25800 -14892 25819 -14858
rect 25881 -14236 26575 -14175
rect 25881 -14270 25942 -14236
rect 25976 -14248 26032 -14236
rect 26066 -14248 26122 -14236
rect 26156 -14248 26212 -14236
rect 25988 -14270 26032 -14248
rect 26088 -14270 26122 -14248
rect 26188 -14270 26212 -14248
rect 26246 -14248 26302 -14236
rect 26246 -14270 26254 -14248
rect 25881 -14282 25954 -14270
rect 25988 -14282 26054 -14270
rect 26088 -14282 26154 -14270
rect 26188 -14282 26254 -14270
rect 26288 -14270 26302 -14248
rect 26336 -14248 26392 -14236
rect 26336 -14270 26354 -14248
rect 26288 -14282 26354 -14270
rect 26388 -14270 26392 -14248
rect 26426 -14248 26482 -14236
rect 26426 -14270 26454 -14248
rect 26516 -14270 26575 -14236
rect 26388 -14282 26454 -14270
rect 26488 -14282 26575 -14270
rect 25881 -14326 26575 -14282
rect 25881 -14360 25942 -14326
rect 25976 -14348 26032 -14326
rect 26066 -14348 26122 -14326
rect 26156 -14348 26212 -14326
rect 25988 -14360 26032 -14348
rect 26088 -14360 26122 -14348
rect 26188 -14360 26212 -14348
rect 26246 -14348 26302 -14326
rect 26246 -14360 26254 -14348
rect 25881 -14382 25954 -14360
rect 25988 -14382 26054 -14360
rect 26088 -14382 26154 -14360
rect 26188 -14382 26254 -14360
rect 26288 -14360 26302 -14348
rect 26336 -14348 26392 -14326
rect 26336 -14360 26354 -14348
rect 26288 -14382 26354 -14360
rect 26388 -14360 26392 -14348
rect 26426 -14348 26482 -14326
rect 26426 -14360 26454 -14348
rect 26516 -14360 26575 -14326
rect 26388 -14382 26454 -14360
rect 26488 -14382 26575 -14360
rect 25881 -14416 26575 -14382
rect 25881 -14450 25942 -14416
rect 25976 -14448 26032 -14416
rect 26066 -14448 26122 -14416
rect 26156 -14448 26212 -14416
rect 25988 -14450 26032 -14448
rect 26088 -14450 26122 -14448
rect 26188 -14450 26212 -14448
rect 26246 -14448 26302 -14416
rect 26246 -14450 26254 -14448
rect 25881 -14482 25954 -14450
rect 25988 -14482 26054 -14450
rect 26088 -14482 26154 -14450
rect 26188 -14482 26254 -14450
rect 26288 -14450 26302 -14448
rect 26336 -14448 26392 -14416
rect 26336 -14450 26354 -14448
rect 26288 -14482 26354 -14450
rect 26388 -14450 26392 -14448
rect 26426 -14448 26482 -14416
rect 26426 -14450 26454 -14448
rect 26516 -14450 26575 -14416
rect 26388 -14482 26454 -14450
rect 26488 -14482 26575 -14450
rect 25881 -14506 26575 -14482
rect 25881 -14540 25942 -14506
rect 25976 -14540 26032 -14506
rect 26066 -14540 26122 -14506
rect 26156 -14540 26212 -14506
rect 26246 -14540 26302 -14506
rect 26336 -14540 26392 -14506
rect 26426 -14540 26482 -14506
rect 26516 -14540 26575 -14506
rect 25881 -14548 26575 -14540
rect 25881 -14582 25954 -14548
rect 25988 -14582 26054 -14548
rect 26088 -14582 26154 -14548
rect 26188 -14582 26254 -14548
rect 26288 -14582 26354 -14548
rect 26388 -14582 26454 -14548
rect 26488 -14582 26575 -14548
rect 25881 -14596 26575 -14582
rect 25881 -14630 25942 -14596
rect 25976 -14630 26032 -14596
rect 26066 -14630 26122 -14596
rect 26156 -14630 26212 -14596
rect 26246 -14630 26302 -14596
rect 26336 -14630 26392 -14596
rect 26426 -14630 26482 -14596
rect 26516 -14630 26575 -14596
rect 25881 -14648 26575 -14630
rect 25881 -14682 25954 -14648
rect 25988 -14682 26054 -14648
rect 26088 -14682 26154 -14648
rect 26188 -14682 26254 -14648
rect 26288 -14682 26354 -14648
rect 26388 -14682 26454 -14648
rect 26488 -14682 26575 -14648
rect 25881 -14686 26575 -14682
rect 25881 -14720 25942 -14686
rect 25976 -14720 26032 -14686
rect 26066 -14720 26122 -14686
rect 26156 -14720 26212 -14686
rect 26246 -14720 26302 -14686
rect 26336 -14720 26392 -14686
rect 26426 -14720 26482 -14686
rect 26516 -14720 26575 -14686
rect 25881 -14748 26575 -14720
rect 25881 -14776 25954 -14748
rect 25988 -14776 26054 -14748
rect 26088 -14776 26154 -14748
rect 26188 -14776 26254 -14748
rect 25881 -14810 25942 -14776
rect 25988 -14782 26032 -14776
rect 26088 -14782 26122 -14776
rect 26188 -14782 26212 -14776
rect 25976 -14810 26032 -14782
rect 26066 -14810 26122 -14782
rect 26156 -14810 26212 -14782
rect 26246 -14782 26254 -14776
rect 26288 -14776 26354 -14748
rect 26288 -14782 26302 -14776
rect 26246 -14810 26302 -14782
rect 26336 -14782 26354 -14776
rect 26388 -14776 26454 -14748
rect 26488 -14776 26575 -14748
rect 26388 -14782 26392 -14776
rect 26336 -14810 26392 -14782
rect 26426 -14782 26454 -14776
rect 26426 -14810 26482 -14782
rect 26516 -14810 26575 -14776
rect 25881 -14869 26575 -14810
rect 26637 -14206 26656 -14172
rect 26690 -14206 26709 -14172
rect 26637 -14262 26709 -14206
rect 26637 -14296 26656 -14262
rect 26690 -14296 26709 -14262
rect 26637 -14352 26709 -14296
rect 26637 -14386 26656 -14352
rect 26690 -14386 26709 -14352
rect 26637 -14442 26709 -14386
rect 26637 -14476 26656 -14442
rect 26690 -14476 26709 -14442
rect 26637 -14532 26709 -14476
rect 26637 -14566 26656 -14532
rect 26690 -14566 26709 -14532
rect 26637 -14622 26709 -14566
rect 26637 -14656 26656 -14622
rect 26690 -14656 26709 -14622
rect 26637 -14712 26709 -14656
rect 26637 -14746 26656 -14712
rect 26690 -14746 26709 -14712
rect 26637 -14802 26709 -14746
rect 26637 -14836 26656 -14802
rect 26690 -14836 26709 -14802
rect 25747 -14931 25819 -14892
rect 26637 -14892 26709 -14836
rect 26637 -14926 26656 -14892
rect 26690 -14926 26709 -14892
rect 26637 -14931 26709 -14926
rect 25747 -14950 26709 -14931
rect 25747 -14984 25860 -14950
rect 25894 -14984 25950 -14950
rect 25984 -14984 26040 -14950
rect 26074 -14984 26130 -14950
rect 26164 -14984 26220 -14950
rect 26254 -14984 26310 -14950
rect 26344 -14984 26400 -14950
rect 26434 -14984 26490 -14950
rect 26524 -14984 26580 -14950
rect 26614 -14984 26709 -14950
rect 25747 -15002 26709 -14984
rect 26773 -14132 26803 -14102
rect 26837 -14132 26872 -14098
rect 26773 -14188 26872 -14132
rect 26773 -14222 26803 -14188
rect 26837 -14222 26872 -14188
rect 26773 -14278 26872 -14222
rect 26773 -14312 26803 -14278
rect 26837 -14312 26872 -14278
rect 26773 -14368 26872 -14312
rect 26773 -14402 26803 -14368
rect 26837 -14402 26872 -14368
rect 26773 -14458 26872 -14402
rect 26773 -14492 26803 -14458
rect 26837 -14492 26872 -14458
rect 26773 -14548 26872 -14492
rect 26773 -14582 26803 -14548
rect 26837 -14582 26872 -14548
rect 26773 -14638 26872 -14582
rect 26773 -14672 26803 -14638
rect 26837 -14672 26872 -14638
rect 26773 -14728 26872 -14672
rect 26773 -14762 26803 -14728
rect 26837 -14762 26872 -14728
rect 26773 -14818 26872 -14762
rect 26773 -14852 26803 -14818
rect 26837 -14852 26872 -14818
rect 26773 -14908 26872 -14852
rect 26773 -14942 26803 -14908
rect 26837 -14942 26872 -14908
rect 26773 -14998 26872 -14942
rect 26773 -15002 26803 -14998
rect 25650 -15032 26803 -15002
rect 26837 -15032 26872 -14998
rect 16568 -15099 26872 -15032
rect 16568 -15133 16684 -15099
rect 16718 -15133 16774 -15099
rect 16808 -15133 16864 -15099
rect 16898 -15133 16954 -15099
rect 16988 -15133 17044 -15099
rect 17078 -15133 17134 -15099
rect 17168 -15133 17224 -15099
rect 17258 -15133 17314 -15099
rect 17348 -15133 17404 -15099
rect 17438 -15133 17494 -15099
rect 17528 -15133 17584 -15099
rect 17618 -15133 17674 -15099
rect 17708 -15133 17764 -15099
rect 17798 -15133 17972 -15099
rect 18006 -15133 18062 -15099
rect 18096 -15133 18152 -15099
rect 18186 -15133 18242 -15099
rect 18276 -15133 18332 -15099
rect 18366 -15133 18422 -15099
rect 18456 -15133 18512 -15099
rect 18546 -15133 18602 -15099
rect 18636 -15133 18692 -15099
rect 18726 -15133 18782 -15099
rect 18816 -15133 18872 -15099
rect 18906 -15133 18962 -15099
rect 18996 -15133 19052 -15099
rect 19086 -15133 19260 -15099
rect 19294 -15133 19350 -15099
rect 19384 -15133 19440 -15099
rect 19474 -15133 19530 -15099
rect 19564 -15133 19620 -15099
rect 19654 -15133 19710 -15099
rect 19744 -15133 19800 -15099
rect 19834 -15133 19890 -15099
rect 19924 -15133 19980 -15099
rect 20014 -15133 20070 -15099
rect 20104 -15133 20160 -15099
rect 20194 -15133 20250 -15099
rect 20284 -15133 20340 -15099
rect 20374 -15133 20548 -15099
rect 20582 -15133 20638 -15099
rect 20672 -15133 20728 -15099
rect 20762 -15133 20818 -15099
rect 20852 -15133 20908 -15099
rect 20942 -15133 20998 -15099
rect 21032 -15133 21088 -15099
rect 21122 -15133 21178 -15099
rect 21212 -15133 21268 -15099
rect 21302 -15133 21358 -15099
rect 21392 -15133 21448 -15099
rect 21482 -15133 21538 -15099
rect 21572 -15133 21628 -15099
rect 21662 -15133 21836 -15099
rect 21870 -15133 21926 -15099
rect 21960 -15133 22016 -15099
rect 22050 -15133 22106 -15099
rect 22140 -15133 22196 -15099
rect 22230 -15133 22286 -15099
rect 22320 -15133 22376 -15099
rect 22410 -15133 22466 -15099
rect 22500 -15133 22556 -15099
rect 22590 -15133 22646 -15099
rect 22680 -15133 22736 -15099
rect 22770 -15133 22826 -15099
rect 22860 -15133 22916 -15099
rect 22950 -15133 23124 -15099
rect 23158 -15133 23214 -15099
rect 23248 -15133 23304 -15099
rect 23338 -15133 23394 -15099
rect 23428 -15133 23484 -15099
rect 23518 -15133 23574 -15099
rect 23608 -15133 23664 -15099
rect 23698 -15133 23754 -15099
rect 23788 -15133 23844 -15099
rect 23878 -15133 23934 -15099
rect 23968 -15133 24024 -15099
rect 24058 -15133 24114 -15099
rect 24148 -15133 24204 -15099
rect 24238 -15133 24412 -15099
rect 24446 -15133 24502 -15099
rect 24536 -15133 24592 -15099
rect 24626 -15133 24682 -15099
rect 24716 -15133 24772 -15099
rect 24806 -15133 24862 -15099
rect 24896 -15133 24952 -15099
rect 24986 -15133 25042 -15099
rect 25076 -15133 25132 -15099
rect 25166 -15133 25222 -15099
rect 25256 -15133 25312 -15099
rect 25346 -15133 25402 -15099
rect 25436 -15133 25492 -15099
rect 25526 -15133 25700 -15099
rect 25734 -15133 25790 -15099
rect 25824 -15133 25880 -15099
rect 25914 -15133 25970 -15099
rect 26004 -15133 26060 -15099
rect 26094 -15133 26150 -15099
rect 26184 -15133 26240 -15099
rect 26274 -15133 26330 -15099
rect 26364 -15133 26420 -15099
rect 26454 -15133 26510 -15099
rect 26544 -15133 26600 -15099
rect 26634 -15133 26690 -15099
rect 26724 -15133 26780 -15099
rect 26814 -15133 26872 -15099
rect 16568 -15200 26872 -15133
rect 16568 -15234 16684 -15200
rect 16718 -15234 16774 -15200
rect 16808 -15234 16864 -15200
rect 16898 -15234 16954 -15200
rect 16988 -15234 17044 -15200
rect 17078 -15234 17134 -15200
rect 17168 -15234 17224 -15200
rect 17258 -15234 17314 -15200
rect 17348 -15234 17404 -15200
rect 17438 -15234 17494 -15200
rect 17528 -15234 17584 -15200
rect 17618 -15234 17674 -15200
rect 17708 -15234 17764 -15200
rect 17798 -15234 17972 -15200
rect 18006 -15234 18062 -15200
rect 18096 -15234 18152 -15200
rect 18186 -15234 18242 -15200
rect 18276 -15234 18332 -15200
rect 18366 -15234 18422 -15200
rect 18456 -15234 18512 -15200
rect 18546 -15234 18602 -15200
rect 18636 -15234 18692 -15200
rect 18726 -15234 18782 -15200
rect 18816 -15234 18872 -15200
rect 18906 -15234 18962 -15200
rect 18996 -15234 19052 -15200
rect 19086 -15234 19260 -15200
rect 19294 -15234 19350 -15200
rect 19384 -15234 19440 -15200
rect 19474 -15234 19530 -15200
rect 19564 -15234 19620 -15200
rect 19654 -15234 19710 -15200
rect 19744 -15234 19800 -15200
rect 19834 -15234 19890 -15200
rect 19924 -15234 19980 -15200
rect 20014 -15234 20070 -15200
rect 20104 -15234 20160 -15200
rect 20194 -15234 20250 -15200
rect 20284 -15234 20340 -15200
rect 20374 -15234 20548 -15200
rect 20582 -15234 20638 -15200
rect 20672 -15234 20728 -15200
rect 20762 -15234 20818 -15200
rect 20852 -15234 20908 -15200
rect 20942 -15234 20998 -15200
rect 21032 -15234 21088 -15200
rect 21122 -15234 21178 -15200
rect 21212 -15234 21268 -15200
rect 21302 -15234 21358 -15200
rect 21392 -15234 21448 -15200
rect 21482 -15234 21538 -15200
rect 21572 -15234 21628 -15200
rect 21662 -15234 21836 -15200
rect 21870 -15234 21926 -15200
rect 21960 -15234 22016 -15200
rect 22050 -15234 22106 -15200
rect 22140 -15234 22196 -15200
rect 22230 -15234 22286 -15200
rect 22320 -15234 22376 -15200
rect 22410 -15234 22466 -15200
rect 22500 -15234 22556 -15200
rect 22590 -15234 22646 -15200
rect 22680 -15234 22736 -15200
rect 22770 -15234 22826 -15200
rect 22860 -15234 22916 -15200
rect 22950 -15234 23124 -15200
rect 23158 -15234 23214 -15200
rect 23248 -15234 23304 -15200
rect 23338 -15234 23394 -15200
rect 23428 -15234 23484 -15200
rect 23518 -15234 23574 -15200
rect 23608 -15234 23664 -15200
rect 23698 -15234 23754 -15200
rect 23788 -15234 23844 -15200
rect 23878 -15234 23934 -15200
rect 23968 -15234 24024 -15200
rect 24058 -15234 24114 -15200
rect 24148 -15234 24204 -15200
rect 24238 -15234 24412 -15200
rect 24446 -15234 24502 -15200
rect 24536 -15234 24592 -15200
rect 24626 -15234 24682 -15200
rect 24716 -15234 24772 -15200
rect 24806 -15234 24862 -15200
rect 24896 -15234 24952 -15200
rect 24986 -15234 25042 -15200
rect 25076 -15234 25132 -15200
rect 25166 -15234 25222 -15200
rect 25256 -15234 25312 -15200
rect 25346 -15234 25402 -15200
rect 25436 -15234 25492 -15200
rect 25526 -15234 25700 -15200
rect 25734 -15234 25790 -15200
rect 25824 -15234 25880 -15200
rect 25914 -15234 25970 -15200
rect 26004 -15234 26060 -15200
rect 26094 -15234 26150 -15200
rect 26184 -15234 26240 -15200
rect 26274 -15234 26330 -15200
rect 26364 -15234 26420 -15200
rect 26454 -15234 26510 -15200
rect 26544 -15234 26600 -15200
rect 26634 -15234 26690 -15200
rect 26724 -15234 26780 -15200
rect 26814 -15234 26872 -15200
rect 16568 -15296 26872 -15234
rect 16568 -15330 16600 -15296
rect 16634 -15330 17787 -15296
rect 17821 -15330 17888 -15296
rect 17922 -15330 19075 -15296
rect 19109 -15330 19176 -15296
rect 19210 -15330 20363 -15296
rect 20397 -15330 20464 -15296
rect 20498 -15330 21651 -15296
rect 21685 -15330 21752 -15296
rect 21786 -15330 22939 -15296
rect 22973 -15330 23040 -15296
rect 23074 -15330 24227 -15296
rect 24261 -15330 24328 -15296
rect 24362 -15330 25515 -15296
rect 25549 -15330 25616 -15296
rect 25650 -15330 26803 -15296
rect 26837 -15330 26872 -15296
rect 16568 -15348 26872 -15330
rect 16568 -15382 16863 -15348
rect 16897 -15382 16953 -15348
rect 16987 -15382 17043 -15348
rect 17077 -15382 17133 -15348
rect 17167 -15382 17223 -15348
rect 17257 -15382 17313 -15348
rect 17347 -15382 17403 -15348
rect 17437 -15382 17493 -15348
rect 17527 -15382 17583 -15348
rect 17617 -15382 18151 -15348
rect 18185 -15382 18241 -15348
rect 18275 -15382 18331 -15348
rect 18365 -15382 18421 -15348
rect 18455 -15382 18511 -15348
rect 18545 -15382 18601 -15348
rect 18635 -15382 18691 -15348
rect 18725 -15382 18781 -15348
rect 18815 -15382 18871 -15348
rect 18905 -15382 19439 -15348
rect 19473 -15382 19529 -15348
rect 19563 -15382 19619 -15348
rect 19653 -15382 19709 -15348
rect 19743 -15382 19799 -15348
rect 19833 -15382 19889 -15348
rect 19923 -15382 19979 -15348
rect 20013 -15382 20069 -15348
rect 20103 -15382 20159 -15348
rect 20193 -15382 20727 -15348
rect 20761 -15382 20817 -15348
rect 20851 -15382 20907 -15348
rect 20941 -15382 20997 -15348
rect 21031 -15382 21087 -15348
rect 21121 -15382 21177 -15348
rect 21211 -15382 21267 -15348
rect 21301 -15382 21357 -15348
rect 21391 -15382 21447 -15348
rect 21481 -15382 22015 -15348
rect 22049 -15382 22105 -15348
rect 22139 -15382 22195 -15348
rect 22229 -15382 22285 -15348
rect 22319 -15382 22375 -15348
rect 22409 -15382 22465 -15348
rect 22499 -15382 22555 -15348
rect 22589 -15382 22645 -15348
rect 22679 -15382 22735 -15348
rect 22769 -15382 23303 -15348
rect 23337 -15382 23393 -15348
rect 23427 -15382 23483 -15348
rect 23517 -15382 23573 -15348
rect 23607 -15382 23663 -15348
rect 23697 -15382 23753 -15348
rect 23787 -15382 23843 -15348
rect 23877 -15382 23933 -15348
rect 23967 -15382 24023 -15348
rect 24057 -15382 24591 -15348
rect 24625 -15382 24681 -15348
rect 24715 -15382 24771 -15348
rect 24805 -15382 24861 -15348
rect 24895 -15382 24951 -15348
rect 24985 -15382 25041 -15348
rect 25075 -15382 25131 -15348
rect 25165 -15382 25221 -15348
rect 25255 -15382 25311 -15348
rect 25345 -15382 25879 -15348
rect 25913 -15382 25969 -15348
rect 26003 -15382 26059 -15348
rect 26093 -15382 26149 -15348
rect 26183 -15382 26239 -15348
rect 26273 -15382 26329 -15348
rect 26363 -15382 26419 -15348
rect 26453 -15382 26509 -15348
rect 26543 -15382 26599 -15348
rect 26633 -15382 26872 -15348
rect 16568 -15386 26872 -15382
rect 16568 -15420 16600 -15386
rect 16634 -15402 17787 -15386
rect 16634 -15420 16667 -15402
rect 16568 -15476 16667 -15420
rect 16568 -15510 16600 -15476
rect 16634 -15510 16667 -15476
rect 16568 -15566 16667 -15510
rect 16568 -15600 16600 -15566
rect 16634 -15600 16667 -15566
rect 16568 -15656 16667 -15600
rect 16568 -15690 16600 -15656
rect 16634 -15690 16667 -15656
rect 16568 -15746 16667 -15690
rect 16568 -15780 16600 -15746
rect 16634 -15780 16667 -15746
rect 16568 -15836 16667 -15780
rect 16568 -15870 16600 -15836
rect 16634 -15870 16667 -15836
rect 16568 -15926 16667 -15870
rect 16568 -15960 16600 -15926
rect 16634 -15960 16667 -15926
rect 16568 -16016 16667 -15960
rect 16568 -16050 16600 -16016
rect 16634 -16050 16667 -16016
rect 16568 -16106 16667 -16050
rect 16568 -16140 16600 -16106
rect 16634 -16140 16667 -16106
rect 16568 -16196 16667 -16140
rect 16568 -16230 16600 -16196
rect 16634 -16202 16667 -16196
rect 16731 -15426 16803 -15402
rect 16731 -15460 16750 -15426
rect 16784 -15460 16803 -15426
rect 16731 -15516 16803 -15460
rect 17621 -15460 17693 -15402
rect 16731 -15550 16750 -15516
rect 16784 -15550 16803 -15516
rect 16731 -15606 16803 -15550
rect 16731 -15640 16750 -15606
rect 16784 -15640 16803 -15606
rect 16731 -15696 16803 -15640
rect 16731 -15730 16750 -15696
rect 16784 -15730 16803 -15696
rect 16731 -15786 16803 -15730
rect 16731 -15820 16750 -15786
rect 16784 -15820 16803 -15786
rect 16731 -15876 16803 -15820
rect 16731 -15910 16750 -15876
rect 16784 -15910 16803 -15876
rect 16731 -15966 16803 -15910
rect 16731 -16000 16750 -15966
rect 16784 -16000 16803 -15966
rect 16731 -16056 16803 -16000
rect 16731 -16090 16750 -16056
rect 16784 -16090 16803 -16056
rect 16731 -16146 16803 -16090
rect 16731 -16180 16750 -16146
rect 16784 -16180 16803 -16146
rect 16865 -15524 17559 -15463
rect 16865 -15558 16926 -15524
rect 16960 -15536 17016 -15524
rect 17050 -15536 17106 -15524
rect 17140 -15536 17196 -15524
rect 16972 -15558 17016 -15536
rect 17072 -15558 17106 -15536
rect 17172 -15558 17196 -15536
rect 17230 -15536 17286 -15524
rect 17230 -15558 17238 -15536
rect 16865 -15570 16938 -15558
rect 16972 -15570 17038 -15558
rect 17072 -15570 17138 -15558
rect 17172 -15570 17238 -15558
rect 17272 -15558 17286 -15536
rect 17320 -15536 17376 -15524
rect 17320 -15558 17338 -15536
rect 17272 -15570 17338 -15558
rect 17372 -15558 17376 -15536
rect 17410 -15536 17466 -15524
rect 17410 -15558 17438 -15536
rect 17500 -15558 17559 -15524
rect 17372 -15570 17438 -15558
rect 17472 -15570 17559 -15558
rect 16865 -15614 17559 -15570
rect 16865 -15648 16926 -15614
rect 16960 -15636 17016 -15614
rect 17050 -15636 17106 -15614
rect 17140 -15636 17196 -15614
rect 16972 -15648 17016 -15636
rect 17072 -15648 17106 -15636
rect 17172 -15648 17196 -15636
rect 17230 -15636 17286 -15614
rect 17230 -15648 17238 -15636
rect 16865 -15670 16938 -15648
rect 16972 -15670 17038 -15648
rect 17072 -15670 17138 -15648
rect 17172 -15670 17238 -15648
rect 17272 -15648 17286 -15636
rect 17320 -15636 17376 -15614
rect 17320 -15648 17338 -15636
rect 17272 -15670 17338 -15648
rect 17372 -15648 17376 -15636
rect 17410 -15636 17466 -15614
rect 17410 -15648 17438 -15636
rect 17500 -15648 17559 -15614
rect 17372 -15670 17438 -15648
rect 17472 -15670 17559 -15648
rect 16865 -15704 17559 -15670
rect 16865 -15738 16926 -15704
rect 16960 -15736 17016 -15704
rect 17050 -15736 17106 -15704
rect 17140 -15736 17196 -15704
rect 16972 -15738 17016 -15736
rect 17072 -15738 17106 -15736
rect 17172 -15738 17196 -15736
rect 17230 -15736 17286 -15704
rect 17230 -15738 17238 -15736
rect 16865 -15770 16938 -15738
rect 16972 -15770 17038 -15738
rect 17072 -15770 17138 -15738
rect 17172 -15770 17238 -15738
rect 17272 -15738 17286 -15736
rect 17320 -15736 17376 -15704
rect 17320 -15738 17338 -15736
rect 17272 -15770 17338 -15738
rect 17372 -15738 17376 -15736
rect 17410 -15736 17466 -15704
rect 17410 -15738 17438 -15736
rect 17500 -15738 17559 -15704
rect 17372 -15770 17438 -15738
rect 17472 -15770 17559 -15738
rect 16865 -15794 17559 -15770
rect 16865 -15828 16926 -15794
rect 16960 -15828 17016 -15794
rect 17050 -15828 17106 -15794
rect 17140 -15828 17196 -15794
rect 17230 -15828 17286 -15794
rect 17320 -15828 17376 -15794
rect 17410 -15828 17466 -15794
rect 17500 -15828 17559 -15794
rect 16865 -15836 17559 -15828
rect 16865 -15870 16938 -15836
rect 16972 -15870 17038 -15836
rect 17072 -15870 17138 -15836
rect 17172 -15870 17238 -15836
rect 17272 -15870 17338 -15836
rect 17372 -15870 17438 -15836
rect 17472 -15870 17559 -15836
rect 16865 -15884 17559 -15870
rect 16865 -15918 16926 -15884
rect 16960 -15918 17016 -15884
rect 17050 -15918 17106 -15884
rect 17140 -15918 17196 -15884
rect 17230 -15918 17286 -15884
rect 17320 -15918 17376 -15884
rect 17410 -15918 17466 -15884
rect 17500 -15918 17559 -15884
rect 16865 -15936 17559 -15918
rect 16865 -15970 16938 -15936
rect 16972 -15970 17038 -15936
rect 17072 -15970 17138 -15936
rect 17172 -15970 17238 -15936
rect 17272 -15970 17338 -15936
rect 17372 -15970 17438 -15936
rect 17472 -15970 17559 -15936
rect 16865 -15974 17559 -15970
rect 16865 -16008 16926 -15974
rect 16960 -16008 17016 -15974
rect 17050 -16008 17106 -15974
rect 17140 -16008 17196 -15974
rect 17230 -16008 17286 -15974
rect 17320 -16008 17376 -15974
rect 17410 -16008 17466 -15974
rect 17500 -16008 17559 -15974
rect 16865 -16036 17559 -16008
rect 16865 -16064 16938 -16036
rect 16972 -16064 17038 -16036
rect 17072 -16064 17138 -16036
rect 17172 -16064 17238 -16036
rect 16865 -16098 16926 -16064
rect 16972 -16070 17016 -16064
rect 17072 -16070 17106 -16064
rect 17172 -16070 17196 -16064
rect 16960 -16098 17016 -16070
rect 17050 -16098 17106 -16070
rect 17140 -16098 17196 -16070
rect 17230 -16070 17238 -16064
rect 17272 -16064 17338 -16036
rect 17272 -16070 17286 -16064
rect 17230 -16098 17286 -16070
rect 17320 -16070 17338 -16064
rect 17372 -16064 17438 -16036
rect 17472 -16064 17559 -16036
rect 17372 -16070 17376 -16064
rect 17320 -16098 17376 -16070
rect 17410 -16070 17438 -16064
rect 17410 -16098 17466 -16070
rect 17500 -16098 17559 -16064
rect 16865 -16157 17559 -16098
rect 17621 -15494 17640 -15460
rect 17674 -15494 17693 -15460
rect 17621 -15550 17693 -15494
rect 17621 -15584 17640 -15550
rect 17674 -15584 17693 -15550
rect 17621 -15640 17693 -15584
rect 17621 -15674 17640 -15640
rect 17674 -15674 17693 -15640
rect 17621 -15730 17693 -15674
rect 17621 -15764 17640 -15730
rect 17674 -15764 17693 -15730
rect 17621 -15820 17693 -15764
rect 17621 -15854 17640 -15820
rect 17674 -15854 17693 -15820
rect 17621 -15910 17693 -15854
rect 17621 -15944 17640 -15910
rect 17674 -15944 17693 -15910
rect 17621 -16000 17693 -15944
rect 17621 -16034 17640 -16000
rect 17674 -16034 17693 -16000
rect 17621 -16090 17693 -16034
rect 17621 -16124 17640 -16090
rect 17674 -16124 17693 -16090
rect 16731 -16202 16803 -16180
rect 17621 -16180 17693 -16124
rect 17621 -16202 17640 -16180
rect 16634 -16214 17640 -16202
rect 17674 -16202 17693 -16180
rect 17757 -15420 17787 -15402
rect 17821 -15420 17888 -15386
rect 17922 -15402 19075 -15386
rect 17922 -15420 17955 -15402
rect 17757 -15476 17955 -15420
rect 17757 -15510 17787 -15476
rect 17821 -15510 17888 -15476
rect 17922 -15510 17955 -15476
rect 17757 -15566 17955 -15510
rect 17757 -15600 17787 -15566
rect 17821 -15600 17888 -15566
rect 17922 -15600 17955 -15566
rect 17757 -15656 17955 -15600
rect 17757 -15690 17787 -15656
rect 17821 -15690 17888 -15656
rect 17922 -15690 17955 -15656
rect 17757 -15746 17955 -15690
rect 17757 -15780 17787 -15746
rect 17821 -15780 17888 -15746
rect 17922 -15780 17955 -15746
rect 17757 -15836 17955 -15780
rect 17757 -15870 17787 -15836
rect 17821 -15870 17888 -15836
rect 17922 -15870 17955 -15836
rect 17757 -15926 17955 -15870
rect 17757 -15960 17787 -15926
rect 17821 -15960 17888 -15926
rect 17922 -15960 17955 -15926
rect 17757 -16016 17955 -15960
rect 17757 -16050 17787 -16016
rect 17821 -16050 17888 -16016
rect 17922 -16050 17955 -16016
rect 17757 -16106 17955 -16050
rect 17757 -16140 17787 -16106
rect 17821 -16140 17888 -16106
rect 17922 -16140 17955 -16106
rect 17757 -16196 17955 -16140
rect 17757 -16202 17787 -16196
rect 17674 -16214 17787 -16202
rect 16634 -16230 17787 -16214
rect 17821 -16230 17888 -16196
rect 17922 -16202 17955 -16196
rect 18019 -15426 18091 -15402
rect 18019 -15460 18038 -15426
rect 18072 -15460 18091 -15426
rect 18019 -15516 18091 -15460
rect 18909 -15460 18981 -15402
rect 18019 -15550 18038 -15516
rect 18072 -15550 18091 -15516
rect 18019 -15606 18091 -15550
rect 18019 -15640 18038 -15606
rect 18072 -15640 18091 -15606
rect 18019 -15696 18091 -15640
rect 18019 -15730 18038 -15696
rect 18072 -15730 18091 -15696
rect 18019 -15786 18091 -15730
rect 18019 -15820 18038 -15786
rect 18072 -15820 18091 -15786
rect 18019 -15876 18091 -15820
rect 18019 -15910 18038 -15876
rect 18072 -15910 18091 -15876
rect 18019 -15966 18091 -15910
rect 18019 -16000 18038 -15966
rect 18072 -16000 18091 -15966
rect 18019 -16056 18091 -16000
rect 18019 -16090 18038 -16056
rect 18072 -16090 18091 -16056
rect 18019 -16146 18091 -16090
rect 18019 -16180 18038 -16146
rect 18072 -16180 18091 -16146
rect 18153 -15524 18847 -15463
rect 18153 -15558 18214 -15524
rect 18248 -15536 18304 -15524
rect 18338 -15536 18394 -15524
rect 18428 -15536 18484 -15524
rect 18260 -15558 18304 -15536
rect 18360 -15558 18394 -15536
rect 18460 -15558 18484 -15536
rect 18518 -15536 18574 -15524
rect 18518 -15558 18526 -15536
rect 18153 -15570 18226 -15558
rect 18260 -15570 18326 -15558
rect 18360 -15570 18426 -15558
rect 18460 -15570 18526 -15558
rect 18560 -15558 18574 -15536
rect 18608 -15536 18664 -15524
rect 18608 -15558 18626 -15536
rect 18560 -15570 18626 -15558
rect 18660 -15558 18664 -15536
rect 18698 -15536 18754 -15524
rect 18698 -15558 18726 -15536
rect 18788 -15558 18847 -15524
rect 18660 -15570 18726 -15558
rect 18760 -15570 18847 -15558
rect 18153 -15614 18847 -15570
rect 18153 -15648 18214 -15614
rect 18248 -15636 18304 -15614
rect 18338 -15636 18394 -15614
rect 18428 -15636 18484 -15614
rect 18260 -15648 18304 -15636
rect 18360 -15648 18394 -15636
rect 18460 -15648 18484 -15636
rect 18518 -15636 18574 -15614
rect 18518 -15648 18526 -15636
rect 18153 -15670 18226 -15648
rect 18260 -15670 18326 -15648
rect 18360 -15670 18426 -15648
rect 18460 -15670 18526 -15648
rect 18560 -15648 18574 -15636
rect 18608 -15636 18664 -15614
rect 18608 -15648 18626 -15636
rect 18560 -15670 18626 -15648
rect 18660 -15648 18664 -15636
rect 18698 -15636 18754 -15614
rect 18698 -15648 18726 -15636
rect 18788 -15648 18847 -15614
rect 18660 -15670 18726 -15648
rect 18760 -15670 18847 -15648
rect 18153 -15704 18847 -15670
rect 18153 -15738 18214 -15704
rect 18248 -15736 18304 -15704
rect 18338 -15736 18394 -15704
rect 18428 -15736 18484 -15704
rect 18260 -15738 18304 -15736
rect 18360 -15738 18394 -15736
rect 18460 -15738 18484 -15736
rect 18518 -15736 18574 -15704
rect 18518 -15738 18526 -15736
rect 18153 -15770 18226 -15738
rect 18260 -15770 18326 -15738
rect 18360 -15770 18426 -15738
rect 18460 -15770 18526 -15738
rect 18560 -15738 18574 -15736
rect 18608 -15736 18664 -15704
rect 18608 -15738 18626 -15736
rect 18560 -15770 18626 -15738
rect 18660 -15738 18664 -15736
rect 18698 -15736 18754 -15704
rect 18698 -15738 18726 -15736
rect 18788 -15738 18847 -15704
rect 18660 -15770 18726 -15738
rect 18760 -15770 18847 -15738
rect 18153 -15794 18847 -15770
rect 18153 -15828 18214 -15794
rect 18248 -15828 18304 -15794
rect 18338 -15828 18394 -15794
rect 18428 -15828 18484 -15794
rect 18518 -15828 18574 -15794
rect 18608 -15828 18664 -15794
rect 18698 -15828 18754 -15794
rect 18788 -15828 18847 -15794
rect 18153 -15836 18847 -15828
rect 18153 -15870 18226 -15836
rect 18260 -15870 18326 -15836
rect 18360 -15870 18426 -15836
rect 18460 -15870 18526 -15836
rect 18560 -15870 18626 -15836
rect 18660 -15870 18726 -15836
rect 18760 -15870 18847 -15836
rect 18153 -15884 18847 -15870
rect 18153 -15918 18214 -15884
rect 18248 -15918 18304 -15884
rect 18338 -15918 18394 -15884
rect 18428 -15918 18484 -15884
rect 18518 -15918 18574 -15884
rect 18608 -15918 18664 -15884
rect 18698 -15918 18754 -15884
rect 18788 -15918 18847 -15884
rect 18153 -15936 18847 -15918
rect 18153 -15970 18226 -15936
rect 18260 -15970 18326 -15936
rect 18360 -15970 18426 -15936
rect 18460 -15970 18526 -15936
rect 18560 -15970 18626 -15936
rect 18660 -15970 18726 -15936
rect 18760 -15970 18847 -15936
rect 18153 -15974 18847 -15970
rect 18153 -16008 18214 -15974
rect 18248 -16008 18304 -15974
rect 18338 -16008 18394 -15974
rect 18428 -16008 18484 -15974
rect 18518 -16008 18574 -15974
rect 18608 -16008 18664 -15974
rect 18698 -16008 18754 -15974
rect 18788 -16008 18847 -15974
rect 18153 -16036 18847 -16008
rect 18153 -16064 18226 -16036
rect 18260 -16064 18326 -16036
rect 18360 -16064 18426 -16036
rect 18460 -16064 18526 -16036
rect 18153 -16098 18214 -16064
rect 18260 -16070 18304 -16064
rect 18360 -16070 18394 -16064
rect 18460 -16070 18484 -16064
rect 18248 -16098 18304 -16070
rect 18338 -16098 18394 -16070
rect 18428 -16098 18484 -16070
rect 18518 -16070 18526 -16064
rect 18560 -16064 18626 -16036
rect 18560 -16070 18574 -16064
rect 18518 -16098 18574 -16070
rect 18608 -16070 18626 -16064
rect 18660 -16064 18726 -16036
rect 18760 -16064 18847 -16036
rect 18660 -16070 18664 -16064
rect 18608 -16098 18664 -16070
rect 18698 -16070 18726 -16064
rect 18698 -16098 18754 -16070
rect 18788 -16098 18847 -16064
rect 18153 -16157 18847 -16098
rect 18909 -15494 18928 -15460
rect 18962 -15494 18981 -15460
rect 18909 -15550 18981 -15494
rect 18909 -15584 18928 -15550
rect 18962 -15584 18981 -15550
rect 18909 -15640 18981 -15584
rect 18909 -15674 18928 -15640
rect 18962 -15674 18981 -15640
rect 18909 -15730 18981 -15674
rect 18909 -15764 18928 -15730
rect 18962 -15764 18981 -15730
rect 18909 -15820 18981 -15764
rect 18909 -15854 18928 -15820
rect 18962 -15854 18981 -15820
rect 18909 -15910 18981 -15854
rect 18909 -15944 18928 -15910
rect 18962 -15944 18981 -15910
rect 18909 -16000 18981 -15944
rect 18909 -16034 18928 -16000
rect 18962 -16034 18981 -16000
rect 18909 -16090 18981 -16034
rect 18909 -16124 18928 -16090
rect 18962 -16124 18981 -16090
rect 18019 -16202 18091 -16180
rect 18909 -16180 18981 -16124
rect 18909 -16202 18928 -16180
rect 17922 -16214 18928 -16202
rect 18962 -16202 18981 -16180
rect 19045 -15420 19075 -15402
rect 19109 -15420 19176 -15386
rect 19210 -15402 20363 -15386
rect 19210 -15420 19243 -15402
rect 19045 -15476 19243 -15420
rect 19045 -15510 19075 -15476
rect 19109 -15510 19176 -15476
rect 19210 -15510 19243 -15476
rect 19045 -15566 19243 -15510
rect 19045 -15600 19075 -15566
rect 19109 -15600 19176 -15566
rect 19210 -15600 19243 -15566
rect 19045 -15656 19243 -15600
rect 19045 -15690 19075 -15656
rect 19109 -15690 19176 -15656
rect 19210 -15690 19243 -15656
rect 19045 -15746 19243 -15690
rect 19045 -15780 19075 -15746
rect 19109 -15780 19176 -15746
rect 19210 -15780 19243 -15746
rect 19045 -15836 19243 -15780
rect 19045 -15870 19075 -15836
rect 19109 -15870 19176 -15836
rect 19210 -15870 19243 -15836
rect 19045 -15926 19243 -15870
rect 19045 -15960 19075 -15926
rect 19109 -15960 19176 -15926
rect 19210 -15960 19243 -15926
rect 19045 -16016 19243 -15960
rect 19045 -16050 19075 -16016
rect 19109 -16050 19176 -16016
rect 19210 -16050 19243 -16016
rect 19045 -16106 19243 -16050
rect 19045 -16140 19075 -16106
rect 19109 -16140 19176 -16106
rect 19210 -16140 19243 -16106
rect 19045 -16196 19243 -16140
rect 19045 -16202 19075 -16196
rect 18962 -16214 19075 -16202
rect 17922 -16230 19075 -16214
rect 19109 -16230 19176 -16196
rect 19210 -16202 19243 -16196
rect 19307 -15426 19379 -15402
rect 19307 -15460 19326 -15426
rect 19360 -15460 19379 -15426
rect 19307 -15516 19379 -15460
rect 20197 -15460 20269 -15402
rect 19307 -15550 19326 -15516
rect 19360 -15550 19379 -15516
rect 19307 -15606 19379 -15550
rect 19307 -15640 19326 -15606
rect 19360 -15640 19379 -15606
rect 19307 -15696 19379 -15640
rect 19307 -15730 19326 -15696
rect 19360 -15730 19379 -15696
rect 19307 -15786 19379 -15730
rect 19307 -15820 19326 -15786
rect 19360 -15820 19379 -15786
rect 19307 -15876 19379 -15820
rect 19307 -15910 19326 -15876
rect 19360 -15910 19379 -15876
rect 19307 -15966 19379 -15910
rect 19307 -16000 19326 -15966
rect 19360 -16000 19379 -15966
rect 19307 -16056 19379 -16000
rect 19307 -16090 19326 -16056
rect 19360 -16090 19379 -16056
rect 19307 -16146 19379 -16090
rect 19307 -16180 19326 -16146
rect 19360 -16180 19379 -16146
rect 19441 -15524 20135 -15463
rect 19441 -15558 19502 -15524
rect 19536 -15536 19592 -15524
rect 19626 -15536 19682 -15524
rect 19716 -15536 19772 -15524
rect 19548 -15558 19592 -15536
rect 19648 -15558 19682 -15536
rect 19748 -15558 19772 -15536
rect 19806 -15536 19862 -15524
rect 19806 -15558 19814 -15536
rect 19441 -15570 19514 -15558
rect 19548 -15570 19614 -15558
rect 19648 -15570 19714 -15558
rect 19748 -15570 19814 -15558
rect 19848 -15558 19862 -15536
rect 19896 -15536 19952 -15524
rect 19896 -15558 19914 -15536
rect 19848 -15570 19914 -15558
rect 19948 -15558 19952 -15536
rect 19986 -15536 20042 -15524
rect 19986 -15558 20014 -15536
rect 20076 -15558 20135 -15524
rect 19948 -15570 20014 -15558
rect 20048 -15570 20135 -15558
rect 19441 -15614 20135 -15570
rect 19441 -15648 19502 -15614
rect 19536 -15636 19592 -15614
rect 19626 -15636 19682 -15614
rect 19716 -15636 19772 -15614
rect 19548 -15648 19592 -15636
rect 19648 -15648 19682 -15636
rect 19748 -15648 19772 -15636
rect 19806 -15636 19862 -15614
rect 19806 -15648 19814 -15636
rect 19441 -15670 19514 -15648
rect 19548 -15670 19614 -15648
rect 19648 -15670 19714 -15648
rect 19748 -15670 19814 -15648
rect 19848 -15648 19862 -15636
rect 19896 -15636 19952 -15614
rect 19896 -15648 19914 -15636
rect 19848 -15670 19914 -15648
rect 19948 -15648 19952 -15636
rect 19986 -15636 20042 -15614
rect 19986 -15648 20014 -15636
rect 20076 -15648 20135 -15614
rect 19948 -15670 20014 -15648
rect 20048 -15670 20135 -15648
rect 19441 -15704 20135 -15670
rect 19441 -15738 19502 -15704
rect 19536 -15736 19592 -15704
rect 19626 -15736 19682 -15704
rect 19716 -15736 19772 -15704
rect 19548 -15738 19592 -15736
rect 19648 -15738 19682 -15736
rect 19748 -15738 19772 -15736
rect 19806 -15736 19862 -15704
rect 19806 -15738 19814 -15736
rect 19441 -15770 19514 -15738
rect 19548 -15770 19614 -15738
rect 19648 -15770 19714 -15738
rect 19748 -15770 19814 -15738
rect 19848 -15738 19862 -15736
rect 19896 -15736 19952 -15704
rect 19896 -15738 19914 -15736
rect 19848 -15770 19914 -15738
rect 19948 -15738 19952 -15736
rect 19986 -15736 20042 -15704
rect 19986 -15738 20014 -15736
rect 20076 -15738 20135 -15704
rect 19948 -15770 20014 -15738
rect 20048 -15770 20135 -15738
rect 19441 -15794 20135 -15770
rect 19441 -15828 19502 -15794
rect 19536 -15828 19592 -15794
rect 19626 -15828 19682 -15794
rect 19716 -15828 19772 -15794
rect 19806 -15828 19862 -15794
rect 19896 -15828 19952 -15794
rect 19986 -15828 20042 -15794
rect 20076 -15828 20135 -15794
rect 19441 -15836 20135 -15828
rect 19441 -15870 19514 -15836
rect 19548 -15870 19614 -15836
rect 19648 -15870 19714 -15836
rect 19748 -15870 19814 -15836
rect 19848 -15870 19914 -15836
rect 19948 -15870 20014 -15836
rect 20048 -15870 20135 -15836
rect 19441 -15884 20135 -15870
rect 19441 -15918 19502 -15884
rect 19536 -15918 19592 -15884
rect 19626 -15918 19682 -15884
rect 19716 -15918 19772 -15884
rect 19806 -15918 19862 -15884
rect 19896 -15918 19952 -15884
rect 19986 -15918 20042 -15884
rect 20076 -15918 20135 -15884
rect 19441 -15936 20135 -15918
rect 19441 -15970 19514 -15936
rect 19548 -15970 19614 -15936
rect 19648 -15970 19714 -15936
rect 19748 -15970 19814 -15936
rect 19848 -15970 19914 -15936
rect 19948 -15970 20014 -15936
rect 20048 -15970 20135 -15936
rect 19441 -15974 20135 -15970
rect 19441 -16008 19502 -15974
rect 19536 -16008 19592 -15974
rect 19626 -16008 19682 -15974
rect 19716 -16008 19772 -15974
rect 19806 -16008 19862 -15974
rect 19896 -16008 19952 -15974
rect 19986 -16008 20042 -15974
rect 20076 -16008 20135 -15974
rect 19441 -16036 20135 -16008
rect 19441 -16064 19514 -16036
rect 19548 -16064 19614 -16036
rect 19648 -16064 19714 -16036
rect 19748 -16064 19814 -16036
rect 19441 -16098 19502 -16064
rect 19548 -16070 19592 -16064
rect 19648 -16070 19682 -16064
rect 19748 -16070 19772 -16064
rect 19536 -16098 19592 -16070
rect 19626 -16098 19682 -16070
rect 19716 -16098 19772 -16070
rect 19806 -16070 19814 -16064
rect 19848 -16064 19914 -16036
rect 19848 -16070 19862 -16064
rect 19806 -16098 19862 -16070
rect 19896 -16070 19914 -16064
rect 19948 -16064 20014 -16036
rect 20048 -16064 20135 -16036
rect 19948 -16070 19952 -16064
rect 19896 -16098 19952 -16070
rect 19986 -16070 20014 -16064
rect 19986 -16098 20042 -16070
rect 20076 -16098 20135 -16064
rect 19441 -16157 20135 -16098
rect 20197 -15494 20216 -15460
rect 20250 -15494 20269 -15460
rect 20197 -15550 20269 -15494
rect 20197 -15584 20216 -15550
rect 20250 -15584 20269 -15550
rect 20197 -15640 20269 -15584
rect 20197 -15674 20216 -15640
rect 20250 -15674 20269 -15640
rect 20197 -15730 20269 -15674
rect 20197 -15764 20216 -15730
rect 20250 -15764 20269 -15730
rect 20197 -15820 20269 -15764
rect 20197 -15854 20216 -15820
rect 20250 -15854 20269 -15820
rect 20197 -15910 20269 -15854
rect 20197 -15944 20216 -15910
rect 20250 -15944 20269 -15910
rect 20197 -16000 20269 -15944
rect 20197 -16034 20216 -16000
rect 20250 -16034 20269 -16000
rect 20197 -16090 20269 -16034
rect 20197 -16124 20216 -16090
rect 20250 -16124 20269 -16090
rect 19307 -16202 19379 -16180
rect 20197 -16180 20269 -16124
rect 20197 -16202 20216 -16180
rect 19210 -16214 20216 -16202
rect 20250 -16202 20269 -16180
rect 20333 -15420 20363 -15402
rect 20397 -15420 20464 -15386
rect 20498 -15402 21651 -15386
rect 20498 -15420 20531 -15402
rect 20333 -15476 20531 -15420
rect 20333 -15510 20363 -15476
rect 20397 -15510 20464 -15476
rect 20498 -15510 20531 -15476
rect 20333 -15566 20531 -15510
rect 20333 -15600 20363 -15566
rect 20397 -15600 20464 -15566
rect 20498 -15600 20531 -15566
rect 20333 -15656 20531 -15600
rect 20333 -15690 20363 -15656
rect 20397 -15690 20464 -15656
rect 20498 -15690 20531 -15656
rect 20333 -15746 20531 -15690
rect 20333 -15780 20363 -15746
rect 20397 -15780 20464 -15746
rect 20498 -15780 20531 -15746
rect 20333 -15836 20531 -15780
rect 20333 -15870 20363 -15836
rect 20397 -15870 20464 -15836
rect 20498 -15870 20531 -15836
rect 20333 -15926 20531 -15870
rect 20333 -15960 20363 -15926
rect 20397 -15960 20464 -15926
rect 20498 -15960 20531 -15926
rect 20333 -16016 20531 -15960
rect 20333 -16050 20363 -16016
rect 20397 -16050 20464 -16016
rect 20498 -16050 20531 -16016
rect 20333 -16106 20531 -16050
rect 20333 -16140 20363 -16106
rect 20397 -16140 20464 -16106
rect 20498 -16140 20531 -16106
rect 20333 -16196 20531 -16140
rect 20333 -16202 20363 -16196
rect 20250 -16214 20363 -16202
rect 19210 -16230 20363 -16214
rect 20397 -16230 20464 -16196
rect 20498 -16202 20531 -16196
rect 20595 -15426 20667 -15402
rect 20595 -15460 20614 -15426
rect 20648 -15460 20667 -15426
rect 20595 -15516 20667 -15460
rect 21485 -15460 21557 -15402
rect 20595 -15550 20614 -15516
rect 20648 -15550 20667 -15516
rect 20595 -15606 20667 -15550
rect 20595 -15640 20614 -15606
rect 20648 -15640 20667 -15606
rect 20595 -15696 20667 -15640
rect 20595 -15730 20614 -15696
rect 20648 -15730 20667 -15696
rect 20595 -15786 20667 -15730
rect 20595 -15820 20614 -15786
rect 20648 -15820 20667 -15786
rect 20595 -15876 20667 -15820
rect 20595 -15910 20614 -15876
rect 20648 -15910 20667 -15876
rect 20595 -15966 20667 -15910
rect 20595 -16000 20614 -15966
rect 20648 -16000 20667 -15966
rect 20595 -16056 20667 -16000
rect 20595 -16090 20614 -16056
rect 20648 -16090 20667 -16056
rect 20595 -16146 20667 -16090
rect 20595 -16180 20614 -16146
rect 20648 -16180 20667 -16146
rect 20729 -15524 21423 -15463
rect 20729 -15558 20790 -15524
rect 20824 -15536 20880 -15524
rect 20914 -15536 20970 -15524
rect 21004 -15536 21060 -15524
rect 20836 -15558 20880 -15536
rect 20936 -15558 20970 -15536
rect 21036 -15558 21060 -15536
rect 21094 -15536 21150 -15524
rect 21094 -15558 21102 -15536
rect 20729 -15570 20802 -15558
rect 20836 -15570 20902 -15558
rect 20936 -15570 21002 -15558
rect 21036 -15570 21102 -15558
rect 21136 -15558 21150 -15536
rect 21184 -15536 21240 -15524
rect 21184 -15558 21202 -15536
rect 21136 -15570 21202 -15558
rect 21236 -15558 21240 -15536
rect 21274 -15536 21330 -15524
rect 21274 -15558 21302 -15536
rect 21364 -15558 21423 -15524
rect 21236 -15570 21302 -15558
rect 21336 -15570 21423 -15558
rect 20729 -15614 21423 -15570
rect 20729 -15648 20790 -15614
rect 20824 -15636 20880 -15614
rect 20914 -15636 20970 -15614
rect 21004 -15636 21060 -15614
rect 20836 -15648 20880 -15636
rect 20936 -15648 20970 -15636
rect 21036 -15648 21060 -15636
rect 21094 -15636 21150 -15614
rect 21094 -15648 21102 -15636
rect 20729 -15670 20802 -15648
rect 20836 -15670 20902 -15648
rect 20936 -15670 21002 -15648
rect 21036 -15670 21102 -15648
rect 21136 -15648 21150 -15636
rect 21184 -15636 21240 -15614
rect 21184 -15648 21202 -15636
rect 21136 -15670 21202 -15648
rect 21236 -15648 21240 -15636
rect 21274 -15636 21330 -15614
rect 21274 -15648 21302 -15636
rect 21364 -15648 21423 -15614
rect 21236 -15670 21302 -15648
rect 21336 -15670 21423 -15648
rect 20729 -15704 21423 -15670
rect 20729 -15738 20790 -15704
rect 20824 -15736 20880 -15704
rect 20914 -15736 20970 -15704
rect 21004 -15736 21060 -15704
rect 20836 -15738 20880 -15736
rect 20936 -15738 20970 -15736
rect 21036 -15738 21060 -15736
rect 21094 -15736 21150 -15704
rect 21094 -15738 21102 -15736
rect 20729 -15770 20802 -15738
rect 20836 -15770 20902 -15738
rect 20936 -15770 21002 -15738
rect 21036 -15770 21102 -15738
rect 21136 -15738 21150 -15736
rect 21184 -15736 21240 -15704
rect 21184 -15738 21202 -15736
rect 21136 -15770 21202 -15738
rect 21236 -15738 21240 -15736
rect 21274 -15736 21330 -15704
rect 21274 -15738 21302 -15736
rect 21364 -15738 21423 -15704
rect 21236 -15770 21302 -15738
rect 21336 -15770 21423 -15738
rect 20729 -15794 21423 -15770
rect 20729 -15828 20790 -15794
rect 20824 -15828 20880 -15794
rect 20914 -15828 20970 -15794
rect 21004 -15828 21060 -15794
rect 21094 -15828 21150 -15794
rect 21184 -15828 21240 -15794
rect 21274 -15828 21330 -15794
rect 21364 -15828 21423 -15794
rect 20729 -15836 21423 -15828
rect 20729 -15870 20802 -15836
rect 20836 -15870 20902 -15836
rect 20936 -15870 21002 -15836
rect 21036 -15870 21102 -15836
rect 21136 -15870 21202 -15836
rect 21236 -15870 21302 -15836
rect 21336 -15870 21423 -15836
rect 20729 -15884 21423 -15870
rect 20729 -15918 20790 -15884
rect 20824 -15918 20880 -15884
rect 20914 -15918 20970 -15884
rect 21004 -15918 21060 -15884
rect 21094 -15918 21150 -15884
rect 21184 -15918 21240 -15884
rect 21274 -15918 21330 -15884
rect 21364 -15918 21423 -15884
rect 20729 -15936 21423 -15918
rect 20729 -15970 20802 -15936
rect 20836 -15970 20902 -15936
rect 20936 -15970 21002 -15936
rect 21036 -15970 21102 -15936
rect 21136 -15970 21202 -15936
rect 21236 -15970 21302 -15936
rect 21336 -15970 21423 -15936
rect 20729 -15974 21423 -15970
rect 20729 -16008 20790 -15974
rect 20824 -16008 20880 -15974
rect 20914 -16008 20970 -15974
rect 21004 -16008 21060 -15974
rect 21094 -16008 21150 -15974
rect 21184 -16008 21240 -15974
rect 21274 -16008 21330 -15974
rect 21364 -16008 21423 -15974
rect 20729 -16036 21423 -16008
rect 20729 -16064 20802 -16036
rect 20836 -16064 20902 -16036
rect 20936 -16064 21002 -16036
rect 21036 -16064 21102 -16036
rect 20729 -16098 20790 -16064
rect 20836 -16070 20880 -16064
rect 20936 -16070 20970 -16064
rect 21036 -16070 21060 -16064
rect 20824 -16098 20880 -16070
rect 20914 -16098 20970 -16070
rect 21004 -16098 21060 -16070
rect 21094 -16070 21102 -16064
rect 21136 -16064 21202 -16036
rect 21136 -16070 21150 -16064
rect 21094 -16098 21150 -16070
rect 21184 -16070 21202 -16064
rect 21236 -16064 21302 -16036
rect 21336 -16064 21423 -16036
rect 21236 -16070 21240 -16064
rect 21184 -16098 21240 -16070
rect 21274 -16070 21302 -16064
rect 21274 -16098 21330 -16070
rect 21364 -16098 21423 -16064
rect 20729 -16157 21423 -16098
rect 21485 -15494 21504 -15460
rect 21538 -15494 21557 -15460
rect 21485 -15550 21557 -15494
rect 21485 -15584 21504 -15550
rect 21538 -15584 21557 -15550
rect 21485 -15640 21557 -15584
rect 21485 -15674 21504 -15640
rect 21538 -15674 21557 -15640
rect 21485 -15730 21557 -15674
rect 21485 -15764 21504 -15730
rect 21538 -15764 21557 -15730
rect 21485 -15820 21557 -15764
rect 21485 -15854 21504 -15820
rect 21538 -15854 21557 -15820
rect 21485 -15910 21557 -15854
rect 21485 -15944 21504 -15910
rect 21538 -15944 21557 -15910
rect 21485 -16000 21557 -15944
rect 21485 -16034 21504 -16000
rect 21538 -16034 21557 -16000
rect 21485 -16090 21557 -16034
rect 21485 -16124 21504 -16090
rect 21538 -16124 21557 -16090
rect 20595 -16202 20667 -16180
rect 21485 -16180 21557 -16124
rect 21485 -16202 21504 -16180
rect 20498 -16214 21504 -16202
rect 21538 -16202 21557 -16180
rect 21621 -15420 21651 -15402
rect 21685 -15420 21752 -15386
rect 21786 -15402 22939 -15386
rect 21786 -15420 21819 -15402
rect 21621 -15476 21819 -15420
rect 21621 -15510 21651 -15476
rect 21685 -15510 21752 -15476
rect 21786 -15510 21819 -15476
rect 21621 -15566 21819 -15510
rect 21621 -15600 21651 -15566
rect 21685 -15600 21752 -15566
rect 21786 -15600 21819 -15566
rect 21621 -15656 21819 -15600
rect 21621 -15690 21651 -15656
rect 21685 -15690 21752 -15656
rect 21786 -15690 21819 -15656
rect 21621 -15746 21819 -15690
rect 21621 -15780 21651 -15746
rect 21685 -15780 21752 -15746
rect 21786 -15780 21819 -15746
rect 21621 -15836 21819 -15780
rect 21621 -15870 21651 -15836
rect 21685 -15870 21752 -15836
rect 21786 -15870 21819 -15836
rect 21621 -15926 21819 -15870
rect 21621 -15960 21651 -15926
rect 21685 -15960 21752 -15926
rect 21786 -15960 21819 -15926
rect 21621 -16016 21819 -15960
rect 21621 -16050 21651 -16016
rect 21685 -16050 21752 -16016
rect 21786 -16050 21819 -16016
rect 21621 -16106 21819 -16050
rect 21621 -16140 21651 -16106
rect 21685 -16140 21752 -16106
rect 21786 -16140 21819 -16106
rect 21621 -16196 21819 -16140
rect 21621 -16202 21651 -16196
rect 21538 -16214 21651 -16202
rect 20498 -16230 21651 -16214
rect 21685 -16230 21752 -16196
rect 21786 -16202 21819 -16196
rect 21883 -15426 21955 -15402
rect 21883 -15460 21902 -15426
rect 21936 -15460 21955 -15426
rect 21883 -15516 21955 -15460
rect 22773 -15460 22845 -15402
rect 21883 -15550 21902 -15516
rect 21936 -15550 21955 -15516
rect 21883 -15606 21955 -15550
rect 21883 -15640 21902 -15606
rect 21936 -15640 21955 -15606
rect 21883 -15696 21955 -15640
rect 21883 -15730 21902 -15696
rect 21936 -15730 21955 -15696
rect 21883 -15786 21955 -15730
rect 21883 -15820 21902 -15786
rect 21936 -15820 21955 -15786
rect 21883 -15876 21955 -15820
rect 21883 -15910 21902 -15876
rect 21936 -15910 21955 -15876
rect 21883 -15966 21955 -15910
rect 21883 -16000 21902 -15966
rect 21936 -16000 21955 -15966
rect 21883 -16056 21955 -16000
rect 21883 -16090 21902 -16056
rect 21936 -16090 21955 -16056
rect 21883 -16146 21955 -16090
rect 21883 -16180 21902 -16146
rect 21936 -16180 21955 -16146
rect 22017 -15524 22711 -15463
rect 22017 -15558 22078 -15524
rect 22112 -15536 22168 -15524
rect 22202 -15536 22258 -15524
rect 22292 -15536 22348 -15524
rect 22124 -15558 22168 -15536
rect 22224 -15558 22258 -15536
rect 22324 -15558 22348 -15536
rect 22382 -15536 22438 -15524
rect 22382 -15558 22390 -15536
rect 22017 -15570 22090 -15558
rect 22124 -15570 22190 -15558
rect 22224 -15570 22290 -15558
rect 22324 -15570 22390 -15558
rect 22424 -15558 22438 -15536
rect 22472 -15536 22528 -15524
rect 22472 -15558 22490 -15536
rect 22424 -15570 22490 -15558
rect 22524 -15558 22528 -15536
rect 22562 -15536 22618 -15524
rect 22562 -15558 22590 -15536
rect 22652 -15558 22711 -15524
rect 22524 -15570 22590 -15558
rect 22624 -15570 22711 -15558
rect 22017 -15614 22711 -15570
rect 22017 -15648 22078 -15614
rect 22112 -15636 22168 -15614
rect 22202 -15636 22258 -15614
rect 22292 -15636 22348 -15614
rect 22124 -15648 22168 -15636
rect 22224 -15648 22258 -15636
rect 22324 -15648 22348 -15636
rect 22382 -15636 22438 -15614
rect 22382 -15648 22390 -15636
rect 22017 -15670 22090 -15648
rect 22124 -15670 22190 -15648
rect 22224 -15670 22290 -15648
rect 22324 -15670 22390 -15648
rect 22424 -15648 22438 -15636
rect 22472 -15636 22528 -15614
rect 22472 -15648 22490 -15636
rect 22424 -15670 22490 -15648
rect 22524 -15648 22528 -15636
rect 22562 -15636 22618 -15614
rect 22562 -15648 22590 -15636
rect 22652 -15648 22711 -15614
rect 22524 -15670 22590 -15648
rect 22624 -15670 22711 -15648
rect 22017 -15704 22711 -15670
rect 22017 -15738 22078 -15704
rect 22112 -15736 22168 -15704
rect 22202 -15736 22258 -15704
rect 22292 -15736 22348 -15704
rect 22124 -15738 22168 -15736
rect 22224 -15738 22258 -15736
rect 22324 -15738 22348 -15736
rect 22382 -15736 22438 -15704
rect 22382 -15738 22390 -15736
rect 22017 -15770 22090 -15738
rect 22124 -15770 22190 -15738
rect 22224 -15770 22290 -15738
rect 22324 -15770 22390 -15738
rect 22424 -15738 22438 -15736
rect 22472 -15736 22528 -15704
rect 22472 -15738 22490 -15736
rect 22424 -15770 22490 -15738
rect 22524 -15738 22528 -15736
rect 22562 -15736 22618 -15704
rect 22562 -15738 22590 -15736
rect 22652 -15738 22711 -15704
rect 22524 -15770 22590 -15738
rect 22624 -15770 22711 -15738
rect 22017 -15794 22711 -15770
rect 22017 -15828 22078 -15794
rect 22112 -15828 22168 -15794
rect 22202 -15828 22258 -15794
rect 22292 -15828 22348 -15794
rect 22382 -15828 22438 -15794
rect 22472 -15828 22528 -15794
rect 22562 -15828 22618 -15794
rect 22652 -15828 22711 -15794
rect 22017 -15836 22711 -15828
rect 22017 -15870 22090 -15836
rect 22124 -15870 22190 -15836
rect 22224 -15870 22290 -15836
rect 22324 -15870 22390 -15836
rect 22424 -15870 22490 -15836
rect 22524 -15870 22590 -15836
rect 22624 -15870 22711 -15836
rect 22017 -15884 22711 -15870
rect 22017 -15918 22078 -15884
rect 22112 -15918 22168 -15884
rect 22202 -15918 22258 -15884
rect 22292 -15918 22348 -15884
rect 22382 -15918 22438 -15884
rect 22472 -15918 22528 -15884
rect 22562 -15918 22618 -15884
rect 22652 -15918 22711 -15884
rect 22017 -15936 22711 -15918
rect 22017 -15970 22090 -15936
rect 22124 -15970 22190 -15936
rect 22224 -15970 22290 -15936
rect 22324 -15970 22390 -15936
rect 22424 -15970 22490 -15936
rect 22524 -15970 22590 -15936
rect 22624 -15970 22711 -15936
rect 22017 -15974 22711 -15970
rect 22017 -16008 22078 -15974
rect 22112 -16008 22168 -15974
rect 22202 -16008 22258 -15974
rect 22292 -16008 22348 -15974
rect 22382 -16008 22438 -15974
rect 22472 -16008 22528 -15974
rect 22562 -16008 22618 -15974
rect 22652 -16008 22711 -15974
rect 22017 -16036 22711 -16008
rect 22017 -16064 22090 -16036
rect 22124 -16064 22190 -16036
rect 22224 -16064 22290 -16036
rect 22324 -16064 22390 -16036
rect 22017 -16098 22078 -16064
rect 22124 -16070 22168 -16064
rect 22224 -16070 22258 -16064
rect 22324 -16070 22348 -16064
rect 22112 -16098 22168 -16070
rect 22202 -16098 22258 -16070
rect 22292 -16098 22348 -16070
rect 22382 -16070 22390 -16064
rect 22424 -16064 22490 -16036
rect 22424 -16070 22438 -16064
rect 22382 -16098 22438 -16070
rect 22472 -16070 22490 -16064
rect 22524 -16064 22590 -16036
rect 22624 -16064 22711 -16036
rect 22524 -16070 22528 -16064
rect 22472 -16098 22528 -16070
rect 22562 -16070 22590 -16064
rect 22562 -16098 22618 -16070
rect 22652 -16098 22711 -16064
rect 22017 -16157 22711 -16098
rect 22773 -15494 22792 -15460
rect 22826 -15494 22845 -15460
rect 22773 -15550 22845 -15494
rect 22773 -15584 22792 -15550
rect 22826 -15584 22845 -15550
rect 22773 -15640 22845 -15584
rect 22773 -15674 22792 -15640
rect 22826 -15674 22845 -15640
rect 22773 -15730 22845 -15674
rect 22773 -15764 22792 -15730
rect 22826 -15764 22845 -15730
rect 22773 -15820 22845 -15764
rect 22773 -15854 22792 -15820
rect 22826 -15854 22845 -15820
rect 22773 -15910 22845 -15854
rect 22773 -15944 22792 -15910
rect 22826 -15944 22845 -15910
rect 22773 -16000 22845 -15944
rect 22773 -16034 22792 -16000
rect 22826 -16034 22845 -16000
rect 22773 -16090 22845 -16034
rect 22773 -16124 22792 -16090
rect 22826 -16124 22845 -16090
rect 21883 -16202 21955 -16180
rect 22773 -16180 22845 -16124
rect 22773 -16202 22792 -16180
rect 21786 -16214 22792 -16202
rect 22826 -16202 22845 -16180
rect 22909 -15420 22939 -15402
rect 22973 -15420 23040 -15386
rect 23074 -15402 24227 -15386
rect 23074 -15420 23107 -15402
rect 22909 -15476 23107 -15420
rect 22909 -15510 22939 -15476
rect 22973 -15510 23040 -15476
rect 23074 -15510 23107 -15476
rect 22909 -15566 23107 -15510
rect 22909 -15600 22939 -15566
rect 22973 -15600 23040 -15566
rect 23074 -15600 23107 -15566
rect 22909 -15656 23107 -15600
rect 22909 -15690 22939 -15656
rect 22973 -15690 23040 -15656
rect 23074 -15690 23107 -15656
rect 22909 -15746 23107 -15690
rect 22909 -15780 22939 -15746
rect 22973 -15780 23040 -15746
rect 23074 -15780 23107 -15746
rect 22909 -15836 23107 -15780
rect 22909 -15870 22939 -15836
rect 22973 -15870 23040 -15836
rect 23074 -15870 23107 -15836
rect 22909 -15926 23107 -15870
rect 22909 -15960 22939 -15926
rect 22973 -15960 23040 -15926
rect 23074 -15960 23107 -15926
rect 22909 -16016 23107 -15960
rect 22909 -16050 22939 -16016
rect 22973 -16050 23040 -16016
rect 23074 -16050 23107 -16016
rect 22909 -16106 23107 -16050
rect 22909 -16140 22939 -16106
rect 22973 -16140 23040 -16106
rect 23074 -16140 23107 -16106
rect 22909 -16196 23107 -16140
rect 22909 -16202 22939 -16196
rect 22826 -16214 22939 -16202
rect 21786 -16230 22939 -16214
rect 22973 -16230 23040 -16196
rect 23074 -16202 23107 -16196
rect 23171 -15426 23243 -15402
rect 23171 -15460 23190 -15426
rect 23224 -15460 23243 -15426
rect 23171 -15516 23243 -15460
rect 24061 -15460 24133 -15402
rect 23171 -15550 23190 -15516
rect 23224 -15550 23243 -15516
rect 23171 -15606 23243 -15550
rect 23171 -15640 23190 -15606
rect 23224 -15640 23243 -15606
rect 23171 -15696 23243 -15640
rect 23171 -15730 23190 -15696
rect 23224 -15730 23243 -15696
rect 23171 -15786 23243 -15730
rect 23171 -15820 23190 -15786
rect 23224 -15820 23243 -15786
rect 23171 -15876 23243 -15820
rect 23171 -15910 23190 -15876
rect 23224 -15910 23243 -15876
rect 23171 -15966 23243 -15910
rect 23171 -16000 23190 -15966
rect 23224 -16000 23243 -15966
rect 23171 -16056 23243 -16000
rect 23171 -16090 23190 -16056
rect 23224 -16090 23243 -16056
rect 23171 -16146 23243 -16090
rect 23171 -16180 23190 -16146
rect 23224 -16180 23243 -16146
rect 23305 -15524 23999 -15463
rect 23305 -15558 23366 -15524
rect 23400 -15536 23456 -15524
rect 23490 -15536 23546 -15524
rect 23580 -15536 23636 -15524
rect 23412 -15558 23456 -15536
rect 23512 -15558 23546 -15536
rect 23612 -15558 23636 -15536
rect 23670 -15536 23726 -15524
rect 23670 -15558 23678 -15536
rect 23305 -15570 23378 -15558
rect 23412 -15570 23478 -15558
rect 23512 -15570 23578 -15558
rect 23612 -15570 23678 -15558
rect 23712 -15558 23726 -15536
rect 23760 -15536 23816 -15524
rect 23760 -15558 23778 -15536
rect 23712 -15570 23778 -15558
rect 23812 -15558 23816 -15536
rect 23850 -15536 23906 -15524
rect 23850 -15558 23878 -15536
rect 23940 -15558 23999 -15524
rect 23812 -15570 23878 -15558
rect 23912 -15570 23999 -15558
rect 23305 -15614 23999 -15570
rect 23305 -15648 23366 -15614
rect 23400 -15636 23456 -15614
rect 23490 -15636 23546 -15614
rect 23580 -15636 23636 -15614
rect 23412 -15648 23456 -15636
rect 23512 -15648 23546 -15636
rect 23612 -15648 23636 -15636
rect 23670 -15636 23726 -15614
rect 23670 -15648 23678 -15636
rect 23305 -15670 23378 -15648
rect 23412 -15670 23478 -15648
rect 23512 -15670 23578 -15648
rect 23612 -15670 23678 -15648
rect 23712 -15648 23726 -15636
rect 23760 -15636 23816 -15614
rect 23760 -15648 23778 -15636
rect 23712 -15670 23778 -15648
rect 23812 -15648 23816 -15636
rect 23850 -15636 23906 -15614
rect 23850 -15648 23878 -15636
rect 23940 -15648 23999 -15614
rect 23812 -15670 23878 -15648
rect 23912 -15670 23999 -15648
rect 23305 -15704 23999 -15670
rect 23305 -15738 23366 -15704
rect 23400 -15736 23456 -15704
rect 23490 -15736 23546 -15704
rect 23580 -15736 23636 -15704
rect 23412 -15738 23456 -15736
rect 23512 -15738 23546 -15736
rect 23612 -15738 23636 -15736
rect 23670 -15736 23726 -15704
rect 23670 -15738 23678 -15736
rect 23305 -15770 23378 -15738
rect 23412 -15770 23478 -15738
rect 23512 -15770 23578 -15738
rect 23612 -15770 23678 -15738
rect 23712 -15738 23726 -15736
rect 23760 -15736 23816 -15704
rect 23760 -15738 23778 -15736
rect 23712 -15770 23778 -15738
rect 23812 -15738 23816 -15736
rect 23850 -15736 23906 -15704
rect 23850 -15738 23878 -15736
rect 23940 -15738 23999 -15704
rect 23812 -15770 23878 -15738
rect 23912 -15770 23999 -15738
rect 23305 -15794 23999 -15770
rect 23305 -15828 23366 -15794
rect 23400 -15828 23456 -15794
rect 23490 -15828 23546 -15794
rect 23580 -15828 23636 -15794
rect 23670 -15828 23726 -15794
rect 23760 -15828 23816 -15794
rect 23850 -15828 23906 -15794
rect 23940 -15828 23999 -15794
rect 23305 -15836 23999 -15828
rect 23305 -15870 23378 -15836
rect 23412 -15870 23478 -15836
rect 23512 -15870 23578 -15836
rect 23612 -15870 23678 -15836
rect 23712 -15870 23778 -15836
rect 23812 -15870 23878 -15836
rect 23912 -15870 23999 -15836
rect 23305 -15884 23999 -15870
rect 23305 -15918 23366 -15884
rect 23400 -15918 23456 -15884
rect 23490 -15918 23546 -15884
rect 23580 -15918 23636 -15884
rect 23670 -15918 23726 -15884
rect 23760 -15918 23816 -15884
rect 23850 -15918 23906 -15884
rect 23940 -15918 23999 -15884
rect 23305 -15936 23999 -15918
rect 23305 -15970 23378 -15936
rect 23412 -15970 23478 -15936
rect 23512 -15970 23578 -15936
rect 23612 -15970 23678 -15936
rect 23712 -15970 23778 -15936
rect 23812 -15970 23878 -15936
rect 23912 -15970 23999 -15936
rect 23305 -15974 23999 -15970
rect 23305 -16008 23366 -15974
rect 23400 -16008 23456 -15974
rect 23490 -16008 23546 -15974
rect 23580 -16008 23636 -15974
rect 23670 -16008 23726 -15974
rect 23760 -16008 23816 -15974
rect 23850 -16008 23906 -15974
rect 23940 -16008 23999 -15974
rect 23305 -16036 23999 -16008
rect 23305 -16064 23378 -16036
rect 23412 -16064 23478 -16036
rect 23512 -16064 23578 -16036
rect 23612 -16064 23678 -16036
rect 23305 -16098 23366 -16064
rect 23412 -16070 23456 -16064
rect 23512 -16070 23546 -16064
rect 23612 -16070 23636 -16064
rect 23400 -16098 23456 -16070
rect 23490 -16098 23546 -16070
rect 23580 -16098 23636 -16070
rect 23670 -16070 23678 -16064
rect 23712 -16064 23778 -16036
rect 23712 -16070 23726 -16064
rect 23670 -16098 23726 -16070
rect 23760 -16070 23778 -16064
rect 23812 -16064 23878 -16036
rect 23912 -16064 23999 -16036
rect 23812 -16070 23816 -16064
rect 23760 -16098 23816 -16070
rect 23850 -16070 23878 -16064
rect 23850 -16098 23906 -16070
rect 23940 -16098 23999 -16064
rect 23305 -16157 23999 -16098
rect 24061 -15494 24080 -15460
rect 24114 -15494 24133 -15460
rect 24061 -15550 24133 -15494
rect 24061 -15584 24080 -15550
rect 24114 -15584 24133 -15550
rect 24061 -15640 24133 -15584
rect 24061 -15674 24080 -15640
rect 24114 -15674 24133 -15640
rect 24061 -15730 24133 -15674
rect 24061 -15764 24080 -15730
rect 24114 -15764 24133 -15730
rect 24061 -15820 24133 -15764
rect 24061 -15854 24080 -15820
rect 24114 -15854 24133 -15820
rect 24061 -15910 24133 -15854
rect 24061 -15944 24080 -15910
rect 24114 -15944 24133 -15910
rect 24061 -16000 24133 -15944
rect 24061 -16034 24080 -16000
rect 24114 -16034 24133 -16000
rect 24061 -16090 24133 -16034
rect 24061 -16124 24080 -16090
rect 24114 -16124 24133 -16090
rect 23171 -16202 23243 -16180
rect 24061 -16180 24133 -16124
rect 24061 -16202 24080 -16180
rect 23074 -16214 24080 -16202
rect 24114 -16202 24133 -16180
rect 24197 -15420 24227 -15402
rect 24261 -15420 24328 -15386
rect 24362 -15402 25515 -15386
rect 24362 -15420 24395 -15402
rect 24197 -15476 24395 -15420
rect 24197 -15510 24227 -15476
rect 24261 -15510 24328 -15476
rect 24362 -15510 24395 -15476
rect 24197 -15566 24395 -15510
rect 24197 -15600 24227 -15566
rect 24261 -15600 24328 -15566
rect 24362 -15600 24395 -15566
rect 24197 -15656 24395 -15600
rect 24197 -15690 24227 -15656
rect 24261 -15690 24328 -15656
rect 24362 -15690 24395 -15656
rect 24197 -15746 24395 -15690
rect 24197 -15780 24227 -15746
rect 24261 -15780 24328 -15746
rect 24362 -15780 24395 -15746
rect 24197 -15836 24395 -15780
rect 24197 -15870 24227 -15836
rect 24261 -15870 24328 -15836
rect 24362 -15870 24395 -15836
rect 24197 -15926 24395 -15870
rect 24197 -15960 24227 -15926
rect 24261 -15960 24328 -15926
rect 24362 -15960 24395 -15926
rect 24197 -16016 24395 -15960
rect 24197 -16050 24227 -16016
rect 24261 -16050 24328 -16016
rect 24362 -16050 24395 -16016
rect 24197 -16106 24395 -16050
rect 24197 -16140 24227 -16106
rect 24261 -16140 24328 -16106
rect 24362 -16140 24395 -16106
rect 24197 -16196 24395 -16140
rect 24197 -16202 24227 -16196
rect 24114 -16214 24227 -16202
rect 23074 -16230 24227 -16214
rect 24261 -16230 24328 -16196
rect 24362 -16202 24395 -16196
rect 24459 -15426 24531 -15402
rect 24459 -15460 24478 -15426
rect 24512 -15460 24531 -15426
rect 24459 -15516 24531 -15460
rect 25349 -15460 25421 -15402
rect 24459 -15550 24478 -15516
rect 24512 -15550 24531 -15516
rect 24459 -15606 24531 -15550
rect 24459 -15640 24478 -15606
rect 24512 -15640 24531 -15606
rect 24459 -15696 24531 -15640
rect 24459 -15730 24478 -15696
rect 24512 -15730 24531 -15696
rect 24459 -15786 24531 -15730
rect 24459 -15820 24478 -15786
rect 24512 -15820 24531 -15786
rect 24459 -15876 24531 -15820
rect 24459 -15910 24478 -15876
rect 24512 -15910 24531 -15876
rect 24459 -15966 24531 -15910
rect 24459 -16000 24478 -15966
rect 24512 -16000 24531 -15966
rect 24459 -16056 24531 -16000
rect 24459 -16090 24478 -16056
rect 24512 -16090 24531 -16056
rect 24459 -16146 24531 -16090
rect 24459 -16180 24478 -16146
rect 24512 -16180 24531 -16146
rect 24593 -15524 25287 -15463
rect 24593 -15558 24654 -15524
rect 24688 -15536 24744 -15524
rect 24778 -15536 24834 -15524
rect 24868 -15536 24924 -15524
rect 24700 -15558 24744 -15536
rect 24800 -15558 24834 -15536
rect 24900 -15558 24924 -15536
rect 24958 -15536 25014 -15524
rect 24958 -15558 24966 -15536
rect 24593 -15570 24666 -15558
rect 24700 -15570 24766 -15558
rect 24800 -15570 24866 -15558
rect 24900 -15570 24966 -15558
rect 25000 -15558 25014 -15536
rect 25048 -15536 25104 -15524
rect 25048 -15558 25066 -15536
rect 25000 -15570 25066 -15558
rect 25100 -15558 25104 -15536
rect 25138 -15536 25194 -15524
rect 25138 -15558 25166 -15536
rect 25228 -15558 25287 -15524
rect 25100 -15570 25166 -15558
rect 25200 -15570 25287 -15558
rect 24593 -15614 25287 -15570
rect 24593 -15648 24654 -15614
rect 24688 -15636 24744 -15614
rect 24778 -15636 24834 -15614
rect 24868 -15636 24924 -15614
rect 24700 -15648 24744 -15636
rect 24800 -15648 24834 -15636
rect 24900 -15648 24924 -15636
rect 24958 -15636 25014 -15614
rect 24958 -15648 24966 -15636
rect 24593 -15670 24666 -15648
rect 24700 -15670 24766 -15648
rect 24800 -15670 24866 -15648
rect 24900 -15670 24966 -15648
rect 25000 -15648 25014 -15636
rect 25048 -15636 25104 -15614
rect 25048 -15648 25066 -15636
rect 25000 -15670 25066 -15648
rect 25100 -15648 25104 -15636
rect 25138 -15636 25194 -15614
rect 25138 -15648 25166 -15636
rect 25228 -15648 25287 -15614
rect 25100 -15670 25166 -15648
rect 25200 -15670 25287 -15648
rect 24593 -15704 25287 -15670
rect 24593 -15738 24654 -15704
rect 24688 -15736 24744 -15704
rect 24778 -15736 24834 -15704
rect 24868 -15736 24924 -15704
rect 24700 -15738 24744 -15736
rect 24800 -15738 24834 -15736
rect 24900 -15738 24924 -15736
rect 24958 -15736 25014 -15704
rect 24958 -15738 24966 -15736
rect 24593 -15770 24666 -15738
rect 24700 -15770 24766 -15738
rect 24800 -15770 24866 -15738
rect 24900 -15770 24966 -15738
rect 25000 -15738 25014 -15736
rect 25048 -15736 25104 -15704
rect 25048 -15738 25066 -15736
rect 25000 -15770 25066 -15738
rect 25100 -15738 25104 -15736
rect 25138 -15736 25194 -15704
rect 25138 -15738 25166 -15736
rect 25228 -15738 25287 -15704
rect 25100 -15770 25166 -15738
rect 25200 -15770 25287 -15738
rect 24593 -15794 25287 -15770
rect 24593 -15828 24654 -15794
rect 24688 -15828 24744 -15794
rect 24778 -15828 24834 -15794
rect 24868 -15828 24924 -15794
rect 24958 -15828 25014 -15794
rect 25048 -15828 25104 -15794
rect 25138 -15828 25194 -15794
rect 25228 -15828 25287 -15794
rect 24593 -15836 25287 -15828
rect 24593 -15870 24666 -15836
rect 24700 -15870 24766 -15836
rect 24800 -15870 24866 -15836
rect 24900 -15870 24966 -15836
rect 25000 -15870 25066 -15836
rect 25100 -15870 25166 -15836
rect 25200 -15870 25287 -15836
rect 24593 -15884 25287 -15870
rect 24593 -15918 24654 -15884
rect 24688 -15918 24744 -15884
rect 24778 -15918 24834 -15884
rect 24868 -15918 24924 -15884
rect 24958 -15918 25014 -15884
rect 25048 -15918 25104 -15884
rect 25138 -15918 25194 -15884
rect 25228 -15918 25287 -15884
rect 24593 -15936 25287 -15918
rect 24593 -15970 24666 -15936
rect 24700 -15970 24766 -15936
rect 24800 -15970 24866 -15936
rect 24900 -15970 24966 -15936
rect 25000 -15970 25066 -15936
rect 25100 -15970 25166 -15936
rect 25200 -15970 25287 -15936
rect 24593 -15974 25287 -15970
rect 24593 -16008 24654 -15974
rect 24688 -16008 24744 -15974
rect 24778 -16008 24834 -15974
rect 24868 -16008 24924 -15974
rect 24958 -16008 25014 -15974
rect 25048 -16008 25104 -15974
rect 25138 -16008 25194 -15974
rect 25228 -16008 25287 -15974
rect 24593 -16036 25287 -16008
rect 24593 -16064 24666 -16036
rect 24700 -16064 24766 -16036
rect 24800 -16064 24866 -16036
rect 24900 -16064 24966 -16036
rect 24593 -16098 24654 -16064
rect 24700 -16070 24744 -16064
rect 24800 -16070 24834 -16064
rect 24900 -16070 24924 -16064
rect 24688 -16098 24744 -16070
rect 24778 -16098 24834 -16070
rect 24868 -16098 24924 -16070
rect 24958 -16070 24966 -16064
rect 25000 -16064 25066 -16036
rect 25000 -16070 25014 -16064
rect 24958 -16098 25014 -16070
rect 25048 -16070 25066 -16064
rect 25100 -16064 25166 -16036
rect 25200 -16064 25287 -16036
rect 25100 -16070 25104 -16064
rect 25048 -16098 25104 -16070
rect 25138 -16070 25166 -16064
rect 25138 -16098 25194 -16070
rect 25228 -16098 25287 -16064
rect 24593 -16157 25287 -16098
rect 25349 -15494 25368 -15460
rect 25402 -15494 25421 -15460
rect 25349 -15550 25421 -15494
rect 25349 -15584 25368 -15550
rect 25402 -15584 25421 -15550
rect 25349 -15640 25421 -15584
rect 25349 -15674 25368 -15640
rect 25402 -15674 25421 -15640
rect 25349 -15730 25421 -15674
rect 25349 -15764 25368 -15730
rect 25402 -15764 25421 -15730
rect 25349 -15820 25421 -15764
rect 25349 -15854 25368 -15820
rect 25402 -15854 25421 -15820
rect 25349 -15910 25421 -15854
rect 25349 -15944 25368 -15910
rect 25402 -15944 25421 -15910
rect 25349 -16000 25421 -15944
rect 25349 -16034 25368 -16000
rect 25402 -16034 25421 -16000
rect 25349 -16090 25421 -16034
rect 25349 -16124 25368 -16090
rect 25402 -16124 25421 -16090
rect 24459 -16202 24531 -16180
rect 25349 -16180 25421 -16124
rect 25349 -16202 25368 -16180
rect 24362 -16214 25368 -16202
rect 25402 -16202 25421 -16180
rect 25485 -15420 25515 -15402
rect 25549 -15420 25616 -15386
rect 25650 -15402 26803 -15386
rect 25650 -15420 25683 -15402
rect 25485 -15476 25683 -15420
rect 25485 -15510 25515 -15476
rect 25549 -15510 25616 -15476
rect 25650 -15510 25683 -15476
rect 25485 -15566 25683 -15510
rect 25485 -15600 25515 -15566
rect 25549 -15600 25616 -15566
rect 25650 -15600 25683 -15566
rect 25485 -15656 25683 -15600
rect 25485 -15690 25515 -15656
rect 25549 -15690 25616 -15656
rect 25650 -15690 25683 -15656
rect 25485 -15746 25683 -15690
rect 25485 -15780 25515 -15746
rect 25549 -15780 25616 -15746
rect 25650 -15780 25683 -15746
rect 25485 -15836 25683 -15780
rect 25485 -15870 25515 -15836
rect 25549 -15870 25616 -15836
rect 25650 -15870 25683 -15836
rect 25485 -15926 25683 -15870
rect 25485 -15960 25515 -15926
rect 25549 -15960 25616 -15926
rect 25650 -15960 25683 -15926
rect 25485 -16016 25683 -15960
rect 25485 -16050 25515 -16016
rect 25549 -16050 25616 -16016
rect 25650 -16050 25683 -16016
rect 25485 -16106 25683 -16050
rect 25485 -16140 25515 -16106
rect 25549 -16140 25616 -16106
rect 25650 -16140 25683 -16106
rect 25485 -16196 25683 -16140
rect 25485 -16202 25515 -16196
rect 25402 -16214 25515 -16202
rect 24362 -16230 25515 -16214
rect 25549 -16230 25616 -16196
rect 25650 -16202 25683 -16196
rect 25747 -15426 25819 -15402
rect 25747 -15460 25766 -15426
rect 25800 -15460 25819 -15426
rect 25747 -15516 25819 -15460
rect 26637 -15460 26709 -15402
rect 25747 -15550 25766 -15516
rect 25800 -15550 25819 -15516
rect 25747 -15606 25819 -15550
rect 25747 -15640 25766 -15606
rect 25800 -15640 25819 -15606
rect 25747 -15696 25819 -15640
rect 25747 -15730 25766 -15696
rect 25800 -15730 25819 -15696
rect 25747 -15786 25819 -15730
rect 25747 -15820 25766 -15786
rect 25800 -15820 25819 -15786
rect 25747 -15876 25819 -15820
rect 25747 -15910 25766 -15876
rect 25800 -15910 25819 -15876
rect 25747 -15966 25819 -15910
rect 25747 -16000 25766 -15966
rect 25800 -16000 25819 -15966
rect 25747 -16056 25819 -16000
rect 25747 -16090 25766 -16056
rect 25800 -16090 25819 -16056
rect 25747 -16146 25819 -16090
rect 25747 -16180 25766 -16146
rect 25800 -16180 25819 -16146
rect 25881 -15524 26575 -15463
rect 25881 -15558 25942 -15524
rect 25976 -15536 26032 -15524
rect 26066 -15536 26122 -15524
rect 26156 -15536 26212 -15524
rect 25988 -15558 26032 -15536
rect 26088 -15558 26122 -15536
rect 26188 -15558 26212 -15536
rect 26246 -15536 26302 -15524
rect 26246 -15558 26254 -15536
rect 25881 -15570 25954 -15558
rect 25988 -15570 26054 -15558
rect 26088 -15570 26154 -15558
rect 26188 -15570 26254 -15558
rect 26288 -15558 26302 -15536
rect 26336 -15536 26392 -15524
rect 26336 -15558 26354 -15536
rect 26288 -15570 26354 -15558
rect 26388 -15558 26392 -15536
rect 26426 -15536 26482 -15524
rect 26426 -15558 26454 -15536
rect 26516 -15558 26575 -15524
rect 26388 -15570 26454 -15558
rect 26488 -15570 26575 -15558
rect 25881 -15614 26575 -15570
rect 25881 -15648 25942 -15614
rect 25976 -15636 26032 -15614
rect 26066 -15636 26122 -15614
rect 26156 -15636 26212 -15614
rect 25988 -15648 26032 -15636
rect 26088 -15648 26122 -15636
rect 26188 -15648 26212 -15636
rect 26246 -15636 26302 -15614
rect 26246 -15648 26254 -15636
rect 25881 -15670 25954 -15648
rect 25988 -15670 26054 -15648
rect 26088 -15670 26154 -15648
rect 26188 -15670 26254 -15648
rect 26288 -15648 26302 -15636
rect 26336 -15636 26392 -15614
rect 26336 -15648 26354 -15636
rect 26288 -15670 26354 -15648
rect 26388 -15648 26392 -15636
rect 26426 -15636 26482 -15614
rect 26426 -15648 26454 -15636
rect 26516 -15648 26575 -15614
rect 26388 -15670 26454 -15648
rect 26488 -15670 26575 -15648
rect 25881 -15704 26575 -15670
rect 25881 -15738 25942 -15704
rect 25976 -15736 26032 -15704
rect 26066 -15736 26122 -15704
rect 26156 -15736 26212 -15704
rect 25988 -15738 26032 -15736
rect 26088 -15738 26122 -15736
rect 26188 -15738 26212 -15736
rect 26246 -15736 26302 -15704
rect 26246 -15738 26254 -15736
rect 25881 -15770 25954 -15738
rect 25988 -15770 26054 -15738
rect 26088 -15770 26154 -15738
rect 26188 -15770 26254 -15738
rect 26288 -15738 26302 -15736
rect 26336 -15736 26392 -15704
rect 26336 -15738 26354 -15736
rect 26288 -15770 26354 -15738
rect 26388 -15738 26392 -15736
rect 26426 -15736 26482 -15704
rect 26426 -15738 26454 -15736
rect 26516 -15738 26575 -15704
rect 26388 -15770 26454 -15738
rect 26488 -15770 26575 -15738
rect 25881 -15794 26575 -15770
rect 25881 -15828 25942 -15794
rect 25976 -15828 26032 -15794
rect 26066 -15828 26122 -15794
rect 26156 -15828 26212 -15794
rect 26246 -15828 26302 -15794
rect 26336 -15828 26392 -15794
rect 26426 -15828 26482 -15794
rect 26516 -15828 26575 -15794
rect 25881 -15836 26575 -15828
rect 25881 -15870 25954 -15836
rect 25988 -15870 26054 -15836
rect 26088 -15870 26154 -15836
rect 26188 -15870 26254 -15836
rect 26288 -15870 26354 -15836
rect 26388 -15870 26454 -15836
rect 26488 -15870 26575 -15836
rect 25881 -15884 26575 -15870
rect 25881 -15918 25942 -15884
rect 25976 -15918 26032 -15884
rect 26066 -15918 26122 -15884
rect 26156 -15918 26212 -15884
rect 26246 -15918 26302 -15884
rect 26336 -15918 26392 -15884
rect 26426 -15918 26482 -15884
rect 26516 -15918 26575 -15884
rect 25881 -15936 26575 -15918
rect 25881 -15970 25954 -15936
rect 25988 -15970 26054 -15936
rect 26088 -15970 26154 -15936
rect 26188 -15970 26254 -15936
rect 26288 -15970 26354 -15936
rect 26388 -15970 26454 -15936
rect 26488 -15970 26575 -15936
rect 25881 -15974 26575 -15970
rect 25881 -16008 25942 -15974
rect 25976 -16008 26032 -15974
rect 26066 -16008 26122 -15974
rect 26156 -16008 26212 -15974
rect 26246 -16008 26302 -15974
rect 26336 -16008 26392 -15974
rect 26426 -16008 26482 -15974
rect 26516 -16008 26575 -15974
rect 25881 -16036 26575 -16008
rect 25881 -16064 25954 -16036
rect 25988 -16064 26054 -16036
rect 26088 -16064 26154 -16036
rect 26188 -16064 26254 -16036
rect 25881 -16098 25942 -16064
rect 25988 -16070 26032 -16064
rect 26088 -16070 26122 -16064
rect 26188 -16070 26212 -16064
rect 25976 -16098 26032 -16070
rect 26066 -16098 26122 -16070
rect 26156 -16098 26212 -16070
rect 26246 -16070 26254 -16064
rect 26288 -16064 26354 -16036
rect 26288 -16070 26302 -16064
rect 26246 -16098 26302 -16070
rect 26336 -16070 26354 -16064
rect 26388 -16064 26454 -16036
rect 26488 -16064 26575 -16036
rect 26388 -16070 26392 -16064
rect 26336 -16098 26392 -16070
rect 26426 -16070 26454 -16064
rect 26426 -16098 26482 -16070
rect 26516 -16098 26575 -16064
rect 25881 -16157 26575 -16098
rect 26637 -15494 26656 -15460
rect 26690 -15494 26709 -15460
rect 26637 -15550 26709 -15494
rect 26637 -15584 26656 -15550
rect 26690 -15584 26709 -15550
rect 26637 -15640 26709 -15584
rect 26637 -15674 26656 -15640
rect 26690 -15674 26709 -15640
rect 26637 -15730 26709 -15674
rect 26637 -15764 26656 -15730
rect 26690 -15764 26709 -15730
rect 26637 -15820 26709 -15764
rect 26637 -15854 26656 -15820
rect 26690 -15854 26709 -15820
rect 26637 -15910 26709 -15854
rect 26637 -15944 26656 -15910
rect 26690 -15944 26709 -15910
rect 26637 -16000 26709 -15944
rect 26637 -16034 26656 -16000
rect 26690 -16034 26709 -16000
rect 26637 -16090 26709 -16034
rect 26637 -16124 26656 -16090
rect 26690 -16124 26709 -16090
rect 25747 -16202 25819 -16180
rect 26637 -16180 26709 -16124
rect 26637 -16202 26656 -16180
rect 25650 -16214 26656 -16202
rect 26690 -16202 26709 -16180
rect 26773 -15420 26803 -15402
rect 26837 -15420 26872 -15386
rect 26773 -15476 26872 -15420
rect 26773 -15510 26803 -15476
rect 26837 -15510 26872 -15476
rect 26773 -15566 26872 -15510
rect 26773 -15600 26803 -15566
rect 26837 -15600 26872 -15566
rect 26773 -15656 26872 -15600
rect 26773 -15690 26803 -15656
rect 26837 -15690 26872 -15656
rect 26773 -15746 26872 -15690
rect 26773 -15780 26803 -15746
rect 26837 -15780 26872 -15746
rect 26773 -15836 26872 -15780
rect 26773 -15870 26803 -15836
rect 26837 -15870 26872 -15836
rect 26773 -15926 26872 -15870
rect 26773 -15960 26803 -15926
rect 26837 -15960 26872 -15926
rect 26773 -16016 26872 -15960
rect 26773 -16050 26803 -16016
rect 26837 -16050 26872 -16016
rect 26773 -16106 26872 -16050
rect 26773 -16140 26803 -16106
rect 26837 -16140 26872 -16106
rect 26773 -16196 26872 -16140
rect 26773 -16202 26803 -16196
rect 26690 -16214 26803 -16202
rect 25650 -16230 26803 -16214
rect 26837 -16202 26872 -16196
rect 26837 -16230 26884 -16202
rect 16568 -16238 26884 -16230
rect 16568 -16272 16844 -16238
rect 16878 -16272 16934 -16238
rect 16968 -16272 17024 -16238
rect 17058 -16272 17114 -16238
rect 17148 -16272 17204 -16238
rect 17238 -16272 17294 -16238
rect 17328 -16272 17384 -16238
rect 17418 -16272 17474 -16238
rect 17508 -16272 17564 -16238
rect 17598 -16272 18132 -16238
rect 18166 -16272 18222 -16238
rect 18256 -16272 18312 -16238
rect 18346 -16272 18402 -16238
rect 18436 -16272 18492 -16238
rect 18526 -16272 18582 -16238
rect 18616 -16272 18672 -16238
rect 18706 -16272 18762 -16238
rect 18796 -16272 18852 -16238
rect 18886 -16272 19420 -16238
rect 19454 -16272 19510 -16238
rect 19544 -16272 19600 -16238
rect 19634 -16272 19690 -16238
rect 19724 -16272 19780 -16238
rect 19814 -16272 19870 -16238
rect 19904 -16272 19960 -16238
rect 19994 -16272 20050 -16238
rect 20084 -16272 20140 -16238
rect 20174 -16272 20708 -16238
rect 20742 -16272 20798 -16238
rect 20832 -16272 20888 -16238
rect 20922 -16272 20978 -16238
rect 21012 -16272 21068 -16238
rect 21102 -16272 21158 -16238
rect 21192 -16272 21248 -16238
rect 21282 -16272 21338 -16238
rect 21372 -16272 21428 -16238
rect 21462 -16272 21996 -16238
rect 22030 -16272 22086 -16238
rect 22120 -16272 22176 -16238
rect 22210 -16272 22266 -16238
rect 22300 -16272 22356 -16238
rect 22390 -16272 22446 -16238
rect 22480 -16272 22536 -16238
rect 22570 -16272 22626 -16238
rect 22660 -16272 22716 -16238
rect 22750 -16272 23284 -16238
rect 23318 -16272 23374 -16238
rect 23408 -16272 23464 -16238
rect 23498 -16272 23554 -16238
rect 23588 -16272 23644 -16238
rect 23678 -16272 23734 -16238
rect 23768 -16272 23824 -16238
rect 23858 -16272 23914 -16238
rect 23948 -16272 24004 -16238
rect 24038 -16272 24572 -16238
rect 24606 -16272 24662 -16238
rect 24696 -16272 24752 -16238
rect 24786 -16272 24842 -16238
rect 24876 -16272 24932 -16238
rect 24966 -16272 25022 -16238
rect 25056 -16272 25112 -16238
rect 25146 -16272 25202 -16238
rect 25236 -16272 25292 -16238
rect 25326 -16272 25860 -16238
rect 25894 -16272 25950 -16238
rect 25984 -16272 26040 -16238
rect 26074 -16272 26130 -16238
rect 26164 -16272 26220 -16238
rect 26254 -16272 26310 -16238
rect 26344 -16272 26400 -16238
rect 26434 -16272 26490 -16238
rect 26524 -16272 26580 -16238
rect 26614 -16272 26884 -16238
rect 16568 -16286 26884 -16272
rect 16568 -16320 16600 -16286
rect 16634 -16320 17787 -16286
rect 17821 -16320 17888 -16286
rect 17922 -16320 19075 -16286
rect 19109 -16320 19176 -16286
rect 19210 -16320 20363 -16286
rect 20397 -16320 20464 -16286
rect 20498 -16320 21651 -16286
rect 21685 -16320 21752 -16286
rect 21786 -16320 22939 -16286
rect 22973 -16320 23040 -16286
rect 23074 -16320 24227 -16286
rect 24261 -16320 24328 -16286
rect 24362 -16320 25515 -16286
rect 25549 -16320 25616 -16286
rect 25650 -16320 26803 -16286
rect 26837 -16320 26884 -16286
rect 16568 -16387 26884 -16320
rect 16568 -16421 16684 -16387
rect 16718 -16421 16774 -16387
rect 16808 -16421 16864 -16387
rect 16898 -16421 16954 -16387
rect 16988 -16421 17044 -16387
rect 17078 -16421 17134 -16387
rect 17168 -16421 17224 -16387
rect 17258 -16421 17314 -16387
rect 17348 -16421 17404 -16387
rect 17438 -16421 17494 -16387
rect 17528 -16421 17584 -16387
rect 17618 -16421 17674 -16387
rect 17708 -16421 17764 -16387
rect 17798 -16421 17972 -16387
rect 18006 -16421 18062 -16387
rect 18096 -16421 18152 -16387
rect 18186 -16421 18242 -16387
rect 18276 -16421 18332 -16387
rect 18366 -16421 18422 -16387
rect 18456 -16421 18512 -16387
rect 18546 -16421 18602 -16387
rect 18636 -16421 18692 -16387
rect 18726 -16421 18782 -16387
rect 18816 -16421 18872 -16387
rect 18906 -16421 18962 -16387
rect 18996 -16421 19052 -16387
rect 19086 -16421 19260 -16387
rect 19294 -16421 19350 -16387
rect 19384 -16421 19440 -16387
rect 19474 -16421 19530 -16387
rect 19564 -16421 19620 -16387
rect 19654 -16421 19710 -16387
rect 19744 -16421 19800 -16387
rect 19834 -16421 19890 -16387
rect 19924 -16421 19980 -16387
rect 20014 -16421 20070 -16387
rect 20104 -16421 20160 -16387
rect 20194 -16421 20250 -16387
rect 20284 -16421 20340 -16387
rect 20374 -16421 20548 -16387
rect 20582 -16421 20638 -16387
rect 20672 -16421 20728 -16387
rect 20762 -16421 20818 -16387
rect 20852 -16421 20908 -16387
rect 20942 -16421 20998 -16387
rect 21032 -16421 21088 -16387
rect 21122 -16421 21178 -16387
rect 21212 -16421 21268 -16387
rect 21302 -16421 21358 -16387
rect 21392 -16421 21448 -16387
rect 21482 -16421 21538 -16387
rect 21572 -16421 21628 -16387
rect 21662 -16421 21836 -16387
rect 21870 -16421 21926 -16387
rect 21960 -16421 22016 -16387
rect 22050 -16421 22106 -16387
rect 22140 -16421 22196 -16387
rect 22230 -16421 22286 -16387
rect 22320 -16421 22376 -16387
rect 22410 -16421 22466 -16387
rect 22500 -16421 22556 -16387
rect 22590 -16421 22646 -16387
rect 22680 -16421 22736 -16387
rect 22770 -16421 22826 -16387
rect 22860 -16421 22916 -16387
rect 22950 -16421 23124 -16387
rect 23158 -16421 23214 -16387
rect 23248 -16421 23304 -16387
rect 23338 -16421 23394 -16387
rect 23428 -16421 23484 -16387
rect 23518 -16421 23574 -16387
rect 23608 -16421 23664 -16387
rect 23698 -16421 23754 -16387
rect 23788 -16421 23844 -16387
rect 23878 -16421 23934 -16387
rect 23968 -16421 24024 -16387
rect 24058 -16421 24114 -16387
rect 24148 -16421 24204 -16387
rect 24238 -16421 24412 -16387
rect 24446 -16421 24502 -16387
rect 24536 -16421 24592 -16387
rect 24626 -16421 24682 -16387
rect 24716 -16421 24772 -16387
rect 24806 -16421 24862 -16387
rect 24896 -16421 24952 -16387
rect 24986 -16421 25042 -16387
rect 25076 -16421 25132 -16387
rect 25166 -16421 25222 -16387
rect 25256 -16421 25312 -16387
rect 25346 -16421 25402 -16387
rect 25436 -16421 25492 -16387
rect 25526 -16421 25700 -16387
rect 25734 -16421 25790 -16387
rect 25824 -16421 25880 -16387
rect 25914 -16421 25970 -16387
rect 26004 -16421 26060 -16387
rect 26094 -16421 26150 -16387
rect 26184 -16421 26240 -16387
rect 26274 -16421 26330 -16387
rect 26364 -16421 26420 -16387
rect 26454 -16421 26510 -16387
rect 26544 -16421 26600 -16387
rect 26634 -16421 26690 -16387
rect 26724 -16421 26780 -16387
rect 26814 -16421 26884 -16387
rect 6870 -16464 7302 -16456
rect 13606 -16464 14038 -16456
rect 6870 -16480 14038 -16464
rect 6870 -17050 7302 -16480
rect 13606 -17050 14038 -16480
rect 6870 -17066 14038 -17050
rect 6870 -17280 7302 -17066
rect 13606 -17280 14038 -17066
rect 16568 -16488 26884 -16421
rect 16568 -16522 16684 -16488
rect 16718 -16522 16774 -16488
rect 16808 -16522 16864 -16488
rect 16898 -16522 16954 -16488
rect 16988 -16522 17044 -16488
rect 17078 -16522 17134 -16488
rect 17168 -16522 17224 -16488
rect 17258 -16522 17314 -16488
rect 17348 -16522 17404 -16488
rect 17438 -16522 17494 -16488
rect 17528 -16522 17584 -16488
rect 17618 -16522 17674 -16488
rect 17708 -16522 17764 -16488
rect 17798 -16522 17972 -16488
rect 18006 -16522 18062 -16488
rect 18096 -16522 18152 -16488
rect 18186 -16522 18242 -16488
rect 18276 -16522 18332 -16488
rect 18366 -16522 18422 -16488
rect 18456 -16522 18512 -16488
rect 18546 -16522 18602 -16488
rect 18636 -16522 18692 -16488
rect 18726 -16522 18782 -16488
rect 18816 -16522 18872 -16488
rect 18906 -16522 18962 -16488
rect 18996 -16522 19052 -16488
rect 19086 -16522 19260 -16488
rect 19294 -16522 19350 -16488
rect 19384 -16522 19440 -16488
rect 19474 -16522 19530 -16488
rect 19564 -16522 19620 -16488
rect 19654 -16522 19710 -16488
rect 19744 -16522 19800 -16488
rect 19834 -16522 19890 -16488
rect 19924 -16522 19980 -16488
rect 20014 -16522 20070 -16488
rect 20104 -16522 20160 -16488
rect 20194 -16522 20250 -16488
rect 20284 -16522 20340 -16488
rect 20374 -16522 20548 -16488
rect 20582 -16522 20638 -16488
rect 20672 -16522 20728 -16488
rect 20762 -16522 20818 -16488
rect 20852 -16522 20908 -16488
rect 20942 -16522 20998 -16488
rect 21032 -16522 21088 -16488
rect 21122 -16522 21178 -16488
rect 21212 -16522 21268 -16488
rect 21302 -16522 21358 -16488
rect 21392 -16522 21448 -16488
rect 21482 -16522 21538 -16488
rect 21572 -16522 21628 -16488
rect 21662 -16522 21836 -16488
rect 21870 -16522 21926 -16488
rect 21960 -16522 22016 -16488
rect 22050 -16522 22106 -16488
rect 22140 -16522 22196 -16488
rect 22230 -16522 22286 -16488
rect 22320 -16522 22376 -16488
rect 22410 -16522 22466 -16488
rect 22500 -16522 22556 -16488
rect 22590 -16522 22646 -16488
rect 22680 -16522 22736 -16488
rect 22770 -16522 22826 -16488
rect 22860 -16522 22916 -16488
rect 22950 -16522 23124 -16488
rect 23158 -16522 23214 -16488
rect 23248 -16522 23304 -16488
rect 23338 -16522 23394 -16488
rect 23428 -16522 23484 -16488
rect 23518 -16522 23574 -16488
rect 23608 -16522 23664 -16488
rect 23698 -16522 23754 -16488
rect 23788 -16522 23844 -16488
rect 23878 -16522 23934 -16488
rect 23968 -16522 24024 -16488
rect 24058 -16522 24114 -16488
rect 24148 -16522 24204 -16488
rect 24238 -16522 24412 -16488
rect 24446 -16522 24502 -16488
rect 24536 -16522 24592 -16488
rect 24626 -16522 24682 -16488
rect 24716 -16522 24772 -16488
rect 24806 -16522 24862 -16488
rect 24896 -16522 24952 -16488
rect 24986 -16522 25042 -16488
rect 25076 -16522 25132 -16488
rect 25166 -16522 25222 -16488
rect 25256 -16522 25312 -16488
rect 25346 -16522 25402 -16488
rect 25436 -16522 25492 -16488
rect 25526 -16522 25700 -16488
rect 25734 -16522 25790 -16488
rect 25824 -16522 25880 -16488
rect 25914 -16522 25970 -16488
rect 26004 -16522 26060 -16488
rect 26094 -16522 26150 -16488
rect 26184 -16522 26240 -16488
rect 26274 -16522 26330 -16488
rect 26364 -16522 26420 -16488
rect 26454 -16522 26510 -16488
rect 26544 -16522 26600 -16488
rect 26634 -16522 26690 -16488
rect 26724 -16522 26780 -16488
rect 26814 -16522 26884 -16488
rect 16568 -16584 26884 -16522
rect 16568 -16618 16600 -16584
rect 16634 -16618 17787 -16584
rect 17821 -16618 17888 -16584
rect 17922 -16618 19075 -16584
rect 19109 -16618 19176 -16584
rect 19210 -16618 20363 -16584
rect 20397 -16618 20464 -16584
rect 20498 -16618 21651 -16584
rect 21685 -16618 21752 -16584
rect 21786 -16618 22939 -16584
rect 22973 -16618 23040 -16584
rect 23074 -16618 24227 -16584
rect 24261 -16618 24328 -16584
rect 24362 -16618 25515 -16584
rect 25549 -16618 25616 -16584
rect 25650 -16618 26803 -16584
rect 26837 -16618 26884 -16584
rect 16568 -16636 26884 -16618
rect 16568 -16670 16863 -16636
rect 16897 -16670 16953 -16636
rect 16987 -16670 17043 -16636
rect 17077 -16670 17133 -16636
rect 17167 -16670 17223 -16636
rect 17257 -16670 17313 -16636
rect 17347 -16670 17403 -16636
rect 17437 -16670 17493 -16636
rect 17527 -16670 17583 -16636
rect 17617 -16670 18151 -16636
rect 18185 -16670 18241 -16636
rect 18275 -16670 18331 -16636
rect 18365 -16670 18421 -16636
rect 18455 -16670 18511 -16636
rect 18545 -16670 18601 -16636
rect 18635 -16670 18691 -16636
rect 18725 -16670 18781 -16636
rect 18815 -16670 18871 -16636
rect 18905 -16670 19439 -16636
rect 19473 -16670 19529 -16636
rect 19563 -16670 19619 -16636
rect 19653 -16670 19709 -16636
rect 19743 -16670 19799 -16636
rect 19833 -16670 19889 -16636
rect 19923 -16670 19979 -16636
rect 20013 -16670 20069 -16636
rect 20103 -16670 20159 -16636
rect 20193 -16670 20727 -16636
rect 20761 -16670 20817 -16636
rect 20851 -16670 20907 -16636
rect 20941 -16670 20997 -16636
rect 21031 -16670 21087 -16636
rect 21121 -16670 21177 -16636
rect 21211 -16670 21267 -16636
rect 21301 -16670 21357 -16636
rect 21391 -16670 21447 -16636
rect 21481 -16670 22015 -16636
rect 22049 -16670 22105 -16636
rect 22139 -16670 22195 -16636
rect 22229 -16670 22285 -16636
rect 22319 -16670 22375 -16636
rect 22409 -16670 22465 -16636
rect 22499 -16670 22555 -16636
rect 22589 -16670 22645 -16636
rect 22679 -16670 22735 -16636
rect 22769 -16670 23303 -16636
rect 23337 -16670 23393 -16636
rect 23427 -16670 23483 -16636
rect 23517 -16670 23573 -16636
rect 23607 -16670 23663 -16636
rect 23697 -16670 23753 -16636
rect 23787 -16670 23843 -16636
rect 23877 -16670 23933 -16636
rect 23967 -16670 24023 -16636
rect 24057 -16670 24591 -16636
rect 24625 -16670 24681 -16636
rect 24715 -16670 24771 -16636
rect 24805 -16670 24861 -16636
rect 24895 -16670 24951 -16636
rect 24985 -16670 25041 -16636
rect 25075 -16670 25131 -16636
rect 25165 -16670 25221 -16636
rect 25255 -16670 25311 -16636
rect 25345 -16670 25879 -16636
rect 25913 -16670 25969 -16636
rect 26003 -16670 26059 -16636
rect 26093 -16670 26149 -16636
rect 26183 -16670 26239 -16636
rect 26273 -16670 26329 -16636
rect 26363 -16670 26419 -16636
rect 26453 -16670 26509 -16636
rect 26543 -16670 26599 -16636
rect 26633 -16670 26884 -16636
rect 16568 -16674 26884 -16670
rect 16568 -16708 16600 -16674
rect 16634 -16702 17787 -16674
rect 16634 -16708 16667 -16702
rect 16568 -16764 16667 -16708
rect 16568 -16798 16600 -16764
rect 16634 -16798 16667 -16764
rect 16568 -16854 16667 -16798
rect 16568 -16888 16600 -16854
rect 16634 -16888 16667 -16854
rect 16568 -16944 16667 -16888
rect 16568 -16978 16600 -16944
rect 16634 -16978 16667 -16944
rect 16568 -17034 16667 -16978
rect 16568 -17068 16600 -17034
rect 16634 -17068 16667 -17034
rect 16568 -17124 16667 -17068
rect 16568 -17158 16600 -17124
rect 16634 -17158 16667 -17124
rect 16568 -17214 16667 -17158
rect 16568 -17248 16600 -17214
rect 16634 -17248 16667 -17214
rect 16568 -17304 16667 -17248
rect 16568 -17338 16600 -17304
rect 16634 -17338 16667 -17304
rect 16568 -17394 16667 -17338
rect 16568 -17428 16600 -17394
rect 16634 -17428 16667 -17394
rect 16568 -17484 16667 -17428
rect 16568 -17518 16600 -17484
rect 16634 -17502 16667 -17484
rect 16731 -16714 16803 -16702
rect 16731 -16748 16750 -16714
rect 16784 -16748 16803 -16714
rect 16731 -16804 16803 -16748
rect 17621 -16748 17693 -16702
rect 16731 -16838 16750 -16804
rect 16784 -16838 16803 -16804
rect 16731 -16894 16803 -16838
rect 16731 -16928 16750 -16894
rect 16784 -16928 16803 -16894
rect 16731 -16984 16803 -16928
rect 16731 -17018 16750 -16984
rect 16784 -17018 16803 -16984
rect 16731 -17074 16803 -17018
rect 16731 -17108 16750 -17074
rect 16784 -17108 16803 -17074
rect 16731 -17164 16803 -17108
rect 16731 -17198 16750 -17164
rect 16784 -17198 16803 -17164
rect 16731 -17254 16803 -17198
rect 16731 -17288 16750 -17254
rect 16784 -17288 16803 -17254
rect 16731 -17344 16803 -17288
rect 16731 -17378 16750 -17344
rect 16784 -17378 16803 -17344
rect 16731 -17434 16803 -17378
rect 16731 -17468 16750 -17434
rect 16784 -17468 16803 -17434
rect 16865 -16812 17559 -16751
rect 16865 -16846 16926 -16812
rect 16960 -16824 17016 -16812
rect 17050 -16824 17106 -16812
rect 17140 -16824 17196 -16812
rect 16972 -16846 17016 -16824
rect 17072 -16846 17106 -16824
rect 17172 -16846 17196 -16824
rect 17230 -16824 17286 -16812
rect 17230 -16846 17238 -16824
rect 16865 -16858 16938 -16846
rect 16972 -16858 17038 -16846
rect 17072 -16858 17138 -16846
rect 17172 -16858 17238 -16846
rect 17272 -16846 17286 -16824
rect 17320 -16824 17376 -16812
rect 17320 -16846 17338 -16824
rect 17272 -16858 17338 -16846
rect 17372 -16846 17376 -16824
rect 17410 -16824 17466 -16812
rect 17410 -16846 17438 -16824
rect 17500 -16846 17559 -16812
rect 17372 -16858 17438 -16846
rect 17472 -16858 17559 -16846
rect 16865 -16902 17559 -16858
rect 16865 -16936 16926 -16902
rect 16960 -16924 17016 -16902
rect 17050 -16924 17106 -16902
rect 17140 -16924 17196 -16902
rect 16972 -16936 17016 -16924
rect 17072 -16936 17106 -16924
rect 17172 -16936 17196 -16924
rect 17230 -16924 17286 -16902
rect 17230 -16936 17238 -16924
rect 16865 -16958 16938 -16936
rect 16972 -16958 17038 -16936
rect 17072 -16958 17138 -16936
rect 17172 -16958 17238 -16936
rect 17272 -16936 17286 -16924
rect 17320 -16924 17376 -16902
rect 17320 -16936 17338 -16924
rect 17272 -16958 17338 -16936
rect 17372 -16936 17376 -16924
rect 17410 -16924 17466 -16902
rect 17410 -16936 17438 -16924
rect 17500 -16936 17559 -16902
rect 17372 -16958 17438 -16936
rect 17472 -16958 17559 -16936
rect 16865 -16992 17559 -16958
rect 16865 -17026 16926 -16992
rect 16960 -17024 17016 -16992
rect 17050 -17024 17106 -16992
rect 17140 -17024 17196 -16992
rect 16972 -17026 17016 -17024
rect 17072 -17026 17106 -17024
rect 17172 -17026 17196 -17024
rect 17230 -17024 17286 -16992
rect 17230 -17026 17238 -17024
rect 16865 -17058 16938 -17026
rect 16972 -17058 17038 -17026
rect 17072 -17058 17138 -17026
rect 17172 -17058 17238 -17026
rect 17272 -17026 17286 -17024
rect 17320 -17024 17376 -16992
rect 17320 -17026 17338 -17024
rect 17272 -17058 17338 -17026
rect 17372 -17026 17376 -17024
rect 17410 -17024 17466 -16992
rect 17410 -17026 17438 -17024
rect 17500 -17026 17559 -16992
rect 17372 -17058 17438 -17026
rect 17472 -17058 17559 -17026
rect 16865 -17082 17559 -17058
rect 16865 -17116 16926 -17082
rect 16960 -17116 17016 -17082
rect 17050 -17116 17106 -17082
rect 17140 -17116 17196 -17082
rect 17230 -17116 17286 -17082
rect 17320 -17116 17376 -17082
rect 17410 -17116 17466 -17082
rect 17500 -17116 17559 -17082
rect 16865 -17124 17559 -17116
rect 16865 -17158 16938 -17124
rect 16972 -17158 17038 -17124
rect 17072 -17158 17138 -17124
rect 17172 -17158 17238 -17124
rect 17272 -17158 17338 -17124
rect 17372 -17158 17438 -17124
rect 17472 -17158 17559 -17124
rect 16865 -17172 17559 -17158
rect 16865 -17206 16926 -17172
rect 16960 -17206 17016 -17172
rect 17050 -17206 17106 -17172
rect 17140 -17206 17196 -17172
rect 17230 -17206 17286 -17172
rect 17320 -17206 17376 -17172
rect 17410 -17206 17466 -17172
rect 17500 -17206 17559 -17172
rect 16865 -17224 17559 -17206
rect 16865 -17258 16938 -17224
rect 16972 -17258 17038 -17224
rect 17072 -17258 17138 -17224
rect 17172 -17258 17238 -17224
rect 17272 -17258 17338 -17224
rect 17372 -17258 17438 -17224
rect 17472 -17258 17559 -17224
rect 16865 -17262 17559 -17258
rect 16865 -17296 16926 -17262
rect 16960 -17296 17016 -17262
rect 17050 -17296 17106 -17262
rect 17140 -17296 17196 -17262
rect 17230 -17296 17286 -17262
rect 17320 -17296 17376 -17262
rect 17410 -17296 17466 -17262
rect 17500 -17296 17559 -17262
rect 16865 -17324 17559 -17296
rect 16865 -17352 16938 -17324
rect 16972 -17352 17038 -17324
rect 17072 -17352 17138 -17324
rect 17172 -17352 17238 -17324
rect 16865 -17386 16926 -17352
rect 16972 -17358 17016 -17352
rect 17072 -17358 17106 -17352
rect 17172 -17358 17196 -17352
rect 16960 -17386 17016 -17358
rect 17050 -17386 17106 -17358
rect 17140 -17386 17196 -17358
rect 17230 -17358 17238 -17352
rect 17272 -17352 17338 -17324
rect 17272 -17358 17286 -17352
rect 17230 -17386 17286 -17358
rect 17320 -17358 17338 -17352
rect 17372 -17352 17438 -17324
rect 17472 -17352 17559 -17324
rect 17372 -17358 17376 -17352
rect 17320 -17386 17376 -17358
rect 17410 -17358 17438 -17352
rect 17410 -17386 17466 -17358
rect 17500 -17386 17559 -17352
rect 16865 -17445 17559 -17386
rect 17621 -16782 17640 -16748
rect 17674 -16782 17693 -16748
rect 17621 -16838 17693 -16782
rect 17621 -16872 17640 -16838
rect 17674 -16872 17693 -16838
rect 17621 -16928 17693 -16872
rect 17621 -16962 17640 -16928
rect 17674 -16962 17693 -16928
rect 17621 -17018 17693 -16962
rect 17621 -17052 17640 -17018
rect 17674 -17052 17693 -17018
rect 17621 -17108 17693 -17052
rect 17621 -17142 17640 -17108
rect 17674 -17142 17693 -17108
rect 17621 -17198 17693 -17142
rect 17621 -17232 17640 -17198
rect 17674 -17232 17693 -17198
rect 17621 -17288 17693 -17232
rect 17621 -17322 17640 -17288
rect 17674 -17322 17693 -17288
rect 17621 -17378 17693 -17322
rect 17621 -17412 17640 -17378
rect 17674 -17412 17693 -17378
rect 16731 -17502 16803 -17468
rect 17621 -17468 17693 -17412
rect 17621 -17502 17640 -17468
rect 17674 -17502 17693 -17468
rect 17757 -16708 17787 -16702
rect 17821 -16708 17888 -16674
rect 17922 -16702 19075 -16674
rect 17922 -16708 17955 -16702
rect 17757 -16764 17955 -16708
rect 17757 -16798 17787 -16764
rect 17821 -16798 17888 -16764
rect 17922 -16798 17955 -16764
rect 17757 -16854 17955 -16798
rect 17757 -16888 17787 -16854
rect 17821 -16888 17888 -16854
rect 17922 -16888 17955 -16854
rect 17757 -16944 17955 -16888
rect 17757 -16978 17787 -16944
rect 17821 -16978 17888 -16944
rect 17922 -16978 17955 -16944
rect 17757 -17034 17955 -16978
rect 17757 -17068 17787 -17034
rect 17821 -17068 17888 -17034
rect 17922 -17068 17955 -17034
rect 17757 -17124 17955 -17068
rect 17757 -17158 17787 -17124
rect 17821 -17158 17888 -17124
rect 17922 -17158 17955 -17124
rect 17757 -17214 17955 -17158
rect 17757 -17248 17787 -17214
rect 17821 -17248 17888 -17214
rect 17922 -17248 17955 -17214
rect 17757 -17304 17955 -17248
rect 17757 -17338 17787 -17304
rect 17821 -17338 17888 -17304
rect 17922 -17338 17955 -17304
rect 17757 -17394 17955 -17338
rect 17757 -17428 17787 -17394
rect 17821 -17428 17888 -17394
rect 17922 -17428 17955 -17394
rect 17757 -17484 17955 -17428
rect 17757 -17502 17787 -17484
rect 16634 -17518 17787 -17502
rect 17821 -17518 17888 -17484
rect 17922 -17502 17955 -17484
rect 18019 -16714 18091 -16702
rect 18019 -16748 18038 -16714
rect 18072 -16748 18091 -16714
rect 18019 -16804 18091 -16748
rect 18909 -16748 18981 -16702
rect 18019 -16838 18038 -16804
rect 18072 -16838 18091 -16804
rect 18019 -16894 18091 -16838
rect 18019 -16928 18038 -16894
rect 18072 -16928 18091 -16894
rect 18019 -16984 18091 -16928
rect 18019 -17018 18038 -16984
rect 18072 -17018 18091 -16984
rect 18019 -17074 18091 -17018
rect 18019 -17108 18038 -17074
rect 18072 -17108 18091 -17074
rect 18019 -17164 18091 -17108
rect 18019 -17198 18038 -17164
rect 18072 -17198 18091 -17164
rect 18019 -17254 18091 -17198
rect 18019 -17288 18038 -17254
rect 18072 -17288 18091 -17254
rect 18019 -17344 18091 -17288
rect 18019 -17378 18038 -17344
rect 18072 -17378 18091 -17344
rect 18019 -17434 18091 -17378
rect 18019 -17468 18038 -17434
rect 18072 -17468 18091 -17434
rect 18153 -16812 18847 -16751
rect 18153 -16846 18214 -16812
rect 18248 -16824 18304 -16812
rect 18338 -16824 18394 -16812
rect 18428 -16824 18484 -16812
rect 18260 -16846 18304 -16824
rect 18360 -16846 18394 -16824
rect 18460 -16846 18484 -16824
rect 18518 -16824 18574 -16812
rect 18518 -16846 18526 -16824
rect 18153 -16858 18226 -16846
rect 18260 -16858 18326 -16846
rect 18360 -16858 18426 -16846
rect 18460 -16858 18526 -16846
rect 18560 -16846 18574 -16824
rect 18608 -16824 18664 -16812
rect 18608 -16846 18626 -16824
rect 18560 -16858 18626 -16846
rect 18660 -16846 18664 -16824
rect 18698 -16824 18754 -16812
rect 18698 -16846 18726 -16824
rect 18788 -16846 18847 -16812
rect 18660 -16858 18726 -16846
rect 18760 -16858 18847 -16846
rect 18153 -16902 18847 -16858
rect 18153 -16936 18214 -16902
rect 18248 -16924 18304 -16902
rect 18338 -16924 18394 -16902
rect 18428 -16924 18484 -16902
rect 18260 -16936 18304 -16924
rect 18360 -16936 18394 -16924
rect 18460 -16936 18484 -16924
rect 18518 -16924 18574 -16902
rect 18518 -16936 18526 -16924
rect 18153 -16958 18226 -16936
rect 18260 -16958 18326 -16936
rect 18360 -16958 18426 -16936
rect 18460 -16958 18526 -16936
rect 18560 -16936 18574 -16924
rect 18608 -16924 18664 -16902
rect 18608 -16936 18626 -16924
rect 18560 -16958 18626 -16936
rect 18660 -16936 18664 -16924
rect 18698 -16924 18754 -16902
rect 18698 -16936 18726 -16924
rect 18788 -16936 18847 -16902
rect 18660 -16958 18726 -16936
rect 18760 -16958 18847 -16936
rect 18153 -16992 18847 -16958
rect 18153 -17026 18214 -16992
rect 18248 -17024 18304 -16992
rect 18338 -17024 18394 -16992
rect 18428 -17024 18484 -16992
rect 18260 -17026 18304 -17024
rect 18360 -17026 18394 -17024
rect 18460 -17026 18484 -17024
rect 18518 -17024 18574 -16992
rect 18518 -17026 18526 -17024
rect 18153 -17058 18226 -17026
rect 18260 -17058 18326 -17026
rect 18360 -17058 18426 -17026
rect 18460 -17058 18526 -17026
rect 18560 -17026 18574 -17024
rect 18608 -17024 18664 -16992
rect 18608 -17026 18626 -17024
rect 18560 -17058 18626 -17026
rect 18660 -17026 18664 -17024
rect 18698 -17024 18754 -16992
rect 18698 -17026 18726 -17024
rect 18788 -17026 18847 -16992
rect 18660 -17058 18726 -17026
rect 18760 -17058 18847 -17026
rect 18153 -17082 18847 -17058
rect 18153 -17116 18214 -17082
rect 18248 -17116 18304 -17082
rect 18338 -17116 18394 -17082
rect 18428 -17116 18484 -17082
rect 18518 -17116 18574 -17082
rect 18608 -17116 18664 -17082
rect 18698 -17116 18754 -17082
rect 18788 -17116 18847 -17082
rect 18153 -17124 18847 -17116
rect 18153 -17158 18226 -17124
rect 18260 -17158 18326 -17124
rect 18360 -17158 18426 -17124
rect 18460 -17158 18526 -17124
rect 18560 -17158 18626 -17124
rect 18660 -17158 18726 -17124
rect 18760 -17158 18847 -17124
rect 18153 -17172 18847 -17158
rect 18153 -17206 18214 -17172
rect 18248 -17206 18304 -17172
rect 18338 -17206 18394 -17172
rect 18428 -17206 18484 -17172
rect 18518 -17206 18574 -17172
rect 18608 -17206 18664 -17172
rect 18698 -17206 18754 -17172
rect 18788 -17206 18847 -17172
rect 18153 -17224 18847 -17206
rect 18153 -17258 18226 -17224
rect 18260 -17258 18326 -17224
rect 18360 -17258 18426 -17224
rect 18460 -17258 18526 -17224
rect 18560 -17258 18626 -17224
rect 18660 -17258 18726 -17224
rect 18760 -17258 18847 -17224
rect 18153 -17262 18847 -17258
rect 18153 -17296 18214 -17262
rect 18248 -17296 18304 -17262
rect 18338 -17296 18394 -17262
rect 18428 -17296 18484 -17262
rect 18518 -17296 18574 -17262
rect 18608 -17296 18664 -17262
rect 18698 -17296 18754 -17262
rect 18788 -17296 18847 -17262
rect 18153 -17324 18847 -17296
rect 18153 -17352 18226 -17324
rect 18260 -17352 18326 -17324
rect 18360 -17352 18426 -17324
rect 18460 -17352 18526 -17324
rect 18153 -17386 18214 -17352
rect 18260 -17358 18304 -17352
rect 18360 -17358 18394 -17352
rect 18460 -17358 18484 -17352
rect 18248 -17386 18304 -17358
rect 18338 -17386 18394 -17358
rect 18428 -17386 18484 -17358
rect 18518 -17358 18526 -17352
rect 18560 -17352 18626 -17324
rect 18560 -17358 18574 -17352
rect 18518 -17386 18574 -17358
rect 18608 -17358 18626 -17352
rect 18660 -17352 18726 -17324
rect 18760 -17352 18847 -17324
rect 18660 -17358 18664 -17352
rect 18608 -17386 18664 -17358
rect 18698 -17358 18726 -17352
rect 18698 -17386 18754 -17358
rect 18788 -17386 18847 -17352
rect 18153 -17445 18847 -17386
rect 18909 -16782 18928 -16748
rect 18962 -16782 18981 -16748
rect 18909 -16838 18981 -16782
rect 18909 -16872 18928 -16838
rect 18962 -16872 18981 -16838
rect 18909 -16928 18981 -16872
rect 18909 -16962 18928 -16928
rect 18962 -16962 18981 -16928
rect 18909 -17018 18981 -16962
rect 18909 -17052 18928 -17018
rect 18962 -17052 18981 -17018
rect 18909 -17108 18981 -17052
rect 18909 -17142 18928 -17108
rect 18962 -17142 18981 -17108
rect 18909 -17198 18981 -17142
rect 18909 -17232 18928 -17198
rect 18962 -17232 18981 -17198
rect 18909 -17288 18981 -17232
rect 18909 -17322 18928 -17288
rect 18962 -17322 18981 -17288
rect 18909 -17378 18981 -17322
rect 18909 -17412 18928 -17378
rect 18962 -17412 18981 -17378
rect 18019 -17502 18091 -17468
rect 18909 -17468 18981 -17412
rect 18909 -17502 18928 -17468
rect 18962 -17502 18981 -17468
rect 19045 -16708 19075 -16702
rect 19109 -16708 19176 -16674
rect 19210 -16702 20363 -16674
rect 19210 -16708 19243 -16702
rect 19045 -16764 19243 -16708
rect 19045 -16798 19075 -16764
rect 19109 -16798 19176 -16764
rect 19210 -16798 19243 -16764
rect 19045 -16854 19243 -16798
rect 19045 -16888 19075 -16854
rect 19109 -16888 19176 -16854
rect 19210 -16888 19243 -16854
rect 19045 -16944 19243 -16888
rect 19045 -16978 19075 -16944
rect 19109 -16978 19176 -16944
rect 19210 -16978 19243 -16944
rect 19045 -17034 19243 -16978
rect 19045 -17068 19075 -17034
rect 19109 -17068 19176 -17034
rect 19210 -17068 19243 -17034
rect 19045 -17124 19243 -17068
rect 19045 -17158 19075 -17124
rect 19109 -17158 19176 -17124
rect 19210 -17158 19243 -17124
rect 19045 -17214 19243 -17158
rect 19045 -17248 19075 -17214
rect 19109 -17248 19176 -17214
rect 19210 -17248 19243 -17214
rect 19045 -17304 19243 -17248
rect 19045 -17338 19075 -17304
rect 19109 -17338 19176 -17304
rect 19210 -17338 19243 -17304
rect 19045 -17394 19243 -17338
rect 19045 -17428 19075 -17394
rect 19109 -17428 19176 -17394
rect 19210 -17428 19243 -17394
rect 19045 -17484 19243 -17428
rect 19045 -17502 19075 -17484
rect 17922 -17518 19075 -17502
rect 19109 -17518 19176 -17484
rect 19210 -17502 19243 -17484
rect 19307 -16714 19379 -16702
rect 19307 -16748 19326 -16714
rect 19360 -16748 19379 -16714
rect 19307 -16804 19379 -16748
rect 20197 -16748 20269 -16702
rect 19307 -16838 19326 -16804
rect 19360 -16838 19379 -16804
rect 19307 -16894 19379 -16838
rect 19307 -16928 19326 -16894
rect 19360 -16928 19379 -16894
rect 19307 -16984 19379 -16928
rect 19307 -17018 19326 -16984
rect 19360 -17018 19379 -16984
rect 19307 -17074 19379 -17018
rect 19307 -17108 19326 -17074
rect 19360 -17108 19379 -17074
rect 19307 -17164 19379 -17108
rect 19307 -17198 19326 -17164
rect 19360 -17198 19379 -17164
rect 19307 -17254 19379 -17198
rect 19307 -17288 19326 -17254
rect 19360 -17288 19379 -17254
rect 19307 -17344 19379 -17288
rect 19307 -17378 19326 -17344
rect 19360 -17378 19379 -17344
rect 19307 -17434 19379 -17378
rect 19307 -17468 19326 -17434
rect 19360 -17468 19379 -17434
rect 19441 -16812 20135 -16751
rect 19441 -16846 19502 -16812
rect 19536 -16824 19592 -16812
rect 19626 -16824 19682 -16812
rect 19716 -16824 19772 -16812
rect 19548 -16846 19592 -16824
rect 19648 -16846 19682 -16824
rect 19748 -16846 19772 -16824
rect 19806 -16824 19862 -16812
rect 19806 -16846 19814 -16824
rect 19441 -16858 19514 -16846
rect 19548 -16858 19614 -16846
rect 19648 -16858 19714 -16846
rect 19748 -16858 19814 -16846
rect 19848 -16846 19862 -16824
rect 19896 -16824 19952 -16812
rect 19896 -16846 19914 -16824
rect 19848 -16858 19914 -16846
rect 19948 -16846 19952 -16824
rect 19986 -16824 20042 -16812
rect 19986 -16846 20014 -16824
rect 20076 -16846 20135 -16812
rect 19948 -16858 20014 -16846
rect 20048 -16858 20135 -16846
rect 19441 -16902 20135 -16858
rect 19441 -16936 19502 -16902
rect 19536 -16924 19592 -16902
rect 19626 -16924 19682 -16902
rect 19716 -16924 19772 -16902
rect 19548 -16936 19592 -16924
rect 19648 -16936 19682 -16924
rect 19748 -16936 19772 -16924
rect 19806 -16924 19862 -16902
rect 19806 -16936 19814 -16924
rect 19441 -16958 19514 -16936
rect 19548 -16958 19614 -16936
rect 19648 -16958 19714 -16936
rect 19748 -16958 19814 -16936
rect 19848 -16936 19862 -16924
rect 19896 -16924 19952 -16902
rect 19896 -16936 19914 -16924
rect 19848 -16958 19914 -16936
rect 19948 -16936 19952 -16924
rect 19986 -16924 20042 -16902
rect 19986 -16936 20014 -16924
rect 20076 -16936 20135 -16902
rect 19948 -16958 20014 -16936
rect 20048 -16958 20135 -16936
rect 19441 -16992 20135 -16958
rect 19441 -17026 19502 -16992
rect 19536 -17024 19592 -16992
rect 19626 -17024 19682 -16992
rect 19716 -17024 19772 -16992
rect 19548 -17026 19592 -17024
rect 19648 -17026 19682 -17024
rect 19748 -17026 19772 -17024
rect 19806 -17024 19862 -16992
rect 19806 -17026 19814 -17024
rect 19441 -17058 19514 -17026
rect 19548 -17058 19614 -17026
rect 19648 -17058 19714 -17026
rect 19748 -17058 19814 -17026
rect 19848 -17026 19862 -17024
rect 19896 -17024 19952 -16992
rect 19896 -17026 19914 -17024
rect 19848 -17058 19914 -17026
rect 19948 -17026 19952 -17024
rect 19986 -17024 20042 -16992
rect 19986 -17026 20014 -17024
rect 20076 -17026 20135 -16992
rect 19948 -17058 20014 -17026
rect 20048 -17058 20135 -17026
rect 19441 -17082 20135 -17058
rect 19441 -17116 19502 -17082
rect 19536 -17116 19592 -17082
rect 19626 -17116 19682 -17082
rect 19716 -17116 19772 -17082
rect 19806 -17116 19862 -17082
rect 19896 -17116 19952 -17082
rect 19986 -17116 20042 -17082
rect 20076 -17116 20135 -17082
rect 19441 -17124 20135 -17116
rect 19441 -17158 19514 -17124
rect 19548 -17158 19614 -17124
rect 19648 -17158 19714 -17124
rect 19748 -17158 19814 -17124
rect 19848 -17158 19914 -17124
rect 19948 -17158 20014 -17124
rect 20048 -17158 20135 -17124
rect 19441 -17172 20135 -17158
rect 19441 -17206 19502 -17172
rect 19536 -17206 19592 -17172
rect 19626 -17206 19682 -17172
rect 19716 -17206 19772 -17172
rect 19806 -17206 19862 -17172
rect 19896 -17206 19952 -17172
rect 19986 -17206 20042 -17172
rect 20076 -17206 20135 -17172
rect 19441 -17224 20135 -17206
rect 19441 -17258 19514 -17224
rect 19548 -17258 19614 -17224
rect 19648 -17258 19714 -17224
rect 19748 -17258 19814 -17224
rect 19848 -17258 19914 -17224
rect 19948 -17258 20014 -17224
rect 20048 -17258 20135 -17224
rect 19441 -17262 20135 -17258
rect 19441 -17296 19502 -17262
rect 19536 -17296 19592 -17262
rect 19626 -17296 19682 -17262
rect 19716 -17296 19772 -17262
rect 19806 -17296 19862 -17262
rect 19896 -17296 19952 -17262
rect 19986 -17296 20042 -17262
rect 20076 -17296 20135 -17262
rect 19441 -17324 20135 -17296
rect 19441 -17352 19514 -17324
rect 19548 -17352 19614 -17324
rect 19648 -17352 19714 -17324
rect 19748 -17352 19814 -17324
rect 19441 -17386 19502 -17352
rect 19548 -17358 19592 -17352
rect 19648 -17358 19682 -17352
rect 19748 -17358 19772 -17352
rect 19536 -17386 19592 -17358
rect 19626 -17386 19682 -17358
rect 19716 -17386 19772 -17358
rect 19806 -17358 19814 -17352
rect 19848 -17352 19914 -17324
rect 19848 -17358 19862 -17352
rect 19806 -17386 19862 -17358
rect 19896 -17358 19914 -17352
rect 19948 -17352 20014 -17324
rect 20048 -17352 20135 -17324
rect 19948 -17358 19952 -17352
rect 19896 -17386 19952 -17358
rect 19986 -17358 20014 -17352
rect 19986 -17386 20042 -17358
rect 20076 -17386 20135 -17352
rect 19441 -17445 20135 -17386
rect 20197 -16782 20216 -16748
rect 20250 -16782 20269 -16748
rect 20197 -16838 20269 -16782
rect 20197 -16872 20216 -16838
rect 20250 -16872 20269 -16838
rect 20197 -16928 20269 -16872
rect 20197 -16962 20216 -16928
rect 20250 -16962 20269 -16928
rect 20197 -17018 20269 -16962
rect 20197 -17052 20216 -17018
rect 20250 -17052 20269 -17018
rect 20197 -17108 20269 -17052
rect 20197 -17142 20216 -17108
rect 20250 -17142 20269 -17108
rect 20197 -17198 20269 -17142
rect 20197 -17232 20216 -17198
rect 20250 -17232 20269 -17198
rect 20197 -17288 20269 -17232
rect 20197 -17322 20216 -17288
rect 20250 -17322 20269 -17288
rect 20197 -17378 20269 -17322
rect 20197 -17412 20216 -17378
rect 20250 -17412 20269 -17378
rect 19307 -17502 19379 -17468
rect 20197 -17468 20269 -17412
rect 20197 -17502 20216 -17468
rect 20250 -17502 20269 -17468
rect 20333 -16708 20363 -16702
rect 20397 -16708 20464 -16674
rect 20498 -16702 21651 -16674
rect 20498 -16708 20531 -16702
rect 20333 -16764 20531 -16708
rect 20333 -16798 20363 -16764
rect 20397 -16798 20464 -16764
rect 20498 -16798 20531 -16764
rect 20333 -16854 20531 -16798
rect 20333 -16888 20363 -16854
rect 20397 -16888 20464 -16854
rect 20498 -16888 20531 -16854
rect 20333 -16944 20531 -16888
rect 20333 -16978 20363 -16944
rect 20397 -16978 20464 -16944
rect 20498 -16978 20531 -16944
rect 20333 -17034 20531 -16978
rect 20333 -17068 20363 -17034
rect 20397 -17068 20464 -17034
rect 20498 -17068 20531 -17034
rect 20333 -17124 20531 -17068
rect 20333 -17158 20363 -17124
rect 20397 -17158 20464 -17124
rect 20498 -17158 20531 -17124
rect 20333 -17214 20531 -17158
rect 20333 -17248 20363 -17214
rect 20397 -17248 20464 -17214
rect 20498 -17248 20531 -17214
rect 20333 -17304 20531 -17248
rect 20333 -17338 20363 -17304
rect 20397 -17338 20464 -17304
rect 20498 -17338 20531 -17304
rect 20333 -17394 20531 -17338
rect 20333 -17428 20363 -17394
rect 20397 -17428 20464 -17394
rect 20498 -17428 20531 -17394
rect 20333 -17484 20531 -17428
rect 20333 -17502 20363 -17484
rect 19210 -17518 20363 -17502
rect 20397 -17518 20464 -17484
rect 20498 -17502 20531 -17484
rect 20595 -16714 20667 -16702
rect 20595 -16748 20614 -16714
rect 20648 -16748 20667 -16714
rect 20595 -16804 20667 -16748
rect 21485 -16748 21557 -16702
rect 20595 -16838 20614 -16804
rect 20648 -16838 20667 -16804
rect 20595 -16894 20667 -16838
rect 20595 -16928 20614 -16894
rect 20648 -16928 20667 -16894
rect 20595 -16984 20667 -16928
rect 20595 -17018 20614 -16984
rect 20648 -17018 20667 -16984
rect 20595 -17074 20667 -17018
rect 20595 -17108 20614 -17074
rect 20648 -17108 20667 -17074
rect 20595 -17164 20667 -17108
rect 20595 -17198 20614 -17164
rect 20648 -17198 20667 -17164
rect 20595 -17254 20667 -17198
rect 20595 -17288 20614 -17254
rect 20648 -17288 20667 -17254
rect 20595 -17344 20667 -17288
rect 20595 -17378 20614 -17344
rect 20648 -17378 20667 -17344
rect 20595 -17434 20667 -17378
rect 20595 -17468 20614 -17434
rect 20648 -17468 20667 -17434
rect 20729 -16812 21423 -16751
rect 20729 -16846 20790 -16812
rect 20824 -16824 20880 -16812
rect 20914 -16824 20970 -16812
rect 21004 -16824 21060 -16812
rect 20836 -16846 20880 -16824
rect 20936 -16846 20970 -16824
rect 21036 -16846 21060 -16824
rect 21094 -16824 21150 -16812
rect 21094 -16846 21102 -16824
rect 20729 -16858 20802 -16846
rect 20836 -16858 20902 -16846
rect 20936 -16858 21002 -16846
rect 21036 -16858 21102 -16846
rect 21136 -16846 21150 -16824
rect 21184 -16824 21240 -16812
rect 21184 -16846 21202 -16824
rect 21136 -16858 21202 -16846
rect 21236 -16846 21240 -16824
rect 21274 -16824 21330 -16812
rect 21274 -16846 21302 -16824
rect 21364 -16846 21423 -16812
rect 21236 -16858 21302 -16846
rect 21336 -16858 21423 -16846
rect 20729 -16902 21423 -16858
rect 20729 -16936 20790 -16902
rect 20824 -16924 20880 -16902
rect 20914 -16924 20970 -16902
rect 21004 -16924 21060 -16902
rect 20836 -16936 20880 -16924
rect 20936 -16936 20970 -16924
rect 21036 -16936 21060 -16924
rect 21094 -16924 21150 -16902
rect 21094 -16936 21102 -16924
rect 20729 -16958 20802 -16936
rect 20836 -16958 20902 -16936
rect 20936 -16958 21002 -16936
rect 21036 -16958 21102 -16936
rect 21136 -16936 21150 -16924
rect 21184 -16924 21240 -16902
rect 21184 -16936 21202 -16924
rect 21136 -16958 21202 -16936
rect 21236 -16936 21240 -16924
rect 21274 -16924 21330 -16902
rect 21274 -16936 21302 -16924
rect 21364 -16936 21423 -16902
rect 21236 -16958 21302 -16936
rect 21336 -16958 21423 -16936
rect 20729 -16992 21423 -16958
rect 20729 -17026 20790 -16992
rect 20824 -17024 20880 -16992
rect 20914 -17024 20970 -16992
rect 21004 -17024 21060 -16992
rect 20836 -17026 20880 -17024
rect 20936 -17026 20970 -17024
rect 21036 -17026 21060 -17024
rect 21094 -17024 21150 -16992
rect 21094 -17026 21102 -17024
rect 20729 -17058 20802 -17026
rect 20836 -17058 20902 -17026
rect 20936 -17058 21002 -17026
rect 21036 -17058 21102 -17026
rect 21136 -17026 21150 -17024
rect 21184 -17024 21240 -16992
rect 21184 -17026 21202 -17024
rect 21136 -17058 21202 -17026
rect 21236 -17026 21240 -17024
rect 21274 -17024 21330 -16992
rect 21274 -17026 21302 -17024
rect 21364 -17026 21423 -16992
rect 21236 -17058 21302 -17026
rect 21336 -17058 21423 -17026
rect 20729 -17082 21423 -17058
rect 20729 -17116 20790 -17082
rect 20824 -17116 20880 -17082
rect 20914 -17116 20970 -17082
rect 21004 -17116 21060 -17082
rect 21094 -17116 21150 -17082
rect 21184 -17116 21240 -17082
rect 21274 -17116 21330 -17082
rect 21364 -17116 21423 -17082
rect 20729 -17124 21423 -17116
rect 20729 -17158 20802 -17124
rect 20836 -17158 20902 -17124
rect 20936 -17158 21002 -17124
rect 21036 -17158 21102 -17124
rect 21136 -17158 21202 -17124
rect 21236 -17158 21302 -17124
rect 21336 -17158 21423 -17124
rect 20729 -17172 21423 -17158
rect 20729 -17206 20790 -17172
rect 20824 -17206 20880 -17172
rect 20914 -17206 20970 -17172
rect 21004 -17206 21060 -17172
rect 21094 -17206 21150 -17172
rect 21184 -17206 21240 -17172
rect 21274 -17206 21330 -17172
rect 21364 -17206 21423 -17172
rect 20729 -17224 21423 -17206
rect 20729 -17258 20802 -17224
rect 20836 -17258 20902 -17224
rect 20936 -17258 21002 -17224
rect 21036 -17258 21102 -17224
rect 21136 -17258 21202 -17224
rect 21236 -17258 21302 -17224
rect 21336 -17258 21423 -17224
rect 20729 -17262 21423 -17258
rect 20729 -17296 20790 -17262
rect 20824 -17296 20880 -17262
rect 20914 -17296 20970 -17262
rect 21004 -17296 21060 -17262
rect 21094 -17296 21150 -17262
rect 21184 -17296 21240 -17262
rect 21274 -17296 21330 -17262
rect 21364 -17296 21423 -17262
rect 20729 -17324 21423 -17296
rect 20729 -17352 20802 -17324
rect 20836 -17352 20902 -17324
rect 20936 -17352 21002 -17324
rect 21036 -17352 21102 -17324
rect 20729 -17386 20790 -17352
rect 20836 -17358 20880 -17352
rect 20936 -17358 20970 -17352
rect 21036 -17358 21060 -17352
rect 20824 -17386 20880 -17358
rect 20914 -17386 20970 -17358
rect 21004 -17386 21060 -17358
rect 21094 -17358 21102 -17352
rect 21136 -17352 21202 -17324
rect 21136 -17358 21150 -17352
rect 21094 -17386 21150 -17358
rect 21184 -17358 21202 -17352
rect 21236 -17352 21302 -17324
rect 21336 -17352 21423 -17324
rect 21236 -17358 21240 -17352
rect 21184 -17386 21240 -17358
rect 21274 -17358 21302 -17352
rect 21274 -17386 21330 -17358
rect 21364 -17386 21423 -17352
rect 20729 -17445 21423 -17386
rect 21485 -16782 21504 -16748
rect 21538 -16782 21557 -16748
rect 21485 -16838 21557 -16782
rect 21485 -16872 21504 -16838
rect 21538 -16872 21557 -16838
rect 21485 -16928 21557 -16872
rect 21485 -16962 21504 -16928
rect 21538 -16962 21557 -16928
rect 21485 -17018 21557 -16962
rect 21485 -17052 21504 -17018
rect 21538 -17052 21557 -17018
rect 21485 -17108 21557 -17052
rect 21485 -17142 21504 -17108
rect 21538 -17142 21557 -17108
rect 21485 -17198 21557 -17142
rect 21485 -17232 21504 -17198
rect 21538 -17232 21557 -17198
rect 21485 -17288 21557 -17232
rect 21485 -17322 21504 -17288
rect 21538 -17322 21557 -17288
rect 21485 -17378 21557 -17322
rect 21485 -17412 21504 -17378
rect 21538 -17412 21557 -17378
rect 20595 -17502 20667 -17468
rect 21485 -17468 21557 -17412
rect 21485 -17502 21504 -17468
rect 21538 -17502 21557 -17468
rect 21621 -16708 21651 -16702
rect 21685 -16708 21752 -16674
rect 21786 -16702 22939 -16674
rect 21786 -16708 21819 -16702
rect 21621 -16764 21819 -16708
rect 21621 -16798 21651 -16764
rect 21685 -16798 21752 -16764
rect 21786 -16798 21819 -16764
rect 21621 -16854 21819 -16798
rect 21621 -16888 21651 -16854
rect 21685 -16888 21752 -16854
rect 21786 -16888 21819 -16854
rect 21621 -16944 21819 -16888
rect 21621 -16978 21651 -16944
rect 21685 -16978 21752 -16944
rect 21786 -16978 21819 -16944
rect 21621 -17034 21819 -16978
rect 21621 -17068 21651 -17034
rect 21685 -17068 21752 -17034
rect 21786 -17068 21819 -17034
rect 21621 -17124 21819 -17068
rect 21621 -17158 21651 -17124
rect 21685 -17158 21752 -17124
rect 21786 -17158 21819 -17124
rect 21621 -17214 21819 -17158
rect 21621 -17248 21651 -17214
rect 21685 -17248 21752 -17214
rect 21786 -17248 21819 -17214
rect 21621 -17304 21819 -17248
rect 21621 -17338 21651 -17304
rect 21685 -17338 21752 -17304
rect 21786 -17338 21819 -17304
rect 21621 -17394 21819 -17338
rect 21621 -17428 21651 -17394
rect 21685 -17428 21752 -17394
rect 21786 -17428 21819 -17394
rect 21621 -17484 21819 -17428
rect 21621 -17502 21651 -17484
rect 20498 -17518 21651 -17502
rect 21685 -17518 21752 -17484
rect 21786 -17502 21819 -17484
rect 21883 -16714 21955 -16702
rect 21883 -16748 21902 -16714
rect 21936 -16748 21955 -16714
rect 21883 -16804 21955 -16748
rect 22773 -16748 22845 -16702
rect 21883 -16838 21902 -16804
rect 21936 -16838 21955 -16804
rect 21883 -16894 21955 -16838
rect 21883 -16928 21902 -16894
rect 21936 -16928 21955 -16894
rect 21883 -16984 21955 -16928
rect 21883 -17018 21902 -16984
rect 21936 -17018 21955 -16984
rect 21883 -17074 21955 -17018
rect 21883 -17108 21902 -17074
rect 21936 -17108 21955 -17074
rect 21883 -17164 21955 -17108
rect 21883 -17198 21902 -17164
rect 21936 -17198 21955 -17164
rect 21883 -17254 21955 -17198
rect 21883 -17288 21902 -17254
rect 21936 -17288 21955 -17254
rect 21883 -17344 21955 -17288
rect 21883 -17378 21902 -17344
rect 21936 -17378 21955 -17344
rect 21883 -17434 21955 -17378
rect 21883 -17468 21902 -17434
rect 21936 -17468 21955 -17434
rect 22017 -16812 22711 -16751
rect 22017 -16846 22078 -16812
rect 22112 -16824 22168 -16812
rect 22202 -16824 22258 -16812
rect 22292 -16824 22348 -16812
rect 22124 -16846 22168 -16824
rect 22224 -16846 22258 -16824
rect 22324 -16846 22348 -16824
rect 22382 -16824 22438 -16812
rect 22382 -16846 22390 -16824
rect 22017 -16858 22090 -16846
rect 22124 -16858 22190 -16846
rect 22224 -16858 22290 -16846
rect 22324 -16858 22390 -16846
rect 22424 -16846 22438 -16824
rect 22472 -16824 22528 -16812
rect 22472 -16846 22490 -16824
rect 22424 -16858 22490 -16846
rect 22524 -16846 22528 -16824
rect 22562 -16824 22618 -16812
rect 22562 -16846 22590 -16824
rect 22652 -16846 22711 -16812
rect 22524 -16858 22590 -16846
rect 22624 -16858 22711 -16846
rect 22017 -16902 22711 -16858
rect 22017 -16936 22078 -16902
rect 22112 -16924 22168 -16902
rect 22202 -16924 22258 -16902
rect 22292 -16924 22348 -16902
rect 22124 -16936 22168 -16924
rect 22224 -16936 22258 -16924
rect 22324 -16936 22348 -16924
rect 22382 -16924 22438 -16902
rect 22382 -16936 22390 -16924
rect 22017 -16958 22090 -16936
rect 22124 -16958 22190 -16936
rect 22224 -16958 22290 -16936
rect 22324 -16958 22390 -16936
rect 22424 -16936 22438 -16924
rect 22472 -16924 22528 -16902
rect 22472 -16936 22490 -16924
rect 22424 -16958 22490 -16936
rect 22524 -16936 22528 -16924
rect 22562 -16924 22618 -16902
rect 22562 -16936 22590 -16924
rect 22652 -16936 22711 -16902
rect 22524 -16958 22590 -16936
rect 22624 -16958 22711 -16936
rect 22017 -16992 22711 -16958
rect 22017 -17026 22078 -16992
rect 22112 -17024 22168 -16992
rect 22202 -17024 22258 -16992
rect 22292 -17024 22348 -16992
rect 22124 -17026 22168 -17024
rect 22224 -17026 22258 -17024
rect 22324 -17026 22348 -17024
rect 22382 -17024 22438 -16992
rect 22382 -17026 22390 -17024
rect 22017 -17058 22090 -17026
rect 22124 -17058 22190 -17026
rect 22224 -17058 22290 -17026
rect 22324 -17058 22390 -17026
rect 22424 -17026 22438 -17024
rect 22472 -17024 22528 -16992
rect 22472 -17026 22490 -17024
rect 22424 -17058 22490 -17026
rect 22524 -17026 22528 -17024
rect 22562 -17024 22618 -16992
rect 22562 -17026 22590 -17024
rect 22652 -17026 22711 -16992
rect 22524 -17058 22590 -17026
rect 22624 -17058 22711 -17026
rect 22017 -17082 22711 -17058
rect 22017 -17116 22078 -17082
rect 22112 -17116 22168 -17082
rect 22202 -17116 22258 -17082
rect 22292 -17116 22348 -17082
rect 22382 -17116 22438 -17082
rect 22472 -17116 22528 -17082
rect 22562 -17116 22618 -17082
rect 22652 -17116 22711 -17082
rect 22017 -17124 22711 -17116
rect 22017 -17158 22090 -17124
rect 22124 -17158 22190 -17124
rect 22224 -17158 22290 -17124
rect 22324 -17158 22390 -17124
rect 22424 -17158 22490 -17124
rect 22524 -17158 22590 -17124
rect 22624 -17158 22711 -17124
rect 22017 -17172 22711 -17158
rect 22017 -17206 22078 -17172
rect 22112 -17206 22168 -17172
rect 22202 -17206 22258 -17172
rect 22292 -17206 22348 -17172
rect 22382 -17206 22438 -17172
rect 22472 -17206 22528 -17172
rect 22562 -17206 22618 -17172
rect 22652 -17206 22711 -17172
rect 22017 -17224 22711 -17206
rect 22017 -17258 22090 -17224
rect 22124 -17258 22190 -17224
rect 22224 -17258 22290 -17224
rect 22324 -17258 22390 -17224
rect 22424 -17258 22490 -17224
rect 22524 -17258 22590 -17224
rect 22624 -17258 22711 -17224
rect 22017 -17262 22711 -17258
rect 22017 -17296 22078 -17262
rect 22112 -17296 22168 -17262
rect 22202 -17296 22258 -17262
rect 22292 -17296 22348 -17262
rect 22382 -17296 22438 -17262
rect 22472 -17296 22528 -17262
rect 22562 -17296 22618 -17262
rect 22652 -17296 22711 -17262
rect 22017 -17324 22711 -17296
rect 22017 -17352 22090 -17324
rect 22124 -17352 22190 -17324
rect 22224 -17352 22290 -17324
rect 22324 -17352 22390 -17324
rect 22017 -17386 22078 -17352
rect 22124 -17358 22168 -17352
rect 22224 -17358 22258 -17352
rect 22324 -17358 22348 -17352
rect 22112 -17386 22168 -17358
rect 22202 -17386 22258 -17358
rect 22292 -17386 22348 -17358
rect 22382 -17358 22390 -17352
rect 22424 -17352 22490 -17324
rect 22424 -17358 22438 -17352
rect 22382 -17386 22438 -17358
rect 22472 -17358 22490 -17352
rect 22524 -17352 22590 -17324
rect 22624 -17352 22711 -17324
rect 22524 -17358 22528 -17352
rect 22472 -17386 22528 -17358
rect 22562 -17358 22590 -17352
rect 22562 -17386 22618 -17358
rect 22652 -17386 22711 -17352
rect 22017 -17445 22711 -17386
rect 22773 -16782 22792 -16748
rect 22826 -16782 22845 -16748
rect 22773 -16838 22845 -16782
rect 22773 -16872 22792 -16838
rect 22826 -16872 22845 -16838
rect 22773 -16928 22845 -16872
rect 22773 -16962 22792 -16928
rect 22826 -16962 22845 -16928
rect 22773 -17018 22845 -16962
rect 22773 -17052 22792 -17018
rect 22826 -17052 22845 -17018
rect 22773 -17108 22845 -17052
rect 22773 -17142 22792 -17108
rect 22826 -17142 22845 -17108
rect 22773 -17198 22845 -17142
rect 22773 -17232 22792 -17198
rect 22826 -17232 22845 -17198
rect 22773 -17288 22845 -17232
rect 22773 -17322 22792 -17288
rect 22826 -17322 22845 -17288
rect 22773 -17378 22845 -17322
rect 22773 -17412 22792 -17378
rect 22826 -17412 22845 -17378
rect 21883 -17502 21955 -17468
rect 22773 -17468 22845 -17412
rect 22773 -17502 22792 -17468
rect 22826 -17502 22845 -17468
rect 22909 -16708 22939 -16702
rect 22973 -16708 23040 -16674
rect 23074 -16702 24227 -16674
rect 23074 -16708 23107 -16702
rect 22909 -16764 23107 -16708
rect 22909 -16798 22939 -16764
rect 22973 -16798 23040 -16764
rect 23074 -16798 23107 -16764
rect 22909 -16854 23107 -16798
rect 22909 -16888 22939 -16854
rect 22973 -16888 23040 -16854
rect 23074 -16888 23107 -16854
rect 22909 -16944 23107 -16888
rect 22909 -16978 22939 -16944
rect 22973 -16978 23040 -16944
rect 23074 -16978 23107 -16944
rect 22909 -17034 23107 -16978
rect 22909 -17068 22939 -17034
rect 22973 -17068 23040 -17034
rect 23074 -17068 23107 -17034
rect 22909 -17124 23107 -17068
rect 22909 -17158 22939 -17124
rect 22973 -17158 23040 -17124
rect 23074 -17158 23107 -17124
rect 22909 -17214 23107 -17158
rect 22909 -17248 22939 -17214
rect 22973 -17248 23040 -17214
rect 23074 -17248 23107 -17214
rect 22909 -17304 23107 -17248
rect 22909 -17338 22939 -17304
rect 22973 -17338 23040 -17304
rect 23074 -17338 23107 -17304
rect 22909 -17394 23107 -17338
rect 22909 -17428 22939 -17394
rect 22973 -17428 23040 -17394
rect 23074 -17428 23107 -17394
rect 22909 -17484 23107 -17428
rect 22909 -17502 22939 -17484
rect 21786 -17518 22939 -17502
rect 22973 -17518 23040 -17484
rect 23074 -17502 23107 -17484
rect 23171 -16714 23243 -16702
rect 23171 -16748 23190 -16714
rect 23224 -16748 23243 -16714
rect 23171 -16804 23243 -16748
rect 24061 -16748 24133 -16702
rect 23171 -16838 23190 -16804
rect 23224 -16838 23243 -16804
rect 23171 -16894 23243 -16838
rect 23171 -16928 23190 -16894
rect 23224 -16928 23243 -16894
rect 23171 -16984 23243 -16928
rect 23171 -17018 23190 -16984
rect 23224 -17018 23243 -16984
rect 23171 -17074 23243 -17018
rect 23171 -17108 23190 -17074
rect 23224 -17108 23243 -17074
rect 23171 -17164 23243 -17108
rect 23171 -17198 23190 -17164
rect 23224 -17198 23243 -17164
rect 23171 -17254 23243 -17198
rect 23171 -17288 23190 -17254
rect 23224 -17288 23243 -17254
rect 23171 -17344 23243 -17288
rect 23171 -17378 23190 -17344
rect 23224 -17378 23243 -17344
rect 23171 -17434 23243 -17378
rect 23171 -17468 23190 -17434
rect 23224 -17468 23243 -17434
rect 23305 -16812 23999 -16751
rect 23305 -16846 23366 -16812
rect 23400 -16824 23456 -16812
rect 23490 -16824 23546 -16812
rect 23580 -16824 23636 -16812
rect 23412 -16846 23456 -16824
rect 23512 -16846 23546 -16824
rect 23612 -16846 23636 -16824
rect 23670 -16824 23726 -16812
rect 23670 -16846 23678 -16824
rect 23305 -16858 23378 -16846
rect 23412 -16858 23478 -16846
rect 23512 -16858 23578 -16846
rect 23612 -16858 23678 -16846
rect 23712 -16846 23726 -16824
rect 23760 -16824 23816 -16812
rect 23760 -16846 23778 -16824
rect 23712 -16858 23778 -16846
rect 23812 -16846 23816 -16824
rect 23850 -16824 23906 -16812
rect 23850 -16846 23878 -16824
rect 23940 -16846 23999 -16812
rect 23812 -16858 23878 -16846
rect 23912 -16858 23999 -16846
rect 23305 -16902 23999 -16858
rect 23305 -16936 23366 -16902
rect 23400 -16924 23456 -16902
rect 23490 -16924 23546 -16902
rect 23580 -16924 23636 -16902
rect 23412 -16936 23456 -16924
rect 23512 -16936 23546 -16924
rect 23612 -16936 23636 -16924
rect 23670 -16924 23726 -16902
rect 23670 -16936 23678 -16924
rect 23305 -16958 23378 -16936
rect 23412 -16958 23478 -16936
rect 23512 -16958 23578 -16936
rect 23612 -16958 23678 -16936
rect 23712 -16936 23726 -16924
rect 23760 -16924 23816 -16902
rect 23760 -16936 23778 -16924
rect 23712 -16958 23778 -16936
rect 23812 -16936 23816 -16924
rect 23850 -16924 23906 -16902
rect 23850 -16936 23878 -16924
rect 23940 -16936 23999 -16902
rect 23812 -16958 23878 -16936
rect 23912 -16958 23999 -16936
rect 23305 -16992 23999 -16958
rect 23305 -17026 23366 -16992
rect 23400 -17024 23456 -16992
rect 23490 -17024 23546 -16992
rect 23580 -17024 23636 -16992
rect 23412 -17026 23456 -17024
rect 23512 -17026 23546 -17024
rect 23612 -17026 23636 -17024
rect 23670 -17024 23726 -16992
rect 23670 -17026 23678 -17024
rect 23305 -17058 23378 -17026
rect 23412 -17058 23478 -17026
rect 23512 -17058 23578 -17026
rect 23612 -17058 23678 -17026
rect 23712 -17026 23726 -17024
rect 23760 -17024 23816 -16992
rect 23760 -17026 23778 -17024
rect 23712 -17058 23778 -17026
rect 23812 -17026 23816 -17024
rect 23850 -17024 23906 -16992
rect 23850 -17026 23878 -17024
rect 23940 -17026 23999 -16992
rect 23812 -17058 23878 -17026
rect 23912 -17058 23999 -17026
rect 23305 -17082 23999 -17058
rect 23305 -17116 23366 -17082
rect 23400 -17116 23456 -17082
rect 23490 -17116 23546 -17082
rect 23580 -17116 23636 -17082
rect 23670 -17116 23726 -17082
rect 23760 -17116 23816 -17082
rect 23850 -17116 23906 -17082
rect 23940 -17116 23999 -17082
rect 23305 -17124 23999 -17116
rect 23305 -17158 23378 -17124
rect 23412 -17158 23478 -17124
rect 23512 -17158 23578 -17124
rect 23612 -17158 23678 -17124
rect 23712 -17158 23778 -17124
rect 23812 -17158 23878 -17124
rect 23912 -17158 23999 -17124
rect 23305 -17172 23999 -17158
rect 23305 -17206 23366 -17172
rect 23400 -17206 23456 -17172
rect 23490 -17206 23546 -17172
rect 23580 -17206 23636 -17172
rect 23670 -17206 23726 -17172
rect 23760 -17206 23816 -17172
rect 23850 -17206 23906 -17172
rect 23940 -17206 23999 -17172
rect 23305 -17224 23999 -17206
rect 23305 -17258 23378 -17224
rect 23412 -17258 23478 -17224
rect 23512 -17258 23578 -17224
rect 23612 -17258 23678 -17224
rect 23712 -17258 23778 -17224
rect 23812 -17258 23878 -17224
rect 23912 -17258 23999 -17224
rect 23305 -17262 23999 -17258
rect 23305 -17296 23366 -17262
rect 23400 -17296 23456 -17262
rect 23490 -17296 23546 -17262
rect 23580 -17296 23636 -17262
rect 23670 -17296 23726 -17262
rect 23760 -17296 23816 -17262
rect 23850 -17296 23906 -17262
rect 23940 -17296 23999 -17262
rect 23305 -17324 23999 -17296
rect 23305 -17352 23378 -17324
rect 23412 -17352 23478 -17324
rect 23512 -17352 23578 -17324
rect 23612 -17352 23678 -17324
rect 23305 -17386 23366 -17352
rect 23412 -17358 23456 -17352
rect 23512 -17358 23546 -17352
rect 23612 -17358 23636 -17352
rect 23400 -17386 23456 -17358
rect 23490 -17386 23546 -17358
rect 23580 -17386 23636 -17358
rect 23670 -17358 23678 -17352
rect 23712 -17352 23778 -17324
rect 23712 -17358 23726 -17352
rect 23670 -17386 23726 -17358
rect 23760 -17358 23778 -17352
rect 23812 -17352 23878 -17324
rect 23912 -17352 23999 -17324
rect 23812 -17358 23816 -17352
rect 23760 -17386 23816 -17358
rect 23850 -17358 23878 -17352
rect 23850 -17386 23906 -17358
rect 23940 -17386 23999 -17352
rect 23305 -17445 23999 -17386
rect 24061 -16782 24080 -16748
rect 24114 -16782 24133 -16748
rect 24061 -16838 24133 -16782
rect 24061 -16872 24080 -16838
rect 24114 -16872 24133 -16838
rect 24061 -16928 24133 -16872
rect 24061 -16962 24080 -16928
rect 24114 -16962 24133 -16928
rect 24061 -17018 24133 -16962
rect 24061 -17052 24080 -17018
rect 24114 -17052 24133 -17018
rect 24061 -17108 24133 -17052
rect 24061 -17142 24080 -17108
rect 24114 -17142 24133 -17108
rect 24061 -17198 24133 -17142
rect 24061 -17232 24080 -17198
rect 24114 -17232 24133 -17198
rect 24061 -17288 24133 -17232
rect 24061 -17322 24080 -17288
rect 24114 -17322 24133 -17288
rect 24061 -17378 24133 -17322
rect 24061 -17412 24080 -17378
rect 24114 -17412 24133 -17378
rect 23171 -17502 23243 -17468
rect 24061 -17468 24133 -17412
rect 24061 -17502 24080 -17468
rect 24114 -17502 24133 -17468
rect 24197 -16708 24227 -16702
rect 24261 -16708 24328 -16674
rect 24362 -16702 25515 -16674
rect 24362 -16708 24395 -16702
rect 24197 -16764 24395 -16708
rect 24197 -16798 24227 -16764
rect 24261 -16798 24328 -16764
rect 24362 -16798 24395 -16764
rect 24197 -16854 24395 -16798
rect 24197 -16888 24227 -16854
rect 24261 -16888 24328 -16854
rect 24362 -16888 24395 -16854
rect 24197 -16944 24395 -16888
rect 24197 -16978 24227 -16944
rect 24261 -16978 24328 -16944
rect 24362 -16978 24395 -16944
rect 24197 -17034 24395 -16978
rect 24197 -17068 24227 -17034
rect 24261 -17068 24328 -17034
rect 24362 -17068 24395 -17034
rect 24197 -17124 24395 -17068
rect 24197 -17158 24227 -17124
rect 24261 -17158 24328 -17124
rect 24362 -17158 24395 -17124
rect 24197 -17214 24395 -17158
rect 24197 -17248 24227 -17214
rect 24261 -17248 24328 -17214
rect 24362 -17248 24395 -17214
rect 24197 -17304 24395 -17248
rect 24197 -17338 24227 -17304
rect 24261 -17338 24328 -17304
rect 24362 -17338 24395 -17304
rect 24197 -17394 24395 -17338
rect 24197 -17428 24227 -17394
rect 24261 -17428 24328 -17394
rect 24362 -17428 24395 -17394
rect 24197 -17484 24395 -17428
rect 24197 -17502 24227 -17484
rect 23074 -17518 24227 -17502
rect 24261 -17518 24328 -17484
rect 24362 -17502 24395 -17484
rect 24459 -16714 24531 -16702
rect 24459 -16748 24478 -16714
rect 24512 -16748 24531 -16714
rect 24459 -16804 24531 -16748
rect 25349 -16748 25421 -16702
rect 24459 -16838 24478 -16804
rect 24512 -16838 24531 -16804
rect 24459 -16894 24531 -16838
rect 24459 -16928 24478 -16894
rect 24512 -16928 24531 -16894
rect 24459 -16984 24531 -16928
rect 24459 -17018 24478 -16984
rect 24512 -17018 24531 -16984
rect 24459 -17074 24531 -17018
rect 24459 -17108 24478 -17074
rect 24512 -17108 24531 -17074
rect 24459 -17164 24531 -17108
rect 24459 -17198 24478 -17164
rect 24512 -17198 24531 -17164
rect 24459 -17254 24531 -17198
rect 24459 -17288 24478 -17254
rect 24512 -17288 24531 -17254
rect 24459 -17344 24531 -17288
rect 24459 -17378 24478 -17344
rect 24512 -17378 24531 -17344
rect 24459 -17434 24531 -17378
rect 24459 -17468 24478 -17434
rect 24512 -17468 24531 -17434
rect 24593 -16812 25287 -16751
rect 24593 -16846 24654 -16812
rect 24688 -16824 24744 -16812
rect 24778 -16824 24834 -16812
rect 24868 -16824 24924 -16812
rect 24700 -16846 24744 -16824
rect 24800 -16846 24834 -16824
rect 24900 -16846 24924 -16824
rect 24958 -16824 25014 -16812
rect 24958 -16846 24966 -16824
rect 24593 -16858 24666 -16846
rect 24700 -16858 24766 -16846
rect 24800 -16858 24866 -16846
rect 24900 -16858 24966 -16846
rect 25000 -16846 25014 -16824
rect 25048 -16824 25104 -16812
rect 25048 -16846 25066 -16824
rect 25000 -16858 25066 -16846
rect 25100 -16846 25104 -16824
rect 25138 -16824 25194 -16812
rect 25138 -16846 25166 -16824
rect 25228 -16846 25287 -16812
rect 25100 -16858 25166 -16846
rect 25200 -16858 25287 -16846
rect 24593 -16902 25287 -16858
rect 24593 -16936 24654 -16902
rect 24688 -16924 24744 -16902
rect 24778 -16924 24834 -16902
rect 24868 -16924 24924 -16902
rect 24700 -16936 24744 -16924
rect 24800 -16936 24834 -16924
rect 24900 -16936 24924 -16924
rect 24958 -16924 25014 -16902
rect 24958 -16936 24966 -16924
rect 24593 -16958 24666 -16936
rect 24700 -16958 24766 -16936
rect 24800 -16958 24866 -16936
rect 24900 -16958 24966 -16936
rect 25000 -16936 25014 -16924
rect 25048 -16924 25104 -16902
rect 25048 -16936 25066 -16924
rect 25000 -16958 25066 -16936
rect 25100 -16936 25104 -16924
rect 25138 -16924 25194 -16902
rect 25138 -16936 25166 -16924
rect 25228 -16936 25287 -16902
rect 25100 -16958 25166 -16936
rect 25200 -16958 25287 -16936
rect 24593 -16992 25287 -16958
rect 24593 -17026 24654 -16992
rect 24688 -17024 24744 -16992
rect 24778 -17024 24834 -16992
rect 24868 -17024 24924 -16992
rect 24700 -17026 24744 -17024
rect 24800 -17026 24834 -17024
rect 24900 -17026 24924 -17024
rect 24958 -17024 25014 -16992
rect 24958 -17026 24966 -17024
rect 24593 -17058 24666 -17026
rect 24700 -17058 24766 -17026
rect 24800 -17058 24866 -17026
rect 24900 -17058 24966 -17026
rect 25000 -17026 25014 -17024
rect 25048 -17024 25104 -16992
rect 25048 -17026 25066 -17024
rect 25000 -17058 25066 -17026
rect 25100 -17026 25104 -17024
rect 25138 -17024 25194 -16992
rect 25138 -17026 25166 -17024
rect 25228 -17026 25287 -16992
rect 25100 -17058 25166 -17026
rect 25200 -17058 25287 -17026
rect 24593 -17082 25287 -17058
rect 24593 -17116 24654 -17082
rect 24688 -17116 24744 -17082
rect 24778 -17116 24834 -17082
rect 24868 -17116 24924 -17082
rect 24958 -17116 25014 -17082
rect 25048 -17116 25104 -17082
rect 25138 -17116 25194 -17082
rect 25228 -17116 25287 -17082
rect 24593 -17124 25287 -17116
rect 24593 -17158 24666 -17124
rect 24700 -17158 24766 -17124
rect 24800 -17158 24866 -17124
rect 24900 -17158 24966 -17124
rect 25000 -17158 25066 -17124
rect 25100 -17158 25166 -17124
rect 25200 -17158 25287 -17124
rect 24593 -17172 25287 -17158
rect 24593 -17206 24654 -17172
rect 24688 -17206 24744 -17172
rect 24778 -17206 24834 -17172
rect 24868 -17206 24924 -17172
rect 24958 -17206 25014 -17172
rect 25048 -17206 25104 -17172
rect 25138 -17206 25194 -17172
rect 25228 -17206 25287 -17172
rect 24593 -17224 25287 -17206
rect 24593 -17258 24666 -17224
rect 24700 -17258 24766 -17224
rect 24800 -17258 24866 -17224
rect 24900 -17258 24966 -17224
rect 25000 -17258 25066 -17224
rect 25100 -17258 25166 -17224
rect 25200 -17258 25287 -17224
rect 24593 -17262 25287 -17258
rect 24593 -17296 24654 -17262
rect 24688 -17296 24744 -17262
rect 24778 -17296 24834 -17262
rect 24868 -17296 24924 -17262
rect 24958 -17296 25014 -17262
rect 25048 -17296 25104 -17262
rect 25138 -17296 25194 -17262
rect 25228 -17296 25287 -17262
rect 24593 -17324 25287 -17296
rect 24593 -17352 24666 -17324
rect 24700 -17352 24766 -17324
rect 24800 -17352 24866 -17324
rect 24900 -17352 24966 -17324
rect 24593 -17386 24654 -17352
rect 24700 -17358 24744 -17352
rect 24800 -17358 24834 -17352
rect 24900 -17358 24924 -17352
rect 24688 -17386 24744 -17358
rect 24778 -17386 24834 -17358
rect 24868 -17386 24924 -17358
rect 24958 -17358 24966 -17352
rect 25000 -17352 25066 -17324
rect 25000 -17358 25014 -17352
rect 24958 -17386 25014 -17358
rect 25048 -17358 25066 -17352
rect 25100 -17352 25166 -17324
rect 25200 -17352 25287 -17324
rect 25100 -17358 25104 -17352
rect 25048 -17386 25104 -17358
rect 25138 -17358 25166 -17352
rect 25138 -17386 25194 -17358
rect 25228 -17386 25287 -17352
rect 24593 -17445 25287 -17386
rect 25349 -16782 25368 -16748
rect 25402 -16782 25421 -16748
rect 25349 -16838 25421 -16782
rect 25349 -16872 25368 -16838
rect 25402 -16872 25421 -16838
rect 25349 -16928 25421 -16872
rect 25349 -16962 25368 -16928
rect 25402 -16962 25421 -16928
rect 25349 -17018 25421 -16962
rect 25349 -17052 25368 -17018
rect 25402 -17052 25421 -17018
rect 25349 -17108 25421 -17052
rect 25349 -17142 25368 -17108
rect 25402 -17142 25421 -17108
rect 25349 -17198 25421 -17142
rect 25349 -17232 25368 -17198
rect 25402 -17232 25421 -17198
rect 25349 -17288 25421 -17232
rect 25349 -17322 25368 -17288
rect 25402 -17322 25421 -17288
rect 25349 -17378 25421 -17322
rect 25349 -17412 25368 -17378
rect 25402 -17412 25421 -17378
rect 24459 -17502 24531 -17468
rect 25349 -17468 25421 -17412
rect 25349 -17502 25368 -17468
rect 25402 -17502 25421 -17468
rect 25485 -16708 25515 -16702
rect 25549 -16708 25616 -16674
rect 25650 -16702 26803 -16674
rect 25650 -16708 25683 -16702
rect 25485 -16764 25683 -16708
rect 25485 -16798 25515 -16764
rect 25549 -16798 25616 -16764
rect 25650 -16798 25683 -16764
rect 25485 -16854 25683 -16798
rect 25485 -16888 25515 -16854
rect 25549 -16888 25616 -16854
rect 25650 -16888 25683 -16854
rect 25485 -16944 25683 -16888
rect 25485 -16978 25515 -16944
rect 25549 -16978 25616 -16944
rect 25650 -16978 25683 -16944
rect 25485 -17034 25683 -16978
rect 25485 -17068 25515 -17034
rect 25549 -17068 25616 -17034
rect 25650 -17068 25683 -17034
rect 25485 -17124 25683 -17068
rect 25485 -17158 25515 -17124
rect 25549 -17158 25616 -17124
rect 25650 -17158 25683 -17124
rect 25485 -17214 25683 -17158
rect 25485 -17248 25515 -17214
rect 25549 -17248 25616 -17214
rect 25650 -17248 25683 -17214
rect 25485 -17304 25683 -17248
rect 25485 -17338 25515 -17304
rect 25549 -17338 25616 -17304
rect 25650 -17338 25683 -17304
rect 25485 -17394 25683 -17338
rect 25485 -17428 25515 -17394
rect 25549 -17428 25616 -17394
rect 25650 -17428 25683 -17394
rect 25485 -17484 25683 -17428
rect 25485 -17502 25515 -17484
rect 24362 -17518 25515 -17502
rect 25549 -17518 25616 -17484
rect 25650 -17502 25683 -17484
rect 25747 -16714 25819 -16702
rect 25747 -16748 25766 -16714
rect 25800 -16748 25819 -16714
rect 25747 -16804 25819 -16748
rect 26637 -16748 26709 -16702
rect 25747 -16838 25766 -16804
rect 25800 -16838 25819 -16804
rect 25747 -16894 25819 -16838
rect 25747 -16928 25766 -16894
rect 25800 -16928 25819 -16894
rect 25747 -16984 25819 -16928
rect 25747 -17018 25766 -16984
rect 25800 -17018 25819 -16984
rect 25747 -17074 25819 -17018
rect 25747 -17108 25766 -17074
rect 25800 -17108 25819 -17074
rect 25747 -17164 25819 -17108
rect 25747 -17198 25766 -17164
rect 25800 -17198 25819 -17164
rect 25747 -17254 25819 -17198
rect 25747 -17288 25766 -17254
rect 25800 -17288 25819 -17254
rect 25747 -17344 25819 -17288
rect 25747 -17378 25766 -17344
rect 25800 -17378 25819 -17344
rect 25747 -17434 25819 -17378
rect 25747 -17468 25766 -17434
rect 25800 -17468 25819 -17434
rect 25881 -16811 26575 -16750
rect 25881 -16846 25942 -16811
rect 25976 -16823 26032 -16811
rect 26066 -16823 26122 -16811
rect 26156 -16823 26212 -16811
rect 25988 -16846 26032 -16823
rect 26088 -16846 26122 -16823
rect 26188 -16846 26212 -16823
rect 26246 -16823 26302 -16811
rect 26246 -16846 26254 -16823
rect 25881 -16858 25954 -16846
rect 25988 -16858 26054 -16846
rect 26088 -16858 26154 -16846
rect 26188 -16858 26254 -16846
rect 26288 -16846 26302 -16823
rect 26336 -16823 26392 -16811
rect 26336 -16846 26354 -16823
rect 26288 -16858 26354 -16846
rect 26388 -16846 26392 -16823
rect 26426 -16823 26482 -16811
rect 26426 -16846 26454 -16823
rect 26516 -16846 26575 -16811
rect 26388 -16858 26454 -16846
rect 26488 -16858 26575 -16846
rect 25881 -16901 26575 -16858
rect 25881 -16936 25942 -16901
rect 25976 -16923 26032 -16901
rect 26066 -16923 26122 -16901
rect 26156 -16923 26212 -16901
rect 25988 -16936 26032 -16923
rect 26088 -16936 26122 -16923
rect 26188 -16936 26212 -16923
rect 26246 -16923 26302 -16901
rect 26246 -16936 26254 -16923
rect 25881 -16958 25954 -16936
rect 25988 -16958 26054 -16936
rect 26088 -16958 26154 -16936
rect 26188 -16958 26254 -16936
rect 26288 -16936 26302 -16923
rect 26336 -16923 26392 -16901
rect 26336 -16936 26354 -16923
rect 26288 -16958 26354 -16936
rect 26388 -16936 26392 -16923
rect 26426 -16923 26482 -16901
rect 26426 -16936 26454 -16923
rect 26516 -16936 26575 -16901
rect 26388 -16958 26454 -16936
rect 26488 -16958 26575 -16936
rect 25881 -16991 26575 -16958
rect 25881 -17026 25942 -16991
rect 25976 -17023 26032 -16991
rect 26066 -17023 26122 -16991
rect 26156 -17023 26212 -16991
rect 25988 -17026 26032 -17023
rect 26088 -17026 26122 -17023
rect 26188 -17026 26212 -17023
rect 26246 -17023 26302 -16991
rect 26246 -17026 26254 -17023
rect 25881 -17058 25954 -17026
rect 25988 -17058 26054 -17026
rect 26088 -17058 26154 -17026
rect 26188 -17058 26254 -17026
rect 26288 -17026 26302 -17023
rect 26336 -17023 26392 -16991
rect 26336 -17026 26354 -17023
rect 26288 -17058 26354 -17026
rect 26388 -17026 26392 -17023
rect 26426 -17023 26482 -16991
rect 26426 -17026 26454 -17023
rect 26516 -17026 26575 -16991
rect 26388 -17058 26454 -17026
rect 26488 -17058 26575 -17026
rect 25881 -17081 26575 -17058
rect 25881 -17116 25942 -17081
rect 25976 -17116 26032 -17081
rect 26066 -17116 26122 -17081
rect 26156 -17116 26212 -17081
rect 26246 -17116 26302 -17081
rect 26336 -17116 26392 -17081
rect 26426 -17116 26482 -17081
rect 26516 -17116 26575 -17081
rect 25881 -17123 26575 -17116
rect 25881 -17158 25954 -17123
rect 25988 -17158 26054 -17123
rect 26088 -17158 26154 -17123
rect 26188 -17158 26254 -17123
rect 26288 -17158 26354 -17123
rect 26388 -17158 26454 -17123
rect 26488 -17158 26575 -17123
rect 25881 -17171 26575 -17158
rect 25881 -17206 25942 -17171
rect 25976 -17206 26032 -17171
rect 26066 -17206 26122 -17171
rect 26156 -17206 26212 -17171
rect 26246 -17206 26302 -17171
rect 26336 -17206 26392 -17171
rect 26426 -17206 26482 -17171
rect 26516 -17206 26575 -17171
rect 25881 -17223 26575 -17206
rect 25881 -17258 25954 -17223
rect 25988 -17258 26054 -17223
rect 26088 -17258 26154 -17223
rect 26188 -17258 26254 -17223
rect 26288 -17258 26354 -17223
rect 26388 -17258 26454 -17223
rect 26488 -17258 26575 -17223
rect 25881 -17261 26575 -17258
rect 25881 -17296 25942 -17261
rect 25976 -17296 26032 -17261
rect 26066 -17296 26122 -17261
rect 26156 -17296 26212 -17261
rect 26246 -17296 26302 -17261
rect 26336 -17296 26392 -17261
rect 26426 -17296 26482 -17261
rect 26516 -17296 26575 -17261
rect 25881 -17323 26575 -17296
rect 25881 -17351 25954 -17323
rect 25988 -17351 26054 -17323
rect 26088 -17351 26154 -17323
rect 26188 -17351 26254 -17323
rect 25881 -17386 25942 -17351
rect 25988 -17358 26032 -17351
rect 26088 -17358 26122 -17351
rect 26188 -17358 26212 -17351
rect 25976 -17386 26032 -17358
rect 26066 -17386 26122 -17358
rect 26156 -17386 26212 -17358
rect 26246 -17358 26254 -17351
rect 26288 -17351 26354 -17323
rect 26288 -17358 26302 -17351
rect 26246 -17386 26302 -17358
rect 26336 -17358 26354 -17351
rect 26388 -17351 26454 -17323
rect 26488 -17351 26575 -17323
rect 26388 -17358 26392 -17351
rect 26336 -17386 26392 -17358
rect 26426 -17358 26454 -17351
rect 26426 -17386 26482 -17358
rect 26516 -17386 26575 -17351
rect 25881 -17445 26575 -17386
rect 26637 -16782 26656 -16748
rect 26690 -16782 26709 -16748
rect 26637 -16838 26709 -16782
rect 26637 -16872 26656 -16838
rect 26690 -16872 26709 -16838
rect 26637 -16928 26709 -16872
rect 26637 -16962 26656 -16928
rect 26690 -16962 26709 -16928
rect 26637 -17018 26709 -16962
rect 26637 -17052 26656 -17018
rect 26690 -17052 26709 -17018
rect 26637 -17108 26709 -17052
rect 26637 -17142 26656 -17108
rect 26690 -17142 26709 -17108
rect 26637 -17198 26709 -17142
rect 26637 -17232 26656 -17198
rect 26690 -17232 26709 -17198
rect 26637 -17288 26709 -17232
rect 26637 -17322 26656 -17288
rect 26690 -17322 26709 -17288
rect 26637 -17378 26709 -17322
rect 26637 -17412 26656 -17378
rect 26690 -17412 26709 -17378
rect 25747 -17502 25819 -17468
rect 26637 -17468 26709 -17412
rect 26637 -17502 26656 -17468
rect 26690 -17502 26709 -17468
rect 26773 -16708 26803 -16702
rect 26837 -16702 26884 -16674
rect 26837 -16708 26872 -16702
rect 26773 -16764 26872 -16708
rect 26773 -16798 26803 -16764
rect 26837 -16798 26872 -16764
rect 26773 -16854 26872 -16798
rect 26773 -16888 26803 -16854
rect 26837 -16888 26872 -16854
rect 26773 -16944 26872 -16888
rect 26773 -16978 26803 -16944
rect 26837 -16978 26872 -16944
rect 26773 -17034 26872 -16978
rect 26773 -17068 26803 -17034
rect 26837 -17068 26872 -17034
rect 26773 -17124 26872 -17068
rect 26773 -17158 26803 -17124
rect 26837 -17158 26872 -17124
rect 26773 -17214 26872 -17158
rect 26773 -17248 26803 -17214
rect 26837 -17248 26872 -17214
rect 26773 -17304 26872 -17248
rect 26773 -17338 26803 -17304
rect 26837 -17338 26872 -17304
rect 26773 -17394 26872 -17338
rect 26773 -17428 26803 -17394
rect 26837 -17428 26872 -17394
rect 26773 -17484 26872 -17428
rect 26773 -17502 26803 -17484
rect 25650 -17518 26803 -17502
rect 26837 -17502 26872 -17484
rect 26837 -17518 26884 -17502
rect 16568 -17526 26884 -17518
rect 16568 -17560 16844 -17526
rect 16878 -17560 16934 -17526
rect 16968 -17560 17024 -17526
rect 17058 -17560 17114 -17526
rect 17148 -17560 17204 -17526
rect 17238 -17560 17294 -17526
rect 17328 -17560 17384 -17526
rect 17418 -17560 17474 -17526
rect 17508 -17560 17564 -17526
rect 17598 -17560 18132 -17526
rect 18166 -17560 18222 -17526
rect 18256 -17560 18312 -17526
rect 18346 -17560 18402 -17526
rect 18436 -17560 18492 -17526
rect 18526 -17560 18582 -17526
rect 18616 -17560 18672 -17526
rect 18706 -17560 18762 -17526
rect 18796 -17560 18852 -17526
rect 18886 -17560 19420 -17526
rect 19454 -17560 19510 -17526
rect 19544 -17560 19600 -17526
rect 19634 -17560 19690 -17526
rect 19724 -17560 19780 -17526
rect 19814 -17560 19870 -17526
rect 19904 -17560 19960 -17526
rect 19994 -17560 20050 -17526
rect 20084 -17560 20140 -17526
rect 20174 -17560 20708 -17526
rect 20742 -17560 20798 -17526
rect 20832 -17560 20888 -17526
rect 20922 -17560 20978 -17526
rect 21012 -17560 21068 -17526
rect 21102 -17560 21158 -17526
rect 21192 -17560 21248 -17526
rect 21282 -17560 21338 -17526
rect 21372 -17560 21428 -17526
rect 21462 -17560 21996 -17526
rect 22030 -17560 22086 -17526
rect 22120 -17560 22176 -17526
rect 22210 -17560 22266 -17526
rect 22300 -17560 22356 -17526
rect 22390 -17560 22446 -17526
rect 22480 -17560 22536 -17526
rect 22570 -17560 22626 -17526
rect 22660 -17560 22716 -17526
rect 22750 -17560 23284 -17526
rect 23318 -17560 23374 -17526
rect 23408 -17560 23464 -17526
rect 23498 -17560 23554 -17526
rect 23588 -17560 23644 -17526
rect 23678 -17560 23734 -17526
rect 23768 -17560 23824 -17526
rect 23858 -17560 23914 -17526
rect 23948 -17560 24004 -17526
rect 24038 -17560 24572 -17526
rect 24606 -17560 24662 -17526
rect 24696 -17560 24752 -17526
rect 24786 -17560 24842 -17526
rect 24876 -17560 24932 -17526
rect 24966 -17560 25022 -17526
rect 25056 -17560 25112 -17526
rect 25146 -17560 25202 -17526
rect 25236 -17560 25292 -17526
rect 25326 -17560 25860 -17526
rect 25894 -17560 25950 -17526
rect 25984 -17560 26040 -17526
rect 26074 -17560 26130 -17526
rect 26164 -17560 26220 -17526
rect 26254 -17560 26310 -17526
rect 26344 -17560 26400 -17526
rect 26434 -17560 26490 -17526
rect 26524 -17560 26580 -17526
rect 26614 -17560 26884 -17526
rect 16568 -17574 26884 -17560
rect 16568 -17608 16600 -17574
rect 16634 -17608 17787 -17574
rect 17821 -17608 17888 -17574
rect 17922 -17608 19075 -17574
rect 19109 -17608 19176 -17574
rect 19210 -17608 20363 -17574
rect 20397 -17608 20464 -17574
rect 20498 -17608 21651 -17574
rect 21685 -17608 21752 -17574
rect 21786 -17608 22939 -17574
rect 22973 -17608 23040 -17574
rect 23074 -17608 24227 -17574
rect 24261 -17608 24328 -17574
rect 24362 -17608 25515 -17574
rect 25549 -17608 25616 -17574
rect 25650 -17608 26803 -17574
rect 26837 -17608 26884 -17574
rect 16568 -17675 26884 -17608
rect 16568 -17709 16684 -17675
rect 16718 -17709 16774 -17675
rect 16808 -17709 16864 -17675
rect 16898 -17709 16954 -17675
rect 16988 -17709 17044 -17675
rect 17078 -17709 17134 -17675
rect 17168 -17709 17224 -17675
rect 17258 -17709 17314 -17675
rect 17348 -17709 17404 -17675
rect 17438 -17709 17494 -17675
rect 17528 -17709 17584 -17675
rect 17618 -17709 17674 -17675
rect 17708 -17709 17764 -17675
rect 17798 -17709 17972 -17675
rect 18006 -17709 18062 -17675
rect 18096 -17709 18152 -17675
rect 18186 -17709 18242 -17675
rect 18276 -17709 18332 -17675
rect 18366 -17709 18422 -17675
rect 18456 -17709 18512 -17675
rect 18546 -17709 18602 -17675
rect 18636 -17709 18692 -17675
rect 18726 -17709 18782 -17675
rect 18816 -17709 18872 -17675
rect 18906 -17709 18962 -17675
rect 18996 -17709 19052 -17675
rect 19086 -17709 19260 -17675
rect 19294 -17709 19350 -17675
rect 19384 -17709 19440 -17675
rect 19474 -17709 19530 -17675
rect 19564 -17709 19620 -17675
rect 19654 -17709 19710 -17675
rect 19744 -17709 19800 -17675
rect 19834 -17709 19890 -17675
rect 19924 -17709 19980 -17675
rect 20014 -17709 20070 -17675
rect 20104 -17709 20160 -17675
rect 20194 -17709 20250 -17675
rect 20284 -17709 20340 -17675
rect 20374 -17709 20548 -17675
rect 20582 -17709 20638 -17675
rect 20672 -17709 20728 -17675
rect 20762 -17709 20818 -17675
rect 20852 -17709 20908 -17675
rect 20942 -17709 20998 -17675
rect 21032 -17709 21088 -17675
rect 21122 -17709 21178 -17675
rect 21212 -17709 21268 -17675
rect 21302 -17709 21358 -17675
rect 21392 -17709 21448 -17675
rect 21482 -17709 21538 -17675
rect 21572 -17709 21628 -17675
rect 21662 -17709 21836 -17675
rect 21870 -17709 21926 -17675
rect 21960 -17709 22016 -17675
rect 22050 -17709 22106 -17675
rect 22140 -17709 22196 -17675
rect 22230 -17709 22286 -17675
rect 22320 -17709 22376 -17675
rect 22410 -17709 22466 -17675
rect 22500 -17709 22556 -17675
rect 22590 -17709 22646 -17675
rect 22680 -17709 22736 -17675
rect 22770 -17709 22826 -17675
rect 22860 -17709 22916 -17675
rect 22950 -17709 23124 -17675
rect 23158 -17709 23214 -17675
rect 23248 -17709 23304 -17675
rect 23338 -17709 23394 -17675
rect 23428 -17709 23484 -17675
rect 23518 -17709 23574 -17675
rect 23608 -17709 23664 -17675
rect 23698 -17709 23754 -17675
rect 23788 -17709 23844 -17675
rect 23878 -17709 23934 -17675
rect 23968 -17709 24024 -17675
rect 24058 -17709 24114 -17675
rect 24148 -17709 24204 -17675
rect 24238 -17709 24412 -17675
rect 24446 -17709 24502 -17675
rect 24536 -17709 24592 -17675
rect 24626 -17709 24682 -17675
rect 24716 -17709 24772 -17675
rect 24806 -17709 24862 -17675
rect 24896 -17709 24952 -17675
rect 24986 -17709 25042 -17675
rect 25076 -17709 25132 -17675
rect 25166 -17709 25222 -17675
rect 25256 -17709 25312 -17675
rect 25346 -17709 25402 -17675
rect 25436 -17709 25492 -17675
rect 25526 -17709 25700 -17675
rect 25734 -17709 25790 -17675
rect 25824 -17709 25880 -17675
rect 25914 -17709 25970 -17675
rect 26004 -17709 26060 -17675
rect 26094 -17709 26150 -17675
rect 26184 -17709 26240 -17675
rect 26274 -17709 26330 -17675
rect 26364 -17709 26420 -17675
rect 26454 -17709 26510 -17675
rect 26544 -17709 26600 -17675
rect 26634 -17709 26690 -17675
rect 26724 -17709 26780 -17675
rect 26814 -17702 26884 -17675
rect 26814 -17709 26872 -17702
rect 16568 -17742 26872 -17709
rect 6808 -30938 6870 -30368
rect 6808 -31152 7302 -30938
rect 13606 -31152 14038 -30938
rect 6808 -31168 14038 -31152
rect 6808 -31738 7302 -31168
rect 13606 -31738 14038 -31168
rect 6808 -31754 14038 -31738
rect 6808 -32822 7302 -31754
rect 7240 -33392 7302 -32822
rect 11540 -32822 12070 -31754
rect 13606 -31762 14038 -31754
rect 11972 -33392 12070 -32822
rect 11540 -33508 12070 -33392
rect 11540 -35276 12070 -35170
rect 11972 -35846 12070 -35276
rect 6808 -36116 7240 -35846
rect 11544 -36112 12070 -35846
rect 12692 -36112 13200 -36102
rect 7286 -36116 13622 -36112
rect 6808 -36128 13622 -36116
rect 6808 -36698 7302 -36128
rect 13606 -36698 13622 -36128
rect 6808 -36714 13622 -36698
rect 6808 -36720 7798 -36714
rect 8194 -36912 8636 -36714
rect 8626 -37482 8636 -36912
rect 11950 -36912 12382 -36714
rect 8194 -37730 8636 -37482
rect 8626 -38300 8636 -37730
rect 8194 -38548 8636 -38300
rect 12692 -38548 13200 -36714
rect 8626 -39118 8636 -38548
rect 12382 -39118 13200 -38548
rect 8194 -39356 8636 -39118
rect 12696 -39356 13200 -39118
rect 7286 -39372 13622 -39356
rect 7286 -39942 7302 -39372
rect 13606 -39942 13622 -39372
rect 7286 -39958 13622 -39942
rect 8194 -39968 8636 -39958
rect 12696 -39962 13200 -39958
<< viali >>
rect 16938 -11694 16960 -11672
rect 16960 -11694 16972 -11672
rect 17038 -11694 17050 -11672
rect 17050 -11694 17072 -11672
rect 17138 -11694 17140 -11672
rect 17140 -11694 17172 -11672
rect 16938 -11706 16972 -11694
rect 17038 -11706 17072 -11694
rect 17138 -11706 17172 -11694
rect 17238 -11706 17272 -11672
rect 17338 -11706 17372 -11672
rect 17438 -11694 17466 -11672
rect 17466 -11694 17472 -11672
rect 17438 -11706 17472 -11694
rect 16938 -11784 16960 -11772
rect 16960 -11784 16972 -11772
rect 17038 -11784 17050 -11772
rect 17050 -11784 17072 -11772
rect 17138 -11784 17140 -11772
rect 17140 -11784 17172 -11772
rect 16938 -11806 16972 -11784
rect 17038 -11806 17072 -11784
rect 17138 -11806 17172 -11784
rect 17238 -11806 17272 -11772
rect 17338 -11806 17372 -11772
rect 17438 -11784 17466 -11772
rect 17466 -11784 17472 -11772
rect 17438 -11806 17472 -11784
rect 16938 -11874 16960 -11872
rect 16960 -11874 16972 -11872
rect 17038 -11874 17050 -11872
rect 17050 -11874 17072 -11872
rect 17138 -11874 17140 -11872
rect 17140 -11874 17172 -11872
rect 16938 -11906 16972 -11874
rect 17038 -11906 17072 -11874
rect 17138 -11906 17172 -11874
rect 17238 -11906 17272 -11872
rect 17338 -11906 17372 -11872
rect 17438 -11874 17466 -11872
rect 17466 -11874 17472 -11872
rect 17438 -11906 17472 -11874
rect 16938 -12006 16972 -11972
rect 17038 -12006 17072 -11972
rect 17138 -12006 17172 -11972
rect 17238 -12006 17272 -11972
rect 17338 -12006 17372 -11972
rect 17438 -12006 17472 -11972
rect 16938 -12106 16972 -12072
rect 17038 -12106 17072 -12072
rect 17138 -12106 17172 -12072
rect 17238 -12106 17272 -12072
rect 17338 -12106 17372 -12072
rect 17438 -12106 17472 -12072
rect 16938 -12200 16972 -12172
rect 17038 -12200 17072 -12172
rect 17138 -12200 17172 -12172
rect 16938 -12206 16960 -12200
rect 16960 -12206 16972 -12200
rect 17038 -12206 17050 -12200
rect 17050 -12206 17072 -12200
rect 17138 -12206 17140 -12200
rect 17140 -12206 17172 -12200
rect 17238 -12206 17272 -12172
rect 17338 -12206 17372 -12172
rect 17438 -12200 17472 -12172
rect 17438 -12206 17466 -12200
rect 17466 -12206 17472 -12200
rect 18226 -11694 18248 -11672
rect 18248 -11694 18260 -11672
rect 18326 -11694 18338 -11672
rect 18338 -11694 18360 -11672
rect 18426 -11694 18428 -11672
rect 18428 -11694 18460 -11672
rect 18226 -11706 18260 -11694
rect 18326 -11706 18360 -11694
rect 18426 -11706 18460 -11694
rect 18526 -11706 18560 -11672
rect 18626 -11706 18660 -11672
rect 18726 -11694 18754 -11672
rect 18754 -11694 18760 -11672
rect 18726 -11706 18760 -11694
rect 18226 -11784 18248 -11772
rect 18248 -11784 18260 -11772
rect 18326 -11784 18338 -11772
rect 18338 -11784 18360 -11772
rect 18426 -11784 18428 -11772
rect 18428 -11784 18460 -11772
rect 18226 -11806 18260 -11784
rect 18326 -11806 18360 -11784
rect 18426 -11806 18460 -11784
rect 18526 -11806 18560 -11772
rect 18626 -11806 18660 -11772
rect 18726 -11784 18754 -11772
rect 18754 -11784 18760 -11772
rect 18726 -11806 18760 -11784
rect 18226 -11874 18248 -11872
rect 18248 -11874 18260 -11872
rect 18326 -11874 18338 -11872
rect 18338 -11874 18360 -11872
rect 18426 -11874 18428 -11872
rect 18428 -11874 18460 -11872
rect 18226 -11906 18260 -11874
rect 18326 -11906 18360 -11874
rect 18426 -11906 18460 -11874
rect 18526 -11906 18560 -11872
rect 18626 -11906 18660 -11872
rect 18726 -11874 18754 -11872
rect 18754 -11874 18760 -11872
rect 18726 -11906 18760 -11874
rect 18226 -12006 18260 -11972
rect 18326 -12006 18360 -11972
rect 18426 -12006 18460 -11972
rect 18526 -12006 18560 -11972
rect 18626 -12006 18660 -11972
rect 18726 -12006 18760 -11972
rect 18226 -12106 18260 -12072
rect 18326 -12106 18360 -12072
rect 18426 -12106 18460 -12072
rect 18526 -12106 18560 -12072
rect 18626 -12106 18660 -12072
rect 18726 -12106 18760 -12072
rect 18226 -12200 18260 -12172
rect 18326 -12200 18360 -12172
rect 18426 -12200 18460 -12172
rect 18226 -12206 18248 -12200
rect 18248 -12206 18260 -12200
rect 18326 -12206 18338 -12200
rect 18338 -12206 18360 -12200
rect 18426 -12206 18428 -12200
rect 18428 -12206 18460 -12200
rect 18526 -12206 18560 -12172
rect 18626 -12206 18660 -12172
rect 18726 -12200 18760 -12172
rect 18726 -12206 18754 -12200
rect 18754 -12206 18760 -12200
rect 19514 -11694 19536 -11672
rect 19536 -11694 19548 -11672
rect 19614 -11694 19626 -11672
rect 19626 -11694 19648 -11672
rect 19714 -11694 19716 -11672
rect 19716 -11694 19748 -11672
rect 19514 -11706 19548 -11694
rect 19614 -11706 19648 -11694
rect 19714 -11706 19748 -11694
rect 19814 -11706 19848 -11672
rect 19914 -11706 19948 -11672
rect 20014 -11694 20042 -11672
rect 20042 -11694 20048 -11672
rect 20014 -11706 20048 -11694
rect 19514 -11784 19536 -11772
rect 19536 -11784 19548 -11772
rect 19614 -11784 19626 -11772
rect 19626 -11784 19648 -11772
rect 19714 -11784 19716 -11772
rect 19716 -11784 19748 -11772
rect 19514 -11806 19548 -11784
rect 19614 -11806 19648 -11784
rect 19714 -11806 19748 -11784
rect 19814 -11806 19848 -11772
rect 19914 -11806 19948 -11772
rect 20014 -11784 20042 -11772
rect 20042 -11784 20048 -11772
rect 20014 -11806 20048 -11784
rect 19514 -11874 19536 -11872
rect 19536 -11874 19548 -11872
rect 19614 -11874 19626 -11872
rect 19626 -11874 19648 -11872
rect 19714 -11874 19716 -11872
rect 19716 -11874 19748 -11872
rect 19514 -11906 19548 -11874
rect 19614 -11906 19648 -11874
rect 19714 -11906 19748 -11874
rect 19814 -11906 19848 -11872
rect 19914 -11906 19948 -11872
rect 20014 -11874 20042 -11872
rect 20042 -11874 20048 -11872
rect 20014 -11906 20048 -11874
rect 19514 -12006 19548 -11972
rect 19614 -12006 19648 -11972
rect 19714 -12006 19748 -11972
rect 19814 -12006 19848 -11972
rect 19914 -12006 19948 -11972
rect 20014 -12006 20048 -11972
rect 19514 -12106 19548 -12072
rect 19614 -12106 19648 -12072
rect 19714 -12106 19748 -12072
rect 19814 -12106 19848 -12072
rect 19914 -12106 19948 -12072
rect 20014 -12106 20048 -12072
rect 19514 -12200 19548 -12172
rect 19614 -12200 19648 -12172
rect 19714 -12200 19748 -12172
rect 19514 -12206 19536 -12200
rect 19536 -12206 19548 -12200
rect 19614 -12206 19626 -12200
rect 19626 -12206 19648 -12200
rect 19714 -12206 19716 -12200
rect 19716 -12206 19748 -12200
rect 19814 -12206 19848 -12172
rect 19914 -12206 19948 -12172
rect 20014 -12200 20048 -12172
rect 20014 -12206 20042 -12200
rect 20042 -12206 20048 -12200
rect 20802 -11694 20824 -11672
rect 20824 -11694 20836 -11672
rect 20902 -11694 20914 -11672
rect 20914 -11694 20936 -11672
rect 21002 -11694 21004 -11672
rect 21004 -11694 21036 -11672
rect 20802 -11706 20836 -11694
rect 20902 -11706 20936 -11694
rect 21002 -11706 21036 -11694
rect 21102 -11706 21136 -11672
rect 21202 -11706 21236 -11672
rect 21302 -11694 21330 -11672
rect 21330 -11694 21336 -11672
rect 21302 -11706 21336 -11694
rect 20802 -11784 20824 -11772
rect 20824 -11784 20836 -11772
rect 20902 -11784 20914 -11772
rect 20914 -11784 20936 -11772
rect 21002 -11784 21004 -11772
rect 21004 -11784 21036 -11772
rect 20802 -11806 20836 -11784
rect 20902 -11806 20936 -11784
rect 21002 -11806 21036 -11784
rect 21102 -11806 21136 -11772
rect 21202 -11806 21236 -11772
rect 21302 -11784 21330 -11772
rect 21330 -11784 21336 -11772
rect 21302 -11806 21336 -11784
rect 20802 -11874 20824 -11872
rect 20824 -11874 20836 -11872
rect 20902 -11874 20914 -11872
rect 20914 -11874 20936 -11872
rect 21002 -11874 21004 -11872
rect 21004 -11874 21036 -11872
rect 20802 -11906 20836 -11874
rect 20902 -11906 20936 -11874
rect 21002 -11906 21036 -11874
rect 21102 -11906 21136 -11872
rect 21202 -11906 21236 -11872
rect 21302 -11874 21330 -11872
rect 21330 -11874 21336 -11872
rect 21302 -11906 21336 -11874
rect 20802 -12006 20836 -11972
rect 20902 -12006 20936 -11972
rect 21002 -12006 21036 -11972
rect 21102 -12006 21136 -11972
rect 21202 -12006 21236 -11972
rect 21302 -12006 21336 -11972
rect 20802 -12106 20836 -12072
rect 20902 -12106 20936 -12072
rect 21002 -12106 21036 -12072
rect 21102 -12106 21136 -12072
rect 21202 -12106 21236 -12072
rect 21302 -12106 21336 -12072
rect 20802 -12200 20836 -12172
rect 20902 -12200 20936 -12172
rect 21002 -12200 21036 -12172
rect 20802 -12206 20824 -12200
rect 20824 -12206 20836 -12200
rect 20902 -12206 20914 -12200
rect 20914 -12206 20936 -12200
rect 21002 -12206 21004 -12200
rect 21004 -12206 21036 -12200
rect 21102 -12206 21136 -12172
rect 21202 -12206 21236 -12172
rect 21302 -12200 21336 -12172
rect 21302 -12206 21330 -12200
rect 21330 -12206 21336 -12200
rect 22090 -11694 22112 -11672
rect 22112 -11694 22124 -11672
rect 22190 -11694 22202 -11672
rect 22202 -11694 22224 -11672
rect 22290 -11694 22292 -11672
rect 22292 -11694 22324 -11672
rect 22090 -11706 22124 -11694
rect 22190 -11706 22224 -11694
rect 22290 -11706 22324 -11694
rect 22390 -11706 22424 -11672
rect 22490 -11706 22524 -11672
rect 22590 -11694 22618 -11672
rect 22618 -11694 22624 -11672
rect 22590 -11706 22624 -11694
rect 22090 -11784 22112 -11772
rect 22112 -11784 22124 -11772
rect 22190 -11784 22202 -11772
rect 22202 -11784 22224 -11772
rect 22290 -11784 22292 -11772
rect 22292 -11784 22324 -11772
rect 22090 -11806 22124 -11784
rect 22190 -11806 22224 -11784
rect 22290 -11806 22324 -11784
rect 22390 -11806 22424 -11772
rect 22490 -11806 22524 -11772
rect 22590 -11784 22618 -11772
rect 22618 -11784 22624 -11772
rect 22590 -11806 22624 -11784
rect 22090 -11874 22112 -11872
rect 22112 -11874 22124 -11872
rect 22190 -11874 22202 -11872
rect 22202 -11874 22224 -11872
rect 22290 -11874 22292 -11872
rect 22292 -11874 22324 -11872
rect 22090 -11906 22124 -11874
rect 22190 -11906 22224 -11874
rect 22290 -11906 22324 -11874
rect 22390 -11906 22424 -11872
rect 22490 -11906 22524 -11872
rect 22590 -11874 22618 -11872
rect 22618 -11874 22624 -11872
rect 22590 -11906 22624 -11874
rect 22090 -12006 22124 -11972
rect 22190 -12006 22224 -11972
rect 22290 -12006 22324 -11972
rect 22390 -12006 22424 -11972
rect 22490 -12006 22524 -11972
rect 22590 -12006 22624 -11972
rect 22090 -12106 22124 -12072
rect 22190 -12106 22224 -12072
rect 22290 -12106 22324 -12072
rect 22390 -12106 22424 -12072
rect 22490 -12106 22524 -12072
rect 22590 -12106 22624 -12072
rect 22090 -12200 22124 -12172
rect 22190 -12200 22224 -12172
rect 22290 -12200 22324 -12172
rect 22090 -12206 22112 -12200
rect 22112 -12206 22124 -12200
rect 22190 -12206 22202 -12200
rect 22202 -12206 22224 -12200
rect 22290 -12206 22292 -12200
rect 22292 -12206 22324 -12200
rect 22390 -12206 22424 -12172
rect 22490 -12206 22524 -12172
rect 22590 -12200 22624 -12172
rect 22590 -12206 22618 -12200
rect 22618 -12206 22624 -12200
rect 23378 -11694 23400 -11672
rect 23400 -11694 23412 -11672
rect 23478 -11694 23490 -11672
rect 23490 -11694 23512 -11672
rect 23578 -11694 23580 -11672
rect 23580 -11694 23612 -11672
rect 23378 -11706 23412 -11694
rect 23478 -11706 23512 -11694
rect 23578 -11706 23612 -11694
rect 23678 -11706 23712 -11672
rect 23778 -11706 23812 -11672
rect 23878 -11694 23906 -11672
rect 23906 -11694 23912 -11672
rect 23878 -11706 23912 -11694
rect 23378 -11784 23400 -11772
rect 23400 -11784 23412 -11772
rect 23478 -11784 23490 -11772
rect 23490 -11784 23512 -11772
rect 23578 -11784 23580 -11772
rect 23580 -11784 23612 -11772
rect 23378 -11806 23412 -11784
rect 23478 -11806 23512 -11784
rect 23578 -11806 23612 -11784
rect 23678 -11806 23712 -11772
rect 23778 -11806 23812 -11772
rect 23878 -11784 23906 -11772
rect 23906 -11784 23912 -11772
rect 23878 -11806 23912 -11784
rect 23378 -11874 23400 -11872
rect 23400 -11874 23412 -11872
rect 23478 -11874 23490 -11872
rect 23490 -11874 23512 -11872
rect 23578 -11874 23580 -11872
rect 23580 -11874 23612 -11872
rect 23378 -11906 23412 -11874
rect 23478 -11906 23512 -11874
rect 23578 -11906 23612 -11874
rect 23678 -11906 23712 -11872
rect 23778 -11906 23812 -11872
rect 23878 -11874 23906 -11872
rect 23906 -11874 23912 -11872
rect 23878 -11906 23912 -11874
rect 23378 -12006 23412 -11972
rect 23478 -12006 23512 -11972
rect 23578 -12006 23612 -11972
rect 23678 -12006 23712 -11972
rect 23778 -12006 23812 -11972
rect 23878 -12006 23912 -11972
rect 23378 -12106 23412 -12072
rect 23478 -12106 23512 -12072
rect 23578 -12106 23612 -12072
rect 23678 -12106 23712 -12072
rect 23778 -12106 23812 -12072
rect 23878 -12106 23912 -12072
rect 23378 -12200 23412 -12172
rect 23478 -12200 23512 -12172
rect 23578 -12200 23612 -12172
rect 23378 -12206 23400 -12200
rect 23400 -12206 23412 -12200
rect 23478 -12206 23490 -12200
rect 23490 -12206 23512 -12200
rect 23578 -12206 23580 -12200
rect 23580 -12206 23612 -12200
rect 23678 -12206 23712 -12172
rect 23778 -12206 23812 -12172
rect 23878 -12200 23912 -12172
rect 23878 -12206 23906 -12200
rect 23906 -12206 23912 -12200
rect 24666 -11694 24688 -11672
rect 24688 -11694 24700 -11672
rect 24766 -11694 24778 -11672
rect 24778 -11694 24800 -11672
rect 24866 -11694 24868 -11672
rect 24868 -11694 24900 -11672
rect 24666 -11706 24700 -11694
rect 24766 -11706 24800 -11694
rect 24866 -11706 24900 -11694
rect 24966 -11706 25000 -11672
rect 25066 -11706 25100 -11672
rect 25166 -11694 25194 -11672
rect 25194 -11694 25200 -11672
rect 25166 -11706 25200 -11694
rect 24666 -11784 24688 -11772
rect 24688 -11784 24700 -11772
rect 24766 -11784 24778 -11772
rect 24778 -11784 24800 -11772
rect 24866 -11784 24868 -11772
rect 24868 -11784 24900 -11772
rect 24666 -11806 24700 -11784
rect 24766 -11806 24800 -11784
rect 24866 -11806 24900 -11784
rect 24966 -11806 25000 -11772
rect 25066 -11806 25100 -11772
rect 25166 -11784 25194 -11772
rect 25194 -11784 25200 -11772
rect 25166 -11806 25200 -11784
rect 24666 -11874 24688 -11872
rect 24688 -11874 24700 -11872
rect 24766 -11874 24778 -11872
rect 24778 -11874 24800 -11872
rect 24866 -11874 24868 -11872
rect 24868 -11874 24900 -11872
rect 24666 -11906 24700 -11874
rect 24766 -11906 24800 -11874
rect 24866 -11906 24900 -11874
rect 24966 -11906 25000 -11872
rect 25066 -11906 25100 -11872
rect 25166 -11874 25194 -11872
rect 25194 -11874 25200 -11872
rect 25166 -11906 25200 -11874
rect 24666 -12006 24700 -11972
rect 24766 -12006 24800 -11972
rect 24866 -12006 24900 -11972
rect 24966 -12006 25000 -11972
rect 25066 -12006 25100 -11972
rect 25166 -12006 25200 -11972
rect 24666 -12106 24700 -12072
rect 24766 -12106 24800 -12072
rect 24866 -12106 24900 -12072
rect 24966 -12106 25000 -12072
rect 25066 -12106 25100 -12072
rect 25166 -12106 25200 -12072
rect 24666 -12200 24700 -12172
rect 24766 -12200 24800 -12172
rect 24866 -12200 24900 -12172
rect 24666 -12206 24688 -12200
rect 24688 -12206 24700 -12200
rect 24766 -12206 24778 -12200
rect 24778 -12206 24800 -12200
rect 24866 -12206 24868 -12200
rect 24868 -12206 24900 -12200
rect 24966 -12206 25000 -12172
rect 25066 -12206 25100 -12172
rect 25166 -12200 25200 -12172
rect 25166 -12206 25194 -12200
rect 25194 -12206 25200 -12200
rect 25954 -11694 25976 -11672
rect 25976 -11694 25988 -11672
rect 26054 -11694 26066 -11672
rect 26066 -11694 26088 -11672
rect 26154 -11694 26156 -11672
rect 26156 -11694 26188 -11672
rect 25954 -11706 25988 -11694
rect 26054 -11706 26088 -11694
rect 26154 -11706 26188 -11694
rect 26254 -11706 26288 -11672
rect 26354 -11706 26388 -11672
rect 26454 -11694 26482 -11672
rect 26482 -11694 26488 -11672
rect 26454 -11706 26488 -11694
rect 25954 -11784 25976 -11772
rect 25976 -11784 25988 -11772
rect 26054 -11784 26066 -11772
rect 26066 -11784 26088 -11772
rect 26154 -11784 26156 -11772
rect 26156 -11784 26188 -11772
rect 25954 -11806 25988 -11784
rect 26054 -11806 26088 -11784
rect 26154 -11806 26188 -11784
rect 26254 -11806 26288 -11772
rect 26354 -11806 26388 -11772
rect 26454 -11784 26482 -11772
rect 26482 -11784 26488 -11772
rect 26454 -11806 26488 -11784
rect 25954 -11874 25976 -11872
rect 25976 -11874 25988 -11872
rect 26054 -11874 26066 -11872
rect 26066 -11874 26088 -11872
rect 26154 -11874 26156 -11872
rect 26156 -11874 26188 -11872
rect 25954 -11906 25988 -11874
rect 26054 -11906 26088 -11874
rect 26154 -11906 26188 -11874
rect 26254 -11906 26288 -11872
rect 26354 -11906 26388 -11872
rect 26454 -11874 26482 -11872
rect 26482 -11874 26488 -11872
rect 26454 -11906 26488 -11874
rect 25954 -12006 25988 -11972
rect 26054 -12006 26088 -11972
rect 26154 -12006 26188 -11972
rect 26254 -12006 26288 -11972
rect 26354 -12006 26388 -11972
rect 26454 -12006 26488 -11972
rect 25954 -12106 25988 -12072
rect 26054 -12106 26088 -12072
rect 26154 -12106 26188 -12072
rect 26254 -12106 26288 -12072
rect 26354 -12106 26388 -12072
rect 26454 -12106 26488 -12072
rect 25954 -12200 25988 -12172
rect 26054 -12200 26088 -12172
rect 26154 -12200 26188 -12172
rect 25954 -12206 25976 -12200
rect 25976 -12206 25988 -12200
rect 26054 -12206 26066 -12200
rect 26066 -12206 26088 -12200
rect 26154 -12206 26156 -12200
rect 26156 -12206 26188 -12200
rect 26254 -12206 26288 -12172
rect 26354 -12206 26388 -12172
rect 26454 -12200 26488 -12172
rect 26454 -12206 26482 -12200
rect 26482 -12206 26488 -12200
rect 16938 -12982 16960 -12960
rect 16960 -12982 16972 -12960
rect 17038 -12982 17050 -12960
rect 17050 -12982 17072 -12960
rect 17138 -12982 17140 -12960
rect 17140 -12982 17172 -12960
rect 16938 -12994 16972 -12982
rect 17038 -12994 17072 -12982
rect 17138 -12994 17172 -12982
rect 17238 -12994 17272 -12960
rect 17338 -12994 17372 -12960
rect 17438 -12982 17466 -12960
rect 17466 -12982 17472 -12960
rect 17438 -12994 17472 -12982
rect 16938 -13072 16960 -13060
rect 16960 -13072 16972 -13060
rect 17038 -13072 17050 -13060
rect 17050 -13072 17072 -13060
rect 17138 -13072 17140 -13060
rect 17140 -13072 17172 -13060
rect 16938 -13094 16972 -13072
rect 17038 -13094 17072 -13072
rect 17138 -13094 17172 -13072
rect 17238 -13094 17272 -13060
rect 17338 -13094 17372 -13060
rect 17438 -13072 17466 -13060
rect 17466 -13072 17472 -13060
rect 17438 -13094 17472 -13072
rect 16938 -13162 16960 -13160
rect 16960 -13162 16972 -13160
rect 17038 -13162 17050 -13160
rect 17050 -13162 17072 -13160
rect 17138 -13162 17140 -13160
rect 17140 -13162 17172 -13160
rect 16938 -13194 16972 -13162
rect 17038 -13194 17072 -13162
rect 17138 -13194 17172 -13162
rect 17238 -13194 17272 -13160
rect 17338 -13194 17372 -13160
rect 17438 -13162 17466 -13160
rect 17466 -13162 17472 -13160
rect 17438 -13194 17472 -13162
rect 16938 -13294 16972 -13260
rect 17038 -13294 17072 -13260
rect 17138 -13294 17172 -13260
rect 17238 -13294 17272 -13260
rect 17338 -13294 17372 -13260
rect 17438 -13294 17472 -13260
rect 16938 -13394 16972 -13360
rect 17038 -13394 17072 -13360
rect 17138 -13394 17172 -13360
rect 17238 -13394 17272 -13360
rect 17338 -13394 17372 -13360
rect 17438 -13394 17472 -13360
rect 16938 -13488 16972 -13460
rect 17038 -13488 17072 -13460
rect 17138 -13488 17172 -13460
rect 16938 -13494 16960 -13488
rect 16960 -13494 16972 -13488
rect 17038 -13494 17050 -13488
rect 17050 -13494 17072 -13488
rect 17138 -13494 17140 -13488
rect 17140 -13494 17172 -13488
rect 17238 -13494 17272 -13460
rect 17338 -13494 17372 -13460
rect 17438 -13488 17472 -13460
rect 17438 -13494 17466 -13488
rect 17466 -13494 17472 -13488
rect 18226 -12982 18248 -12960
rect 18248 -12982 18260 -12960
rect 18326 -12982 18338 -12960
rect 18338 -12982 18360 -12960
rect 18426 -12982 18428 -12960
rect 18428 -12982 18460 -12960
rect 18226 -12994 18260 -12982
rect 18326 -12994 18360 -12982
rect 18426 -12994 18460 -12982
rect 18526 -12994 18560 -12960
rect 18626 -12994 18660 -12960
rect 18726 -12982 18754 -12960
rect 18754 -12982 18760 -12960
rect 18726 -12994 18760 -12982
rect 18226 -13072 18248 -13060
rect 18248 -13072 18260 -13060
rect 18326 -13072 18338 -13060
rect 18338 -13072 18360 -13060
rect 18426 -13072 18428 -13060
rect 18428 -13072 18460 -13060
rect 18226 -13094 18260 -13072
rect 18326 -13094 18360 -13072
rect 18426 -13094 18460 -13072
rect 18526 -13094 18560 -13060
rect 18626 -13094 18660 -13060
rect 18726 -13072 18754 -13060
rect 18754 -13072 18760 -13060
rect 18726 -13094 18760 -13072
rect 18226 -13162 18248 -13160
rect 18248 -13162 18260 -13160
rect 18326 -13162 18338 -13160
rect 18338 -13162 18360 -13160
rect 18426 -13162 18428 -13160
rect 18428 -13162 18460 -13160
rect 18226 -13194 18260 -13162
rect 18326 -13194 18360 -13162
rect 18426 -13194 18460 -13162
rect 18526 -13194 18560 -13160
rect 18626 -13194 18660 -13160
rect 18726 -13162 18754 -13160
rect 18754 -13162 18760 -13160
rect 18726 -13194 18760 -13162
rect 18226 -13294 18260 -13260
rect 18326 -13294 18360 -13260
rect 18426 -13294 18460 -13260
rect 18526 -13294 18560 -13260
rect 18626 -13294 18660 -13260
rect 18726 -13294 18760 -13260
rect 18226 -13394 18260 -13360
rect 18326 -13394 18360 -13360
rect 18426 -13394 18460 -13360
rect 18526 -13394 18560 -13360
rect 18626 -13394 18660 -13360
rect 18726 -13394 18760 -13360
rect 18226 -13488 18260 -13460
rect 18326 -13488 18360 -13460
rect 18426 -13488 18460 -13460
rect 18226 -13494 18248 -13488
rect 18248 -13494 18260 -13488
rect 18326 -13494 18338 -13488
rect 18338 -13494 18360 -13488
rect 18426 -13494 18428 -13488
rect 18428 -13494 18460 -13488
rect 18526 -13494 18560 -13460
rect 18626 -13494 18660 -13460
rect 18726 -13488 18760 -13460
rect 18726 -13494 18754 -13488
rect 18754 -13494 18760 -13488
rect 19514 -12982 19536 -12960
rect 19536 -12982 19548 -12960
rect 19614 -12982 19626 -12960
rect 19626 -12982 19648 -12960
rect 19714 -12982 19716 -12960
rect 19716 -12982 19748 -12960
rect 19514 -12994 19548 -12982
rect 19614 -12994 19648 -12982
rect 19714 -12994 19748 -12982
rect 19814 -12994 19848 -12960
rect 19914 -12994 19948 -12960
rect 20014 -12982 20042 -12960
rect 20042 -12982 20048 -12960
rect 20014 -12994 20048 -12982
rect 19514 -13072 19536 -13060
rect 19536 -13072 19548 -13060
rect 19614 -13072 19626 -13060
rect 19626 -13072 19648 -13060
rect 19714 -13072 19716 -13060
rect 19716 -13072 19748 -13060
rect 19514 -13094 19548 -13072
rect 19614 -13094 19648 -13072
rect 19714 -13094 19748 -13072
rect 19814 -13094 19848 -13060
rect 19914 -13094 19948 -13060
rect 20014 -13072 20042 -13060
rect 20042 -13072 20048 -13060
rect 20014 -13094 20048 -13072
rect 19514 -13162 19536 -13160
rect 19536 -13162 19548 -13160
rect 19614 -13162 19626 -13160
rect 19626 -13162 19648 -13160
rect 19714 -13162 19716 -13160
rect 19716 -13162 19748 -13160
rect 19514 -13194 19548 -13162
rect 19614 -13194 19648 -13162
rect 19714 -13194 19748 -13162
rect 19814 -13194 19848 -13160
rect 19914 -13194 19948 -13160
rect 20014 -13162 20042 -13160
rect 20042 -13162 20048 -13160
rect 20014 -13194 20048 -13162
rect 19514 -13294 19548 -13260
rect 19614 -13294 19648 -13260
rect 19714 -13294 19748 -13260
rect 19814 -13294 19848 -13260
rect 19914 -13294 19948 -13260
rect 20014 -13294 20048 -13260
rect 19514 -13394 19548 -13360
rect 19614 -13394 19648 -13360
rect 19714 -13394 19748 -13360
rect 19814 -13394 19848 -13360
rect 19914 -13394 19948 -13360
rect 20014 -13394 20048 -13360
rect 19514 -13488 19548 -13460
rect 19614 -13488 19648 -13460
rect 19714 -13488 19748 -13460
rect 19514 -13494 19536 -13488
rect 19536 -13494 19548 -13488
rect 19614 -13494 19626 -13488
rect 19626 -13494 19648 -13488
rect 19714 -13494 19716 -13488
rect 19716 -13494 19748 -13488
rect 19814 -13494 19848 -13460
rect 19914 -13494 19948 -13460
rect 20014 -13488 20048 -13460
rect 20014 -13494 20042 -13488
rect 20042 -13494 20048 -13488
rect 20802 -12982 20824 -12960
rect 20824 -12982 20836 -12960
rect 20902 -12982 20914 -12960
rect 20914 -12982 20936 -12960
rect 21002 -12982 21004 -12960
rect 21004 -12982 21036 -12960
rect 20802 -12994 20836 -12982
rect 20902 -12994 20936 -12982
rect 21002 -12994 21036 -12982
rect 21102 -12994 21136 -12960
rect 21202 -12994 21236 -12960
rect 21302 -12982 21330 -12960
rect 21330 -12982 21336 -12960
rect 21302 -12994 21336 -12982
rect 20802 -13072 20824 -13060
rect 20824 -13072 20836 -13060
rect 20902 -13072 20914 -13060
rect 20914 -13072 20936 -13060
rect 21002 -13072 21004 -13060
rect 21004 -13072 21036 -13060
rect 20802 -13094 20836 -13072
rect 20902 -13094 20936 -13072
rect 21002 -13094 21036 -13072
rect 21102 -13094 21136 -13060
rect 21202 -13094 21236 -13060
rect 21302 -13072 21330 -13060
rect 21330 -13072 21336 -13060
rect 21302 -13094 21336 -13072
rect 20802 -13162 20824 -13160
rect 20824 -13162 20836 -13160
rect 20902 -13162 20914 -13160
rect 20914 -13162 20936 -13160
rect 21002 -13162 21004 -13160
rect 21004 -13162 21036 -13160
rect 20802 -13194 20836 -13162
rect 20902 -13194 20936 -13162
rect 21002 -13194 21036 -13162
rect 21102 -13194 21136 -13160
rect 21202 -13194 21236 -13160
rect 21302 -13162 21330 -13160
rect 21330 -13162 21336 -13160
rect 21302 -13194 21336 -13162
rect 20802 -13294 20836 -13260
rect 20902 -13294 20936 -13260
rect 21002 -13294 21036 -13260
rect 21102 -13294 21136 -13260
rect 21202 -13294 21236 -13260
rect 21302 -13294 21336 -13260
rect 20802 -13394 20836 -13360
rect 20902 -13394 20936 -13360
rect 21002 -13394 21036 -13360
rect 21102 -13394 21136 -13360
rect 21202 -13394 21236 -13360
rect 21302 -13394 21336 -13360
rect 20802 -13488 20836 -13460
rect 20902 -13488 20936 -13460
rect 21002 -13488 21036 -13460
rect 20802 -13494 20824 -13488
rect 20824 -13494 20836 -13488
rect 20902 -13494 20914 -13488
rect 20914 -13494 20936 -13488
rect 21002 -13494 21004 -13488
rect 21004 -13494 21036 -13488
rect 21102 -13494 21136 -13460
rect 21202 -13494 21236 -13460
rect 21302 -13488 21336 -13460
rect 21302 -13494 21330 -13488
rect 21330 -13494 21336 -13488
rect 22090 -12982 22112 -12960
rect 22112 -12982 22124 -12960
rect 22190 -12982 22202 -12960
rect 22202 -12982 22224 -12960
rect 22290 -12982 22292 -12960
rect 22292 -12982 22324 -12960
rect 22090 -12994 22124 -12982
rect 22190 -12994 22224 -12982
rect 22290 -12994 22324 -12982
rect 22390 -12994 22424 -12960
rect 22490 -12994 22524 -12960
rect 22590 -12982 22618 -12960
rect 22618 -12982 22624 -12960
rect 22590 -12994 22624 -12982
rect 22090 -13072 22112 -13060
rect 22112 -13072 22124 -13060
rect 22190 -13072 22202 -13060
rect 22202 -13072 22224 -13060
rect 22290 -13072 22292 -13060
rect 22292 -13072 22324 -13060
rect 22090 -13094 22124 -13072
rect 22190 -13094 22224 -13072
rect 22290 -13094 22324 -13072
rect 22390 -13094 22424 -13060
rect 22490 -13094 22524 -13060
rect 22590 -13072 22618 -13060
rect 22618 -13072 22624 -13060
rect 22590 -13094 22624 -13072
rect 22090 -13162 22112 -13160
rect 22112 -13162 22124 -13160
rect 22190 -13162 22202 -13160
rect 22202 -13162 22224 -13160
rect 22290 -13162 22292 -13160
rect 22292 -13162 22324 -13160
rect 22090 -13194 22124 -13162
rect 22190 -13194 22224 -13162
rect 22290 -13194 22324 -13162
rect 22390 -13194 22424 -13160
rect 22490 -13194 22524 -13160
rect 22590 -13162 22618 -13160
rect 22618 -13162 22624 -13160
rect 22590 -13194 22624 -13162
rect 22090 -13294 22124 -13260
rect 22190 -13294 22224 -13260
rect 22290 -13294 22324 -13260
rect 22390 -13294 22424 -13260
rect 22490 -13294 22524 -13260
rect 22590 -13294 22624 -13260
rect 22090 -13394 22124 -13360
rect 22190 -13394 22224 -13360
rect 22290 -13394 22324 -13360
rect 22390 -13394 22424 -13360
rect 22490 -13394 22524 -13360
rect 22590 -13394 22624 -13360
rect 22090 -13488 22124 -13460
rect 22190 -13488 22224 -13460
rect 22290 -13488 22324 -13460
rect 22090 -13494 22112 -13488
rect 22112 -13494 22124 -13488
rect 22190 -13494 22202 -13488
rect 22202 -13494 22224 -13488
rect 22290 -13494 22292 -13488
rect 22292 -13494 22324 -13488
rect 22390 -13494 22424 -13460
rect 22490 -13494 22524 -13460
rect 22590 -13488 22624 -13460
rect 22590 -13494 22618 -13488
rect 22618 -13494 22624 -13488
rect 23378 -12982 23400 -12960
rect 23400 -12982 23412 -12960
rect 23478 -12982 23490 -12960
rect 23490 -12982 23512 -12960
rect 23578 -12982 23580 -12960
rect 23580 -12982 23612 -12960
rect 23378 -12994 23412 -12982
rect 23478 -12994 23512 -12982
rect 23578 -12994 23612 -12982
rect 23678 -12994 23712 -12960
rect 23778 -12994 23812 -12960
rect 23878 -12982 23906 -12960
rect 23906 -12982 23912 -12960
rect 23878 -12994 23912 -12982
rect 23378 -13072 23400 -13060
rect 23400 -13072 23412 -13060
rect 23478 -13072 23490 -13060
rect 23490 -13072 23512 -13060
rect 23578 -13072 23580 -13060
rect 23580 -13072 23612 -13060
rect 23378 -13094 23412 -13072
rect 23478 -13094 23512 -13072
rect 23578 -13094 23612 -13072
rect 23678 -13094 23712 -13060
rect 23778 -13094 23812 -13060
rect 23878 -13072 23906 -13060
rect 23906 -13072 23912 -13060
rect 23878 -13094 23912 -13072
rect 23378 -13162 23400 -13160
rect 23400 -13162 23412 -13160
rect 23478 -13162 23490 -13160
rect 23490 -13162 23512 -13160
rect 23578 -13162 23580 -13160
rect 23580 -13162 23612 -13160
rect 23378 -13194 23412 -13162
rect 23478 -13194 23512 -13162
rect 23578 -13194 23612 -13162
rect 23678 -13194 23712 -13160
rect 23778 -13194 23812 -13160
rect 23878 -13162 23906 -13160
rect 23906 -13162 23912 -13160
rect 23878 -13194 23912 -13162
rect 23378 -13294 23412 -13260
rect 23478 -13294 23512 -13260
rect 23578 -13294 23612 -13260
rect 23678 -13294 23712 -13260
rect 23778 -13294 23812 -13260
rect 23878 -13294 23912 -13260
rect 23378 -13394 23412 -13360
rect 23478 -13394 23512 -13360
rect 23578 -13394 23612 -13360
rect 23678 -13394 23712 -13360
rect 23778 -13394 23812 -13360
rect 23878 -13394 23912 -13360
rect 23378 -13488 23412 -13460
rect 23478 -13488 23512 -13460
rect 23578 -13488 23612 -13460
rect 23378 -13494 23400 -13488
rect 23400 -13494 23412 -13488
rect 23478 -13494 23490 -13488
rect 23490 -13494 23512 -13488
rect 23578 -13494 23580 -13488
rect 23580 -13494 23612 -13488
rect 23678 -13494 23712 -13460
rect 23778 -13494 23812 -13460
rect 23878 -13488 23912 -13460
rect 23878 -13494 23906 -13488
rect 23906 -13494 23912 -13488
rect 24666 -12982 24688 -12960
rect 24688 -12982 24700 -12960
rect 24766 -12982 24778 -12960
rect 24778 -12982 24800 -12960
rect 24866 -12982 24868 -12960
rect 24868 -12982 24900 -12960
rect 24666 -12994 24700 -12982
rect 24766 -12994 24800 -12982
rect 24866 -12994 24900 -12982
rect 24966 -12994 25000 -12960
rect 25066 -12994 25100 -12960
rect 25166 -12982 25194 -12960
rect 25194 -12982 25200 -12960
rect 25166 -12994 25200 -12982
rect 24666 -13072 24688 -13060
rect 24688 -13072 24700 -13060
rect 24766 -13072 24778 -13060
rect 24778 -13072 24800 -13060
rect 24866 -13072 24868 -13060
rect 24868 -13072 24900 -13060
rect 24666 -13094 24700 -13072
rect 24766 -13094 24800 -13072
rect 24866 -13094 24900 -13072
rect 24966 -13094 25000 -13060
rect 25066 -13094 25100 -13060
rect 25166 -13072 25194 -13060
rect 25194 -13072 25200 -13060
rect 25166 -13094 25200 -13072
rect 24666 -13162 24688 -13160
rect 24688 -13162 24700 -13160
rect 24766 -13162 24778 -13160
rect 24778 -13162 24800 -13160
rect 24866 -13162 24868 -13160
rect 24868 -13162 24900 -13160
rect 24666 -13194 24700 -13162
rect 24766 -13194 24800 -13162
rect 24866 -13194 24900 -13162
rect 24966 -13194 25000 -13160
rect 25066 -13194 25100 -13160
rect 25166 -13162 25194 -13160
rect 25194 -13162 25200 -13160
rect 25166 -13194 25200 -13162
rect 24666 -13294 24700 -13260
rect 24766 -13294 24800 -13260
rect 24866 -13294 24900 -13260
rect 24966 -13294 25000 -13260
rect 25066 -13294 25100 -13260
rect 25166 -13294 25200 -13260
rect 24666 -13394 24700 -13360
rect 24766 -13394 24800 -13360
rect 24866 -13394 24900 -13360
rect 24966 -13394 25000 -13360
rect 25066 -13394 25100 -13360
rect 25166 -13394 25200 -13360
rect 24666 -13488 24700 -13460
rect 24766 -13488 24800 -13460
rect 24866 -13488 24900 -13460
rect 24666 -13494 24688 -13488
rect 24688 -13494 24700 -13488
rect 24766 -13494 24778 -13488
rect 24778 -13494 24800 -13488
rect 24866 -13494 24868 -13488
rect 24868 -13494 24900 -13488
rect 24966 -13494 25000 -13460
rect 25066 -13494 25100 -13460
rect 25166 -13488 25200 -13460
rect 25166 -13494 25194 -13488
rect 25194 -13494 25200 -13488
rect 25954 -12982 25976 -12960
rect 25976 -12982 25988 -12960
rect 26054 -12982 26066 -12960
rect 26066 -12982 26088 -12960
rect 26154 -12982 26156 -12960
rect 26156 -12982 26188 -12960
rect 25954 -12994 25988 -12982
rect 26054 -12994 26088 -12982
rect 26154 -12994 26188 -12982
rect 26254 -12994 26288 -12960
rect 26354 -12994 26388 -12960
rect 26454 -12982 26482 -12960
rect 26482 -12982 26488 -12960
rect 26454 -12994 26488 -12982
rect 25954 -13072 25976 -13060
rect 25976 -13072 25988 -13060
rect 26054 -13072 26066 -13060
rect 26066 -13072 26088 -13060
rect 26154 -13072 26156 -13060
rect 26156 -13072 26188 -13060
rect 25954 -13094 25988 -13072
rect 26054 -13094 26088 -13072
rect 26154 -13094 26188 -13072
rect 26254 -13094 26288 -13060
rect 26354 -13094 26388 -13060
rect 26454 -13072 26482 -13060
rect 26482 -13072 26488 -13060
rect 26454 -13094 26488 -13072
rect 25954 -13162 25976 -13160
rect 25976 -13162 25988 -13160
rect 26054 -13162 26066 -13160
rect 26066 -13162 26088 -13160
rect 26154 -13162 26156 -13160
rect 26156 -13162 26188 -13160
rect 25954 -13194 25988 -13162
rect 26054 -13194 26088 -13162
rect 26154 -13194 26188 -13162
rect 26254 -13194 26288 -13160
rect 26354 -13194 26388 -13160
rect 26454 -13162 26482 -13160
rect 26482 -13162 26488 -13160
rect 26454 -13194 26488 -13162
rect 25954 -13294 25988 -13260
rect 26054 -13294 26088 -13260
rect 26154 -13294 26188 -13260
rect 26254 -13294 26288 -13260
rect 26354 -13294 26388 -13260
rect 26454 -13294 26488 -13260
rect 25954 -13394 25988 -13360
rect 26054 -13394 26088 -13360
rect 26154 -13394 26188 -13360
rect 26254 -13394 26288 -13360
rect 26354 -13394 26388 -13360
rect 26454 -13394 26488 -13360
rect 25954 -13488 25988 -13460
rect 26054 -13488 26088 -13460
rect 26154 -13488 26188 -13460
rect 25954 -13494 25976 -13488
rect 25976 -13494 25988 -13488
rect 26054 -13494 26066 -13488
rect 26066 -13494 26088 -13488
rect 26154 -13494 26156 -13488
rect 26156 -13494 26188 -13488
rect 26254 -13494 26288 -13460
rect 26354 -13494 26388 -13460
rect 26454 -13488 26488 -13460
rect 26454 -13494 26482 -13488
rect 26482 -13494 26488 -13488
rect 16938 -14270 16960 -14248
rect 16960 -14270 16972 -14248
rect 17038 -14270 17050 -14248
rect 17050 -14270 17072 -14248
rect 17138 -14270 17140 -14248
rect 17140 -14270 17172 -14248
rect 16938 -14282 16972 -14270
rect 17038 -14282 17072 -14270
rect 17138 -14282 17172 -14270
rect 17238 -14282 17272 -14248
rect 17338 -14282 17372 -14248
rect 17438 -14270 17466 -14248
rect 17466 -14270 17472 -14248
rect 17438 -14282 17472 -14270
rect 16938 -14360 16960 -14348
rect 16960 -14360 16972 -14348
rect 17038 -14360 17050 -14348
rect 17050 -14360 17072 -14348
rect 17138 -14360 17140 -14348
rect 17140 -14360 17172 -14348
rect 16938 -14382 16972 -14360
rect 17038 -14382 17072 -14360
rect 17138 -14382 17172 -14360
rect 17238 -14382 17272 -14348
rect 17338 -14382 17372 -14348
rect 17438 -14360 17466 -14348
rect 17466 -14360 17472 -14348
rect 17438 -14382 17472 -14360
rect 16938 -14450 16960 -14448
rect 16960 -14450 16972 -14448
rect 17038 -14450 17050 -14448
rect 17050 -14450 17072 -14448
rect 17138 -14450 17140 -14448
rect 17140 -14450 17172 -14448
rect 16938 -14482 16972 -14450
rect 17038 -14482 17072 -14450
rect 17138 -14482 17172 -14450
rect 17238 -14482 17272 -14448
rect 17338 -14482 17372 -14448
rect 17438 -14450 17466 -14448
rect 17466 -14450 17472 -14448
rect 17438 -14482 17472 -14450
rect 16938 -14582 16972 -14548
rect 17038 -14582 17072 -14548
rect 17138 -14582 17172 -14548
rect 17238 -14582 17272 -14548
rect 17338 -14582 17372 -14548
rect 17438 -14582 17472 -14548
rect 16938 -14682 16972 -14648
rect 17038 -14682 17072 -14648
rect 17138 -14682 17172 -14648
rect 17238 -14682 17272 -14648
rect 17338 -14682 17372 -14648
rect 17438 -14682 17472 -14648
rect 16938 -14776 16972 -14748
rect 17038 -14776 17072 -14748
rect 17138 -14776 17172 -14748
rect 16938 -14782 16960 -14776
rect 16960 -14782 16972 -14776
rect 17038 -14782 17050 -14776
rect 17050 -14782 17072 -14776
rect 17138 -14782 17140 -14776
rect 17140 -14782 17172 -14776
rect 17238 -14782 17272 -14748
rect 17338 -14782 17372 -14748
rect 17438 -14776 17472 -14748
rect 17438 -14782 17466 -14776
rect 17466 -14782 17472 -14776
rect 18226 -14270 18248 -14248
rect 18248 -14270 18260 -14248
rect 18326 -14270 18338 -14248
rect 18338 -14270 18360 -14248
rect 18426 -14270 18428 -14248
rect 18428 -14270 18460 -14248
rect 18226 -14282 18260 -14270
rect 18326 -14282 18360 -14270
rect 18426 -14282 18460 -14270
rect 18526 -14282 18560 -14248
rect 18626 -14282 18660 -14248
rect 18726 -14270 18754 -14248
rect 18754 -14270 18760 -14248
rect 18726 -14282 18760 -14270
rect 18226 -14360 18248 -14348
rect 18248 -14360 18260 -14348
rect 18326 -14360 18338 -14348
rect 18338 -14360 18360 -14348
rect 18426 -14360 18428 -14348
rect 18428 -14360 18460 -14348
rect 18226 -14382 18260 -14360
rect 18326 -14382 18360 -14360
rect 18426 -14382 18460 -14360
rect 18526 -14382 18560 -14348
rect 18626 -14382 18660 -14348
rect 18726 -14360 18754 -14348
rect 18754 -14360 18760 -14348
rect 18726 -14382 18760 -14360
rect 18226 -14450 18248 -14448
rect 18248 -14450 18260 -14448
rect 18326 -14450 18338 -14448
rect 18338 -14450 18360 -14448
rect 18426 -14450 18428 -14448
rect 18428 -14450 18460 -14448
rect 18226 -14482 18260 -14450
rect 18326 -14482 18360 -14450
rect 18426 -14482 18460 -14450
rect 18526 -14482 18560 -14448
rect 18626 -14482 18660 -14448
rect 18726 -14450 18754 -14448
rect 18754 -14450 18760 -14448
rect 18726 -14482 18760 -14450
rect 18226 -14582 18260 -14548
rect 18326 -14582 18360 -14548
rect 18426 -14582 18460 -14548
rect 18526 -14582 18560 -14548
rect 18626 -14582 18660 -14548
rect 18726 -14582 18760 -14548
rect 18226 -14682 18260 -14648
rect 18326 -14682 18360 -14648
rect 18426 -14682 18460 -14648
rect 18526 -14682 18560 -14648
rect 18626 -14682 18660 -14648
rect 18726 -14682 18760 -14648
rect 18226 -14776 18260 -14748
rect 18326 -14776 18360 -14748
rect 18426 -14776 18460 -14748
rect 18226 -14782 18248 -14776
rect 18248 -14782 18260 -14776
rect 18326 -14782 18338 -14776
rect 18338 -14782 18360 -14776
rect 18426 -14782 18428 -14776
rect 18428 -14782 18460 -14776
rect 18526 -14782 18560 -14748
rect 18626 -14782 18660 -14748
rect 18726 -14776 18760 -14748
rect 18726 -14782 18754 -14776
rect 18754 -14782 18760 -14776
rect 19514 -14270 19536 -14248
rect 19536 -14270 19548 -14248
rect 19614 -14270 19626 -14248
rect 19626 -14270 19648 -14248
rect 19714 -14270 19716 -14248
rect 19716 -14270 19748 -14248
rect 19514 -14282 19548 -14270
rect 19614 -14282 19648 -14270
rect 19714 -14282 19748 -14270
rect 19814 -14282 19848 -14248
rect 19914 -14282 19948 -14248
rect 20014 -14270 20042 -14248
rect 20042 -14270 20048 -14248
rect 20014 -14282 20048 -14270
rect 19514 -14360 19536 -14348
rect 19536 -14360 19548 -14348
rect 19614 -14360 19626 -14348
rect 19626 -14360 19648 -14348
rect 19714 -14360 19716 -14348
rect 19716 -14360 19748 -14348
rect 19514 -14382 19548 -14360
rect 19614 -14382 19648 -14360
rect 19714 -14382 19748 -14360
rect 19814 -14382 19848 -14348
rect 19914 -14382 19948 -14348
rect 20014 -14360 20042 -14348
rect 20042 -14360 20048 -14348
rect 20014 -14382 20048 -14360
rect 19514 -14450 19536 -14448
rect 19536 -14450 19548 -14448
rect 19614 -14450 19626 -14448
rect 19626 -14450 19648 -14448
rect 19714 -14450 19716 -14448
rect 19716 -14450 19748 -14448
rect 19514 -14482 19548 -14450
rect 19614 -14482 19648 -14450
rect 19714 -14482 19748 -14450
rect 19814 -14482 19848 -14448
rect 19914 -14482 19948 -14448
rect 20014 -14450 20042 -14448
rect 20042 -14450 20048 -14448
rect 20014 -14482 20048 -14450
rect 19514 -14582 19548 -14548
rect 19614 -14582 19648 -14548
rect 19714 -14582 19748 -14548
rect 19814 -14582 19848 -14548
rect 19914 -14582 19948 -14548
rect 20014 -14582 20048 -14548
rect 19514 -14682 19548 -14648
rect 19614 -14682 19648 -14648
rect 19714 -14682 19748 -14648
rect 19814 -14682 19848 -14648
rect 19914 -14682 19948 -14648
rect 20014 -14682 20048 -14648
rect 19514 -14776 19548 -14748
rect 19614 -14776 19648 -14748
rect 19714 -14776 19748 -14748
rect 19514 -14782 19536 -14776
rect 19536 -14782 19548 -14776
rect 19614 -14782 19626 -14776
rect 19626 -14782 19648 -14776
rect 19714 -14782 19716 -14776
rect 19716 -14782 19748 -14776
rect 19814 -14782 19848 -14748
rect 19914 -14782 19948 -14748
rect 20014 -14776 20048 -14748
rect 20014 -14782 20042 -14776
rect 20042 -14782 20048 -14776
rect 20802 -14270 20824 -14248
rect 20824 -14270 20836 -14248
rect 20902 -14270 20914 -14248
rect 20914 -14270 20936 -14248
rect 21002 -14270 21004 -14248
rect 21004 -14270 21036 -14248
rect 20802 -14282 20836 -14270
rect 20902 -14282 20936 -14270
rect 21002 -14282 21036 -14270
rect 21102 -14282 21136 -14248
rect 21202 -14282 21236 -14248
rect 21302 -14270 21330 -14248
rect 21330 -14270 21336 -14248
rect 21302 -14282 21336 -14270
rect 20802 -14360 20824 -14348
rect 20824 -14360 20836 -14348
rect 20902 -14360 20914 -14348
rect 20914 -14360 20936 -14348
rect 21002 -14360 21004 -14348
rect 21004 -14360 21036 -14348
rect 20802 -14382 20836 -14360
rect 20902 -14382 20936 -14360
rect 21002 -14382 21036 -14360
rect 21102 -14382 21136 -14348
rect 21202 -14382 21236 -14348
rect 21302 -14360 21330 -14348
rect 21330 -14360 21336 -14348
rect 21302 -14382 21336 -14360
rect 20802 -14450 20824 -14448
rect 20824 -14450 20836 -14448
rect 20902 -14450 20914 -14448
rect 20914 -14450 20936 -14448
rect 21002 -14450 21004 -14448
rect 21004 -14450 21036 -14448
rect 20802 -14482 20836 -14450
rect 20902 -14482 20936 -14450
rect 21002 -14482 21036 -14450
rect 21102 -14482 21136 -14448
rect 21202 -14482 21236 -14448
rect 21302 -14450 21330 -14448
rect 21330 -14450 21336 -14448
rect 21302 -14482 21336 -14450
rect 20802 -14582 20836 -14548
rect 20902 -14582 20936 -14548
rect 21002 -14582 21036 -14548
rect 21102 -14582 21136 -14548
rect 21202 -14582 21236 -14548
rect 21302 -14582 21336 -14548
rect 20802 -14682 20836 -14648
rect 20902 -14682 20936 -14648
rect 21002 -14682 21036 -14648
rect 21102 -14682 21136 -14648
rect 21202 -14682 21236 -14648
rect 21302 -14682 21336 -14648
rect 20802 -14776 20836 -14748
rect 20902 -14776 20936 -14748
rect 21002 -14776 21036 -14748
rect 20802 -14782 20824 -14776
rect 20824 -14782 20836 -14776
rect 20902 -14782 20914 -14776
rect 20914 -14782 20936 -14776
rect 21002 -14782 21004 -14776
rect 21004 -14782 21036 -14776
rect 21102 -14782 21136 -14748
rect 21202 -14782 21236 -14748
rect 21302 -14776 21336 -14748
rect 21302 -14782 21330 -14776
rect 21330 -14782 21336 -14776
rect 22090 -14270 22112 -14248
rect 22112 -14270 22124 -14248
rect 22190 -14270 22202 -14248
rect 22202 -14270 22224 -14248
rect 22290 -14270 22292 -14248
rect 22292 -14270 22324 -14248
rect 22090 -14282 22124 -14270
rect 22190 -14282 22224 -14270
rect 22290 -14282 22324 -14270
rect 22390 -14282 22424 -14248
rect 22490 -14282 22524 -14248
rect 22590 -14270 22618 -14248
rect 22618 -14270 22624 -14248
rect 22590 -14282 22624 -14270
rect 22090 -14360 22112 -14348
rect 22112 -14360 22124 -14348
rect 22190 -14360 22202 -14348
rect 22202 -14360 22224 -14348
rect 22290 -14360 22292 -14348
rect 22292 -14360 22324 -14348
rect 22090 -14382 22124 -14360
rect 22190 -14382 22224 -14360
rect 22290 -14382 22324 -14360
rect 22390 -14382 22424 -14348
rect 22490 -14382 22524 -14348
rect 22590 -14360 22618 -14348
rect 22618 -14360 22624 -14348
rect 22590 -14382 22624 -14360
rect 22090 -14450 22112 -14448
rect 22112 -14450 22124 -14448
rect 22190 -14450 22202 -14448
rect 22202 -14450 22224 -14448
rect 22290 -14450 22292 -14448
rect 22292 -14450 22324 -14448
rect 22090 -14482 22124 -14450
rect 22190 -14482 22224 -14450
rect 22290 -14482 22324 -14450
rect 22390 -14482 22424 -14448
rect 22490 -14482 22524 -14448
rect 22590 -14450 22618 -14448
rect 22618 -14450 22624 -14448
rect 22590 -14482 22624 -14450
rect 22090 -14582 22124 -14548
rect 22190 -14582 22224 -14548
rect 22290 -14582 22324 -14548
rect 22390 -14582 22424 -14548
rect 22490 -14582 22524 -14548
rect 22590 -14582 22624 -14548
rect 22090 -14682 22124 -14648
rect 22190 -14682 22224 -14648
rect 22290 -14682 22324 -14648
rect 22390 -14682 22424 -14648
rect 22490 -14682 22524 -14648
rect 22590 -14682 22624 -14648
rect 22090 -14776 22124 -14748
rect 22190 -14776 22224 -14748
rect 22290 -14776 22324 -14748
rect 22090 -14782 22112 -14776
rect 22112 -14782 22124 -14776
rect 22190 -14782 22202 -14776
rect 22202 -14782 22224 -14776
rect 22290 -14782 22292 -14776
rect 22292 -14782 22324 -14776
rect 22390 -14782 22424 -14748
rect 22490 -14782 22524 -14748
rect 22590 -14776 22624 -14748
rect 22590 -14782 22618 -14776
rect 22618 -14782 22624 -14776
rect 23378 -14270 23400 -14248
rect 23400 -14270 23412 -14248
rect 23478 -14270 23490 -14248
rect 23490 -14270 23512 -14248
rect 23578 -14270 23580 -14248
rect 23580 -14270 23612 -14248
rect 23378 -14282 23412 -14270
rect 23478 -14282 23512 -14270
rect 23578 -14282 23612 -14270
rect 23678 -14282 23712 -14248
rect 23778 -14282 23812 -14248
rect 23878 -14270 23906 -14248
rect 23906 -14270 23912 -14248
rect 23878 -14282 23912 -14270
rect 23378 -14360 23400 -14348
rect 23400 -14360 23412 -14348
rect 23478 -14360 23490 -14348
rect 23490 -14360 23512 -14348
rect 23578 -14360 23580 -14348
rect 23580 -14360 23612 -14348
rect 23378 -14382 23412 -14360
rect 23478 -14382 23512 -14360
rect 23578 -14382 23612 -14360
rect 23678 -14382 23712 -14348
rect 23778 -14382 23812 -14348
rect 23878 -14360 23906 -14348
rect 23906 -14360 23912 -14348
rect 23878 -14382 23912 -14360
rect 23378 -14450 23400 -14448
rect 23400 -14450 23412 -14448
rect 23478 -14450 23490 -14448
rect 23490 -14450 23512 -14448
rect 23578 -14450 23580 -14448
rect 23580 -14450 23612 -14448
rect 23378 -14482 23412 -14450
rect 23478 -14482 23512 -14450
rect 23578 -14482 23612 -14450
rect 23678 -14482 23712 -14448
rect 23778 -14482 23812 -14448
rect 23878 -14450 23906 -14448
rect 23906 -14450 23912 -14448
rect 23878 -14482 23912 -14450
rect 23378 -14582 23412 -14548
rect 23478 -14582 23512 -14548
rect 23578 -14582 23612 -14548
rect 23678 -14582 23712 -14548
rect 23778 -14582 23812 -14548
rect 23878 -14582 23912 -14548
rect 23378 -14682 23412 -14648
rect 23478 -14682 23512 -14648
rect 23578 -14682 23612 -14648
rect 23678 -14682 23712 -14648
rect 23778 -14682 23812 -14648
rect 23878 -14682 23912 -14648
rect 23378 -14776 23412 -14748
rect 23478 -14776 23512 -14748
rect 23578 -14776 23612 -14748
rect 23378 -14782 23400 -14776
rect 23400 -14782 23412 -14776
rect 23478 -14782 23490 -14776
rect 23490 -14782 23512 -14776
rect 23578 -14782 23580 -14776
rect 23580 -14782 23612 -14776
rect 23678 -14782 23712 -14748
rect 23778 -14782 23812 -14748
rect 23878 -14776 23912 -14748
rect 23878 -14782 23906 -14776
rect 23906 -14782 23912 -14776
rect 24666 -14270 24688 -14248
rect 24688 -14270 24700 -14248
rect 24766 -14270 24778 -14248
rect 24778 -14270 24800 -14248
rect 24866 -14270 24868 -14248
rect 24868 -14270 24900 -14248
rect 24666 -14282 24700 -14270
rect 24766 -14282 24800 -14270
rect 24866 -14282 24900 -14270
rect 24966 -14282 25000 -14248
rect 25066 -14282 25100 -14248
rect 25166 -14270 25194 -14248
rect 25194 -14270 25200 -14248
rect 25166 -14282 25200 -14270
rect 24666 -14360 24688 -14348
rect 24688 -14360 24700 -14348
rect 24766 -14360 24778 -14348
rect 24778 -14360 24800 -14348
rect 24866 -14360 24868 -14348
rect 24868 -14360 24900 -14348
rect 24666 -14382 24700 -14360
rect 24766 -14382 24800 -14360
rect 24866 -14382 24900 -14360
rect 24966 -14382 25000 -14348
rect 25066 -14382 25100 -14348
rect 25166 -14360 25194 -14348
rect 25194 -14360 25200 -14348
rect 25166 -14382 25200 -14360
rect 24666 -14450 24688 -14448
rect 24688 -14450 24700 -14448
rect 24766 -14450 24778 -14448
rect 24778 -14450 24800 -14448
rect 24866 -14450 24868 -14448
rect 24868 -14450 24900 -14448
rect 24666 -14482 24700 -14450
rect 24766 -14482 24800 -14450
rect 24866 -14482 24900 -14450
rect 24966 -14482 25000 -14448
rect 25066 -14482 25100 -14448
rect 25166 -14450 25194 -14448
rect 25194 -14450 25200 -14448
rect 25166 -14482 25200 -14450
rect 24666 -14582 24700 -14548
rect 24766 -14582 24800 -14548
rect 24866 -14582 24900 -14548
rect 24966 -14582 25000 -14548
rect 25066 -14582 25100 -14548
rect 25166 -14582 25200 -14548
rect 24666 -14682 24700 -14648
rect 24766 -14682 24800 -14648
rect 24866 -14682 24900 -14648
rect 24966 -14682 25000 -14648
rect 25066 -14682 25100 -14648
rect 25166 -14682 25200 -14648
rect 24666 -14776 24700 -14748
rect 24766 -14776 24800 -14748
rect 24866 -14776 24900 -14748
rect 24666 -14782 24688 -14776
rect 24688 -14782 24700 -14776
rect 24766 -14782 24778 -14776
rect 24778 -14782 24800 -14776
rect 24866 -14782 24868 -14776
rect 24868 -14782 24900 -14776
rect 24966 -14782 25000 -14748
rect 25066 -14782 25100 -14748
rect 25166 -14776 25200 -14748
rect 25166 -14782 25194 -14776
rect 25194 -14782 25200 -14776
rect 25954 -14270 25976 -14248
rect 25976 -14270 25988 -14248
rect 26054 -14270 26066 -14248
rect 26066 -14270 26088 -14248
rect 26154 -14270 26156 -14248
rect 26156 -14270 26188 -14248
rect 25954 -14282 25988 -14270
rect 26054 -14282 26088 -14270
rect 26154 -14282 26188 -14270
rect 26254 -14282 26288 -14248
rect 26354 -14282 26388 -14248
rect 26454 -14270 26482 -14248
rect 26482 -14270 26488 -14248
rect 26454 -14282 26488 -14270
rect 25954 -14360 25976 -14348
rect 25976 -14360 25988 -14348
rect 26054 -14360 26066 -14348
rect 26066 -14360 26088 -14348
rect 26154 -14360 26156 -14348
rect 26156 -14360 26188 -14348
rect 25954 -14382 25988 -14360
rect 26054 -14382 26088 -14360
rect 26154 -14382 26188 -14360
rect 26254 -14382 26288 -14348
rect 26354 -14382 26388 -14348
rect 26454 -14360 26482 -14348
rect 26482 -14360 26488 -14348
rect 26454 -14382 26488 -14360
rect 25954 -14450 25976 -14448
rect 25976 -14450 25988 -14448
rect 26054 -14450 26066 -14448
rect 26066 -14450 26088 -14448
rect 26154 -14450 26156 -14448
rect 26156 -14450 26188 -14448
rect 25954 -14482 25988 -14450
rect 26054 -14482 26088 -14450
rect 26154 -14482 26188 -14450
rect 26254 -14482 26288 -14448
rect 26354 -14482 26388 -14448
rect 26454 -14450 26482 -14448
rect 26482 -14450 26488 -14448
rect 26454 -14482 26488 -14450
rect 25954 -14582 25988 -14548
rect 26054 -14582 26088 -14548
rect 26154 -14582 26188 -14548
rect 26254 -14582 26288 -14548
rect 26354 -14582 26388 -14548
rect 26454 -14582 26488 -14548
rect 25954 -14682 25988 -14648
rect 26054 -14682 26088 -14648
rect 26154 -14682 26188 -14648
rect 26254 -14682 26288 -14648
rect 26354 -14682 26388 -14648
rect 26454 -14682 26488 -14648
rect 25954 -14776 25988 -14748
rect 26054 -14776 26088 -14748
rect 26154 -14776 26188 -14748
rect 25954 -14782 25976 -14776
rect 25976 -14782 25988 -14776
rect 26054 -14782 26066 -14776
rect 26066 -14782 26088 -14776
rect 26154 -14782 26156 -14776
rect 26156 -14782 26188 -14776
rect 26254 -14782 26288 -14748
rect 26354 -14782 26388 -14748
rect 26454 -14776 26488 -14748
rect 26454 -14782 26482 -14776
rect 26482 -14782 26488 -14776
rect 16938 -15558 16960 -15536
rect 16960 -15558 16972 -15536
rect 17038 -15558 17050 -15536
rect 17050 -15558 17072 -15536
rect 17138 -15558 17140 -15536
rect 17140 -15558 17172 -15536
rect 16938 -15570 16972 -15558
rect 17038 -15570 17072 -15558
rect 17138 -15570 17172 -15558
rect 17238 -15570 17272 -15536
rect 17338 -15570 17372 -15536
rect 17438 -15558 17466 -15536
rect 17466 -15558 17472 -15536
rect 17438 -15570 17472 -15558
rect 16938 -15648 16960 -15636
rect 16960 -15648 16972 -15636
rect 17038 -15648 17050 -15636
rect 17050 -15648 17072 -15636
rect 17138 -15648 17140 -15636
rect 17140 -15648 17172 -15636
rect 16938 -15670 16972 -15648
rect 17038 -15670 17072 -15648
rect 17138 -15670 17172 -15648
rect 17238 -15670 17272 -15636
rect 17338 -15670 17372 -15636
rect 17438 -15648 17466 -15636
rect 17466 -15648 17472 -15636
rect 17438 -15670 17472 -15648
rect 16938 -15738 16960 -15736
rect 16960 -15738 16972 -15736
rect 17038 -15738 17050 -15736
rect 17050 -15738 17072 -15736
rect 17138 -15738 17140 -15736
rect 17140 -15738 17172 -15736
rect 16938 -15770 16972 -15738
rect 17038 -15770 17072 -15738
rect 17138 -15770 17172 -15738
rect 17238 -15770 17272 -15736
rect 17338 -15770 17372 -15736
rect 17438 -15738 17466 -15736
rect 17466 -15738 17472 -15736
rect 17438 -15770 17472 -15738
rect 16938 -15870 16972 -15836
rect 17038 -15870 17072 -15836
rect 17138 -15870 17172 -15836
rect 17238 -15870 17272 -15836
rect 17338 -15870 17372 -15836
rect 17438 -15870 17472 -15836
rect 16938 -15970 16972 -15936
rect 17038 -15970 17072 -15936
rect 17138 -15970 17172 -15936
rect 17238 -15970 17272 -15936
rect 17338 -15970 17372 -15936
rect 17438 -15970 17472 -15936
rect 16938 -16064 16972 -16036
rect 17038 -16064 17072 -16036
rect 17138 -16064 17172 -16036
rect 16938 -16070 16960 -16064
rect 16960 -16070 16972 -16064
rect 17038 -16070 17050 -16064
rect 17050 -16070 17072 -16064
rect 17138 -16070 17140 -16064
rect 17140 -16070 17172 -16064
rect 17238 -16070 17272 -16036
rect 17338 -16070 17372 -16036
rect 17438 -16064 17472 -16036
rect 17438 -16070 17466 -16064
rect 17466 -16070 17472 -16064
rect 18226 -15558 18248 -15536
rect 18248 -15558 18260 -15536
rect 18326 -15558 18338 -15536
rect 18338 -15558 18360 -15536
rect 18426 -15558 18428 -15536
rect 18428 -15558 18460 -15536
rect 18226 -15570 18260 -15558
rect 18326 -15570 18360 -15558
rect 18426 -15570 18460 -15558
rect 18526 -15570 18560 -15536
rect 18626 -15570 18660 -15536
rect 18726 -15558 18754 -15536
rect 18754 -15558 18760 -15536
rect 18726 -15570 18760 -15558
rect 18226 -15648 18248 -15636
rect 18248 -15648 18260 -15636
rect 18326 -15648 18338 -15636
rect 18338 -15648 18360 -15636
rect 18426 -15648 18428 -15636
rect 18428 -15648 18460 -15636
rect 18226 -15670 18260 -15648
rect 18326 -15670 18360 -15648
rect 18426 -15670 18460 -15648
rect 18526 -15670 18560 -15636
rect 18626 -15670 18660 -15636
rect 18726 -15648 18754 -15636
rect 18754 -15648 18760 -15636
rect 18726 -15670 18760 -15648
rect 18226 -15738 18248 -15736
rect 18248 -15738 18260 -15736
rect 18326 -15738 18338 -15736
rect 18338 -15738 18360 -15736
rect 18426 -15738 18428 -15736
rect 18428 -15738 18460 -15736
rect 18226 -15770 18260 -15738
rect 18326 -15770 18360 -15738
rect 18426 -15770 18460 -15738
rect 18526 -15770 18560 -15736
rect 18626 -15770 18660 -15736
rect 18726 -15738 18754 -15736
rect 18754 -15738 18760 -15736
rect 18726 -15770 18760 -15738
rect 18226 -15870 18260 -15836
rect 18326 -15870 18360 -15836
rect 18426 -15870 18460 -15836
rect 18526 -15870 18560 -15836
rect 18626 -15870 18660 -15836
rect 18726 -15870 18760 -15836
rect 18226 -15970 18260 -15936
rect 18326 -15970 18360 -15936
rect 18426 -15970 18460 -15936
rect 18526 -15970 18560 -15936
rect 18626 -15970 18660 -15936
rect 18726 -15970 18760 -15936
rect 18226 -16064 18260 -16036
rect 18326 -16064 18360 -16036
rect 18426 -16064 18460 -16036
rect 18226 -16070 18248 -16064
rect 18248 -16070 18260 -16064
rect 18326 -16070 18338 -16064
rect 18338 -16070 18360 -16064
rect 18426 -16070 18428 -16064
rect 18428 -16070 18460 -16064
rect 18526 -16070 18560 -16036
rect 18626 -16070 18660 -16036
rect 18726 -16064 18760 -16036
rect 18726 -16070 18754 -16064
rect 18754 -16070 18760 -16064
rect 19514 -15558 19536 -15536
rect 19536 -15558 19548 -15536
rect 19614 -15558 19626 -15536
rect 19626 -15558 19648 -15536
rect 19714 -15558 19716 -15536
rect 19716 -15558 19748 -15536
rect 19514 -15570 19548 -15558
rect 19614 -15570 19648 -15558
rect 19714 -15570 19748 -15558
rect 19814 -15570 19848 -15536
rect 19914 -15570 19948 -15536
rect 20014 -15558 20042 -15536
rect 20042 -15558 20048 -15536
rect 20014 -15570 20048 -15558
rect 19514 -15648 19536 -15636
rect 19536 -15648 19548 -15636
rect 19614 -15648 19626 -15636
rect 19626 -15648 19648 -15636
rect 19714 -15648 19716 -15636
rect 19716 -15648 19748 -15636
rect 19514 -15670 19548 -15648
rect 19614 -15670 19648 -15648
rect 19714 -15670 19748 -15648
rect 19814 -15670 19848 -15636
rect 19914 -15670 19948 -15636
rect 20014 -15648 20042 -15636
rect 20042 -15648 20048 -15636
rect 20014 -15670 20048 -15648
rect 19514 -15738 19536 -15736
rect 19536 -15738 19548 -15736
rect 19614 -15738 19626 -15736
rect 19626 -15738 19648 -15736
rect 19714 -15738 19716 -15736
rect 19716 -15738 19748 -15736
rect 19514 -15770 19548 -15738
rect 19614 -15770 19648 -15738
rect 19714 -15770 19748 -15738
rect 19814 -15770 19848 -15736
rect 19914 -15770 19948 -15736
rect 20014 -15738 20042 -15736
rect 20042 -15738 20048 -15736
rect 20014 -15770 20048 -15738
rect 19514 -15870 19548 -15836
rect 19614 -15870 19648 -15836
rect 19714 -15870 19748 -15836
rect 19814 -15870 19848 -15836
rect 19914 -15870 19948 -15836
rect 20014 -15870 20048 -15836
rect 19514 -15970 19548 -15936
rect 19614 -15970 19648 -15936
rect 19714 -15970 19748 -15936
rect 19814 -15970 19848 -15936
rect 19914 -15970 19948 -15936
rect 20014 -15970 20048 -15936
rect 19514 -16064 19548 -16036
rect 19614 -16064 19648 -16036
rect 19714 -16064 19748 -16036
rect 19514 -16070 19536 -16064
rect 19536 -16070 19548 -16064
rect 19614 -16070 19626 -16064
rect 19626 -16070 19648 -16064
rect 19714 -16070 19716 -16064
rect 19716 -16070 19748 -16064
rect 19814 -16070 19848 -16036
rect 19914 -16070 19948 -16036
rect 20014 -16064 20048 -16036
rect 20014 -16070 20042 -16064
rect 20042 -16070 20048 -16064
rect 20802 -15558 20824 -15536
rect 20824 -15558 20836 -15536
rect 20902 -15558 20914 -15536
rect 20914 -15558 20936 -15536
rect 21002 -15558 21004 -15536
rect 21004 -15558 21036 -15536
rect 20802 -15570 20836 -15558
rect 20902 -15570 20936 -15558
rect 21002 -15570 21036 -15558
rect 21102 -15570 21136 -15536
rect 21202 -15570 21236 -15536
rect 21302 -15558 21330 -15536
rect 21330 -15558 21336 -15536
rect 21302 -15570 21336 -15558
rect 20802 -15648 20824 -15636
rect 20824 -15648 20836 -15636
rect 20902 -15648 20914 -15636
rect 20914 -15648 20936 -15636
rect 21002 -15648 21004 -15636
rect 21004 -15648 21036 -15636
rect 20802 -15670 20836 -15648
rect 20902 -15670 20936 -15648
rect 21002 -15670 21036 -15648
rect 21102 -15670 21136 -15636
rect 21202 -15670 21236 -15636
rect 21302 -15648 21330 -15636
rect 21330 -15648 21336 -15636
rect 21302 -15670 21336 -15648
rect 20802 -15738 20824 -15736
rect 20824 -15738 20836 -15736
rect 20902 -15738 20914 -15736
rect 20914 -15738 20936 -15736
rect 21002 -15738 21004 -15736
rect 21004 -15738 21036 -15736
rect 20802 -15770 20836 -15738
rect 20902 -15770 20936 -15738
rect 21002 -15770 21036 -15738
rect 21102 -15770 21136 -15736
rect 21202 -15770 21236 -15736
rect 21302 -15738 21330 -15736
rect 21330 -15738 21336 -15736
rect 21302 -15770 21336 -15738
rect 20802 -15870 20836 -15836
rect 20902 -15870 20936 -15836
rect 21002 -15870 21036 -15836
rect 21102 -15870 21136 -15836
rect 21202 -15870 21236 -15836
rect 21302 -15870 21336 -15836
rect 20802 -15970 20836 -15936
rect 20902 -15970 20936 -15936
rect 21002 -15970 21036 -15936
rect 21102 -15970 21136 -15936
rect 21202 -15970 21236 -15936
rect 21302 -15970 21336 -15936
rect 20802 -16064 20836 -16036
rect 20902 -16064 20936 -16036
rect 21002 -16064 21036 -16036
rect 20802 -16070 20824 -16064
rect 20824 -16070 20836 -16064
rect 20902 -16070 20914 -16064
rect 20914 -16070 20936 -16064
rect 21002 -16070 21004 -16064
rect 21004 -16070 21036 -16064
rect 21102 -16070 21136 -16036
rect 21202 -16070 21236 -16036
rect 21302 -16064 21336 -16036
rect 21302 -16070 21330 -16064
rect 21330 -16070 21336 -16064
rect 22090 -15558 22112 -15536
rect 22112 -15558 22124 -15536
rect 22190 -15558 22202 -15536
rect 22202 -15558 22224 -15536
rect 22290 -15558 22292 -15536
rect 22292 -15558 22324 -15536
rect 22090 -15570 22124 -15558
rect 22190 -15570 22224 -15558
rect 22290 -15570 22324 -15558
rect 22390 -15570 22424 -15536
rect 22490 -15570 22524 -15536
rect 22590 -15558 22618 -15536
rect 22618 -15558 22624 -15536
rect 22590 -15570 22624 -15558
rect 22090 -15648 22112 -15636
rect 22112 -15648 22124 -15636
rect 22190 -15648 22202 -15636
rect 22202 -15648 22224 -15636
rect 22290 -15648 22292 -15636
rect 22292 -15648 22324 -15636
rect 22090 -15670 22124 -15648
rect 22190 -15670 22224 -15648
rect 22290 -15670 22324 -15648
rect 22390 -15670 22424 -15636
rect 22490 -15670 22524 -15636
rect 22590 -15648 22618 -15636
rect 22618 -15648 22624 -15636
rect 22590 -15670 22624 -15648
rect 22090 -15738 22112 -15736
rect 22112 -15738 22124 -15736
rect 22190 -15738 22202 -15736
rect 22202 -15738 22224 -15736
rect 22290 -15738 22292 -15736
rect 22292 -15738 22324 -15736
rect 22090 -15770 22124 -15738
rect 22190 -15770 22224 -15738
rect 22290 -15770 22324 -15738
rect 22390 -15770 22424 -15736
rect 22490 -15770 22524 -15736
rect 22590 -15738 22618 -15736
rect 22618 -15738 22624 -15736
rect 22590 -15770 22624 -15738
rect 22090 -15870 22124 -15836
rect 22190 -15870 22224 -15836
rect 22290 -15870 22324 -15836
rect 22390 -15870 22424 -15836
rect 22490 -15870 22524 -15836
rect 22590 -15870 22624 -15836
rect 22090 -15970 22124 -15936
rect 22190 -15970 22224 -15936
rect 22290 -15970 22324 -15936
rect 22390 -15970 22424 -15936
rect 22490 -15970 22524 -15936
rect 22590 -15970 22624 -15936
rect 22090 -16064 22124 -16036
rect 22190 -16064 22224 -16036
rect 22290 -16064 22324 -16036
rect 22090 -16070 22112 -16064
rect 22112 -16070 22124 -16064
rect 22190 -16070 22202 -16064
rect 22202 -16070 22224 -16064
rect 22290 -16070 22292 -16064
rect 22292 -16070 22324 -16064
rect 22390 -16070 22424 -16036
rect 22490 -16070 22524 -16036
rect 22590 -16064 22624 -16036
rect 22590 -16070 22618 -16064
rect 22618 -16070 22624 -16064
rect 23378 -15558 23400 -15536
rect 23400 -15558 23412 -15536
rect 23478 -15558 23490 -15536
rect 23490 -15558 23512 -15536
rect 23578 -15558 23580 -15536
rect 23580 -15558 23612 -15536
rect 23378 -15570 23412 -15558
rect 23478 -15570 23512 -15558
rect 23578 -15570 23612 -15558
rect 23678 -15570 23712 -15536
rect 23778 -15570 23812 -15536
rect 23878 -15558 23906 -15536
rect 23906 -15558 23912 -15536
rect 23878 -15570 23912 -15558
rect 23378 -15648 23400 -15636
rect 23400 -15648 23412 -15636
rect 23478 -15648 23490 -15636
rect 23490 -15648 23512 -15636
rect 23578 -15648 23580 -15636
rect 23580 -15648 23612 -15636
rect 23378 -15670 23412 -15648
rect 23478 -15670 23512 -15648
rect 23578 -15670 23612 -15648
rect 23678 -15670 23712 -15636
rect 23778 -15670 23812 -15636
rect 23878 -15648 23906 -15636
rect 23906 -15648 23912 -15636
rect 23878 -15670 23912 -15648
rect 23378 -15738 23400 -15736
rect 23400 -15738 23412 -15736
rect 23478 -15738 23490 -15736
rect 23490 -15738 23512 -15736
rect 23578 -15738 23580 -15736
rect 23580 -15738 23612 -15736
rect 23378 -15770 23412 -15738
rect 23478 -15770 23512 -15738
rect 23578 -15770 23612 -15738
rect 23678 -15770 23712 -15736
rect 23778 -15770 23812 -15736
rect 23878 -15738 23906 -15736
rect 23906 -15738 23912 -15736
rect 23878 -15770 23912 -15738
rect 23378 -15870 23412 -15836
rect 23478 -15870 23512 -15836
rect 23578 -15870 23612 -15836
rect 23678 -15870 23712 -15836
rect 23778 -15870 23812 -15836
rect 23878 -15870 23912 -15836
rect 23378 -15970 23412 -15936
rect 23478 -15970 23512 -15936
rect 23578 -15970 23612 -15936
rect 23678 -15970 23712 -15936
rect 23778 -15970 23812 -15936
rect 23878 -15970 23912 -15936
rect 23378 -16064 23412 -16036
rect 23478 -16064 23512 -16036
rect 23578 -16064 23612 -16036
rect 23378 -16070 23400 -16064
rect 23400 -16070 23412 -16064
rect 23478 -16070 23490 -16064
rect 23490 -16070 23512 -16064
rect 23578 -16070 23580 -16064
rect 23580 -16070 23612 -16064
rect 23678 -16070 23712 -16036
rect 23778 -16070 23812 -16036
rect 23878 -16064 23912 -16036
rect 23878 -16070 23906 -16064
rect 23906 -16070 23912 -16064
rect 24666 -15558 24688 -15536
rect 24688 -15558 24700 -15536
rect 24766 -15558 24778 -15536
rect 24778 -15558 24800 -15536
rect 24866 -15558 24868 -15536
rect 24868 -15558 24900 -15536
rect 24666 -15570 24700 -15558
rect 24766 -15570 24800 -15558
rect 24866 -15570 24900 -15558
rect 24966 -15570 25000 -15536
rect 25066 -15570 25100 -15536
rect 25166 -15558 25194 -15536
rect 25194 -15558 25200 -15536
rect 25166 -15570 25200 -15558
rect 24666 -15648 24688 -15636
rect 24688 -15648 24700 -15636
rect 24766 -15648 24778 -15636
rect 24778 -15648 24800 -15636
rect 24866 -15648 24868 -15636
rect 24868 -15648 24900 -15636
rect 24666 -15670 24700 -15648
rect 24766 -15670 24800 -15648
rect 24866 -15670 24900 -15648
rect 24966 -15670 25000 -15636
rect 25066 -15670 25100 -15636
rect 25166 -15648 25194 -15636
rect 25194 -15648 25200 -15636
rect 25166 -15670 25200 -15648
rect 24666 -15738 24688 -15736
rect 24688 -15738 24700 -15736
rect 24766 -15738 24778 -15736
rect 24778 -15738 24800 -15736
rect 24866 -15738 24868 -15736
rect 24868 -15738 24900 -15736
rect 24666 -15770 24700 -15738
rect 24766 -15770 24800 -15738
rect 24866 -15770 24900 -15738
rect 24966 -15770 25000 -15736
rect 25066 -15770 25100 -15736
rect 25166 -15738 25194 -15736
rect 25194 -15738 25200 -15736
rect 25166 -15770 25200 -15738
rect 24666 -15870 24700 -15836
rect 24766 -15870 24800 -15836
rect 24866 -15870 24900 -15836
rect 24966 -15870 25000 -15836
rect 25066 -15870 25100 -15836
rect 25166 -15870 25200 -15836
rect 24666 -15970 24700 -15936
rect 24766 -15970 24800 -15936
rect 24866 -15970 24900 -15936
rect 24966 -15970 25000 -15936
rect 25066 -15970 25100 -15936
rect 25166 -15970 25200 -15936
rect 24666 -16064 24700 -16036
rect 24766 -16064 24800 -16036
rect 24866 -16064 24900 -16036
rect 24666 -16070 24688 -16064
rect 24688 -16070 24700 -16064
rect 24766 -16070 24778 -16064
rect 24778 -16070 24800 -16064
rect 24866 -16070 24868 -16064
rect 24868 -16070 24900 -16064
rect 24966 -16070 25000 -16036
rect 25066 -16070 25100 -16036
rect 25166 -16064 25200 -16036
rect 25166 -16070 25194 -16064
rect 25194 -16070 25200 -16064
rect 25954 -15558 25976 -15536
rect 25976 -15558 25988 -15536
rect 26054 -15558 26066 -15536
rect 26066 -15558 26088 -15536
rect 26154 -15558 26156 -15536
rect 26156 -15558 26188 -15536
rect 25954 -15570 25988 -15558
rect 26054 -15570 26088 -15558
rect 26154 -15570 26188 -15558
rect 26254 -15570 26288 -15536
rect 26354 -15570 26388 -15536
rect 26454 -15558 26482 -15536
rect 26482 -15558 26488 -15536
rect 26454 -15570 26488 -15558
rect 25954 -15648 25976 -15636
rect 25976 -15648 25988 -15636
rect 26054 -15648 26066 -15636
rect 26066 -15648 26088 -15636
rect 26154 -15648 26156 -15636
rect 26156 -15648 26188 -15636
rect 25954 -15670 25988 -15648
rect 26054 -15670 26088 -15648
rect 26154 -15670 26188 -15648
rect 26254 -15670 26288 -15636
rect 26354 -15670 26388 -15636
rect 26454 -15648 26482 -15636
rect 26482 -15648 26488 -15636
rect 26454 -15670 26488 -15648
rect 25954 -15738 25976 -15736
rect 25976 -15738 25988 -15736
rect 26054 -15738 26066 -15736
rect 26066 -15738 26088 -15736
rect 26154 -15738 26156 -15736
rect 26156 -15738 26188 -15736
rect 25954 -15770 25988 -15738
rect 26054 -15770 26088 -15738
rect 26154 -15770 26188 -15738
rect 26254 -15770 26288 -15736
rect 26354 -15770 26388 -15736
rect 26454 -15738 26482 -15736
rect 26482 -15738 26488 -15736
rect 26454 -15770 26488 -15738
rect 25954 -15870 25988 -15836
rect 26054 -15870 26088 -15836
rect 26154 -15870 26188 -15836
rect 26254 -15870 26288 -15836
rect 26354 -15870 26388 -15836
rect 26454 -15870 26488 -15836
rect 25954 -15970 25988 -15936
rect 26054 -15970 26088 -15936
rect 26154 -15970 26188 -15936
rect 26254 -15970 26288 -15936
rect 26354 -15970 26388 -15936
rect 26454 -15970 26488 -15936
rect 25954 -16064 25988 -16036
rect 26054 -16064 26088 -16036
rect 26154 -16064 26188 -16036
rect 25954 -16070 25976 -16064
rect 25976 -16070 25988 -16064
rect 26054 -16070 26066 -16064
rect 26066 -16070 26088 -16064
rect 26154 -16070 26156 -16064
rect 26156 -16070 26188 -16064
rect 26254 -16070 26288 -16036
rect 26354 -16070 26388 -16036
rect 26454 -16064 26488 -16036
rect 26454 -16070 26482 -16064
rect 26482 -16070 26488 -16064
rect 6888 -17834 7285 -17296
rect 13623 -17834 14020 -17296
rect 16938 -16846 16960 -16824
rect 16960 -16846 16972 -16824
rect 17038 -16846 17050 -16824
rect 17050 -16846 17072 -16824
rect 17138 -16846 17140 -16824
rect 17140 -16846 17172 -16824
rect 16938 -16858 16972 -16846
rect 17038 -16858 17072 -16846
rect 17138 -16858 17172 -16846
rect 17238 -16858 17272 -16824
rect 17338 -16858 17372 -16824
rect 17438 -16846 17466 -16824
rect 17466 -16846 17472 -16824
rect 17438 -16858 17472 -16846
rect 16938 -16936 16960 -16924
rect 16960 -16936 16972 -16924
rect 17038 -16936 17050 -16924
rect 17050 -16936 17072 -16924
rect 17138 -16936 17140 -16924
rect 17140 -16936 17172 -16924
rect 16938 -16958 16972 -16936
rect 17038 -16958 17072 -16936
rect 17138 -16958 17172 -16936
rect 17238 -16958 17272 -16924
rect 17338 -16958 17372 -16924
rect 17438 -16936 17466 -16924
rect 17466 -16936 17472 -16924
rect 17438 -16958 17472 -16936
rect 16938 -17026 16960 -17024
rect 16960 -17026 16972 -17024
rect 17038 -17026 17050 -17024
rect 17050 -17026 17072 -17024
rect 17138 -17026 17140 -17024
rect 17140 -17026 17172 -17024
rect 16938 -17058 16972 -17026
rect 17038 -17058 17072 -17026
rect 17138 -17058 17172 -17026
rect 17238 -17058 17272 -17024
rect 17338 -17058 17372 -17024
rect 17438 -17026 17466 -17024
rect 17466 -17026 17472 -17024
rect 17438 -17058 17472 -17026
rect 16938 -17158 16972 -17124
rect 17038 -17158 17072 -17124
rect 17138 -17158 17172 -17124
rect 17238 -17158 17272 -17124
rect 17338 -17158 17372 -17124
rect 17438 -17158 17472 -17124
rect 16938 -17258 16972 -17224
rect 17038 -17258 17072 -17224
rect 17138 -17258 17172 -17224
rect 17238 -17258 17272 -17224
rect 17338 -17258 17372 -17224
rect 17438 -17258 17472 -17224
rect 16938 -17352 16972 -17324
rect 17038 -17352 17072 -17324
rect 17138 -17352 17172 -17324
rect 16938 -17358 16960 -17352
rect 16960 -17358 16972 -17352
rect 17038 -17358 17050 -17352
rect 17050 -17358 17072 -17352
rect 17138 -17358 17140 -17352
rect 17140 -17358 17172 -17352
rect 17238 -17358 17272 -17324
rect 17338 -17358 17372 -17324
rect 17438 -17352 17472 -17324
rect 17438 -17358 17466 -17352
rect 17466 -17358 17472 -17352
rect 18226 -16846 18248 -16824
rect 18248 -16846 18260 -16824
rect 18326 -16846 18338 -16824
rect 18338 -16846 18360 -16824
rect 18426 -16846 18428 -16824
rect 18428 -16846 18460 -16824
rect 18226 -16858 18260 -16846
rect 18326 -16858 18360 -16846
rect 18426 -16858 18460 -16846
rect 18526 -16858 18560 -16824
rect 18626 -16858 18660 -16824
rect 18726 -16846 18754 -16824
rect 18754 -16846 18760 -16824
rect 18726 -16858 18760 -16846
rect 18226 -16936 18248 -16924
rect 18248 -16936 18260 -16924
rect 18326 -16936 18338 -16924
rect 18338 -16936 18360 -16924
rect 18426 -16936 18428 -16924
rect 18428 -16936 18460 -16924
rect 18226 -16958 18260 -16936
rect 18326 -16958 18360 -16936
rect 18426 -16958 18460 -16936
rect 18526 -16958 18560 -16924
rect 18626 -16958 18660 -16924
rect 18726 -16936 18754 -16924
rect 18754 -16936 18760 -16924
rect 18726 -16958 18760 -16936
rect 18226 -17026 18248 -17024
rect 18248 -17026 18260 -17024
rect 18326 -17026 18338 -17024
rect 18338 -17026 18360 -17024
rect 18426 -17026 18428 -17024
rect 18428 -17026 18460 -17024
rect 18226 -17058 18260 -17026
rect 18326 -17058 18360 -17026
rect 18426 -17058 18460 -17026
rect 18526 -17058 18560 -17024
rect 18626 -17058 18660 -17024
rect 18726 -17026 18754 -17024
rect 18754 -17026 18760 -17024
rect 18726 -17058 18760 -17026
rect 18226 -17158 18260 -17124
rect 18326 -17158 18360 -17124
rect 18426 -17158 18460 -17124
rect 18526 -17158 18560 -17124
rect 18626 -17158 18660 -17124
rect 18726 -17158 18760 -17124
rect 18226 -17258 18260 -17224
rect 18326 -17258 18360 -17224
rect 18426 -17258 18460 -17224
rect 18526 -17258 18560 -17224
rect 18626 -17258 18660 -17224
rect 18726 -17258 18760 -17224
rect 18226 -17352 18260 -17324
rect 18326 -17352 18360 -17324
rect 18426 -17352 18460 -17324
rect 18226 -17358 18248 -17352
rect 18248 -17358 18260 -17352
rect 18326 -17358 18338 -17352
rect 18338 -17358 18360 -17352
rect 18426 -17358 18428 -17352
rect 18428 -17358 18460 -17352
rect 18526 -17358 18560 -17324
rect 18626 -17358 18660 -17324
rect 18726 -17352 18760 -17324
rect 18726 -17358 18754 -17352
rect 18754 -17358 18760 -17352
rect 19514 -16846 19536 -16824
rect 19536 -16846 19548 -16824
rect 19614 -16846 19626 -16824
rect 19626 -16846 19648 -16824
rect 19714 -16846 19716 -16824
rect 19716 -16846 19748 -16824
rect 19514 -16858 19548 -16846
rect 19614 -16858 19648 -16846
rect 19714 -16858 19748 -16846
rect 19814 -16858 19848 -16824
rect 19914 -16858 19948 -16824
rect 20014 -16846 20042 -16824
rect 20042 -16846 20048 -16824
rect 20014 -16858 20048 -16846
rect 19514 -16936 19536 -16924
rect 19536 -16936 19548 -16924
rect 19614 -16936 19626 -16924
rect 19626 -16936 19648 -16924
rect 19714 -16936 19716 -16924
rect 19716 -16936 19748 -16924
rect 19514 -16958 19548 -16936
rect 19614 -16958 19648 -16936
rect 19714 -16958 19748 -16936
rect 19814 -16958 19848 -16924
rect 19914 -16958 19948 -16924
rect 20014 -16936 20042 -16924
rect 20042 -16936 20048 -16924
rect 20014 -16958 20048 -16936
rect 19514 -17026 19536 -17024
rect 19536 -17026 19548 -17024
rect 19614 -17026 19626 -17024
rect 19626 -17026 19648 -17024
rect 19714 -17026 19716 -17024
rect 19716 -17026 19748 -17024
rect 19514 -17058 19548 -17026
rect 19614 -17058 19648 -17026
rect 19714 -17058 19748 -17026
rect 19814 -17058 19848 -17024
rect 19914 -17058 19948 -17024
rect 20014 -17026 20042 -17024
rect 20042 -17026 20048 -17024
rect 20014 -17058 20048 -17026
rect 19514 -17158 19548 -17124
rect 19614 -17158 19648 -17124
rect 19714 -17158 19748 -17124
rect 19814 -17158 19848 -17124
rect 19914 -17158 19948 -17124
rect 20014 -17158 20048 -17124
rect 19514 -17258 19548 -17224
rect 19614 -17258 19648 -17224
rect 19714 -17258 19748 -17224
rect 19814 -17258 19848 -17224
rect 19914 -17258 19948 -17224
rect 20014 -17258 20048 -17224
rect 19514 -17352 19548 -17324
rect 19614 -17352 19648 -17324
rect 19714 -17352 19748 -17324
rect 19514 -17358 19536 -17352
rect 19536 -17358 19548 -17352
rect 19614 -17358 19626 -17352
rect 19626 -17358 19648 -17352
rect 19714 -17358 19716 -17352
rect 19716 -17358 19748 -17352
rect 19814 -17358 19848 -17324
rect 19914 -17358 19948 -17324
rect 20014 -17352 20048 -17324
rect 20014 -17358 20042 -17352
rect 20042 -17358 20048 -17352
rect 20802 -16846 20824 -16824
rect 20824 -16846 20836 -16824
rect 20902 -16846 20914 -16824
rect 20914 -16846 20936 -16824
rect 21002 -16846 21004 -16824
rect 21004 -16846 21036 -16824
rect 20802 -16858 20836 -16846
rect 20902 -16858 20936 -16846
rect 21002 -16858 21036 -16846
rect 21102 -16858 21136 -16824
rect 21202 -16858 21236 -16824
rect 21302 -16846 21330 -16824
rect 21330 -16846 21336 -16824
rect 21302 -16858 21336 -16846
rect 20802 -16936 20824 -16924
rect 20824 -16936 20836 -16924
rect 20902 -16936 20914 -16924
rect 20914 -16936 20936 -16924
rect 21002 -16936 21004 -16924
rect 21004 -16936 21036 -16924
rect 20802 -16958 20836 -16936
rect 20902 -16958 20936 -16936
rect 21002 -16958 21036 -16936
rect 21102 -16958 21136 -16924
rect 21202 -16958 21236 -16924
rect 21302 -16936 21330 -16924
rect 21330 -16936 21336 -16924
rect 21302 -16958 21336 -16936
rect 20802 -17026 20824 -17024
rect 20824 -17026 20836 -17024
rect 20902 -17026 20914 -17024
rect 20914 -17026 20936 -17024
rect 21002 -17026 21004 -17024
rect 21004 -17026 21036 -17024
rect 20802 -17058 20836 -17026
rect 20902 -17058 20936 -17026
rect 21002 -17058 21036 -17026
rect 21102 -17058 21136 -17024
rect 21202 -17058 21236 -17024
rect 21302 -17026 21330 -17024
rect 21330 -17026 21336 -17024
rect 21302 -17058 21336 -17026
rect 20802 -17158 20836 -17124
rect 20902 -17158 20936 -17124
rect 21002 -17158 21036 -17124
rect 21102 -17158 21136 -17124
rect 21202 -17158 21236 -17124
rect 21302 -17158 21336 -17124
rect 20802 -17258 20836 -17224
rect 20902 -17258 20936 -17224
rect 21002 -17258 21036 -17224
rect 21102 -17258 21136 -17224
rect 21202 -17258 21236 -17224
rect 21302 -17258 21336 -17224
rect 20802 -17352 20836 -17324
rect 20902 -17352 20936 -17324
rect 21002 -17352 21036 -17324
rect 20802 -17358 20824 -17352
rect 20824 -17358 20836 -17352
rect 20902 -17358 20914 -17352
rect 20914 -17358 20936 -17352
rect 21002 -17358 21004 -17352
rect 21004 -17358 21036 -17352
rect 21102 -17358 21136 -17324
rect 21202 -17358 21236 -17324
rect 21302 -17352 21336 -17324
rect 21302 -17358 21330 -17352
rect 21330 -17358 21336 -17352
rect 22090 -16846 22112 -16824
rect 22112 -16846 22124 -16824
rect 22190 -16846 22202 -16824
rect 22202 -16846 22224 -16824
rect 22290 -16846 22292 -16824
rect 22292 -16846 22324 -16824
rect 22090 -16858 22124 -16846
rect 22190 -16858 22224 -16846
rect 22290 -16858 22324 -16846
rect 22390 -16858 22424 -16824
rect 22490 -16858 22524 -16824
rect 22590 -16846 22618 -16824
rect 22618 -16846 22624 -16824
rect 22590 -16858 22624 -16846
rect 22090 -16936 22112 -16924
rect 22112 -16936 22124 -16924
rect 22190 -16936 22202 -16924
rect 22202 -16936 22224 -16924
rect 22290 -16936 22292 -16924
rect 22292 -16936 22324 -16924
rect 22090 -16958 22124 -16936
rect 22190 -16958 22224 -16936
rect 22290 -16958 22324 -16936
rect 22390 -16958 22424 -16924
rect 22490 -16958 22524 -16924
rect 22590 -16936 22618 -16924
rect 22618 -16936 22624 -16924
rect 22590 -16958 22624 -16936
rect 22090 -17026 22112 -17024
rect 22112 -17026 22124 -17024
rect 22190 -17026 22202 -17024
rect 22202 -17026 22224 -17024
rect 22290 -17026 22292 -17024
rect 22292 -17026 22324 -17024
rect 22090 -17058 22124 -17026
rect 22190 -17058 22224 -17026
rect 22290 -17058 22324 -17026
rect 22390 -17058 22424 -17024
rect 22490 -17058 22524 -17024
rect 22590 -17026 22618 -17024
rect 22618 -17026 22624 -17024
rect 22590 -17058 22624 -17026
rect 22090 -17158 22124 -17124
rect 22190 -17158 22224 -17124
rect 22290 -17158 22324 -17124
rect 22390 -17158 22424 -17124
rect 22490 -17158 22524 -17124
rect 22590 -17158 22624 -17124
rect 22090 -17258 22124 -17224
rect 22190 -17258 22224 -17224
rect 22290 -17258 22324 -17224
rect 22390 -17258 22424 -17224
rect 22490 -17258 22524 -17224
rect 22590 -17258 22624 -17224
rect 22090 -17352 22124 -17324
rect 22190 -17352 22224 -17324
rect 22290 -17352 22324 -17324
rect 22090 -17358 22112 -17352
rect 22112 -17358 22124 -17352
rect 22190 -17358 22202 -17352
rect 22202 -17358 22224 -17352
rect 22290 -17358 22292 -17352
rect 22292 -17358 22324 -17352
rect 22390 -17358 22424 -17324
rect 22490 -17358 22524 -17324
rect 22590 -17352 22624 -17324
rect 22590 -17358 22618 -17352
rect 22618 -17358 22624 -17352
rect 23378 -16846 23400 -16824
rect 23400 -16846 23412 -16824
rect 23478 -16846 23490 -16824
rect 23490 -16846 23512 -16824
rect 23578 -16846 23580 -16824
rect 23580 -16846 23612 -16824
rect 23378 -16858 23412 -16846
rect 23478 -16858 23512 -16846
rect 23578 -16858 23612 -16846
rect 23678 -16858 23712 -16824
rect 23778 -16858 23812 -16824
rect 23878 -16846 23906 -16824
rect 23906 -16846 23912 -16824
rect 23878 -16858 23912 -16846
rect 23378 -16936 23400 -16924
rect 23400 -16936 23412 -16924
rect 23478 -16936 23490 -16924
rect 23490 -16936 23512 -16924
rect 23578 -16936 23580 -16924
rect 23580 -16936 23612 -16924
rect 23378 -16958 23412 -16936
rect 23478 -16958 23512 -16936
rect 23578 -16958 23612 -16936
rect 23678 -16958 23712 -16924
rect 23778 -16958 23812 -16924
rect 23878 -16936 23906 -16924
rect 23906 -16936 23912 -16924
rect 23878 -16958 23912 -16936
rect 23378 -17026 23400 -17024
rect 23400 -17026 23412 -17024
rect 23478 -17026 23490 -17024
rect 23490 -17026 23512 -17024
rect 23578 -17026 23580 -17024
rect 23580 -17026 23612 -17024
rect 23378 -17058 23412 -17026
rect 23478 -17058 23512 -17026
rect 23578 -17058 23612 -17026
rect 23678 -17058 23712 -17024
rect 23778 -17058 23812 -17024
rect 23878 -17026 23906 -17024
rect 23906 -17026 23912 -17024
rect 23878 -17058 23912 -17026
rect 23378 -17158 23412 -17124
rect 23478 -17158 23512 -17124
rect 23578 -17158 23612 -17124
rect 23678 -17158 23712 -17124
rect 23778 -17158 23812 -17124
rect 23878 -17158 23912 -17124
rect 23378 -17258 23412 -17224
rect 23478 -17258 23512 -17224
rect 23578 -17258 23612 -17224
rect 23678 -17258 23712 -17224
rect 23778 -17258 23812 -17224
rect 23878 -17258 23912 -17224
rect 23378 -17352 23412 -17324
rect 23478 -17352 23512 -17324
rect 23578 -17352 23612 -17324
rect 23378 -17358 23400 -17352
rect 23400 -17358 23412 -17352
rect 23478 -17358 23490 -17352
rect 23490 -17358 23512 -17352
rect 23578 -17358 23580 -17352
rect 23580 -17358 23612 -17352
rect 23678 -17358 23712 -17324
rect 23778 -17358 23812 -17324
rect 23878 -17352 23912 -17324
rect 23878 -17358 23906 -17352
rect 23906 -17358 23912 -17352
rect 24666 -16846 24688 -16824
rect 24688 -16846 24700 -16824
rect 24766 -16846 24778 -16824
rect 24778 -16846 24800 -16824
rect 24866 -16846 24868 -16824
rect 24868 -16846 24900 -16824
rect 24666 -16858 24700 -16846
rect 24766 -16858 24800 -16846
rect 24866 -16858 24900 -16846
rect 24966 -16858 25000 -16824
rect 25066 -16858 25100 -16824
rect 25166 -16846 25194 -16824
rect 25194 -16846 25200 -16824
rect 25166 -16858 25200 -16846
rect 24666 -16936 24688 -16924
rect 24688 -16936 24700 -16924
rect 24766 -16936 24778 -16924
rect 24778 -16936 24800 -16924
rect 24866 -16936 24868 -16924
rect 24868 -16936 24900 -16924
rect 24666 -16958 24700 -16936
rect 24766 -16958 24800 -16936
rect 24866 -16958 24900 -16936
rect 24966 -16958 25000 -16924
rect 25066 -16958 25100 -16924
rect 25166 -16936 25194 -16924
rect 25194 -16936 25200 -16924
rect 25166 -16958 25200 -16936
rect 24666 -17026 24688 -17024
rect 24688 -17026 24700 -17024
rect 24766 -17026 24778 -17024
rect 24778 -17026 24800 -17024
rect 24866 -17026 24868 -17024
rect 24868 -17026 24900 -17024
rect 24666 -17058 24700 -17026
rect 24766 -17058 24800 -17026
rect 24866 -17058 24900 -17026
rect 24966 -17058 25000 -17024
rect 25066 -17058 25100 -17024
rect 25166 -17026 25194 -17024
rect 25194 -17026 25200 -17024
rect 25166 -17058 25200 -17026
rect 24666 -17158 24700 -17124
rect 24766 -17158 24800 -17124
rect 24866 -17158 24900 -17124
rect 24966 -17158 25000 -17124
rect 25066 -17158 25100 -17124
rect 25166 -17158 25200 -17124
rect 24666 -17258 24700 -17224
rect 24766 -17258 24800 -17224
rect 24866 -17258 24900 -17224
rect 24966 -17258 25000 -17224
rect 25066 -17258 25100 -17224
rect 25166 -17258 25200 -17224
rect 24666 -17352 24700 -17324
rect 24766 -17352 24800 -17324
rect 24866 -17352 24900 -17324
rect 24666 -17358 24688 -17352
rect 24688 -17358 24700 -17352
rect 24766 -17358 24778 -17352
rect 24778 -17358 24800 -17352
rect 24866 -17358 24868 -17352
rect 24868 -17358 24900 -17352
rect 24966 -17358 25000 -17324
rect 25066 -17358 25100 -17324
rect 25166 -17352 25200 -17324
rect 25166 -17358 25194 -17352
rect 25194 -17358 25200 -17352
rect 25954 -16846 25976 -16823
rect 25976 -16846 25988 -16823
rect 26054 -16846 26066 -16823
rect 26066 -16846 26088 -16823
rect 26154 -16846 26156 -16823
rect 26156 -16846 26188 -16823
rect 25954 -16858 25988 -16846
rect 26054 -16858 26088 -16846
rect 26154 -16858 26188 -16846
rect 26254 -16858 26288 -16823
rect 26354 -16858 26388 -16823
rect 26454 -16846 26482 -16823
rect 26482 -16846 26488 -16823
rect 26454 -16858 26488 -16846
rect 25954 -16936 25976 -16923
rect 25976 -16936 25988 -16923
rect 26054 -16936 26066 -16923
rect 26066 -16936 26088 -16923
rect 26154 -16936 26156 -16923
rect 26156 -16936 26188 -16923
rect 25954 -16958 25988 -16936
rect 26054 -16958 26088 -16936
rect 26154 -16958 26188 -16936
rect 26254 -16958 26288 -16923
rect 26354 -16958 26388 -16923
rect 26454 -16936 26482 -16923
rect 26482 -16936 26488 -16923
rect 26454 -16958 26488 -16936
rect 25954 -17026 25976 -17023
rect 25976 -17026 25988 -17023
rect 26054 -17026 26066 -17023
rect 26066 -17026 26088 -17023
rect 26154 -17026 26156 -17023
rect 26156 -17026 26188 -17023
rect 25954 -17058 25988 -17026
rect 26054 -17058 26088 -17026
rect 26154 -17058 26188 -17026
rect 26254 -17058 26288 -17023
rect 26354 -17058 26388 -17023
rect 26454 -17026 26482 -17023
rect 26482 -17026 26488 -17023
rect 26454 -17058 26488 -17026
rect 25954 -17158 25988 -17123
rect 26054 -17158 26088 -17123
rect 26154 -17158 26188 -17123
rect 26254 -17158 26288 -17123
rect 26354 -17158 26388 -17123
rect 26454 -17158 26488 -17123
rect 25954 -17258 25988 -17223
rect 26054 -17258 26088 -17223
rect 26154 -17258 26188 -17223
rect 26254 -17258 26288 -17223
rect 26354 -17258 26388 -17223
rect 26454 -17258 26488 -17223
rect 25954 -17351 25988 -17323
rect 26054 -17351 26088 -17323
rect 26154 -17351 26188 -17323
rect 25954 -17358 25976 -17351
rect 25976 -17358 25988 -17351
rect 26054 -17358 26066 -17351
rect 26066 -17358 26088 -17351
rect 26154 -17358 26156 -17351
rect 26156 -17358 26188 -17351
rect 26254 -17358 26288 -17323
rect 26354 -17358 26388 -17323
rect 26454 -17351 26488 -17323
rect 26454 -17358 26482 -17351
rect 26482 -17358 26488 -17351
rect 6888 -18652 7285 -18114
rect 13623 -18652 14020 -18114
rect 6888 -19470 7285 -18932
rect 13623 -19470 14020 -18932
rect 6888 -20288 7285 -19750
rect 13623 -20288 14020 -19750
rect 6888 -21106 7285 -20568
rect 13623 -21106 14020 -20568
rect 6888 -21924 7285 -21386
rect 13623 -21924 14021 -21386
rect 6888 -22742 7285 -22204
rect 13623 -22742 14020 -22204
rect 6888 -23560 7285 -23022
rect 13623 -23560 14020 -23022
rect 6888 -24378 7285 -23840
rect 13623 -24378 14020 -23840
rect 6888 -25196 7285 -24658
rect 13623 -25196 14021 -24658
rect 6888 -26014 7285 -25476
rect 13623 -26014 14020 -25476
rect 6888 -26832 7285 -26294
rect 13623 -26832 14020 -26294
rect 6888 -27650 7285 -27112
rect 13623 -27650 14021 -27112
rect 6888 -28468 7285 -27930
rect 13623 -28468 14020 -27930
rect 6888 -29286 7285 -28748
rect 13623 -29286 14020 -28748
rect 6888 -30104 7285 -29566
rect 13623 -30104 14021 -29566
rect 6888 -30922 7285 -30384
rect 13623 -30922 14020 -30384
rect 11570 -31694 12622 -31182
rect 6826 -33376 7223 -32838
rect 11557 -33376 11954 -32838
rect 6826 -34194 7223 -33656
rect 11557 -34194 11954 -33656
rect 6826 -35012 7223 -34474
rect 11557 -35012 11954 -34474
rect 6826 -35830 7223 -35292
rect 11557 -35830 11954 -35292
rect 11568 -36646 12634 -36152
rect 8212 -37466 8609 -36928
rect 11967 -37466 12364 -36928
rect 8212 -38284 8609 -37746
rect 11967 -38284 12364 -37746
rect 8212 -39102 8609 -38564
rect 11967 -39102 12364 -38564
<< metal1 >>
rect 16884 -11672 26584 -11602
rect 16884 -11706 16938 -11672
rect 16972 -11706 17038 -11672
rect 17072 -11706 17138 -11672
rect 17172 -11706 17238 -11672
rect 17272 -11706 17338 -11672
rect 17372 -11706 17438 -11672
rect 17472 -11706 18226 -11672
rect 18260 -11706 18326 -11672
rect 18360 -11706 18426 -11672
rect 18460 -11706 18526 -11672
rect 18560 -11706 18626 -11672
rect 18660 -11706 18726 -11672
rect 18760 -11706 19514 -11672
rect 19548 -11706 19614 -11672
rect 19648 -11706 19714 -11672
rect 19748 -11706 19814 -11672
rect 19848 -11706 19914 -11672
rect 19948 -11706 20014 -11672
rect 20048 -11706 20802 -11672
rect 20836 -11706 20902 -11672
rect 20936 -11706 21002 -11672
rect 21036 -11706 21102 -11672
rect 21136 -11706 21202 -11672
rect 21236 -11706 21302 -11672
rect 21336 -11706 22090 -11672
rect 22124 -11706 22190 -11672
rect 22224 -11706 22290 -11672
rect 22324 -11706 22390 -11672
rect 22424 -11706 22490 -11672
rect 22524 -11706 22590 -11672
rect 22624 -11706 23378 -11672
rect 23412 -11706 23478 -11672
rect 23512 -11706 23578 -11672
rect 23612 -11706 23678 -11672
rect 23712 -11706 23778 -11672
rect 23812 -11706 23878 -11672
rect 23912 -11706 24666 -11672
rect 24700 -11706 24766 -11672
rect 24800 -11706 24866 -11672
rect 24900 -11706 24966 -11672
rect 25000 -11706 25066 -11672
rect 25100 -11706 25166 -11672
rect 25200 -11706 25954 -11672
rect 25988 -11706 26054 -11672
rect 26088 -11706 26154 -11672
rect 26188 -11706 26254 -11672
rect 26288 -11706 26354 -11672
rect 26388 -11706 26454 -11672
rect 26488 -11706 26584 -11672
rect 16884 -11772 26584 -11706
rect 16884 -11806 16938 -11772
rect 16972 -11806 17038 -11772
rect 17072 -11806 17138 -11772
rect 17172 -11806 17238 -11772
rect 17272 -11806 17338 -11772
rect 17372 -11806 17438 -11772
rect 17472 -11806 18226 -11772
rect 18260 -11806 18326 -11772
rect 18360 -11806 18426 -11772
rect 18460 -11806 18526 -11772
rect 18560 -11806 18626 -11772
rect 18660 -11806 18726 -11772
rect 18760 -11806 19514 -11772
rect 19548 -11806 19614 -11772
rect 19648 -11806 19714 -11772
rect 19748 -11806 19814 -11772
rect 19848 -11806 19914 -11772
rect 19948 -11806 20014 -11772
rect 20048 -11806 20802 -11772
rect 20836 -11806 20902 -11772
rect 20936 -11806 21002 -11772
rect 21036 -11806 21102 -11772
rect 21136 -11806 21202 -11772
rect 21236 -11806 21302 -11772
rect 21336 -11806 22090 -11772
rect 22124 -11806 22190 -11772
rect 22224 -11806 22290 -11772
rect 22324 -11806 22390 -11772
rect 22424 -11806 22490 -11772
rect 22524 -11806 22590 -11772
rect 22624 -11806 23378 -11772
rect 23412 -11806 23478 -11772
rect 23512 -11806 23578 -11772
rect 23612 -11806 23678 -11772
rect 23712 -11806 23778 -11772
rect 23812 -11806 23878 -11772
rect 23912 -11806 24666 -11772
rect 24700 -11806 24766 -11772
rect 24800 -11806 24866 -11772
rect 24900 -11806 24966 -11772
rect 25000 -11806 25066 -11772
rect 25100 -11806 25166 -11772
rect 25200 -11806 25954 -11772
rect 25988 -11806 26054 -11772
rect 26088 -11806 26154 -11772
rect 26188 -11806 26254 -11772
rect 26288 -11806 26354 -11772
rect 26388 -11806 26454 -11772
rect 26488 -11806 26584 -11772
rect 16884 -11872 26584 -11806
rect 16884 -11906 16938 -11872
rect 16972 -11906 17038 -11872
rect 17072 -11906 17138 -11872
rect 17172 -11906 17238 -11872
rect 17272 -11906 17338 -11872
rect 17372 -11906 17438 -11872
rect 17472 -11906 18226 -11872
rect 18260 -11906 18326 -11872
rect 18360 -11906 18426 -11872
rect 18460 -11906 18526 -11872
rect 18560 -11906 18626 -11872
rect 18660 -11906 18726 -11872
rect 18760 -11906 19514 -11872
rect 19548 -11906 19614 -11872
rect 19648 -11906 19714 -11872
rect 19748 -11906 19814 -11872
rect 19848 -11906 19914 -11872
rect 19948 -11906 20014 -11872
rect 20048 -11906 20802 -11872
rect 20836 -11906 20902 -11872
rect 20936 -11906 21002 -11872
rect 21036 -11906 21102 -11872
rect 21136 -11906 21202 -11872
rect 21236 -11906 21302 -11872
rect 21336 -11906 22090 -11872
rect 22124 -11906 22190 -11872
rect 22224 -11906 22290 -11872
rect 22324 -11906 22390 -11872
rect 22424 -11906 22490 -11872
rect 22524 -11906 22590 -11872
rect 22624 -11906 23378 -11872
rect 23412 -11906 23478 -11872
rect 23512 -11906 23578 -11872
rect 23612 -11906 23678 -11872
rect 23712 -11906 23778 -11872
rect 23812 -11906 23878 -11872
rect 23912 -11906 24666 -11872
rect 24700 -11906 24766 -11872
rect 24800 -11906 24866 -11872
rect 24900 -11906 24966 -11872
rect 25000 -11906 25066 -11872
rect 25100 -11906 25166 -11872
rect 25200 -11906 25954 -11872
rect 25988 -11906 26054 -11872
rect 26088 -11906 26154 -11872
rect 26188 -11906 26254 -11872
rect 26288 -11906 26354 -11872
rect 26388 -11906 26454 -11872
rect 26488 -11906 26584 -11872
rect 16884 -11972 26584 -11906
rect 16884 -12006 16938 -11972
rect 16972 -12006 17038 -11972
rect 17072 -12006 17138 -11972
rect 17172 -12006 17238 -11972
rect 17272 -12006 17338 -11972
rect 17372 -12006 17438 -11972
rect 17472 -12006 18226 -11972
rect 18260 -12006 18326 -11972
rect 18360 -12006 18426 -11972
rect 18460 -12006 18526 -11972
rect 18560 -12006 18626 -11972
rect 18660 -12006 18726 -11972
rect 18760 -12006 19514 -11972
rect 19548 -12006 19614 -11972
rect 19648 -12006 19714 -11972
rect 19748 -12006 19814 -11972
rect 19848 -12006 19914 -11972
rect 19948 -12006 20014 -11972
rect 20048 -12006 20802 -11972
rect 20836 -12006 20902 -11972
rect 20936 -12006 21002 -11972
rect 21036 -12006 21102 -11972
rect 21136 -12006 21202 -11972
rect 21236 -12006 21302 -11972
rect 21336 -12006 22090 -11972
rect 22124 -12006 22190 -11972
rect 22224 -12006 22290 -11972
rect 22324 -12006 22390 -11972
rect 22424 -12006 22490 -11972
rect 22524 -12006 22590 -11972
rect 22624 -12006 23378 -11972
rect 23412 -12006 23478 -11972
rect 23512 -12006 23578 -11972
rect 23612 -12006 23678 -11972
rect 23712 -12006 23778 -11972
rect 23812 -12006 23878 -11972
rect 23912 -12006 24666 -11972
rect 24700 -12006 24766 -11972
rect 24800 -12006 24866 -11972
rect 24900 -12006 24966 -11972
rect 25000 -12006 25066 -11972
rect 25100 -12006 25166 -11972
rect 25200 -12006 25954 -11972
rect 25988 -12006 26054 -11972
rect 26088 -12006 26154 -11972
rect 26188 -12006 26254 -11972
rect 26288 -12006 26354 -11972
rect 26388 -12006 26454 -11972
rect 26488 -12006 26584 -11972
rect 16884 -12072 26584 -12006
rect 16884 -12106 16938 -12072
rect 16972 -12106 17038 -12072
rect 17072 -12106 17138 -12072
rect 17172 -12106 17238 -12072
rect 17272 -12106 17338 -12072
rect 17372 -12106 17438 -12072
rect 17472 -12106 18226 -12072
rect 18260 -12106 18326 -12072
rect 18360 -12106 18426 -12072
rect 18460 -12106 18526 -12072
rect 18560 -12106 18626 -12072
rect 18660 -12106 18726 -12072
rect 18760 -12106 19514 -12072
rect 19548 -12106 19614 -12072
rect 19648 -12106 19714 -12072
rect 19748 -12106 19814 -12072
rect 19848 -12106 19914 -12072
rect 19948 -12106 20014 -12072
rect 20048 -12106 20802 -12072
rect 20836 -12106 20902 -12072
rect 20936 -12106 21002 -12072
rect 21036 -12106 21102 -12072
rect 21136 -12106 21202 -12072
rect 21236 -12106 21302 -12072
rect 21336 -12106 22090 -12072
rect 22124 -12106 22190 -12072
rect 22224 -12106 22290 -12072
rect 22324 -12106 22390 -12072
rect 22424 -12106 22490 -12072
rect 22524 -12106 22590 -12072
rect 22624 -12106 23378 -12072
rect 23412 -12106 23478 -12072
rect 23512 -12106 23578 -12072
rect 23612 -12106 23678 -12072
rect 23712 -12106 23778 -12072
rect 23812 -12106 23878 -12072
rect 23912 -12106 24666 -12072
rect 24700 -12106 24766 -12072
rect 24800 -12106 24866 -12072
rect 24900 -12106 24966 -12072
rect 25000 -12106 25066 -12072
rect 25100 -12106 25166 -12072
rect 25200 -12106 25954 -12072
rect 25988 -12106 26054 -12072
rect 26088 -12106 26154 -12072
rect 26188 -12106 26254 -12072
rect 26288 -12106 26354 -12072
rect 26388 -12106 26454 -12072
rect 26488 -12106 26584 -12072
rect 16884 -12172 26584 -12106
rect 16884 -12206 16938 -12172
rect 16972 -12206 17038 -12172
rect 17072 -12206 17138 -12172
rect 17172 -12206 17238 -12172
rect 17272 -12206 17338 -12172
rect 17372 -12206 17438 -12172
rect 17472 -12206 18226 -12172
rect 18260 -12206 18326 -12172
rect 18360 -12206 18426 -12172
rect 18460 -12206 18526 -12172
rect 18560 -12206 18626 -12172
rect 18660 -12206 18726 -12172
rect 18760 -12206 19514 -12172
rect 19548 -12206 19614 -12172
rect 19648 -12206 19714 -12172
rect 19748 -12206 19814 -12172
rect 19848 -12206 19914 -12172
rect 19948 -12206 20014 -12172
rect 20048 -12206 20802 -12172
rect 20836 -12206 20902 -12172
rect 20936 -12206 21002 -12172
rect 21036 -12206 21102 -12172
rect 21136 -12206 21202 -12172
rect 21236 -12206 21302 -12172
rect 21336 -12206 22090 -12172
rect 22124 -12206 22190 -12172
rect 22224 -12206 22290 -12172
rect 22324 -12206 22390 -12172
rect 22424 -12206 22490 -12172
rect 22524 -12206 22590 -12172
rect 22624 -12206 23378 -12172
rect 23412 -12206 23478 -12172
rect 23512 -12206 23578 -12172
rect 23612 -12206 23678 -12172
rect 23712 -12206 23778 -12172
rect 23812 -12206 23878 -12172
rect 23912 -12206 24666 -12172
rect 24700 -12206 24766 -12172
rect 24800 -12206 24866 -12172
rect 24900 -12206 24966 -12172
rect 25000 -12206 25066 -12172
rect 25100 -12206 25166 -12172
rect 25200 -12206 25954 -12172
rect 25988 -12206 26054 -12172
rect 26088 -12206 26154 -12172
rect 26188 -12206 26254 -12172
rect 26288 -12206 26354 -12172
rect 26388 -12206 26454 -12172
rect 26488 -12206 26584 -12172
rect 16884 -12960 26584 -12206
rect 16884 -12994 16938 -12960
rect 16972 -12994 17038 -12960
rect 17072 -12994 17138 -12960
rect 17172 -12994 17238 -12960
rect 17272 -12994 17338 -12960
rect 17372 -12994 17438 -12960
rect 17472 -12994 18226 -12960
rect 18260 -12994 18326 -12960
rect 18360 -12994 18426 -12960
rect 18460 -12994 18526 -12960
rect 18560 -12994 18626 -12960
rect 18660 -12994 18726 -12960
rect 18760 -12994 19514 -12960
rect 19548 -12994 19614 -12960
rect 19648 -12994 19714 -12960
rect 19748 -12994 19814 -12960
rect 19848 -12994 19914 -12960
rect 19948 -12994 20014 -12960
rect 20048 -12994 20802 -12960
rect 20836 -12994 20902 -12960
rect 20936 -12994 21002 -12960
rect 21036 -12994 21102 -12960
rect 21136 -12994 21202 -12960
rect 21236 -12994 21302 -12960
rect 21336 -12994 22090 -12960
rect 22124 -12994 22190 -12960
rect 22224 -12994 22290 -12960
rect 22324 -12994 22390 -12960
rect 22424 -12994 22490 -12960
rect 22524 -12994 22590 -12960
rect 22624 -12994 23378 -12960
rect 23412 -12994 23478 -12960
rect 23512 -12994 23578 -12960
rect 23612 -12994 23678 -12960
rect 23712 -12994 23778 -12960
rect 23812 -12994 23878 -12960
rect 23912 -12994 24666 -12960
rect 24700 -12994 24766 -12960
rect 24800 -12994 24866 -12960
rect 24900 -12994 24966 -12960
rect 25000 -12994 25066 -12960
rect 25100 -12994 25166 -12960
rect 25200 -12994 25954 -12960
rect 25988 -12994 26054 -12960
rect 26088 -12994 26154 -12960
rect 26188 -12994 26254 -12960
rect 26288 -12994 26354 -12960
rect 26388 -12994 26454 -12960
rect 26488 -12994 26584 -12960
rect 16884 -13060 26584 -12994
rect 16884 -13094 16938 -13060
rect 16972 -13094 17038 -13060
rect 17072 -13094 17138 -13060
rect 17172 -13094 17238 -13060
rect 17272 -13094 17338 -13060
rect 17372 -13094 17438 -13060
rect 17472 -13094 18226 -13060
rect 18260 -13094 18326 -13060
rect 18360 -13094 18426 -13060
rect 18460 -13094 18526 -13060
rect 18560 -13094 18626 -13060
rect 18660 -13094 18726 -13060
rect 18760 -13094 19514 -13060
rect 19548 -13094 19614 -13060
rect 19648 -13094 19714 -13060
rect 19748 -13094 19814 -13060
rect 19848 -13094 19914 -13060
rect 19948 -13094 20014 -13060
rect 20048 -13094 20802 -13060
rect 20836 -13094 20902 -13060
rect 20936 -13094 21002 -13060
rect 21036 -13094 21102 -13060
rect 21136 -13094 21202 -13060
rect 21236 -13094 21302 -13060
rect 21336 -13094 22090 -13060
rect 22124 -13094 22190 -13060
rect 22224 -13094 22290 -13060
rect 22324 -13094 22390 -13060
rect 22424 -13094 22490 -13060
rect 22524 -13094 22590 -13060
rect 22624 -13094 23378 -13060
rect 23412 -13094 23478 -13060
rect 23512 -13094 23578 -13060
rect 23612 -13094 23678 -13060
rect 23712 -13094 23778 -13060
rect 23812 -13094 23878 -13060
rect 23912 -13094 24666 -13060
rect 24700 -13094 24766 -13060
rect 24800 -13094 24866 -13060
rect 24900 -13094 24966 -13060
rect 25000 -13094 25066 -13060
rect 25100 -13094 25166 -13060
rect 25200 -13094 25954 -13060
rect 25988 -13094 26054 -13060
rect 26088 -13094 26154 -13060
rect 26188 -13094 26254 -13060
rect 26288 -13094 26354 -13060
rect 26388 -13094 26454 -13060
rect 26488 -13094 26584 -13060
rect 16884 -13160 26584 -13094
rect 16884 -13194 16938 -13160
rect 16972 -13194 17038 -13160
rect 17072 -13194 17138 -13160
rect 17172 -13194 17238 -13160
rect 17272 -13194 17338 -13160
rect 17372 -13194 17438 -13160
rect 17472 -13194 18226 -13160
rect 18260 -13194 18326 -13160
rect 18360 -13194 18426 -13160
rect 18460 -13194 18526 -13160
rect 18560 -13194 18626 -13160
rect 18660 -13194 18726 -13160
rect 18760 -13194 19514 -13160
rect 19548 -13194 19614 -13160
rect 19648 -13194 19714 -13160
rect 19748 -13194 19814 -13160
rect 19848 -13194 19914 -13160
rect 19948 -13194 20014 -13160
rect 20048 -13194 20802 -13160
rect 20836 -13194 20902 -13160
rect 20936 -13194 21002 -13160
rect 21036 -13194 21102 -13160
rect 21136 -13194 21202 -13160
rect 21236 -13194 21302 -13160
rect 21336 -13194 22090 -13160
rect 22124 -13194 22190 -13160
rect 22224 -13194 22290 -13160
rect 22324 -13194 22390 -13160
rect 22424 -13194 22490 -13160
rect 22524 -13194 22590 -13160
rect 22624 -13194 23378 -13160
rect 23412 -13194 23478 -13160
rect 23512 -13194 23578 -13160
rect 23612 -13194 23678 -13160
rect 23712 -13194 23778 -13160
rect 23812 -13194 23878 -13160
rect 23912 -13194 24666 -13160
rect 24700 -13194 24766 -13160
rect 24800 -13194 24866 -13160
rect 24900 -13194 24966 -13160
rect 25000 -13194 25066 -13160
rect 25100 -13194 25166 -13160
rect 25200 -13194 25954 -13160
rect 25988 -13194 26054 -13160
rect 26088 -13194 26154 -13160
rect 26188 -13194 26254 -13160
rect 26288 -13194 26354 -13160
rect 26388 -13194 26454 -13160
rect 26488 -13194 26584 -13160
rect 16884 -13260 26584 -13194
rect 16884 -13294 16938 -13260
rect 16972 -13294 17038 -13260
rect 17072 -13294 17138 -13260
rect 17172 -13294 17238 -13260
rect 17272 -13294 17338 -13260
rect 17372 -13294 17438 -13260
rect 17472 -13294 18226 -13260
rect 18260 -13294 18326 -13260
rect 18360 -13294 18426 -13260
rect 18460 -13294 18526 -13260
rect 18560 -13294 18626 -13260
rect 18660 -13294 18726 -13260
rect 18760 -13294 19514 -13260
rect 19548 -13294 19614 -13260
rect 19648 -13294 19714 -13260
rect 19748 -13294 19814 -13260
rect 19848 -13294 19914 -13260
rect 19948 -13294 20014 -13260
rect 20048 -13294 20802 -13260
rect 20836 -13294 20902 -13260
rect 20936 -13294 21002 -13260
rect 21036 -13294 21102 -13260
rect 21136 -13294 21202 -13260
rect 21236 -13294 21302 -13260
rect 21336 -13294 22090 -13260
rect 22124 -13294 22190 -13260
rect 22224 -13294 22290 -13260
rect 22324 -13294 22390 -13260
rect 22424 -13294 22490 -13260
rect 22524 -13294 22590 -13260
rect 22624 -13294 23378 -13260
rect 23412 -13294 23478 -13260
rect 23512 -13294 23578 -13260
rect 23612 -13294 23678 -13260
rect 23712 -13294 23778 -13260
rect 23812 -13294 23878 -13260
rect 23912 -13294 24666 -13260
rect 24700 -13294 24766 -13260
rect 24800 -13294 24866 -13260
rect 24900 -13294 24966 -13260
rect 25000 -13294 25066 -13260
rect 25100 -13294 25166 -13260
rect 25200 -13294 25954 -13260
rect 25988 -13294 26054 -13260
rect 26088 -13294 26154 -13260
rect 26188 -13294 26254 -13260
rect 26288 -13294 26354 -13260
rect 26388 -13294 26454 -13260
rect 26488 -13294 26584 -13260
rect 16884 -13360 26584 -13294
rect 16884 -13394 16938 -13360
rect 16972 -13394 17038 -13360
rect 17072 -13394 17138 -13360
rect 17172 -13394 17238 -13360
rect 17272 -13394 17338 -13360
rect 17372 -13394 17438 -13360
rect 17472 -13394 18226 -13360
rect 18260 -13394 18326 -13360
rect 18360 -13394 18426 -13360
rect 18460 -13394 18526 -13360
rect 18560 -13394 18626 -13360
rect 18660 -13394 18726 -13360
rect 18760 -13394 19514 -13360
rect 19548 -13394 19614 -13360
rect 19648 -13394 19714 -13360
rect 19748 -13394 19814 -13360
rect 19848 -13394 19914 -13360
rect 19948 -13394 20014 -13360
rect 20048 -13394 20802 -13360
rect 20836 -13394 20902 -13360
rect 20936 -13394 21002 -13360
rect 21036 -13394 21102 -13360
rect 21136 -13394 21202 -13360
rect 21236 -13394 21302 -13360
rect 21336 -13394 22090 -13360
rect 22124 -13394 22190 -13360
rect 22224 -13394 22290 -13360
rect 22324 -13394 22390 -13360
rect 22424 -13394 22490 -13360
rect 22524 -13394 22590 -13360
rect 22624 -13394 23378 -13360
rect 23412 -13394 23478 -13360
rect 23512 -13394 23578 -13360
rect 23612 -13394 23678 -13360
rect 23712 -13394 23778 -13360
rect 23812 -13394 23878 -13360
rect 23912 -13394 24666 -13360
rect 24700 -13394 24766 -13360
rect 24800 -13394 24866 -13360
rect 24900 -13394 24966 -13360
rect 25000 -13394 25066 -13360
rect 25100 -13394 25166 -13360
rect 25200 -13394 25954 -13360
rect 25988 -13394 26054 -13360
rect 26088 -13394 26154 -13360
rect 26188 -13394 26254 -13360
rect 26288 -13394 26354 -13360
rect 26388 -13394 26454 -13360
rect 26488 -13394 26584 -13360
rect 16884 -13460 26584 -13394
rect 16884 -13494 16938 -13460
rect 16972 -13494 17038 -13460
rect 17072 -13494 17138 -13460
rect 17172 -13494 17238 -13460
rect 17272 -13494 17338 -13460
rect 17372 -13494 17438 -13460
rect 17472 -13494 18226 -13460
rect 18260 -13494 18326 -13460
rect 18360 -13494 18426 -13460
rect 18460 -13494 18526 -13460
rect 18560 -13494 18626 -13460
rect 18660 -13494 18726 -13460
rect 18760 -13494 19514 -13460
rect 19548 -13494 19614 -13460
rect 19648 -13494 19714 -13460
rect 19748 -13494 19814 -13460
rect 19848 -13494 19914 -13460
rect 19948 -13494 20014 -13460
rect 20048 -13494 20802 -13460
rect 20836 -13494 20902 -13460
rect 20936 -13494 21002 -13460
rect 21036 -13494 21102 -13460
rect 21136 -13494 21202 -13460
rect 21236 -13494 21302 -13460
rect 21336 -13494 22090 -13460
rect 22124 -13494 22190 -13460
rect 22224 -13494 22290 -13460
rect 22324 -13494 22390 -13460
rect 22424 -13494 22490 -13460
rect 22524 -13494 22590 -13460
rect 22624 -13494 23378 -13460
rect 23412 -13494 23478 -13460
rect 23512 -13494 23578 -13460
rect 23612 -13494 23678 -13460
rect 23712 -13494 23778 -13460
rect 23812 -13494 23878 -13460
rect 23912 -13494 24666 -13460
rect 24700 -13494 24766 -13460
rect 24800 -13494 24866 -13460
rect 24900 -13494 24966 -13460
rect 25000 -13494 25066 -13460
rect 25100 -13494 25166 -13460
rect 25200 -13494 25954 -13460
rect 25988 -13494 26054 -13460
rect 26088 -13494 26154 -13460
rect 26188 -13494 26254 -13460
rect 26288 -13494 26354 -13460
rect 26388 -13494 26454 -13460
rect 26488 -13494 26584 -13460
rect 16884 -14112 26584 -13494
rect 16884 -14248 20666 -14112
rect 16884 -14282 16938 -14248
rect 16972 -14282 17038 -14248
rect 17072 -14282 17138 -14248
rect 17172 -14282 17238 -14248
rect 17272 -14282 17338 -14248
rect 17372 -14282 17438 -14248
rect 17472 -14282 18226 -14248
rect 18260 -14282 18326 -14248
rect 18360 -14282 18426 -14248
rect 18460 -14282 18526 -14248
rect 18560 -14282 18626 -14248
rect 18660 -14282 18726 -14248
rect 18760 -14282 19514 -14248
rect 19548 -14282 19614 -14248
rect 19648 -14282 19714 -14248
rect 19748 -14282 19814 -14248
rect 19848 -14282 19914 -14248
rect 19948 -14282 20014 -14248
rect 20048 -14282 20666 -14248
rect 16884 -14348 20666 -14282
rect 16884 -14382 16938 -14348
rect 16972 -14382 17038 -14348
rect 17072 -14382 17138 -14348
rect 17172 -14382 17238 -14348
rect 17272 -14382 17338 -14348
rect 17372 -14382 17438 -14348
rect 17472 -14382 18226 -14348
rect 18260 -14382 18326 -14348
rect 18360 -14382 18426 -14348
rect 18460 -14382 18526 -14348
rect 18560 -14382 18626 -14348
rect 18660 -14382 18726 -14348
rect 18760 -14382 19514 -14348
rect 19548 -14382 19614 -14348
rect 19648 -14382 19714 -14348
rect 19748 -14382 19814 -14348
rect 19848 -14382 19914 -14348
rect 19948 -14382 20014 -14348
rect 20048 -14382 20666 -14348
rect 16884 -14448 20666 -14382
rect 16884 -14482 16938 -14448
rect 16972 -14482 17038 -14448
rect 17072 -14482 17138 -14448
rect 17172 -14482 17238 -14448
rect 17272 -14482 17338 -14448
rect 17372 -14482 17438 -14448
rect 17472 -14482 18226 -14448
rect 18260 -14482 18326 -14448
rect 18360 -14482 18426 -14448
rect 18460 -14482 18526 -14448
rect 18560 -14482 18626 -14448
rect 18660 -14482 18726 -14448
rect 18760 -14482 19514 -14448
rect 19548 -14482 19614 -14448
rect 19648 -14482 19714 -14448
rect 19748 -14482 19814 -14448
rect 19848 -14482 19914 -14448
rect 19948 -14482 20014 -14448
rect 20048 -14482 20666 -14448
rect 16884 -14548 20666 -14482
rect 16884 -14582 16938 -14548
rect 16972 -14582 17038 -14548
rect 17072 -14582 17138 -14548
rect 17172 -14582 17238 -14548
rect 17272 -14582 17338 -14548
rect 17372 -14582 17438 -14548
rect 17472 -14582 18226 -14548
rect 18260 -14582 18326 -14548
rect 18360 -14582 18426 -14548
rect 18460 -14582 18526 -14548
rect 18560 -14582 18626 -14548
rect 18660 -14582 18726 -14548
rect 18760 -14582 19514 -14548
rect 19548 -14582 19614 -14548
rect 19648 -14582 19714 -14548
rect 19748 -14582 19814 -14548
rect 19848 -14582 19914 -14548
rect 19948 -14582 20014 -14548
rect 20048 -14582 20666 -14548
rect 16884 -14648 20666 -14582
rect 16884 -14682 16938 -14648
rect 16972 -14682 17038 -14648
rect 17072 -14682 17138 -14648
rect 17172 -14682 17238 -14648
rect 17272 -14682 17338 -14648
rect 17372 -14682 17438 -14648
rect 17472 -14682 18226 -14648
rect 18260 -14682 18326 -14648
rect 18360 -14682 18426 -14648
rect 18460 -14682 18526 -14648
rect 18560 -14682 18626 -14648
rect 18660 -14682 18726 -14648
rect 18760 -14682 19514 -14648
rect 19548 -14682 19614 -14648
rect 19648 -14682 19714 -14648
rect 19748 -14682 19814 -14648
rect 19848 -14682 19914 -14648
rect 19948 -14682 20014 -14648
rect 20048 -14682 20666 -14648
rect 16884 -14748 20666 -14682
rect 16884 -14782 16938 -14748
rect 16972 -14782 17038 -14748
rect 17072 -14782 17138 -14748
rect 17172 -14782 17238 -14748
rect 17272 -14782 17338 -14748
rect 17372 -14782 17438 -14748
rect 17472 -14782 18226 -14748
rect 18260 -14782 18326 -14748
rect 18360 -14782 18426 -14748
rect 18460 -14782 18526 -14748
rect 18560 -14782 18626 -14748
rect 18660 -14782 18726 -14748
rect 18760 -14782 19514 -14748
rect 19548 -14782 19614 -14748
rect 19648 -14782 19714 -14748
rect 19748 -14782 19814 -14748
rect 19848 -14782 19914 -14748
rect 19948 -14782 20014 -14748
rect 20048 -14782 20666 -14748
rect 16884 -14932 20666 -14782
rect 20724 -14176 21428 -14170
rect 20724 -14868 20730 -14176
rect 21422 -14868 21428 -14176
rect 20724 -14874 21428 -14868
rect 21484 -14248 26584 -14112
rect 21484 -14282 22090 -14248
rect 22124 -14282 22190 -14248
rect 22224 -14282 22290 -14248
rect 22324 -14282 22390 -14248
rect 22424 -14282 22490 -14248
rect 22524 -14282 22590 -14248
rect 22624 -14282 23378 -14248
rect 23412 -14282 23478 -14248
rect 23512 -14282 23578 -14248
rect 23612 -14282 23678 -14248
rect 23712 -14282 23778 -14248
rect 23812 -14282 23878 -14248
rect 23912 -14282 24666 -14248
rect 24700 -14282 24766 -14248
rect 24800 -14282 24866 -14248
rect 24900 -14282 24966 -14248
rect 25000 -14282 25066 -14248
rect 25100 -14282 25166 -14248
rect 25200 -14282 25954 -14248
rect 25988 -14282 26054 -14248
rect 26088 -14282 26154 -14248
rect 26188 -14282 26254 -14248
rect 26288 -14282 26354 -14248
rect 26388 -14282 26454 -14248
rect 26488 -14282 26584 -14248
rect 21484 -14348 26584 -14282
rect 21484 -14382 22090 -14348
rect 22124 -14382 22190 -14348
rect 22224 -14382 22290 -14348
rect 22324 -14382 22390 -14348
rect 22424 -14382 22490 -14348
rect 22524 -14382 22590 -14348
rect 22624 -14382 23378 -14348
rect 23412 -14382 23478 -14348
rect 23512 -14382 23578 -14348
rect 23612 -14382 23678 -14348
rect 23712 -14382 23778 -14348
rect 23812 -14382 23878 -14348
rect 23912 -14382 24666 -14348
rect 24700 -14382 24766 -14348
rect 24800 -14382 24866 -14348
rect 24900 -14382 24966 -14348
rect 25000 -14382 25066 -14348
rect 25100 -14382 25166 -14348
rect 25200 -14382 25954 -14348
rect 25988 -14382 26054 -14348
rect 26088 -14382 26154 -14348
rect 26188 -14382 26254 -14348
rect 26288 -14382 26354 -14348
rect 26388 -14382 26454 -14348
rect 26488 -14382 26584 -14348
rect 21484 -14448 26584 -14382
rect 21484 -14482 22090 -14448
rect 22124 -14482 22190 -14448
rect 22224 -14482 22290 -14448
rect 22324 -14482 22390 -14448
rect 22424 -14482 22490 -14448
rect 22524 -14482 22590 -14448
rect 22624 -14482 23378 -14448
rect 23412 -14482 23478 -14448
rect 23512 -14482 23578 -14448
rect 23612 -14482 23678 -14448
rect 23712 -14482 23778 -14448
rect 23812 -14482 23878 -14448
rect 23912 -14482 24666 -14448
rect 24700 -14482 24766 -14448
rect 24800 -14482 24866 -14448
rect 24900 -14482 24966 -14448
rect 25000 -14482 25066 -14448
rect 25100 -14482 25166 -14448
rect 25200 -14482 25954 -14448
rect 25988 -14482 26054 -14448
rect 26088 -14482 26154 -14448
rect 26188 -14482 26254 -14448
rect 26288 -14482 26354 -14448
rect 26388 -14482 26454 -14448
rect 26488 -14482 26584 -14448
rect 21484 -14548 26584 -14482
rect 21484 -14582 22090 -14548
rect 22124 -14582 22190 -14548
rect 22224 -14582 22290 -14548
rect 22324 -14582 22390 -14548
rect 22424 -14582 22490 -14548
rect 22524 -14582 22590 -14548
rect 22624 -14582 23378 -14548
rect 23412 -14582 23478 -14548
rect 23512 -14582 23578 -14548
rect 23612 -14582 23678 -14548
rect 23712 -14582 23778 -14548
rect 23812 -14582 23878 -14548
rect 23912 -14582 24666 -14548
rect 24700 -14582 24766 -14548
rect 24800 -14582 24866 -14548
rect 24900 -14582 24966 -14548
rect 25000 -14582 25066 -14548
rect 25100 -14582 25166 -14548
rect 25200 -14582 25954 -14548
rect 25988 -14582 26054 -14548
rect 26088 -14582 26154 -14548
rect 26188 -14582 26254 -14548
rect 26288 -14582 26354 -14548
rect 26388 -14582 26454 -14548
rect 26488 -14582 26584 -14548
rect 21484 -14648 26584 -14582
rect 21484 -14682 22090 -14648
rect 22124 -14682 22190 -14648
rect 22224 -14682 22290 -14648
rect 22324 -14682 22390 -14648
rect 22424 -14682 22490 -14648
rect 22524 -14682 22590 -14648
rect 22624 -14682 23378 -14648
rect 23412 -14682 23478 -14648
rect 23512 -14682 23578 -14648
rect 23612 -14682 23678 -14648
rect 23712 -14682 23778 -14648
rect 23812 -14682 23878 -14648
rect 23912 -14682 24666 -14648
rect 24700 -14682 24766 -14648
rect 24800 -14682 24866 -14648
rect 24900 -14682 24966 -14648
rect 25000 -14682 25066 -14648
rect 25100 -14682 25166 -14648
rect 25200 -14682 25954 -14648
rect 25988 -14682 26054 -14648
rect 26088 -14682 26154 -14648
rect 26188 -14682 26254 -14648
rect 26288 -14682 26354 -14648
rect 26388 -14682 26454 -14648
rect 26488 -14682 26584 -14648
rect 21484 -14748 26584 -14682
rect 21484 -14782 22090 -14748
rect 22124 -14782 22190 -14748
rect 22224 -14782 22290 -14748
rect 22324 -14782 22390 -14748
rect 22424 -14782 22490 -14748
rect 22524 -14782 22590 -14748
rect 22624 -14782 23378 -14748
rect 23412 -14782 23478 -14748
rect 23512 -14782 23578 -14748
rect 23612 -14782 23678 -14748
rect 23712 -14782 23778 -14748
rect 23812 -14782 23878 -14748
rect 23912 -14782 24666 -14748
rect 24700 -14782 24766 -14748
rect 24800 -14782 24866 -14748
rect 24900 -14782 24966 -14748
rect 25000 -14782 25066 -14748
rect 25100 -14782 25166 -14748
rect 25200 -14782 25954 -14748
rect 25988 -14782 26054 -14748
rect 26088 -14782 26154 -14748
rect 26188 -14782 26254 -14748
rect 26288 -14782 26354 -14748
rect 26388 -14782 26454 -14748
rect 26488 -14782 26584 -14748
rect 21484 -14932 26584 -14782
rect 16884 -15464 26584 -14932
rect 16884 -15536 25882 -15464
rect 16884 -15570 16938 -15536
rect 16972 -15570 17038 -15536
rect 17072 -15570 17138 -15536
rect 17172 -15570 17238 -15536
rect 17272 -15570 17338 -15536
rect 17372 -15570 17438 -15536
rect 17472 -15570 18226 -15536
rect 18260 -15570 18326 -15536
rect 18360 -15570 18426 -15536
rect 18460 -15570 18526 -15536
rect 18560 -15570 18626 -15536
rect 18660 -15570 18726 -15536
rect 18760 -15570 19514 -15536
rect 19548 -15570 19614 -15536
rect 19648 -15570 19714 -15536
rect 19748 -15570 19814 -15536
rect 19848 -15570 19914 -15536
rect 19948 -15570 20014 -15536
rect 20048 -15570 20802 -15536
rect 20836 -15570 20902 -15536
rect 20936 -15570 21002 -15536
rect 21036 -15570 21102 -15536
rect 21136 -15570 21202 -15536
rect 21236 -15570 21302 -15536
rect 21336 -15570 22090 -15536
rect 22124 -15570 22190 -15536
rect 22224 -15570 22290 -15536
rect 22324 -15570 22390 -15536
rect 22424 -15570 22490 -15536
rect 22524 -15570 22590 -15536
rect 22624 -15570 23378 -15536
rect 23412 -15570 23478 -15536
rect 23512 -15570 23578 -15536
rect 23612 -15570 23678 -15536
rect 23712 -15570 23778 -15536
rect 23812 -15570 23878 -15536
rect 23912 -15570 24666 -15536
rect 24700 -15570 24766 -15536
rect 24800 -15570 24866 -15536
rect 24900 -15570 24966 -15536
rect 25000 -15570 25066 -15536
rect 25100 -15570 25166 -15536
rect 25200 -15570 25882 -15536
rect 16884 -15636 25882 -15570
rect 16884 -15670 16938 -15636
rect 16972 -15670 17038 -15636
rect 17072 -15670 17138 -15636
rect 17172 -15670 17238 -15636
rect 17272 -15670 17338 -15636
rect 17372 -15670 17438 -15636
rect 17472 -15670 18226 -15636
rect 18260 -15670 18326 -15636
rect 18360 -15670 18426 -15636
rect 18460 -15670 18526 -15636
rect 18560 -15670 18626 -15636
rect 18660 -15670 18726 -15636
rect 18760 -15670 19514 -15636
rect 19548 -15670 19614 -15636
rect 19648 -15670 19714 -15636
rect 19748 -15670 19814 -15636
rect 19848 -15670 19914 -15636
rect 19948 -15670 20014 -15636
rect 20048 -15670 20802 -15636
rect 20836 -15670 20902 -15636
rect 20936 -15670 21002 -15636
rect 21036 -15670 21102 -15636
rect 21136 -15670 21202 -15636
rect 21236 -15670 21302 -15636
rect 21336 -15670 22090 -15636
rect 22124 -15670 22190 -15636
rect 22224 -15670 22290 -15636
rect 22324 -15670 22390 -15636
rect 22424 -15670 22490 -15636
rect 22524 -15670 22590 -15636
rect 22624 -15670 23378 -15636
rect 23412 -15670 23478 -15636
rect 23512 -15670 23578 -15636
rect 23612 -15670 23678 -15636
rect 23712 -15670 23778 -15636
rect 23812 -15670 23878 -15636
rect 23912 -15670 24666 -15636
rect 24700 -15670 24766 -15636
rect 24800 -15670 24866 -15636
rect 24900 -15670 24966 -15636
rect 25000 -15670 25066 -15636
rect 25100 -15670 25166 -15636
rect 25200 -15670 25882 -15636
rect 16884 -15736 25882 -15670
rect 16884 -15770 16938 -15736
rect 16972 -15770 17038 -15736
rect 17072 -15770 17138 -15736
rect 17172 -15770 17238 -15736
rect 17272 -15770 17338 -15736
rect 17372 -15770 17438 -15736
rect 17472 -15770 18226 -15736
rect 18260 -15770 18326 -15736
rect 18360 -15770 18426 -15736
rect 18460 -15770 18526 -15736
rect 18560 -15770 18626 -15736
rect 18660 -15770 18726 -15736
rect 18760 -15770 19514 -15736
rect 19548 -15770 19614 -15736
rect 19648 -15770 19714 -15736
rect 19748 -15770 19814 -15736
rect 19848 -15770 19914 -15736
rect 19948 -15770 20014 -15736
rect 20048 -15770 20802 -15736
rect 20836 -15770 20902 -15736
rect 20936 -15770 21002 -15736
rect 21036 -15770 21102 -15736
rect 21136 -15770 21202 -15736
rect 21236 -15770 21302 -15736
rect 21336 -15770 22090 -15736
rect 22124 -15770 22190 -15736
rect 22224 -15770 22290 -15736
rect 22324 -15770 22390 -15736
rect 22424 -15770 22490 -15736
rect 22524 -15770 22590 -15736
rect 22624 -15770 23378 -15736
rect 23412 -15770 23478 -15736
rect 23512 -15770 23578 -15736
rect 23612 -15770 23678 -15736
rect 23712 -15770 23778 -15736
rect 23812 -15770 23878 -15736
rect 23912 -15770 24666 -15736
rect 24700 -15770 24766 -15736
rect 24800 -15770 24866 -15736
rect 24900 -15770 24966 -15736
rect 25000 -15770 25066 -15736
rect 25100 -15770 25166 -15736
rect 25200 -15770 25882 -15736
rect 16884 -15836 25882 -15770
rect 16884 -15870 16938 -15836
rect 16972 -15870 17038 -15836
rect 17072 -15870 17138 -15836
rect 17172 -15870 17238 -15836
rect 17272 -15870 17338 -15836
rect 17372 -15870 17438 -15836
rect 17472 -15870 18226 -15836
rect 18260 -15870 18326 -15836
rect 18360 -15870 18426 -15836
rect 18460 -15870 18526 -15836
rect 18560 -15870 18626 -15836
rect 18660 -15870 18726 -15836
rect 18760 -15870 19514 -15836
rect 19548 -15870 19614 -15836
rect 19648 -15870 19714 -15836
rect 19748 -15870 19814 -15836
rect 19848 -15870 19914 -15836
rect 19948 -15870 20014 -15836
rect 20048 -15870 20802 -15836
rect 20836 -15870 20902 -15836
rect 20936 -15870 21002 -15836
rect 21036 -15870 21102 -15836
rect 21136 -15870 21202 -15836
rect 21236 -15870 21302 -15836
rect 21336 -15870 22090 -15836
rect 22124 -15870 22190 -15836
rect 22224 -15870 22290 -15836
rect 22324 -15870 22390 -15836
rect 22424 -15870 22490 -15836
rect 22524 -15870 22590 -15836
rect 22624 -15870 23378 -15836
rect 23412 -15870 23478 -15836
rect 23512 -15870 23578 -15836
rect 23612 -15870 23678 -15836
rect 23712 -15870 23778 -15836
rect 23812 -15870 23878 -15836
rect 23912 -15870 24666 -15836
rect 24700 -15870 24766 -15836
rect 24800 -15870 24866 -15836
rect 24900 -15870 24966 -15836
rect 25000 -15870 25066 -15836
rect 25100 -15870 25166 -15836
rect 25200 -15870 25882 -15836
rect 16884 -15936 25882 -15870
rect 16884 -15970 16938 -15936
rect 16972 -15970 17038 -15936
rect 17072 -15970 17138 -15936
rect 17172 -15970 17238 -15936
rect 17272 -15970 17338 -15936
rect 17372 -15970 17438 -15936
rect 17472 -15970 18226 -15936
rect 18260 -15970 18326 -15936
rect 18360 -15970 18426 -15936
rect 18460 -15970 18526 -15936
rect 18560 -15970 18626 -15936
rect 18660 -15970 18726 -15936
rect 18760 -15970 19514 -15936
rect 19548 -15970 19614 -15936
rect 19648 -15970 19714 -15936
rect 19748 -15970 19814 -15936
rect 19848 -15970 19914 -15936
rect 19948 -15970 20014 -15936
rect 20048 -15970 20802 -15936
rect 20836 -15970 20902 -15936
rect 20936 -15970 21002 -15936
rect 21036 -15970 21102 -15936
rect 21136 -15970 21202 -15936
rect 21236 -15970 21302 -15936
rect 21336 -15970 22090 -15936
rect 22124 -15970 22190 -15936
rect 22224 -15970 22290 -15936
rect 22324 -15970 22390 -15936
rect 22424 -15970 22490 -15936
rect 22524 -15970 22590 -15936
rect 22624 -15970 23378 -15936
rect 23412 -15970 23478 -15936
rect 23512 -15970 23578 -15936
rect 23612 -15970 23678 -15936
rect 23712 -15970 23778 -15936
rect 23812 -15970 23878 -15936
rect 23912 -15970 24666 -15936
rect 24700 -15970 24766 -15936
rect 24800 -15970 24866 -15936
rect 24900 -15970 24966 -15936
rect 25000 -15970 25066 -15936
rect 25100 -15970 25166 -15936
rect 25200 -15970 25882 -15936
rect 16884 -16036 25882 -15970
rect 16884 -16070 16938 -16036
rect 16972 -16070 17038 -16036
rect 17072 -16070 17138 -16036
rect 17172 -16070 17238 -16036
rect 17272 -16070 17338 -16036
rect 17372 -16070 17438 -16036
rect 17472 -16070 18226 -16036
rect 18260 -16070 18326 -16036
rect 18360 -16070 18426 -16036
rect 18460 -16070 18526 -16036
rect 18560 -16070 18626 -16036
rect 18660 -16070 18726 -16036
rect 18760 -16070 19514 -16036
rect 19548 -16070 19614 -16036
rect 19648 -16070 19714 -16036
rect 19748 -16070 19814 -16036
rect 19848 -16070 19914 -16036
rect 19948 -16070 20014 -16036
rect 20048 -16070 20802 -16036
rect 20836 -16070 20902 -16036
rect 20936 -16070 21002 -16036
rect 21036 -16070 21102 -16036
rect 21136 -16070 21202 -16036
rect 21236 -16070 21302 -16036
rect 21336 -16070 22090 -16036
rect 22124 -16070 22190 -16036
rect 22224 -16070 22290 -16036
rect 22324 -16070 22390 -16036
rect 22424 -16070 22490 -16036
rect 22524 -16070 22590 -16036
rect 22624 -16070 23378 -16036
rect 23412 -16070 23478 -16036
rect 23512 -16070 23578 -16036
rect 23612 -16070 23678 -16036
rect 23712 -16070 23778 -16036
rect 23812 -16070 23878 -16036
rect 23912 -16070 24666 -16036
rect 24700 -16070 24766 -16036
rect 24800 -16070 24866 -16036
rect 24900 -16070 24966 -16036
rect 25000 -16070 25066 -16036
rect 25100 -16070 25166 -16036
rect 25200 -16070 25882 -16036
rect 16884 -16156 25882 -16070
rect 26574 -16156 26584 -15464
rect 16884 -16751 26584 -16156
rect 16884 -16824 25882 -16751
rect 16884 -16858 16938 -16824
rect 16972 -16858 17038 -16824
rect 17072 -16858 17138 -16824
rect 17172 -16858 17238 -16824
rect 17272 -16858 17338 -16824
rect 17372 -16858 17438 -16824
rect 17472 -16858 18226 -16824
rect 18260 -16858 18326 -16824
rect 18360 -16858 18426 -16824
rect 18460 -16858 18526 -16824
rect 18560 -16858 18626 -16824
rect 18660 -16858 18726 -16824
rect 18760 -16858 19514 -16824
rect 19548 -16858 19614 -16824
rect 19648 -16858 19714 -16824
rect 19748 -16858 19814 -16824
rect 19848 -16858 19914 -16824
rect 19948 -16858 20014 -16824
rect 20048 -16858 20802 -16824
rect 20836 -16858 20902 -16824
rect 20936 -16858 21002 -16824
rect 21036 -16858 21102 -16824
rect 21136 -16858 21202 -16824
rect 21236 -16858 21302 -16824
rect 21336 -16858 22090 -16824
rect 22124 -16858 22190 -16824
rect 22224 -16858 22290 -16824
rect 22324 -16858 22390 -16824
rect 22424 -16858 22490 -16824
rect 22524 -16858 22590 -16824
rect 22624 -16858 23378 -16824
rect 23412 -16858 23478 -16824
rect 23512 -16858 23578 -16824
rect 23612 -16858 23678 -16824
rect 23712 -16858 23778 -16824
rect 23812 -16858 23878 -16824
rect 23912 -16858 24666 -16824
rect 24700 -16858 24766 -16824
rect 24800 -16858 24866 -16824
rect 24900 -16858 24966 -16824
rect 25000 -16858 25066 -16824
rect 25100 -16858 25166 -16824
rect 25200 -16858 25882 -16824
rect 16884 -16924 25882 -16858
rect 16884 -16958 16938 -16924
rect 16972 -16958 17038 -16924
rect 17072 -16958 17138 -16924
rect 17172 -16958 17238 -16924
rect 17272 -16958 17338 -16924
rect 17372 -16958 17438 -16924
rect 17472 -16958 18226 -16924
rect 18260 -16958 18326 -16924
rect 18360 -16958 18426 -16924
rect 18460 -16958 18526 -16924
rect 18560 -16958 18626 -16924
rect 18660 -16958 18726 -16924
rect 18760 -16958 19514 -16924
rect 19548 -16958 19614 -16924
rect 19648 -16958 19714 -16924
rect 19748 -16958 19814 -16924
rect 19848 -16958 19914 -16924
rect 19948 -16958 20014 -16924
rect 20048 -16958 20802 -16924
rect 20836 -16958 20902 -16924
rect 20936 -16958 21002 -16924
rect 21036 -16958 21102 -16924
rect 21136 -16958 21202 -16924
rect 21236 -16958 21302 -16924
rect 21336 -16958 22090 -16924
rect 22124 -16958 22190 -16924
rect 22224 -16958 22290 -16924
rect 22324 -16958 22390 -16924
rect 22424 -16958 22490 -16924
rect 22524 -16958 22590 -16924
rect 22624 -16958 23378 -16924
rect 23412 -16958 23478 -16924
rect 23512 -16958 23578 -16924
rect 23612 -16958 23678 -16924
rect 23712 -16958 23778 -16924
rect 23812 -16958 23878 -16924
rect 23912 -16958 24666 -16924
rect 24700 -16958 24766 -16924
rect 24800 -16958 24866 -16924
rect 24900 -16958 24966 -16924
rect 25000 -16958 25066 -16924
rect 25100 -16958 25166 -16924
rect 25200 -16958 25882 -16924
rect 16884 -17024 25882 -16958
rect 16884 -17058 16938 -17024
rect 16972 -17058 17038 -17024
rect 17072 -17058 17138 -17024
rect 17172 -17058 17238 -17024
rect 17272 -17058 17338 -17024
rect 17372 -17058 17438 -17024
rect 17472 -17058 18226 -17024
rect 18260 -17058 18326 -17024
rect 18360 -17058 18426 -17024
rect 18460 -17058 18526 -17024
rect 18560 -17058 18626 -17024
rect 18660 -17058 18726 -17024
rect 18760 -17058 19514 -17024
rect 19548 -17058 19614 -17024
rect 19648 -17058 19714 -17024
rect 19748 -17058 19814 -17024
rect 19848 -17058 19914 -17024
rect 19948 -17058 20014 -17024
rect 20048 -17058 20802 -17024
rect 20836 -17058 20902 -17024
rect 20936 -17058 21002 -17024
rect 21036 -17058 21102 -17024
rect 21136 -17058 21202 -17024
rect 21236 -17058 21302 -17024
rect 21336 -17058 22090 -17024
rect 22124 -17058 22190 -17024
rect 22224 -17058 22290 -17024
rect 22324 -17058 22390 -17024
rect 22424 -17058 22490 -17024
rect 22524 -17058 22590 -17024
rect 22624 -17058 23378 -17024
rect 23412 -17058 23478 -17024
rect 23512 -17058 23578 -17024
rect 23612 -17058 23678 -17024
rect 23712 -17058 23778 -17024
rect 23812 -17058 23878 -17024
rect 23912 -17058 24666 -17024
rect 24700 -17058 24766 -17024
rect 24800 -17058 24866 -17024
rect 24900 -17058 24966 -17024
rect 25000 -17058 25066 -17024
rect 25100 -17058 25166 -17024
rect 25200 -17058 25882 -17024
rect 16884 -17124 25882 -17058
rect 16884 -17158 16938 -17124
rect 16972 -17158 17038 -17124
rect 17072 -17158 17138 -17124
rect 17172 -17158 17238 -17124
rect 17272 -17158 17338 -17124
rect 17372 -17158 17438 -17124
rect 17472 -17158 18226 -17124
rect 18260 -17158 18326 -17124
rect 18360 -17158 18426 -17124
rect 18460 -17158 18526 -17124
rect 18560 -17158 18626 -17124
rect 18660 -17158 18726 -17124
rect 18760 -17158 19514 -17124
rect 19548 -17158 19614 -17124
rect 19648 -17158 19714 -17124
rect 19748 -17158 19814 -17124
rect 19848 -17158 19914 -17124
rect 19948 -17158 20014 -17124
rect 20048 -17158 20802 -17124
rect 20836 -17158 20902 -17124
rect 20936 -17158 21002 -17124
rect 21036 -17158 21102 -17124
rect 21136 -17158 21202 -17124
rect 21236 -17158 21302 -17124
rect 21336 -17158 22090 -17124
rect 22124 -17158 22190 -17124
rect 22224 -17158 22290 -17124
rect 22324 -17158 22390 -17124
rect 22424 -17158 22490 -17124
rect 22524 -17158 22590 -17124
rect 22624 -17158 23378 -17124
rect 23412 -17158 23478 -17124
rect 23512 -17158 23578 -17124
rect 23612 -17158 23678 -17124
rect 23712 -17158 23778 -17124
rect 23812 -17158 23878 -17124
rect 23912 -17158 24666 -17124
rect 24700 -17158 24766 -17124
rect 24800 -17158 24866 -17124
rect 24900 -17158 24966 -17124
rect 25000 -17158 25066 -17124
rect 25100 -17158 25166 -17124
rect 25200 -17158 25882 -17124
rect 16884 -17224 25882 -17158
rect 16884 -17258 16938 -17224
rect 16972 -17258 17038 -17224
rect 17072 -17258 17138 -17224
rect 17172 -17258 17238 -17224
rect 17272 -17258 17338 -17224
rect 17372 -17258 17438 -17224
rect 17472 -17258 18226 -17224
rect 18260 -17258 18326 -17224
rect 18360 -17258 18426 -17224
rect 18460 -17258 18526 -17224
rect 18560 -17258 18626 -17224
rect 18660 -17258 18726 -17224
rect 18760 -17258 19514 -17224
rect 19548 -17258 19614 -17224
rect 19648 -17258 19714 -17224
rect 19748 -17258 19814 -17224
rect 19848 -17258 19914 -17224
rect 19948 -17258 20014 -17224
rect 20048 -17258 20802 -17224
rect 20836 -17258 20902 -17224
rect 20936 -17258 21002 -17224
rect 21036 -17258 21102 -17224
rect 21136 -17258 21202 -17224
rect 21236 -17258 21302 -17224
rect 21336 -17258 22090 -17224
rect 22124 -17258 22190 -17224
rect 22224 -17258 22290 -17224
rect 22324 -17258 22390 -17224
rect 22424 -17258 22490 -17224
rect 22524 -17258 22590 -17224
rect 22624 -17258 23378 -17224
rect 23412 -17258 23478 -17224
rect 23512 -17258 23578 -17224
rect 23612 -17258 23678 -17224
rect 23712 -17258 23778 -17224
rect 23812 -17258 23878 -17224
rect 23912 -17258 24666 -17224
rect 24700 -17258 24766 -17224
rect 24800 -17258 24866 -17224
rect 24900 -17258 24966 -17224
rect 25000 -17258 25066 -17224
rect 25100 -17258 25166 -17224
rect 25200 -17258 25882 -17224
rect 6882 -17296 7291 -17284
rect 6882 -17834 6888 -17296
rect 7285 -17834 7291 -17296
rect 6882 -17846 7291 -17834
rect 13617 -17296 14026 -17284
rect 13617 -17834 13623 -17296
rect 14020 -17834 14026 -17296
rect 16884 -17324 25882 -17258
rect 16884 -17358 16938 -17324
rect 16972 -17358 17038 -17324
rect 17072 -17358 17138 -17324
rect 17172 -17358 17238 -17324
rect 17272 -17358 17338 -17324
rect 17372 -17358 17438 -17324
rect 17472 -17358 18226 -17324
rect 18260 -17358 18326 -17324
rect 18360 -17358 18426 -17324
rect 18460 -17358 18526 -17324
rect 18560 -17358 18626 -17324
rect 18660 -17358 18726 -17324
rect 18760 -17358 19514 -17324
rect 19548 -17358 19614 -17324
rect 19648 -17358 19714 -17324
rect 19748 -17358 19814 -17324
rect 19848 -17358 19914 -17324
rect 19948 -17358 20014 -17324
rect 20048 -17358 20802 -17324
rect 20836 -17358 20902 -17324
rect 20936 -17358 21002 -17324
rect 21036 -17358 21102 -17324
rect 21136 -17358 21202 -17324
rect 21236 -17358 21302 -17324
rect 21336 -17358 22090 -17324
rect 22124 -17358 22190 -17324
rect 22224 -17358 22290 -17324
rect 22324 -17358 22390 -17324
rect 22424 -17358 22490 -17324
rect 22524 -17358 22590 -17324
rect 22624 -17358 23378 -17324
rect 23412 -17358 23478 -17324
rect 23512 -17358 23578 -17324
rect 23612 -17358 23678 -17324
rect 23712 -17358 23778 -17324
rect 23812 -17358 23878 -17324
rect 23912 -17358 24666 -17324
rect 24700 -17358 24766 -17324
rect 24800 -17358 24866 -17324
rect 24900 -17358 24966 -17324
rect 25000 -17358 25066 -17324
rect 25100 -17358 25166 -17324
rect 25200 -17358 25882 -17324
rect 16884 -17443 25882 -17358
rect 26574 -17443 26584 -16751
rect 16884 -17446 26584 -17443
rect 25876 -17449 26580 -17446
rect 13617 -17846 14026 -17834
rect 13606 -18048 14304 -18042
rect 6070 -18104 6640 -18098
rect 6070 -18662 6076 -18104
rect 6634 -18662 6640 -18104
rect 5270 -19740 5840 -19728
rect 5270 -20298 5276 -19740
rect 5834 -20298 5840 -19740
rect 5270 -22194 5840 -20298
rect 6070 -20558 6640 -18662
rect 6870 -18104 7302 -18098
rect 6870 -18662 6876 -18104
rect 7296 -18662 7302 -18104
rect 6870 -18668 7302 -18662
rect 13606 -18740 13612 -18048
rect 13606 -18746 14304 -18740
rect 13606 -18866 21430 -18860
rect 6870 -18922 7302 -18916
rect 6870 -19480 6876 -18922
rect 7296 -19480 7302 -18922
rect 6870 -19486 7302 -19480
rect 7532 -18922 8102 -18916
rect 7532 -19480 7538 -18922
rect 8096 -19480 8102 -18922
rect 6870 -19740 7302 -19734
rect 6870 -20298 6876 -19740
rect 7296 -20298 7302 -19740
rect 6870 -20304 7302 -20298
rect 6070 -21116 6076 -20558
rect 6634 -21116 6640 -20558
rect 6070 -21236 6640 -21116
rect 6870 -20558 7302 -20552
rect 6870 -21116 6876 -20558
rect 7296 -21116 7302 -20558
rect 6870 -21122 7302 -21116
rect 6870 -21376 7302 -21370
rect 6870 -21934 6876 -21376
rect 7296 -21934 7302 -21376
rect 6870 -21940 7302 -21934
rect 7532 -21376 8102 -19480
rect 13606 -19558 13612 -18866
rect 14304 -19558 20730 -18866
rect 21422 -19558 21430 -18866
rect 13606 -19564 21430 -19558
rect 13606 -19684 14310 -19678
rect 13606 -20376 13612 -19684
rect 14304 -20376 14310 -19684
rect 13606 -20382 14310 -20376
rect 16156 -19966 26582 -19960
rect 7532 -21934 7538 -21376
rect 8096 -21934 8102 -21376
rect 7532 -21940 8102 -21934
rect 12006 -20558 12576 -20552
rect 12006 -21116 12012 -20558
rect 12570 -21116 12576 -20558
rect 5270 -22752 5276 -22194
rect 5834 -22752 5840 -22194
rect 5270 -22926 5840 -22752
rect 6870 -22194 7302 -22188
rect 6870 -22752 6876 -22194
rect 7296 -22752 7302 -22194
rect 6870 -22758 7302 -22752
rect 6070 -23012 6640 -23006
rect 6070 -23570 6076 -23012
rect 6634 -23570 6640 -23012
rect 6070 -25466 6640 -23570
rect 6870 -23012 7302 -23006
rect 6870 -23570 6876 -23012
rect 7296 -23570 7302 -23012
rect 12006 -23012 12576 -21116
rect 13606 -20558 14038 -20552
rect 13606 -21116 13612 -20558
rect 14032 -21116 14038 -20558
rect 16156 -20900 16162 -19966
rect 16680 -20900 25640 -19966
rect 16156 -20902 25640 -20900
rect 26576 -20902 26582 -19966
rect 16156 -20906 26582 -20902
rect 16680 -20908 26582 -20906
rect 13606 -21122 14038 -21116
rect 13606 -21376 14038 -21370
rect 13606 -21934 13612 -21376
rect 14032 -21934 14038 -21376
rect 13606 -21940 14038 -21934
rect 14268 -21376 14838 -21370
rect 14268 -21934 14274 -21376
rect 14832 -21934 14838 -21376
rect 12006 -23570 12012 -23012
rect 12570 -23570 12576 -23012
rect 12806 -22194 13376 -22188
rect 12806 -22752 12812 -22194
rect 13370 -22752 13376 -22194
rect 6870 -23576 7302 -23570
rect 6870 -23830 7302 -23824
rect 6870 -24388 6876 -23830
rect 7296 -24388 7302 -23830
rect 6870 -24394 7302 -24388
rect 6870 -24648 7302 -24642
rect 6870 -25206 6876 -24648
rect 7296 -25206 7302 -24648
rect 6870 -25212 7302 -25206
rect 7532 -24648 8102 -24642
rect 7532 -25206 7538 -24648
rect 8096 -25206 8102 -24648
rect 6070 -26024 6076 -25466
rect 6634 -26024 6640 -25466
rect 6070 -26152 6640 -26024
rect 6870 -25466 7302 -25460
rect 6870 -26024 6876 -25466
rect 7296 -26024 7302 -25466
rect 6870 -26030 7302 -26024
rect 5270 -26284 5840 -26278
rect 5270 -26842 5276 -26284
rect 5834 -26842 5840 -26284
rect 5270 -27908 5840 -26842
rect 6870 -26284 7302 -26278
rect 6870 -26842 6876 -26284
rect 7296 -26842 7302 -26284
rect 6870 -26848 7302 -26842
rect 6870 -27102 7302 -27096
rect 6870 -27660 6876 -27102
rect 7296 -27660 7302 -27102
rect 6870 -27666 7302 -27660
rect 7532 -27102 8102 -25206
rect 7532 -27660 7538 -27102
rect 8096 -27660 8102 -27102
rect 7532 -27666 8102 -27660
rect 12006 -25466 12576 -25460
rect 12006 -26024 12012 -25466
rect 12570 -26024 12576 -25466
rect 5270 -28466 5276 -27908
rect 5834 -28466 5840 -27908
rect 5270 -28472 5840 -28466
rect 6870 -27920 7302 -27914
rect 6870 -28478 6876 -27920
rect 7296 -28478 7302 -27920
rect 6870 -28484 7302 -28478
rect 6070 -28738 6640 -28732
rect 6070 -29296 6076 -28738
rect 6634 -29296 6640 -28738
rect 6070 -34464 6640 -29296
rect 6870 -28738 7302 -28732
rect 6870 -29296 6876 -28738
rect 7296 -29296 7302 -28738
rect 6870 -29302 7302 -29296
rect 12006 -28738 12576 -26024
rect 12806 -26284 13376 -22752
rect 13606 -22194 14038 -22188
rect 13606 -22752 13612 -22194
rect 14032 -22752 14038 -22194
rect 13606 -22758 14038 -22752
rect 13606 -23012 14038 -23006
rect 13606 -23570 13612 -23012
rect 14032 -23570 14038 -23012
rect 13606 -23576 14038 -23570
rect 13606 -23774 14162 -23768
rect 13606 -23830 13644 -23774
rect 13606 -24388 13612 -23830
rect 13606 -24466 13644 -24388
rect 13606 -24472 14162 -24466
rect 13606 -24648 14038 -24642
rect 13606 -25206 13612 -24648
rect 14032 -25206 14038 -24648
rect 13606 -25212 14038 -25206
rect 14268 -24648 14838 -21934
rect 14268 -25206 14274 -24648
rect 14832 -25206 14838 -24648
rect 14268 -25212 14838 -25206
rect 13606 -25466 14038 -25460
rect 13606 -26024 13612 -25466
rect 14032 -26024 14038 -25466
rect 13606 -26030 14038 -26024
rect 12806 -26842 12812 -26284
rect 13370 -26842 13376 -26284
rect 12806 -26848 13376 -26842
rect 13606 -26284 14038 -26278
rect 13606 -26842 13612 -26284
rect 14032 -26842 14038 -26284
rect 13606 -26848 14038 -26842
rect 13606 -27102 14038 -27096
rect 13606 -27660 13612 -27102
rect 14032 -27660 14038 -27102
rect 13606 -27666 14038 -27660
rect 14268 -27102 14838 -27096
rect 14268 -27660 14274 -27102
rect 14832 -27660 14838 -27102
rect 12006 -29296 12012 -28738
rect 12570 -29296 12576 -28738
rect 12006 -29302 12576 -29296
rect 12806 -27920 13376 -27914
rect 12806 -28478 12812 -27920
rect 13370 -28478 13376 -27920
rect 6870 -29556 7302 -29550
rect 6870 -30114 6876 -29556
rect 7296 -30114 7302 -29556
rect 6870 -30120 7302 -30114
rect 7532 -29556 8102 -29550
rect 7532 -30114 7538 -29556
rect 8096 -30114 8102 -29556
rect 6882 -30384 7291 -30372
rect 6882 -30922 6888 -30384
rect 7285 -30922 7291 -30384
rect 6882 -30934 7291 -30922
rect 6820 -32838 7229 -32826
rect 6820 -33376 6826 -32838
rect 7223 -33376 7229 -32838
rect 6820 -33388 7229 -33376
rect 6808 -33646 7240 -33640
rect 6808 -34204 6814 -33646
rect 7234 -34204 7240 -33646
rect 6808 -34210 7240 -34204
rect 7532 -33646 8102 -30114
rect 7532 -34204 7538 -33646
rect 8030 -34204 8102 -33646
rect 7532 -34212 8102 -34204
rect 11540 -31182 12676 -31172
rect 11540 -31694 11570 -31182
rect 12622 -31694 12676 -31182
rect 11540 -32838 12676 -31694
rect 11540 -33376 11557 -32838
rect 11954 -33376 12676 -32838
rect 11540 -33656 12676 -33376
rect 11540 -34194 11557 -33656
rect 11954 -34194 12676 -33656
rect 6070 -35022 6076 -34464
rect 6634 -35022 6640 -34464
rect 6070 -35028 6640 -35022
rect 6808 -34464 7240 -34458
rect 6808 -35022 6814 -34464
rect 7234 -35022 7240 -34464
rect 6808 -35028 7240 -35022
rect 11540 -34474 12676 -34194
rect 11540 -35012 11557 -34474
rect 11954 -35012 12676 -34474
rect 6820 -35292 7229 -35280
rect 6820 -35830 6826 -35292
rect 7223 -35830 7229 -35292
rect 6820 -35842 7229 -35830
rect 11540 -35292 12676 -35012
rect 11540 -35830 11557 -35292
rect 11954 -35830 12676 -35292
rect 11540 -36152 12676 -35830
rect 11540 -36646 11568 -36152
rect 12634 -36646 12676 -36152
rect 11540 -36668 12676 -36646
rect 8206 -36928 8615 -36916
rect 8206 -37466 8212 -36928
rect 8609 -37466 8615 -36928
rect 8206 -37478 8615 -37466
rect 11961 -36928 12370 -36916
rect 11961 -37466 11967 -36928
rect 12364 -37466 12370 -36928
rect 11961 -37478 12370 -37466
rect 12806 -37730 13376 -28478
rect 13606 -27920 14038 -27914
rect 13606 -28478 13612 -27920
rect 14032 -28478 14038 -27920
rect 13606 -28484 14038 -28478
rect 13606 -28738 14038 -28732
rect 13606 -29296 13612 -28738
rect 14032 -29296 14038 -28738
rect 13606 -29302 14038 -29296
rect 13606 -29556 14038 -29550
rect 13606 -30114 13612 -29556
rect 14032 -30114 14038 -29556
rect 13606 -30120 14038 -30114
rect 14268 -29556 14838 -27660
rect 14268 -30114 14274 -29556
rect 14832 -30114 14838 -29556
rect 14268 -30120 14838 -30114
rect 13617 -30384 14026 -30372
rect 13617 -30922 13623 -30384
rect 14020 -30922 14026 -30384
rect 13617 -30934 14026 -30922
rect 8206 -37746 8615 -37734
rect 8206 -38284 8212 -37746
rect 8609 -38284 8615 -37746
rect 8206 -38296 8615 -38284
rect 11950 -37746 13376 -37730
rect 11950 -38284 11967 -37746
rect 12364 -38284 13376 -37746
rect 11950 -38300 13376 -38284
rect 8206 -38564 8615 -38552
rect 8206 -39102 8212 -38564
rect 8609 -39102 8615 -38564
rect 8206 -39114 8615 -39102
rect 11961 -38564 12370 -38552
rect 11961 -39102 11967 -38564
rect 12364 -39102 12370 -38564
rect 11961 -39114 12370 -39102
<< via1 >>
rect 20730 -14248 21422 -14176
rect 20730 -14282 20802 -14248
rect 20802 -14282 20836 -14248
rect 20836 -14282 20902 -14248
rect 20902 -14282 20936 -14248
rect 20936 -14282 21002 -14248
rect 21002 -14282 21036 -14248
rect 21036 -14282 21102 -14248
rect 21102 -14282 21136 -14248
rect 21136 -14282 21202 -14248
rect 21202 -14282 21236 -14248
rect 21236 -14282 21302 -14248
rect 21302 -14282 21336 -14248
rect 21336 -14282 21422 -14248
rect 20730 -14348 21422 -14282
rect 20730 -14382 20802 -14348
rect 20802 -14382 20836 -14348
rect 20836 -14382 20902 -14348
rect 20902 -14382 20936 -14348
rect 20936 -14382 21002 -14348
rect 21002 -14382 21036 -14348
rect 21036 -14382 21102 -14348
rect 21102 -14382 21136 -14348
rect 21136 -14382 21202 -14348
rect 21202 -14382 21236 -14348
rect 21236 -14382 21302 -14348
rect 21302 -14382 21336 -14348
rect 21336 -14382 21422 -14348
rect 20730 -14448 21422 -14382
rect 20730 -14482 20802 -14448
rect 20802 -14482 20836 -14448
rect 20836 -14482 20902 -14448
rect 20902 -14482 20936 -14448
rect 20936 -14482 21002 -14448
rect 21002 -14482 21036 -14448
rect 21036 -14482 21102 -14448
rect 21102 -14482 21136 -14448
rect 21136 -14482 21202 -14448
rect 21202 -14482 21236 -14448
rect 21236 -14482 21302 -14448
rect 21302 -14482 21336 -14448
rect 21336 -14482 21422 -14448
rect 20730 -14548 21422 -14482
rect 20730 -14582 20802 -14548
rect 20802 -14582 20836 -14548
rect 20836 -14582 20902 -14548
rect 20902 -14582 20936 -14548
rect 20936 -14582 21002 -14548
rect 21002 -14582 21036 -14548
rect 21036 -14582 21102 -14548
rect 21102 -14582 21136 -14548
rect 21136 -14582 21202 -14548
rect 21202 -14582 21236 -14548
rect 21236 -14582 21302 -14548
rect 21302 -14582 21336 -14548
rect 21336 -14582 21422 -14548
rect 20730 -14648 21422 -14582
rect 20730 -14682 20802 -14648
rect 20802 -14682 20836 -14648
rect 20836 -14682 20902 -14648
rect 20902 -14682 20936 -14648
rect 20936 -14682 21002 -14648
rect 21002 -14682 21036 -14648
rect 21036 -14682 21102 -14648
rect 21102 -14682 21136 -14648
rect 21136 -14682 21202 -14648
rect 21202 -14682 21236 -14648
rect 21236 -14682 21302 -14648
rect 21302 -14682 21336 -14648
rect 21336 -14682 21422 -14648
rect 20730 -14748 21422 -14682
rect 20730 -14782 20802 -14748
rect 20802 -14782 20836 -14748
rect 20836 -14782 20902 -14748
rect 20902 -14782 20936 -14748
rect 20936 -14782 21002 -14748
rect 21002 -14782 21036 -14748
rect 21036 -14782 21102 -14748
rect 21102 -14782 21136 -14748
rect 21136 -14782 21202 -14748
rect 21202 -14782 21236 -14748
rect 21236 -14782 21302 -14748
rect 21302 -14782 21336 -14748
rect 21336 -14782 21422 -14748
rect 20730 -14868 21422 -14782
rect 25882 -15536 26574 -15464
rect 25882 -15570 25954 -15536
rect 25954 -15570 25988 -15536
rect 25988 -15570 26054 -15536
rect 26054 -15570 26088 -15536
rect 26088 -15570 26154 -15536
rect 26154 -15570 26188 -15536
rect 26188 -15570 26254 -15536
rect 26254 -15570 26288 -15536
rect 26288 -15570 26354 -15536
rect 26354 -15570 26388 -15536
rect 26388 -15570 26454 -15536
rect 26454 -15570 26488 -15536
rect 26488 -15570 26574 -15536
rect 25882 -15636 26574 -15570
rect 25882 -15670 25954 -15636
rect 25954 -15670 25988 -15636
rect 25988 -15670 26054 -15636
rect 26054 -15670 26088 -15636
rect 26088 -15670 26154 -15636
rect 26154 -15670 26188 -15636
rect 26188 -15670 26254 -15636
rect 26254 -15670 26288 -15636
rect 26288 -15670 26354 -15636
rect 26354 -15670 26388 -15636
rect 26388 -15670 26454 -15636
rect 26454 -15670 26488 -15636
rect 26488 -15670 26574 -15636
rect 25882 -15736 26574 -15670
rect 25882 -15770 25954 -15736
rect 25954 -15770 25988 -15736
rect 25988 -15770 26054 -15736
rect 26054 -15770 26088 -15736
rect 26088 -15770 26154 -15736
rect 26154 -15770 26188 -15736
rect 26188 -15770 26254 -15736
rect 26254 -15770 26288 -15736
rect 26288 -15770 26354 -15736
rect 26354 -15770 26388 -15736
rect 26388 -15770 26454 -15736
rect 26454 -15770 26488 -15736
rect 26488 -15770 26574 -15736
rect 25882 -15836 26574 -15770
rect 25882 -15870 25954 -15836
rect 25954 -15870 25988 -15836
rect 25988 -15870 26054 -15836
rect 26054 -15870 26088 -15836
rect 26088 -15870 26154 -15836
rect 26154 -15870 26188 -15836
rect 26188 -15870 26254 -15836
rect 26254 -15870 26288 -15836
rect 26288 -15870 26354 -15836
rect 26354 -15870 26388 -15836
rect 26388 -15870 26454 -15836
rect 26454 -15870 26488 -15836
rect 26488 -15870 26574 -15836
rect 25882 -15936 26574 -15870
rect 25882 -15970 25954 -15936
rect 25954 -15970 25988 -15936
rect 25988 -15970 26054 -15936
rect 26054 -15970 26088 -15936
rect 26088 -15970 26154 -15936
rect 26154 -15970 26188 -15936
rect 26188 -15970 26254 -15936
rect 26254 -15970 26288 -15936
rect 26288 -15970 26354 -15936
rect 26354 -15970 26388 -15936
rect 26388 -15970 26454 -15936
rect 26454 -15970 26488 -15936
rect 26488 -15970 26574 -15936
rect 25882 -16036 26574 -15970
rect 25882 -16070 25954 -16036
rect 25954 -16070 25988 -16036
rect 25988 -16070 26054 -16036
rect 26054 -16070 26088 -16036
rect 26088 -16070 26154 -16036
rect 26154 -16070 26188 -16036
rect 26188 -16070 26254 -16036
rect 26254 -16070 26288 -16036
rect 26288 -16070 26354 -16036
rect 26354 -16070 26388 -16036
rect 26388 -16070 26454 -16036
rect 26454 -16070 26488 -16036
rect 26488 -16070 26574 -16036
rect 25882 -16156 26574 -16070
rect 25882 -16823 26574 -16751
rect 25882 -16858 25954 -16823
rect 25954 -16858 25988 -16823
rect 25988 -16858 26054 -16823
rect 26054 -16858 26088 -16823
rect 26088 -16858 26154 -16823
rect 26154 -16858 26188 -16823
rect 26188 -16858 26254 -16823
rect 26254 -16858 26288 -16823
rect 26288 -16858 26354 -16823
rect 26354 -16858 26388 -16823
rect 26388 -16858 26454 -16823
rect 26454 -16858 26488 -16823
rect 26488 -16858 26574 -16823
rect 25882 -16923 26574 -16858
rect 25882 -16958 25954 -16923
rect 25954 -16958 25988 -16923
rect 25988 -16958 26054 -16923
rect 26054 -16958 26088 -16923
rect 26088 -16958 26154 -16923
rect 26154 -16958 26188 -16923
rect 26188 -16958 26254 -16923
rect 26254 -16958 26288 -16923
rect 26288 -16958 26354 -16923
rect 26354 -16958 26388 -16923
rect 26388 -16958 26454 -16923
rect 26454 -16958 26488 -16923
rect 26488 -16958 26574 -16923
rect 25882 -17023 26574 -16958
rect 25882 -17058 25954 -17023
rect 25954 -17058 25988 -17023
rect 25988 -17058 26054 -17023
rect 26054 -17058 26088 -17023
rect 26088 -17058 26154 -17023
rect 26154 -17058 26188 -17023
rect 26188 -17058 26254 -17023
rect 26254 -17058 26288 -17023
rect 26288 -17058 26354 -17023
rect 26354 -17058 26388 -17023
rect 26388 -17058 26454 -17023
rect 26454 -17058 26488 -17023
rect 26488 -17058 26574 -17023
rect 25882 -17123 26574 -17058
rect 25882 -17158 25954 -17123
rect 25954 -17158 25988 -17123
rect 25988 -17158 26054 -17123
rect 26054 -17158 26088 -17123
rect 26088 -17158 26154 -17123
rect 26154 -17158 26188 -17123
rect 26188 -17158 26254 -17123
rect 26254 -17158 26288 -17123
rect 26288 -17158 26354 -17123
rect 26354 -17158 26388 -17123
rect 26388 -17158 26454 -17123
rect 26454 -17158 26488 -17123
rect 26488 -17158 26574 -17123
rect 25882 -17223 26574 -17158
rect 25882 -17258 25954 -17223
rect 25954 -17258 25988 -17223
rect 25988 -17258 26054 -17223
rect 26054 -17258 26088 -17223
rect 26088 -17258 26154 -17223
rect 26154 -17258 26188 -17223
rect 26188 -17258 26254 -17223
rect 26254 -17258 26288 -17223
rect 26288 -17258 26354 -17223
rect 26354 -17258 26388 -17223
rect 26388 -17258 26454 -17223
rect 26454 -17258 26488 -17223
rect 26488 -17258 26574 -17223
rect 25882 -17323 26574 -17258
rect 25882 -17358 25954 -17323
rect 25954 -17358 25988 -17323
rect 25988 -17358 26054 -17323
rect 26054 -17358 26088 -17323
rect 26088 -17358 26154 -17323
rect 26154 -17358 26188 -17323
rect 26188 -17358 26254 -17323
rect 26254 -17358 26288 -17323
rect 26288 -17358 26354 -17323
rect 26354 -17358 26388 -17323
rect 26388 -17358 26454 -17323
rect 26454 -17358 26488 -17323
rect 26488 -17358 26574 -17323
rect 25882 -17443 26574 -17358
rect 6076 -18662 6634 -18104
rect 5276 -20298 5834 -19740
rect 6876 -18114 7296 -18104
rect 6876 -18652 6888 -18114
rect 6888 -18652 7285 -18114
rect 7285 -18652 7296 -18114
rect 6876 -18662 7296 -18652
rect 13612 -18114 14304 -18048
rect 13612 -18652 13623 -18114
rect 13623 -18652 14020 -18114
rect 14020 -18652 14304 -18114
rect 13612 -18740 14304 -18652
rect 6876 -18932 7296 -18922
rect 6876 -19470 6888 -18932
rect 6888 -19470 7285 -18932
rect 7285 -19470 7296 -18932
rect 6876 -19480 7296 -19470
rect 7538 -19480 8096 -18922
rect 6876 -19750 7296 -19740
rect 6876 -20288 6888 -19750
rect 6888 -20288 7285 -19750
rect 7285 -20288 7296 -19750
rect 6876 -20298 7296 -20288
rect 6076 -21116 6634 -20558
rect 6876 -20568 7296 -20558
rect 6876 -21106 6888 -20568
rect 6888 -21106 7285 -20568
rect 7285 -21106 7296 -20568
rect 6876 -21116 7296 -21106
rect 6876 -21386 7296 -21376
rect 6876 -21924 6888 -21386
rect 6888 -21924 7285 -21386
rect 7285 -21924 7296 -21386
rect 6876 -21934 7296 -21924
rect 13612 -18932 14304 -18866
rect 13612 -19470 13623 -18932
rect 13623 -19470 14020 -18932
rect 14020 -19470 14304 -18932
rect 13612 -19558 14304 -19470
rect 20730 -19558 21422 -18866
rect 13612 -19750 14304 -19684
rect 13612 -20288 13623 -19750
rect 13623 -20288 14020 -19750
rect 14020 -20288 14304 -19750
rect 13612 -20376 14304 -20288
rect 7538 -21934 8096 -21376
rect 12012 -21116 12570 -20558
rect 5276 -22752 5834 -22194
rect 6876 -22204 7296 -22194
rect 6876 -22742 6888 -22204
rect 6888 -22742 7285 -22204
rect 7285 -22742 7296 -22204
rect 6876 -22752 7296 -22742
rect 6076 -23570 6634 -23012
rect 6876 -23022 7296 -23012
rect 6876 -23560 6888 -23022
rect 6888 -23560 7285 -23022
rect 7285 -23560 7296 -23022
rect 6876 -23570 7296 -23560
rect 13612 -20568 14032 -20558
rect 13612 -21106 13623 -20568
rect 13623 -21106 14020 -20568
rect 14020 -21106 14032 -20568
rect 13612 -21116 14032 -21106
rect 16162 -20900 16680 -19966
rect 25640 -20902 26576 -19966
rect 13612 -21386 14032 -21376
rect 13612 -21924 13623 -21386
rect 13623 -21924 14021 -21386
rect 14021 -21924 14032 -21386
rect 13612 -21934 14032 -21924
rect 14274 -21934 14832 -21376
rect 12012 -23570 12570 -23012
rect 12812 -22752 13370 -22194
rect 6876 -23840 7296 -23830
rect 6876 -24378 6888 -23840
rect 6888 -24378 7285 -23840
rect 7285 -24378 7296 -23840
rect 6876 -24388 7296 -24378
rect 6876 -24658 7296 -24648
rect 6876 -25196 6888 -24658
rect 6888 -25196 7285 -24658
rect 7285 -25196 7296 -24658
rect 6876 -25206 7296 -25196
rect 7538 -25206 8096 -24648
rect 6076 -26024 6634 -25466
rect 6876 -25476 7296 -25466
rect 6876 -26014 6888 -25476
rect 6888 -26014 7285 -25476
rect 7285 -26014 7296 -25476
rect 6876 -26024 7296 -26014
rect 5276 -26842 5834 -26284
rect 6876 -26294 7296 -26284
rect 6876 -26832 6888 -26294
rect 6888 -26832 7285 -26294
rect 7285 -26832 7296 -26294
rect 6876 -26842 7296 -26832
rect 6876 -27112 7296 -27102
rect 6876 -27650 6888 -27112
rect 6888 -27650 7285 -27112
rect 7285 -27650 7296 -27112
rect 6876 -27660 7296 -27650
rect 7538 -27660 8096 -27102
rect 12012 -26024 12570 -25466
rect 5276 -28466 5834 -27908
rect 6876 -27930 7296 -27920
rect 6876 -28468 6888 -27930
rect 6888 -28468 7285 -27930
rect 7285 -28468 7296 -27930
rect 6876 -28478 7296 -28468
rect 6076 -29296 6634 -28738
rect 6876 -28748 7296 -28738
rect 6876 -29286 6888 -28748
rect 6888 -29286 7285 -28748
rect 7285 -29286 7296 -28748
rect 6876 -29296 7296 -29286
rect 13612 -22204 14032 -22194
rect 13612 -22742 13623 -22204
rect 13623 -22742 14020 -22204
rect 14020 -22742 14032 -22204
rect 13612 -22752 14032 -22742
rect 13612 -23022 14032 -23012
rect 13612 -23560 13623 -23022
rect 13623 -23560 14020 -23022
rect 14020 -23560 14032 -23022
rect 13612 -23570 14032 -23560
rect 13644 -23830 14162 -23774
rect 13612 -23840 14162 -23830
rect 13612 -24378 13623 -23840
rect 13623 -24378 14020 -23840
rect 14020 -24378 14162 -23840
rect 13612 -24388 14162 -24378
rect 13644 -24466 14162 -24388
rect 13612 -24658 14032 -24648
rect 13612 -25196 13623 -24658
rect 13623 -25196 14021 -24658
rect 14021 -25196 14032 -24658
rect 13612 -25206 14032 -25196
rect 14274 -25206 14832 -24648
rect 13612 -25476 14032 -25466
rect 13612 -26014 13623 -25476
rect 13623 -26014 14020 -25476
rect 14020 -26014 14032 -25476
rect 13612 -26024 14032 -26014
rect 12812 -26842 13370 -26284
rect 13612 -26294 14032 -26284
rect 13612 -26832 13623 -26294
rect 13623 -26832 14020 -26294
rect 14020 -26832 14032 -26294
rect 13612 -26842 14032 -26832
rect 13612 -27112 14032 -27102
rect 13612 -27650 13623 -27112
rect 13623 -27650 14021 -27112
rect 14021 -27650 14032 -27112
rect 13612 -27660 14032 -27650
rect 14274 -27660 14832 -27102
rect 12012 -29296 12570 -28738
rect 12812 -28478 13370 -27920
rect 6876 -29566 7296 -29556
rect 6876 -30104 6888 -29566
rect 6888 -30104 7285 -29566
rect 7285 -30104 7296 -29566
rect 6876 -30114 7296 -30104
rect 7538 -30114 8096 -29556
rect 6814 -33656 7234 -33646
rect 6814 -34194 6826 -33656
rect 6826 -34194 7223 -33656
rect 7223 -34194 7234 -33656
rect 6814 -34204 7234 -34194
rect 7538 -34204 8030 -33646
rect 6076 -35022 6634 -34464
rect 6814 -34474 7234 -34464
rect 6814 -35012 6826 -34474
rect 6826 -35012 7223 -34474
rect 7223 -35012 7234 -34474
rect 6814 -35022 7234 -35012
rect 13612 -27930 14032 -27920
rect 13612 -28468 13623 -27930
rect 13623 -28468 14020 -27930
rect 14020 -28468 14032 -27930
rect 13612 -28478 14032 -28468
rect 13612 -28748 14032 -28738
rect 13612 -29286 13623 -28748
rect 13623 -29286 14020 -28748
rect 14020 -29286 14032 -28748
rect 13612 -29296 14032 -29286
rect 13612 -29566 14032 -29556
rect 13612 -30104 13623 -29566
rect 13623 -30104 14021 -29566
rect 14021 -30104 14032 -29566
rect 13612 -30114 14032 -30104
rect 14274 -30114 14832 -29556
<< metal2 >>
rect 20724 -14176 21428 -14170
rect 20724 -14868 20730 -14176
rect 21422 -14868 21428 -14176
rect 13606 -18048 14310 -18042
rect 6070 -18104 7302 -18098
rect 6070 -18662 6076 -18104
rect 6634 -18662 6876 -18104
rect 7296 -18662 7302 -18104
rect 13606 -18110 13612 -18048
rect 6070 -18668 7302 -18662
rect 9732 -18680 13612 -18110
rect 6870 -18922 8102 -18916
rect 6870 -19480 6876 -18922
rect 7296 -19480 7538 -18922
rect 8096 -19480 8102 -18922
rect 6870 -19486 8102 -19480
rect 5270 -19740 7302 -19734
rect 5270 -20298 5276 -19740
rect 5834 -20298 6876 -19740
rect 7296 -20298 7302 -19740
rect 5840 -20304 7302 -20298
rect 6070 -20558 7302 -20552
rect 6070 -21116 6076 -20558
rect 6634 -21116 6876 -20558
rect 7296 -21116 7302 -20558
rect 6070 -21122 7302 -21116
rect 6870 -21376 8102 -21370
rect 6870 -21934 6876 -21376
rect 7296 -21934 7538 -21376
rect 8096 -21934 8102 -21376
rect 6870 -21940 8102 -21934
rect 5270 -22194 7302 -22188
rect 5270 -22752 5276 -22194
rect 5834 -22752 6876 -22194
rect 7296 -22752 7302 -22194
rect 5270 -22758 7302 -22752
rect 6070 -23012 7302 -23006
rect 6070 -23570 6076 -23012
rect 6634 -23570 6876 -23012
rect 7296 -23570 7302 -23012
rect 6070 -23576 7302 -23570
rect 9732 -23824 10302 -18680
rect 13606 -18740 13612 -18680
rect 14304 -18740 14310 -18048
rect 13606 -18746 14310 -18740
rect 13606 -18866 14304 -18860
rect 13606 -19558 13612 -18866
rect 13606 -19564 14304 -19558
rect 20724 -18866 21428 -14868
rect 25876 -15464 26580 -15458
rect 25876 -16156 25882 -15464
rect 26574 -15470 26580 -15464
rect 26574 -16156 26582 -15470
rect 25876 -16162 26582 -16156
rect 25902 -16745 26582 -16162
rect 25876 -16751 26582 -16745
rect 25876 -17443 25882 -16751
rect 26574 -17443 26582 -16751
rect 25876 -17449 26582 -17443
rect 20724 -19558 20730 -18866
rect 21422 -19558 21428 -18866
rect 20724 -19564 21428 -19558
rect 13606 -19684 14310 -19678
rect 13606 -20376 13612 -19684
rect 14304 -20376 14310 -19684
rect 13606 -20382 14310 -20376
rect 16156 -19966 16686 -19960
rect 25902 -19966 26582 -17449
rect 12006 -20558 14038 -20552
rect 12006 -21116 12012 -20558
rect 12570 -21116 13612 -20558
rect 14032 -21116 14038 -20558
rect 12006 -21122 14038 -21116
rect 16156 -20900 16162 -19966
rect 16680 -20900 16686 -19966
rect 13606 -21376 14838 -21370
rect 13606 -21934 13612 -21376
rect 14032 -21934 14274 -21376
rect 14832 -21934 14838 -21376
rect 13606 -21940 14838 -21934
rect 12806 -22194 14038 -22188
rect 12806 -22752 12812 -22194
rect 13370 -22752 13612 -22194
rect 14032 -22752 14038 -22194
rect 12806 -22758 14038 -22752
rect 12006 -23012 14038 -23006
rect 12006 -23570 12012 -23012
rect 12570 -23570 13612 -23012
rect 14032 -23570 14038 -23012
rect 12006 -23576 14038 -23570
rect 13644 -23770 14910 -23768
rect 16156 -23770 16686 -20900
rect 25634 -20902 25640 -19966
rect 26576 -20902 26582 -19966
rect 25634 -20908 26582 -20902
rect 13644 -23774 16686 -23770
rect 6870 -23830 10302 -23824
rect 6870 -24388 6876 -23830
rect 7296 -24388 10302 -23830
rect 6870 -24394 10302 -24388
rect 13606 -23830 13644 -23824
rect 13606 -24388 13612 -23830
rect 13606 -24394 13644 -24388
rect 14162 -24466 16686 -23774
rect 13644 -24472 16686 -24466
rect 6870 -24648 8102 -24642
rect 6870 -25206 6876 -24648
rect 7296 -25206 7538 -24648
rect 8096 -25206 8102 -24648
rect 6870 -25212 8102 -25206
rect 13606 -24648 14832 -24642
rect 13606 -25206 13612 -24648
rect 14032 -25206 14274 -24648
rect 14832 -25206 14838 -24648
rect 13606 -25212 14838 -25206
rect 6070 -25466 7302 -25460
rect 6070 -26024 6076 -25466
rect 6634 -26024 6876 -25466
rect 7296 -26024 7302 -25466
rect 6070 -26030 7302 -26024
rect 12006 -25466 14038 -25460
rect 12006 -26024 12012 -25466
rect 12570 -26024 13612 -25466
rect 14032 -26024 14038 -25466
rect 12006 -26030 14038 -26024
rect 5270 -26284 7302 -26278
rect 5270 -26842 5276 -26284
rect 5834 -26842 6876 -26284
rect 7296 -26842 7302 -26284
rect 5270 -26848 7302 -26842
rect 12806 -26284 14038 -26278
rect 12806 -26842 12812 -26284
rect 13370 -26842 13612 -26284
rect 14032 -26842 14038 -26284
rect 12806 -26848 14038 -26842
rect 6870 -27102 8102 -27096
rect 6870 -27660 6876 -27102
rect 7296 -27660 7538 -27102
rect 8096 -27660 8102 -27102
rect 6870 -27666 8102 -27660
rect 13606 -27102 14832 -27096
rect 13606 -27660 13612 -27102
rect 14032 -27660 14274 -27102
rect 14832 -27660 14838 -27102
rect 13606 -27666 14838 -27660
rect 5270 -27908 7284 -27902
rect 5270 -28466 5276 -27908
rect 5834 -27914 7284 -27908
rect 5834 -27920 7302 -27914
rect 5834 -28466 6876 -27920
rect 5270 -28472 6876 -28466
rect 6870 -28478 6876 -28472
rect 7296 -28478 7302 -27920
rect 6870 -28484 7302 -28478
rect 12806 -27920 14038 -27914
rect 12806 -28478 12812 -27920
rect 13370 -28478 13612 -27920
rect 14032 -28478 14038 -27920
rect 12806 -28484 14038 -28478
rect 6070 -28738 7302 -28732
rect 6070 -29296 6076 -28738
rect 6634 -29296 6876 -28738
rect 7296 -29296 7302 -28738
rect 6070 -29302 7302 -29296
rect 12006 -28738 14038 -28732
rect 12006 -29296 12012 -28738
rect 12570 -29296 13612 -28738
rect 14032 -29296 14038 -28738
rect 12006 -29302 14038 -29296
rect 6870 -29556 8102 -29550
rect 6870 -30114 6876 -29556
rect 7296 -30114 7538 -29556
rect 8096 -30114 8102 -29556
rect 6870 -30120 8102 -30114
rect 13606 -29556 14832 -29550
rect 13606 -30114 13612 -29556
rect 14032 -30114 14274 -29556
rect 14832 -30114 14838 -29556
rect 13606 -30120 14838 -30114
rect 6808 -33646 8040 -33640
rect 6808 -34204 6814 -33646
rect 7234 -34204 7538 -33646
rect 8030 -34204 8040 -33646
rect 6808 -34210 8040 -34204
rect 6070 -34464 7240 -34458
rect 6070 -35022 6076 -34464
rect 6634 -35022 6814 -34464
rect 7234 -35022 7240 -34464
rect 6070 -35028 7240 -35022
<< res2p85 >>
rect 7300 -17852 13608 -17278
rect 7300 -18670 13608 -18096
rect 7300 -19488 13608 -18914
rect 7300 -20306 13608 -19732
rect 7300 -21124 13608 -20550
rect 7300 -21942 13608 -21368
rect 7300 -22760 13608 -22186
rect 7300 -23578 13608 -23004
rect 7300 -24396 13608 -23822
rect 7300 -25214 13608 -24640
rect 7300 -26032 13608 -25458
rect 7300 -26850 13608 -26276
rect 7300 -27668 13608 -27094
rect 7300 -28486 13608 -27912
rect 7300 -29304 13608 -28730
rect 7300 -30122 13608 -29548
rect 7300 -30940 13608 -30366
rect 7238 -33394 11542 -32820
rect 7238 -34212 11542 -33638
rect 7238 -35030 11542 -34456
rect 7238 -35848 11542 -35274
rect 8624 -37484 11952 -36910
rect 8624 -38302 11952 -37728
rect 8624 -39120 11952 -38546
<< labels >>
flabel metal2 6870 -29302 7302 -28732 7 FreeSans 800 90 0 0 VbEnd
flabel metal2 13606 -28484 14038 -27914 7 FreeSans 800 90 0 0 VbgEnd
flabel metal2 6870 -30120 8102 -29550 7 FreeSans 800 90 0 0 VaEnd
flabel metal2 13612 -20376 14304 -19684 7 FreeSans 1600 90 0 0 Vbg
port 3 n
flabel metal2 13606 -18746 14310 -18042 7 FreeSans 1600 90 0 0 Vb
port 1 n
flabel metal1 14304 -19564 14876 -18860 1 FreeSans 1600 0 0 0 Va
port 5 n
flabel metal1 12028 -35032 12470 -33566 1 FreeSans 1600 0 0 0 GND!
port 6 n
flabel locali 17168 -12078 17272 -11830 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,0]/Emitter
flabel locali 17794 -11990 17843 -11889 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,0]/Collector
flabel locali 17644 -11984 17684 -11866 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,0]/Base
flabel locali 17168 -13366 17272 -13118 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,1]/Emitter
flabel locali 17794 -13278 17843 -13177 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,1]/Collector
flabel locali 17644 -13272 17684 -13154 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,1]/Base
flabel locali 17168 -14654 17272 -14406 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,2]/Emitter
flabel locali 17794 -14566 17843 -14465 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,2]/Collector
flabel locali 17644 -14560 17684 -14442 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,2]/Base
flabel locali 17168 -15942 17272 -15694 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,3]/Emitter
flabel locali 17794 -15854 17843 -15753 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,3]/Collector
flabel locali 17644 -15848 17684 -15730 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,3]/Base
flabel locali 17168 -17230 17272 -16982 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,4]/Emitter
flabel locali 17794 -17142 17843 -17041 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,4]/Collector
flabel locali 17644 -17136 17684 -17018 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,4]/Base
flabel locali 18456 -12078 18560 -11830 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,0]/Emitter
flabel locali 19082 -11990 19131 -11889 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,0]/Collector
flabel locali 18932 -11984 18972 -11866 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,0]/Base
flabel locali 18456 -13366 18560 -13118 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,1]/Emitter
flabel locali 19082 -13278 19131 -13177 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,1]/Collector
flabel locali 18932 -13272 18972 -13154 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,1]/Base
flabel locali 18456 -14654 18560 -14406 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,2]/Emitter
flabel locali 19082 -14566 19131 -14465 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,2]/Collector
flabel locali 18932 -14560 18972 -14442 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,2]/Base
flabel locali 18456 -15942 18560 -15694 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,3]/Emitter
flabel locali 19082 -15854 19131 -15753 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,3]/Collector
flabel locali 18932 -15848 18972 -15730 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,3]/Base
flabel locali 18456 -17230 18560 -16982 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,4]/Emitter
flabel locali 19082 -17142 19131 -17041 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,4]/Collector
flabel locali 18932 -17136 18972 -17018 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,4]/Base
flabel locali 19744 -12078 19848 -11830 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,0]/Emitter
flabel locali 20370 -11990 20419 -11889 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,0]/Collector
flabel locali 20220 -11984 20260 -11866 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,0]/Base
flabel locali 19744 -13366 19848 -13118 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,1]/Emitter
flabel locali 20370 -13278 20419 -13177 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,1]/Collector
flabel locali 20220 -13272 20260 -13154 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,1]/Base
flabel locali 19744 -14654 19848 -14406 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,2]/Emitter
flabel locali 20370 -14566 20419 -14465 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,2]/Collector
flabel locali 20220 -14560 20260 -14442 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,2]/Base
flabel locali 19744 -15942 19848 -15694 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,3]/Emitter
flabel locali 20370 -15854 20419 -15753 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,3]/Collector
flabel locali 20220 -15848 20260 -15730 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,3]/Base
flabel locali 19744 -17230 19848 -16982 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,4]/Emitter
flabel locali 20370 -17142 20419 -17041 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,4]/Collector
flabel locali 20220 -17136 20260 -17018 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,4]/Base
flabel locali 21032 -12078 21136 -11830 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,0]/Emitter
flabel locali 21658 -11990 21707 -11889 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,0]/Collector
flabel locali 21508 -11984 21548 -11866 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,0]/Base
flabel locali 21032 -13366 21136 -13118 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,1]/Emitter
flabel locali 21658 -13278 21707 -13177 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,1]/Collector
flabel locali 21508 -13272 21548 -13154 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,1]/Base
flabel locali 21032 -14654 21136 -14406 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,2]/Emitter
flabel locali 21658 -14566 21707 -14465 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,2]/Collector
flabel locali 21508 -14560 21548 -14442 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,2]/Base
flabel locali 21032 -15942 21136 -15694 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,3]/Emitter
flabel locali 21658 -15854 21707 -15753 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,3]/Collector
flabel locali 21508 -15848 21548 -15730 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,3]/Base
flabel locali 21032 -17230 21136 -16982 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,4]/Emitter
flabel locali 21658 -17142 21707 -17041 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,4]/Collector
flabel locali 21508 -17136 21548 -17018 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,4]/Base
flabel locali 22320 -12078 22424 -11830 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,0]/Emitter
flabel locali 22946 -11990 22995 -11889 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,0]/Collector
flabel locali 22796 -11984 22836 -11866 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,0]/Base
flabel locali 22320 -13366 22424 -13118 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,1]/Emitter
flabel locali 22946 -13278 22995 -13177 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,1]/Collector
flabel locali 22796 -13272 22836 -13154 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,1]/Base
flabel locali 22320 -14654 22424 -14406 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,2]/Emitter
flabel locali 22946 -14566 22995 -14465 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,2]/Collector
flabel locali 22796 -14560 22836 -14442 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,2]/Base
flabel locali 22320 -15942 22424 -15694 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,3]/Emitter
flabel locali 22946 -15854 22995 -15753 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,3]/Collector
flabel locali 22796 -15848 22836 -15730 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,3]/Base
flabel locali 22320 -17230 22424 -16982 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,4]/Emitter
flabel locali 22946 -17142 22995 -17041 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,4]/Collector
flabel locali 22796 -17136 22836 -17018 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,4]/Base
flabel locali 23608 -12078 23712 -11830 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,0]/Emitter
flabel locali 24234 -11990 24283 -11889 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,0]/Collector
flabel locali 24084 -11984 24124 -11866 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,0]/Base
flabel locali 23608 -13366 23712 -13118 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,1]/Emitter
flabel locali 24234 -13278 24283 -13177 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,1]/Collector
flabel locali 24084 -13272 24124 -13154 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,1]/Base
flabel locali 23608 -14654 23712 -14406 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,2]/Emitter
flabel locali 24234 -14566 24283 -14465 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,2]/Collector
flabel locali 24084 -14560 24124 -14442 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,2]/Base
flabel locali 23608 -15942 23712 -15694 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,3]/Emitter
flabel locali 24234 -15854 24283 -15753 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,3]/Collector
flabel locali 24084 -15848 24124 -15730 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,3]/Base
flabel locali 23608 -17230 23712 -16982 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,4]/Emitter
flabel locali 24234 -17142 24283 -17041 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,4]/Collector
flabel locali 24084 -17136 24124 -17018 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,4]/Base
flabel locali 24896 -12078 25000 -11830 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,0]/Emitter
flabel locali 25522 -11990 25571 -11889 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,0]/Collector
flabel locali 25372 -11984 25412 -11866 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,0]/Base
flabel locali 24896 -13366 25000 -13118 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,1]/Emitter
flabel locali 25522 -13278 25571 -13177 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,1]/Collector
flabel locali 25372 -13272 25412 -13154 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,1]/Base
flabel locali 24896 -14654 25000 -14406 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,2]/Emitter
flabel locali 25522 -14566 25571 -14465 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,2]/Collector
flabel locali 25372 -14560 25412 -14442 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,2]/Base
flabel locali 24896 -15942 25000 -15694 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,3]/Emitter
flabel locali 25522 -15854 25571 -15753 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,3]/Collector
flabel locali 25372 -15848 25412 -15730 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,3]/Base
flabel locali 24896 -17230 25000 -16982 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,4]/Emitter
flabel locali 25522 -17142 25571 -17041 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,4]/Collector
flabel locali 25372 -17136 25412 -17018 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,4]/Base
flabel locali 26184 -12078 26288 -11830 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,0]/Emitter
flabel locali 26810 -11990 26859 -11889 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,0]/Collector
flabel locali 26660 -11984 26700 -11866 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,0]/Base
flabel locali 26184 -13366 26288 -13118 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,1]/Emitter
flabel locali 26810 -13278 26859 -13177 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,1]/Collector
flabel locali 26660 -13272 26700 -13154 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,1]/Base
flabel locali 26184 -14654 26288 -14406 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,2]/Emitter
flabel locali 26810 -14566 26859 -14465 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,2]/Collector
flabel locali 26660 -14560 26700 -14442 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,2]/Base
flabel locali 26184 -15942 26288 -15694 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,3]/Emitter
flabel locali 26810 -15854 26859 -15753 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,3]/Collector
flabel locali 26660 -15848 26700 -15730 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,3]/Base
flabel locali 26184 -17230 26288 -16982 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,4]/Emitter
flabel locali 26810 -17142 26859 -17041 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,4]/Collector
flabel locali 26660 -17136 26700 -17018 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,4]/Base
flabel locali 26184 -17229 26288 -16981 0 FreeSans 400 0 0 0 sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,3]/Emitter
flabel metal2 25902 -19966 26582 -17443 1 FreeSans 1600 0 0 0 Vbneg
<< end >>
