magic
tech sky130A
magscale 1 2
timestamp 1620938299
<< psubdiff >>
rect 12480 6690 12998 6714
rect 12480 6504 12504 6690
rect 12974 6504 12998 6690
rect 12480 6480 12998 6504
<< psubdiffcont >>
rect 12504 6504 12974 6690
<< xpolycontact >>
rect 8502 6600 8572 7032
rect 9302 6600 9372 7032
rect 10102 6600 10172 7032
rect 10502 6600 10572 7032
rect 10902 6600 10972 7032
rect 12102 6600 12172 7032
<< viali >>
rect 8518 6618 8556 7015
rect 9318 6618 9356 7015
rect 10118 6618 10156 7015
rect 10518 6618 10556 7015
rect 10918 6618 10956 7015
rect 12118 6618 12156 7015
rect 12488 6690 12990 6706
rect 12488 6504 12504 6690
rect 12504 6504 12974 6690
rect 12974 6504 12990 6690
rect 12488 6488 12990 6504
<< metal1 >>
rect 8102 8196 8172 8216
rect 8102 8144 8108 8196
rect 8160 8144 8172 8196
rect 8102 7784 8172 8144
rect 8502 7864 8572 8216
rect 8502 7812 8508 7864
rect 8560 7812 8572 7864
rect 8502 7784 8572 7812
rect 8902 8196 8972 8216
rect 8902 8144 8908 8196
rect 8960 8144 8972 8196
rect 8902 7784 8972 8144
rect 9302 7864 9372 8216
rect 9302 7812 9308 7864
rect 9360 7812 9372 7864
rect 9302 7784 9372 7812
rect 9702 8196 9772 8216
rect 9702 8144 9708 8196
rect 9760 8144 9772 8196
rect 9702 7784 9772 8144
rect 10102 7864 10172 8216
rect 10102 7812 10108 7864
rect 10160 7812 10172 7864
rect 10102 7784 10172 7812
rect 10502 8196 10572 8216
rect 10502 8144 10508 8196
rect 10560 8144 10572 8196
rect 10502 7784 10572 8144
rect 10902 7864 10972 8216
rect 10902 7812 10908 7864
rect 10960 7812 10972 7864
rect 10902 7784 10972 7812
rect 8502 7448 8572 7468
rect 8502 7396 8510 7448
rect 8562 7396 8572 7448
rect 8102 5900 8172 7032
rect 8502 7015 8572 7396
rect 11302 7448 11372 8216
rect 11702 8196 11772 8216
rect 11702 8144 11708 8196
rect 11760 8144 11772 8196
rect 11702 7784 11772 8144
rect 12102 7864 12172 8216
rect 12102 7812 12108 7864
rect 12160 7812 12172 7864
rect 12102 7784 12172 7812
rect 12504 8196 12574 8202
rect 12504 8144 12510 8196
rect 12562 8144 12574 8196
rect 12504 7754 12574 8144
rect 12904 7864 12974 8186
rect 12904 7812 12910 7864
rect 12962 7812 12974 7864
rect 12904 7754 12974 7812
rect 11302 7396 11308 7448
rect 11360 7396 11372 7448
rect 11302 7368 11372 7396
rect 12504 7032 12974 7248
rect 8502 6618 8518 7015
rect 8556 6618 8572 7015
rect 8502 6492 8572 6618
rect 8902 6680 8972 7032
rect 8902 6628 8908 6680
rect 8960 6628 8972 6680
rect 8902 6600 8972 6628
rect 9302 7015 9372 7032
rect 9302 7012 9318 7015
rect 9356 7012 9372 7015
rect 9302 6952 9308 7012
rect 9360 6952 9372 7012
rect 9302 6618 9318 6952
rect 9356 6618 9372 6952
rect 9302 6600 9372 6618
rect 9702 6680 9772 7032
rect 9702 6628 9708 6680
rect 9760 6628 9772 6680
rect 9702 6600 9772 6628
rect 10102 7015 10172 7032
rect 10102 7012 10118 7015
rect 10156 7012 10172 7015
rect 10102 6960 10108 7012
rect 10160 6960 10172 7012
rect 10102 6618 10118 6960
rect 10156 6618 10172 6960
rect 10102 6600 10172 6618
rect 10502 7015 10572 7032
rect 10502 6672 10518 7015
rect 10556 6672 10572 7015
rect 10502 6620 10508 6672
rect 10560 6620 10572 6672
rect 10502 6618 10518 6620
rect 10556 6618 10572 6620
rect 10502 6600 10572 6618
rect 10902 7015 10972 7032
rect 10902 7012 10918 7015
rect 10956 7012 10972 7015
rect 10902 6960 10908 7012
rect 10960 6960 10972 7012
rect 10902 6618 10918 6960
rect 10956 6618 10972 6960
rect 10902 6600 10972 6618
rect 11302 6500 11372 7032
rect 11702 6680 11772 7032
rect 11702 6628 11708 6680
rect 11760 6628 11772 6680
rect 11702 6600 11772 6628
rect 12102 7015 12172 7032
rect 12102 7012 12118 7015
rect 12156 7012 12172 7015
rect 12102 6960 12108 7012
rect 12160 6960 12172 7012
rect 12102 6618 12118 6960
rect 12156 6618 12172 6960
rect 12504 6720 13272 7032
rect 12102 6600 12172 6618
rect 12474 6706 13272 6720
rect 8444 6486 8630 6492
rect 8444 6300 8450 6486
rect 8624 6300 8630 6486
rect 8444 6294 8630 6300
rect 8102 5686 9400 5900
rect 8102 5500 8450 5686
rect 8624 5500 9400 5686
rect 8102 5302 9400 5500
rect 11000 5302 11700 6500
rect 12474 6488 12488 6706
rect 12990 6600 13272 6706
rect 12990 6488 13004 6600
rect 12474 6474 13004 6488
<< via1 >>
rect 8108 8144 8160 8196
rect 8508 7812 8560 7864
rect 8908 8144 8960 8196
rect 9308 7812 9360 7864
rect 9708 8144 9760 8196
rect 10108 7812 10160 7864
rect 10508 8144 10560 8196
rect 10908 7812 10960 7864
rect 8510 7396 8562 7448
rect 11708 8144 11760 8196
rect 12108 7812 12160 7864
rect 12510 8144 12562 8196
rect 12910 7812 12962 7864
rect 11308 7396 11360 7448
rect 8908 6628 8960 6680
rect 9308 6952 9318 7012
rect 9318 6952 9356 7012
rect 9356 6952 9360 7012
rect 9708 6628 9760 6680
rect 10108 6960 10118 7012
rect 10118 6960 10156 7012
rect 10156 6960 10160 7012
rect 10508 6620 10518 6672
rect 10518 6620 10556 6672
rect 10556 6620 10560 6672
rect 10908 6960 10918 7012
rect 10918 6960 10956 7012
rect 10956 6960 10960 7012
rect 11708 6628 11760 6680
rect 12108 6960 12118 7012
rect 12118 6960 12156 7012
rect 12156 6960 12160 7012
rect 8450 6300 8624 6486
rect 8450 5500 8624 5686
<< metal2 >>
rect 8090 8196 8990 8216
rect 8090 8144 8108 8196
rect 8160 8144 8908 8196
rect 8960 8144 8990 8196
rect 8090 8116 8990 8144
rect 9690 8196 10590 8216
rect 9690 8144 9708 8196
rect 9760 8144 10508 8196
rect 10560 8144 10590 8196
rect 9690 8116 10590 8144
rect 11690 8196 12574 8216
rect 11690 8144 11708 8196
rect 11760 8144 12510 8196
rect 12562 8144 12574 8196
rect 11690 8116 12574 8144
rect 8490 7864 9390 7884
rect 8490 7812 8508 7864
rect 8560 7812 9308 7864
rect 9360 7812 9390 7864
rect 8490 7784 9390 7812
rect 10090 7864 10990 7884
rect 10090 7812 10108 7864
rect 10160 7812 10908 7864
rect 10960 7812 10990 7864
rect 10090 7784 10990 7812
rect 12090 7864 12974 7884
rect 12090 7812 12108 7864
rect 12160 7812 12910 7864
rect 12962 7812 12974 7864
rect 12090 7784 12974 7812
rect 8500 7448 11390 7468
rect 8500 7396 8510 7448
rect 8562 7396 11308 7448
rect 11360 7396 11390 7448
rect 8500 7368 11390 7396
rect 9290 7012 10190 7032
rect 9290 6952 9308 7012
rect 9360 6960 10108 7012
rect 10160 6960 10190 7012
rect 9360 6952 10190 6960
rect 9290 6932 10190 6952
rect 10890 7012 12190 7032
rect 10890 6960 10908 7012
rect 10960 6960 12108 7012
rect 12160 6960 12190 7012
rect 10890 6932 12190 6960
rect 8890 6680 9790 6700
rect 8890 6628 8908 6680
rect 8960 6628 9708 6680
rect 9760 6628 9790 6680
rect 8890 6600 9790 6628
rect 10502 6680 11790 6700
rect 10502 6672 11708 6680
rect 10502 6620 10508 6672
rect 10560 6628 11708 6672
rect 11760 6628 11790 6680
rect 10560 6620 11790 6628
rect 10502 6600 11790 6620
rect 8444 6486 8630 6492
rect 8444 6300 8450 6486
rect 8624 6300 8630 6486
rect 8444 6294 8630 6300
rect 8444 5686 8630 5692
rect 8444 5500 8450 5686
rect 8624 5500 8630 5686
rect 8444 5494 8630 5500
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_2
timestamp 1620883575
transform 1 0 8937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_3
timestamp 1620883575
transform 1 0 9337 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_3LWQVB  sky130_fd_pr__res_xhigh_po_0p35_3LWQVB_0
timestamp 1620936259
transform 1 0 8537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_3LWQVB  sky130_fd_pr__res_xhigh_po_0p35_3LWQVB_1
timestamp 1620936259
transform 1 0 8137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_5
timestamp 1620883575
transform 1 0 10137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_7
timestamp 1620883575
transform 1 0 10937 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_6
timestamp 1620883575
transform 1 0 10537 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_4
timestamp 1620883575
transform 1 0 9737 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_10
timestamp 1620883575
transform 1 0 12137 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_5SLMZ4  sky130_fd_pr__res_xhigh_po_0p35_5SLMZ4_1
timestamp 1620886403
transform 1 0 12939 0 1 7493
box -37 -677 37 677
use sky130_fd_pr__res_xhigh_po_0p35_5SLMZ4  sky130_fd_pr__res_xhigh_po_0p35_5SLMZ4_0
timestamp 1620886403
transform 1 0 12539 0 1 7493
box -37 -677 37 677
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_8
timestamp 1620883575
transform 1 0 11337 0 1 7408
box -37 -808 37 808
use sky130_fd_pr__res_xhigh_po_0p35_BNSLGU  sky130_fd_pr__res_xhigh_po_0p35_BNSLGU_9
timestamp 1620883575
transform 1 0 11737 0 1 7408
box -37 -808 37 808
<< labels >>
flabel metal1 8700 5500 9000 5800 1 FreeSans 1600 0 0 0 Va
port 1 n
flabel via1 8458 6304 8606 6468 1 FreeSans 1600 0 0 0 Vb
port 0 n
flabel metal1 11240 5360 11440 5580 1 FreeSans 800 0 0 0 Vbneg
flabel metal1 13056 6674 13196 6820 1 FreeSans 800 0 0 0 GND!
port 2 n
<< end >>
