magic
tech sky130A
timestamp 1621277573
<< error_p >>
rect -2359 1495 -2249 1725
rect -2800 1425 -2249 1495
rect -2239 1495 -2129 1725
rect -1798 1495 -1688 1725
rect -2239 1425 -1688 1495
rect -1678 1495 -1568 1725
rect -1237 1495 -1127 1725
rect -1678 1425 -1127 1495
rect -1117 1495 -1007 1725
rect -676 1495 -566 1725
rect -1117 1425 -566 1495
rect -556 1495 -446 1725
rect -115 1495 -5 1725
rect -556 1425 -5 1495
rect 5 1495 115 1725
rect 446 1495 556 1725
rect 5 1425 556 1495
rect 566 1495 676 1725
rect 1007 1495 1117 1725
rect 566 1425 1117 1495
rect 1127 1495 1237 1725
rect 1568 1495 1678 1725
rect 1127 1425 1678 1495
rect 1688 1495 1798 1725
rect 2129 1495 2239 1725
rect 1688 1425 2239 1495
rect 2249 1495 2359 1725
rect 2249 1425 2800 1495
rect -2800 1305 -2249 1375
rect -2359 1145 -2249 1305
rect -2800 1075 -2249 1145
rect -2239 1305 -1688 1375
rect -2239 1145 -2129 1305
rect -1798 1145 -1688 1305
rect -2239 1075 -1688 1145
rect -1678 1305 -1127 1375
rect -1678 1145 -1568 1305
rect -1237 1145 -1127 1305
rect -1678 1075 -1127 1145
rect -1117 1305 -566 1375
rect -1117 1145 -1007 1305
rect -676 1145 -566 1305
rect -1117 1075 -566 1145
rect -556 1305 -5 1375
rect -556 1145 -446 1305
rect -115 1145 -5 1305
rect -556 1075 -5 1145
rect 5 1305 556 1375
rect 5 1145 115 1305
rect 446 1145 556 1305
rect 5 1075 556 1145
rect 566 1305 1117 1375
rect 566 1145 676 1305
rect 1007 1145 1117 1305
rect 566 1075 1117 1145
rect 1127 1305 1678 1375
rect 1127 1145 1237 1305
rect 1568 1145 1678 1305
rect 1127 1075 1678 1145
rect 1688 1305 2239 1375
rect 1688 1145 1798 1305
rect 2129 1145 2239 1305
rect 1688 1075 2239 1145
rect 2249 1305 2800 1375
rect 2249 1145 2359 1305
rect 2249 1075 2800 1145
rect -2800 955 -2249 1025
rect -2359 795 -2249 955
rect -2800 725 -2249 795
rect -2239 955 -1688 1025
rect -2239 795 -2129 955
rect -1798 795 -1688 955
rect -2239 725 -1688 795
rect -1678 955 -1127 1025
rect -1678 795 -1568 955
rect -1237 795 -1127 955
rect -1678 725 -1127 795
rect -1117 955 -566 1025
rect -1117 795 -1007 955
rect -676 795 -566 955
rect -1117 725 -566 795
rect -556 955 -5 1025
rect -556 795 -446 955
rect -115 795 -5 955
rect -556 725 -5 795
rect 5 955 556 1025
rect 5 795 115 955
rect 446 795 556 955
rect 5 725 556 795
rect 566 955 1117 1025
rect 566 795 676 955
rect 1007 795 1117 955
rect 566 725 1117 795
rect 1127 955 1678 1025
rect 1127 795 1237 955
rect 1568 795 1678 955
rect 1127 725 1678 795
rect 1688 955 2239 1025
rect 1688 795 1798 955
rect 2129 795 2239 955
rect 1688 725 2239 795
rect 2249 955 2800 1025
rect 2249 795 2359 955
rect 2249 725 2800 795
rect -2800 605 -2249 675
rect -2359 445 -2249 605
rect -2800 375 -2249 445
rect -2239 605 -1688 675
rect -2239 445 -2129 605
rect -1798 445 -1688 605
rect -2239 375 -1688 445
rect -1678 605 -1127 675
rect -1678 445 -1568 605
rect -1237 445 -1127 605
rect -1678 375 -1127 445
rect -1117 605 -566 675
rect -1117 445 -1007 605
rect -676 445 -566 605
rect -1117 375 -566 445
rect -556 605 -5 675
rect -556 445 -446 605
rect -115 445 -5 605
rect -556 375 -5 445
rect 5 605 556 675
rect 5 445 115 605
rect 446 445 556 605
rect 5 375 556 445
rect 566 605 1117 675
rect 566 445 676 605
rect 1007 445 1117 605
rect 566 375 1117 445
rect 1127 605 1678 675
rect 1127 445 1237 605
rect 1568 445 1678 605
rect 1127 375 1678 445
rect 1688 605 2239 675
rect 1688 445 1798 605
rect 2129 445 2239 605
rect 1688 375 2239 445
rect 2249 605 2800 675
rect 2249 445 2359 605
rect 2249 375 2800 445
rect -2800 255 -2249 325
rect -2359 95 -2249 255
rect -2800 25 -2249 95
rect -2239 255 -1688 325
rect -2239 95 -2129 255
rect -1798 95 -1688 255
rect -2239 25 -1688 95
rect -1678 255 -1127 325
rect -1678 95 -1568 255
rect -1237 95 -1127 255
rect -1678 25 -1127 95
rect -1117 255 -566 325
rect -1117 95 -1007 255
rect -676 95 -566 255
rect -1117 25 -566 95
rect -556 255 -5 325
rect -556 95 -446 255
rect -115 95 -5 255
rect -556 25 -5 95
rect 5 255 556 325
rect 5 95 115 255
rect 446 95 556 255
rect 5 25 556 95
rect 566 255 1117 325
rect 566 95 676 255
rect 1007 95 1117 255
rect 566 25 1117 95
rect 1127 255 1678 325
rect 1127 95 1237 255
rect 1568 95 1678 255
rect 1127 25 1678 95
rect 1688 255 2239 325
rect 1688 95 1798 255
rect 2129 95 2239 255
rect 1688 25 2239 95
rect 2249 255 2800 325
rect 2249 95 2359 255
rect 2249 25 2800 95
rect -2800 -95 -2249 -25
rect -2359 -255 -2249 -95
rect -2800 -325 -2249 -255
rect -2239 -95 -1688 -25
rect -2239 -255 -2129 -95
rect -1798 -255 -1688 -95
rect -2239 -325 -1688 -255
rect -1678 -95 -1127 -25
rect -1678 -255 -1568 -95
rect -1237 -255 -1127 -95
rect -1678 -325 -1127 -255
rect -1117 -95 -566 -25
rect -1117 -255 -1007 -95
rect -676 -255 -566 -95
rect -1117 -325 -566 -255
rect -556 -95 -5 -25
rect -556 -255 -446 -95
rect -115 -255 -5 -95
rect -556 -325 -5 -255
rect 5 -95 556 -25
rect 5 -255 115 -95
rect 446 -255 556 -95
rect 5 -325 556 -255
rect 566 -95 1117 -25
rect 566 -255 676 -95
rect 1007 -255 1117 -95
rect 566 -325 1117 -255
rect 1127 -95 1678 -25
rect 1127 -255 1237 -95
rect 1568 -255 1678 -95
rect 1127 -325 1678 -255
rect 1688 -95 2239 -25
rect 1688 -255 1798 -95
rect 2129 -255 2239 -95
rect 1688 -325 2239 -255
rect 2249 -95 2800 -25
rect 2249 -255 2359 -95
rect 2249 -325 2800 -255
rect -2800 -445 -2249 -375
rect -2359 -605 -2249 -445
rect -2800 -675 -2249 -605
rect -2239 -445 -1688 -375
rect -2239 -605 -2129 -445
rect -1798 -605 -1688 -445
rect -2239 -675 -1688 -605
rect -1678 -445 -1127 -375
rect -1678 -605 -1568 -445
rect -1237 -605 -1127 -445
rect -1678 -675 -1127 -605
rect -1117 -445 -566 -375
rect -1117 -605 -1007 -445
rect -676 -605 -566 -445
rect -1117 -675 -566 -605
rect -556 -445 -5 -375
rect -556 -605 -446 -445
rect -115 -605 -5 -445
rect -556 -675 -5 -605
rect 5 -445 556 -375
rect 5 -605 115 -445
rect 446 -605 556 -445
rect 5 -675 556 -605
rect 566 -445 1117 -375
rect 566 -605 676 -445
rect 1007 -605 1117 -445
rect 566 -675 1117 -605
rect 1127 -445 1678 -375
rect 1127 -605 1237 -445
rect 1568 -605 1678 -445
rect 1127 -675 1678 -605
rect 1688 -445 2239 -375
rect 1688 -605 1798 -445
rect 2129 -605 2239 -445
rect 1688 -675 2239 -605
rect 2249 -445 2800 -375
rect 2249 -605 2359 -445
rect 2249 -675 2800 -605
rect -2800 -795 -2249 -725
rect -2359 -955 -2249 -795
rect -2800 -1025 -2249 -955
rect -2239 -795 -1688 -725
rect -2239 -955 -2129 -795
rect -1798 -955 -1688 -795
rect -2239 -1025 -1688 -955
rect -1678 -795 -1127 -725
rect -1678 -955 -1568 -795
rect -1237 -955 -1127 -795
rect -1678 -1025 -1127 -955
rect -1117 -795 -566 -725
rect -1117 -955 -1007 -795
rect -676 -955 -566 -795
rect -1117 -1025 -566 -955
rect -556 -795 -5 -725
rect -556 -955 -446 -795
rect -115 -955 -5 -795
rect -556 -1025 -5 -955
rect 5 -795 556 -725
rect 5 -955 115 -795
rect 446 -955 556 -795
rect 5 -1025 556 -955
rect 566 -795 1117 -725
rect 566 -955 676 -795
rect 1007 -955 1117 -795
rect 566 -1025 1117 -955
rect 1127 -795 1678 -725
rect 1127 -955 1237 -795
rect 1568 -955 1678 -795
rect 1127 -1025 1678 -955
rect 1688 -795 2239 -725
rect 1688 -955 1798 -795
rect 2129 -955 2239 -795
rect 1688 -1025 2239 -955
rect 2249 -795 2800 -725
rect 2249 -955 2359 -795
rect 2249 -1025 2800 -955
rect -2800 -1145 -2249 -1075
rect -2359 -1305 -2249 -1145
rect -2800 -1375 -2249 -1305
rect -2239 -1145 -1688 -1075
rect -2239 -1305 -2129 -1145
rect -1798 -1305 -1688 -1145
rect -2239 -1375 -1688 -1305
rect -1678 -1145 -1127 -1075
rect -1678 -1305 -1568 -1145
rect -1237 -1305 -1127 -1145
rect -1678 -1375 -1127 -1305
rect -1117 -1145 -566 -1075
rect -1117 -1305 -1007 -1145
rect -676 -1305 -566 -1145
rect -1117 -1375 -566 -1305
rect -556 -1145 -5 -1075
rect -556 -1305 -446 -1145
rect -115 -1305 -5 -1145
rect -556 -1375 -5 -1305
rect 5 -1145 556 -1075
rect 5 -1305 115 -1145
rect 446 -1305 556 -1145
rect 5 -1375 556 -1305
rect 566 -1145 1117 -1075
rect 566 -1305 676 -1145
rect 1007 -1305 1117 -1145
rect 566 -1375 1117 -1305
rect 1127 -1145 1678 -1075
rect 1127 -1305 1237 -1145
rect 1568 -1305 1678 -1145
rect 1127 -1375 1678 -1305
rect 1688 -1145 2239 -1075
rect 1688 -1305 1798 -1145
rect 2129 -1305 2239 -1145
rect 1688 -1375 2239 -1305
rect 2249 -1145 2800 -1075
rect 2249 -1305 2359 -1145
rect 2249 -1375 2800 -1305
rect -2800 -1495 -2249 -1425
rect -2359 -1725 -2249 -1495
rect -2239 -1495 -1688 -1425
rect -2239 -1725 -2129 -1495
rect -1798 -1725 -1688 -1495
rect -1678 -1495 -1127 -1425
rect -1678 -1725 -1568 -1495
rect -1237 -1725 -1127 -1495
rect -1117 -1495 -566 -1425
rect -1117 -1725 -1007 -1495
rect -676 -1725 -566 -1495
rect -556 -1495 -5 -1425
rect -556 -1725 -446 -1495
rect -115 -1725 -5 -1495
rect 5 -1495 556 -1425
rect 5 -1725 115 -1495
rect 446 -1725 556 -1495
rect 566 -1495 1117 -1425
rect 566 -1725 676 -1495
rect 1007 -1725 1117 -1495
rect 1127 -1495 1678 -1425
rect 1127 -1725 1237 -1495
rect 1568 -1725 1678 -1495
rect 1688 -1495 2239 -1425
rect 1688 -1725 1798 -1495
rect 2129 -1725 2239 -1495
rect 2249 -1495 2800 -1425
rect 2249 -1725 2359 -1495
<< metal4 >>
rect -2800 1425 -2249 1725
rect -2239 1425 -1688 1725
rect -1678 1425 -1127 1725
rect -1117 1425 -566 1725
rect -556 1425 -5 1725
rect 5 1425 556 1725
rect 566 1425 1117 1725
rect 1127 1425 1678 1725
rect 1688 1425 2239 1725
rect 2249 1425 2800 1725
rect -2800 1075 -2249 1375
rect -2239 1075 -1688 1375
rect -1678 1075 -1127 1375
rect -1117 1075 -566 1375
rect -556 1075 -5 1375
rect 5 1075 556 1375
rect 566 1075 1117 1375
rect 1127 1075 1678 1375
rect 1688 1075 2239 1375
rect 2249 1075 2800 1375
rect -2800 725 -2249 1025
rect -2239 725 -1688 1025
rect -1678 725 -1127 1025
rect -1117 725 -566 1025
rect -556 725 -5 1025
rect 5 725 556 1025
rect 566 725 1117 1025
rect 1127 725 1678 1025
rect 1688 725 2239 1025
rect 2249 725 2800 1025
rect -2800 375 -2249 675
rect -2239 375 -1688 675
rect -1678 375 -1127 675
rect -1117 375 -566 675
rect -556 375 -5 675
rect 5 375 556 675
rect 566 375 1117 675
rect 1127 375 1678 675
rect 1688 375 2239 675
rect 2249 375 2800 675
rect -2800 25 -2249 325
rect -2239 25 -1688 325
rect -1678 25 -1127 325
rect -1117 25 -566 325
rect -556 25 -5 325
rect 5 25 556 325
rect 566 25 1117 325
rect 1127 25 1678 325
rect 1688 25 2239 325
rect 2249 25 2800 325
rect -2800 -325 -2249 -25
rect -2239 -325 -1688 -25
rect -1678 -325 -1127 -25
rect -1117 -325 -566 -25
rect -556 -325 -5 -25
rect 5 -325 556 -25
rect 566 -325 1117 -25
rect 1127 -325 1678 -25
rect 1688 -325 2239 -25
rect 2249 -325 2800 -25
rect -2800 -675 -2249 -375
rect -2239 -675 -1688 -375
rect -1678 -675 -1127 -375
rect -1117 -675 -566 -375
rect -556 -675 -5 -375
rect 5 -675 556 -375
rect 566 -675 1117 -375
rect 1127 -675 1678 -375
rect 1688 -675 2239 -375
rect 2249 -675 2800 -375
rect -2800 -1025 -2249 -725
rect -2239 -1025 -1688 -725
rect -1678 -1025 -1127 -725
rect -1117 -1025 -566 -725
rect -556 -1025 -5 -725
rect 5 -1025 556 -725
rect 566 -1025 1117 -725
rect 1127 -1025 1678 -725
rect 1688 -1025 2239 -725
rect 2249 -1025 2800 -725
rect -2800 -1375 -2249 -1075
rect -2239 -1375 -1688 -1075
rect -1678 -1375 -1127 -1075
rect -1117 -1375 -566 -1075
rect -556 -1375 -5 -1075
rect 5 -1375 556 -1075
rect 566 -1375 1117 -1075
rect 1127 -1375 1678 -1075
rect 1688 -1375 2239 -1075
rect 2249 -1375 2800 -1075
rect -2800 -1725 -2249 -1425
rect -2239 -1725 -1688 -1425
rect -1678 -1725 -1127 -1425
rect -1117 -1725 -566 -1425
rect -556 -1725 -5 -1425
rect 5 -1725 556 -1425
rect 566 -1725 1117 -1425
rect 1127 -1725 1678 -1425
rect 1688 -1725 2239 -1425
rect 2249 -1725 2800 -1425
<< mimcap2 >>
rect -2750 1655 -2550 1675
rect -2750 1495 -2730 1655
rect -2570 1495 -2550 1655
rect -2750 1475 -2550 1495
rect -2189 1655 -1989 1675
rect -2189 1495 -2169 1655
rect -2009 1495 -1989 1655
rect -2189 1475 -1989 1495
rect -1628 1655 -1428 1675
rect -1628 1495 -1608 1655
rect -1448 1495 -1428 1655
rect -1628 1475 -1428 1495
rect -1067 1655 -867 1675
rect -1067 1495 -1047 1655
rect -887 1495 -867 1655
rect -1067 1475 -867 1495
rect -506 1655 -306 1675
rect -506 1495 -486 1655
rect -326 1495 -306 1655
rect -506 1475 -306 1495
rect 55 1655 255 1675
rect 55 1495 75 1655
rect 235 1495 255 1655
rect 55 1475 255 1495
rect 616 1655 816 1675
rect 616 1495 636 1655
rect 796 1495 816 1655
rect 616 1475 816 1495
rect 1177 1655 1377 1675
rect 1177 1495 1197 1655
rect 1357 1495 1377 1655
rect 1177 1475 1377 1495
rect 1738 1655 1938 1675
rect 1738 1495 1758 1655
rect 1918 1495 1938 1655
rect 1738 1475 1938 1495
rect 2299 1655 2499 1675
rect 2299 1495 2319 1655
rect 2479 1495 2499 1655
rect 2299 1475 2499 1495
rect -2750 1305 -2550 1325
rect -2750 1145 -2730 1305
rect -2570 1145 -2550 1305
rect -2750 1125 -2550 1145
rect -2189 1305 -1989 1325
rect -2189 1145 -2169 1305
rect -2009 1145 -1989 1305
rect -2189 1125 -1989 1145
rect -1628 1305 -1428 1325
rect -1628 1145 -1608 1305
rect -1448 1145 -1428 1305
rect -1628 1125 -1428 1145
rect -1067 1305 -867 1325
rect -1067 1145 -1047 1305
rect -887 1145 -867 1305
rect -1067 1125 -867 1145
rect -506 1305 -306 1325
rect -506 1145 -486 1305
rect -326 1145 -306 1305
rect -506 1125 -306 1145
rect 55 1305 255 1325
rect 55 1145 75 1305
rect 235 1145 255 1305
rect 55 1125 255 1145
rect 616 1305 816 1325
rect 616 1145 636 1305
rect 796 1145 816 1305
rect 616 1125 816 1145
rect 1177 1305 1377 1325
rect 1177 1145 1197 1305
rect 1357 1145 1377 1305
rect 1177 1125 1377 1145
rect 1738 1305 1938 1325
rect 1738 1145 1758 1305
rect 1918 1145 1938 1305
rect 1738 1125 1938 1145
rect 2299 1305 2499 1325
rect 2299 1145 2319 1305
rect 2479 1145 2499 1305
rect 2299 1125 2499 1145
rect -2750 955 -2550 975
rect -2750 795 -2730 955
rect -2570 795 -2550 955
rect -2750 775 -2550 795
rect -2189 955 -1989 975
rect -2189 795 -2169 955
rect -2009 795 -1989 955
rect -2189 775 -1989 795
rect -1628 955 -1428 975
rect -1628 795 -1608 955
rect -1448 795 -1428 955
rect -1628 775 -1428 795
rect -1067 955 -867 975
rect -1067 795 -1047 955
rect -887 795 -867 955
rect -1067 775 -867 795
rect -506 955 -306 975
rect -506 795 -486 955
rect -326 795 -306 955
rect -506 775 -306 795
rect 55 955 255 975
rect 55 795 75 955
rect 235 795 255 955
rect 55 775 255 795
rect 616 955 816 975
rect 616 795 636 955
rect 796 795 816 955
rect 616 775 816 795
rect 1177 955 1377 975
rect 1177 795 1197 955
rect 1357 795 1377 955
rect 1177 775 1377 795
rect 1738 955 1938 975
rect 1738 795 1758 955
rect 1918 795 1938 955
rect 1738 775 1938 795
rect 2299 955 2499 975
rect 2299 795 2319 955
rect 2479 795 2499 955
rect 2299 775 2499 795
rect -2750 605 -2550 625
rect -2750 445 -2730 605
rect -2570 445 -2550 605
rect -2750 425 -2550 445
rect -2189 605 -1989 625
rect -2189 445 -2169 605
rect -2009 445 -1989 605
rect -2189 425 -1989 445
rect -1628 605 -1428 625
rect -1628 445 -1608 605
rect -1448 445 -1428 605
rect -1628 425 -1428 445
rect -1067 605 -867 625
rect -1067 445 -1047 605
rect -887 445 -867 605
rect -1067 425 -867 445
rect -506 605 -306 625
rect -506 445 -486 605
rect -326 445 -306 605
rect -506 425 -306 445
rect 55 605 255 625
rect 55 445 75 605
rect 235 445 255 605
rect 55 425 255 445
rect 616 605 816 625
rect 616 445 636 605
rect 796 445 816 605
rect 616 425 816 445
rect 1177 605 1377 625
rect 1177 445 1197 605
rect 1357 445 1377 605
rect 1177 425 1377 445
rect 1738 605 1938 625
rect 1738 445 1758 605
rect 1918 445 1938 605
rect 1738 425 1938 445
rect 2299 605 2499 625
rect 2299 445 2319 605
rect 2479 445 2499 605
rect 2299 425 2499 445
rect -2750 255 -2550 275
rect -2750 95 -2730 255
rect -2570 95 -2550 255
rect -2750 75 -2550 95
rect -2189 255 -1989 275
rect -2189 95 -2169 255
rect -2009 95 -1989 255
rect -2189 75 -1989 95
rect -1628 255 -1428 275
rect -1628 95 -1608 255
rect -1448 95 -1428 255
rect -1628 75 -1428 95
rect -1067 255 -867 275
rect -1067 95 -1047 255
rect -887 95 -867 255
rect -1067 75 -867 95
rect -506 255 -306 275
rect -506 95 -486 255
rect -326 95 -306 255
rect -506 75 -306 95
rect 55 255 255 275
rect 55 95 75 255
rect 235 95 255 255
rect 55 75 255 95
rect 616 255 816 275
rect 616 95 636 255
rect 796 95 816 255
rect 616 75 816 95
rect 1177 255 1377 275
rect 1177 95 1197 255
rect 1357 95 1377 255
rect 1177 75 1377 95
rect 1738 255 1938 275
rect 1738 95 1758 255
rect 1918 95 1938 255
rect 1738 75 1938 95
rect 2299 255 2499 275
rect 2299 95 2319 255
rect 2479 95 2499 255
rect 2299 75 2499 95
rect -2750 -95 -2550 -75
rect -2750 -255 -2730 -95
rect -2570 -255 -2550 -95
rect -2750 -275 -2550 -255
rect -2189 -95 -1989 -75
rect -2189 -255 -2169 -95
rect -2009 -255 -1989 -95
rect -2189 -275 -1989 -255
rect -1628 -95 -1428 -75
rect -1628 -255 -1608 -95
rect -1448 -255 -1428 -95
rect -1628 -275 -1428 -255
rect -1067 -95 -867 -75
rect -1067 -255 -1047 -95
rect -887 -255 -867 -95
rect -1067 -275 -867 -255
rect -506 -95 -306 -75
rect -506 -255 -486 -95
rect -326 -255 -306 -95
rect -506 -275 -306 -255
rect 55 -95 255 -75
rect 55 -255 75 -95
rect 235 -255 255 -95
rect 55 -275 255 -255
rect 616 -95 816 -75
rect 616 -255 636 -95
rect 796 -255 816 -95
rect 616 -275 816 -255
rect 1177 -95 1377 -75
rect 1177 -255 1197 -95
rect 1357 -255 1377 -95
rect 1177 -275 1377 -255
rect 1738 -95 1938 -75
rect 1738 -255 1758 -95
rect 1918 -255 1938 -95
rect 1738 -275 1938 -255
rect 2299 -95 2499 -75
rect 2299 -255 2319 -95
rect 2479 -255 2499 -95
rect 2299 -275 2499 -255
rect -2750 -445 -2550 -425
rect -2750 -605 -2730 -445
rect -2570 -605 -2550 -445
rect -2750 -625 -2550 -605
rect -2189 -445 -1989 -425
rect -2189 -605 -2169 -445
rect -2009 -605 -1989 -445
rect -2189 -625 -1989 -605
rect -1628 -445 -1428 -425
rect -1628 -605 -1608 -445
rect -1448 -605 -1428 -445
rect -1628 -625 -1428 -605
rect -1067 -445 -867 -425
rect -1067 -605 -1047 -445
rect -887 -605 -867 -445
rect -1067 -625 -867 -605
rect -506 -445 -306 -425
rect -506 -605 -486 -445
rect -326 -605 -306 -445
rect -506 -625 -306 -605
rect 55 -445 255 -425
rect 55 -605 75 -445
rect 235 -605 255 -445
rect 55 -625 255 -605
rect 616 -445 816 -425
rect 616 -605 636 -445
rect 796 -605 816 -445
rect 616 -625 816 -605
rect 1177 -445 1377 -425
rect 1177 -605 1197 -445
rect 1357 -605 1377 -445
rect 1177 -625 1377 -605
rect 1738 -445 1938 -425
rect 1738 -605 1758 -445
rect 1918 -605 1938 -445
rect 1738 -625 1938 -605
rect 2299 -445 2499 -425
rect 2299 -605 2319 -445
rect 2479 -605 2499 -445
rect 2299 -625 2499 -605
rect -2750 -795 -2550 -775
rect -2750 -955 -2730 -795
rect -2570 -955 -2550 -795
rect -2750 -975 -2550 -955
rect -2189 -795 -1989 -775
rect -2189 -955 -2169 -795
rect -2009 -955 -1989 -795
rect -2189 -975 -1989 -955
rect -1628 -795 -1428 -775
rect -1628 -955 -1608 -795
rect -1448 -955 -1428 -795
rect -1628 -975 -1428 -955
rect -1067 -795 -867 -775
rect -1067 -955 -1047 -795
rect -887 -955 -867 -795
rect -1067 -975 -867 -955
rect -506 -795 -306 -775
rect -506 -955 -486 -795
rect -326 -955 -306 -795
rect -506 -975 -306 -955
rect 55 -795 255 -775
rect 55 -955 75 -795
rect 235 -955 255 -795
rect 55 -975 255 -955
rect 616 -795 816 -775
rect 616 -955 636 -795
rect 796 -955 816 -795
rect 616 -975 816 -955
rect 1177 -795 1377 -775
rect 1177 -955 1197 -795
rect 1357 -955 1377 -795
rect 1177 -975 1377 -955
rect 1738 -795 1938 -775
rect 1738 -955 1758 -795
rect 1918 -955 1938 -795
rect 1738 -975 1938 -955
rect 2299 -795 2499 -775
rect 2299 -955 2319 -795
rect 2479 -955 2499 -795
rect 2299 -975 2499 -955
rect -2750 -1145 -2550 -1125
rect -2750 -1305 -2730 -1145
rect -2570 -1305 -2550 -1145
rect -2750 -1325 -2550 -1305
rect -2189 -1145 -1989 -1125
rect -2189 -1305 -2169 -1145
rect -2009 -1305 -1989 -1145
rect -2189 -1325 -1989 -1305
rect -1628 -1145 -1428 -1125
rect -1628 -1305 -1608 -1145
rect -1448 -1305 -1428 -1145
rect -1628 -1325 -1428 -1305
rect -1067 -1145 -867 -1125
rect -1067 -1305 -1047 -1145
rect -887 -1305 -867 -1145
rect -1067 -1325 -867 -1305
rect -506 -1145 -306 -1125
rect -506 -1305 -486 -1145
rect -326 -1305 -306 -1145
rect -506 -1325 -306 -1305
rect 55 -1145 255 -1125
rect 55 -1305 75 -1145
rect 235 -1305 255 -1145
rect 55 -1325 255 -1305
rect 616 -1145 816 -1125
rect 616 -1305 636 -1145
rect 796 -1305 816 -1145
rect 616 -1325 816 -1305
rect 1177 -1145 1377 -1125
rect 1177 -1305 1197 -1145
rect 1357 -1305 1377 -1145
rect 1177 -1325 1377 -1305
rect 1738 -1145 1938 -1125
rect 1738 -1305 1758 -1145
rect 1918 -1305 1938 -1145
rect 1738 -1325 1938 -1305
rect 2299 -1145 2499 -1125
rect 2299 -1305 2319 -1145
rect 2479 -1305 2499 -1145
rect 2299 -1325 2499 -1305
rect -2750 -1495 -2550 -1475
rect -2750 -1655 -2730 -1495
rect -2570 -1655 -2550 -1495
rect -2750 -1675 -2550 -1655
rect -2189 -1495 -1989 -1475
rect -2189 -1655 -2169 -1495
rect -2009 -1655 -1989 -1495
rect -2189 -1675 -1989 -1655
rect -1628 -1495 -1428 -1475
rect -1628 -1655 -1608 -1495
rect -1448 -1655 -1428 -1495
rect -1628 -1675 -1428 -1655
rect -1067 -1495 -867 -1475
rect -1067 -1655 -1047 -1495
rect -887 -1655 -867 -1495
rect -1067 -1675 -867 -1655
rect -506 -1495 -306 -1475
rect -506 -1655 -486 -1495
rect -326 -1655 -306 -1495
rect -506 -1675 -306 -1655
rect 55 -1495 255 -1475
rect 55 -1655 75 -1495
rect 235 -1655 255 -1495
rect 55 -1675 255 -1655
rect 616 -1495 816 -1475
rect 616 -1655 636 -1495
rect 796 -1655 816 -1495
rect 616 -1675 816 -1655
rect 1177 -1495 1377 -1475
rect 1177 -1655 1197 -1495
rect 1357 -1655 1377 -1495
rect 1177 -1675 1377 -1655
rect 1738 -1495 1938 -1475
rect 1738 -1655 1758 -1495
rect 1918 -1655 1938 -1495
rect 1738 -1675 1938 -1655
rect 2299 -1495 2499 -1475
rect 2299 -1655 2319 -1495
rect 2479 -1655 2499 -1495
rect 2299 -1675 2499 -1655
<< mimcap2contact >>
rect -2730 1495 -2570 1655
rect -2169 1495 -2009 1655
rect -1608 1495 -1448 1655
rect -1047 1495 -887 1655
rect -486 1495 -326 1655
rect 75 1495 235 1655
rect 636 1495 796 1655
rect 1197 1495 1357 1655
rect 1758 1495 1918 1655
rect 2319 1495 2479 1655
rect -2730 1145 -2570 1305
rect -2169 1145 -2009 1305
rect -1608 1145 -1448 1305
rect -1047 1145 -887 1305
rect -486 1145 -326 1305
rect 75 1145 235 1305
rect 636 1145 796 1305
rect 1197 1145 1357 1305
rect 1758 1145 1918 1305
rect 2319 1145 2479 1305
rect -2730 795 -2570 955
rect -2169 795 -2009 955
rect -1608 795 -1448 955
rect -1047 795 -887 955
rect -486 795 -326 955
rect 75 795 235 955
rect 636 795 796 955
rect 1197 795 1357 955
rect 1758 795 1918 955
rect 2319 795 2479 955
rect -2730 445 -2570 605
rect -2169 445 -2009 605
rect -1608 445 -1448 605
rect -1047 445 -887 605
rect -486 445 -326 605
rect 75 445 235 605
rect 636 445 796 605
rect 1197 445 1357 605
rect 1758 445 1918 605
rect 2319 445 2479 605
rect -2730 95 -2570 255
rect -2169 95 -2009 255
rect -1608 95 -1448 255
rect -1047 95 -887 255
rect -486 95 -326 255
rect 75 95 235 255
rect 636 95 796 255
rect 1197 95 1357 255
rect 1758 95 1918 255
rect 2319 95 2479 255
rect -2730 -255 -2570 -95
rect -2169 -255 -2009 -95
rect -1608 -255 -1448 -95
rect -1047 -255 -887 -95
rect -486 -255 -326 -95
rect 75 -255 235 -95
rect 636 -255 796 -95
rect 1197 -255 1357 -95
rect 1758 -255 1918 -95
rect 2319 -255 2479 -95
rect -2730 -605 -2570 -445
rect -2169 -605 -2009 -445
rect -1608 -605 -1448 -445
rect -1047 -605 -887 -445
rect -486 -605 -326 -445
rect 75 -605 235 -445
rect 636 -605 796 -445
rect 1197 -605 1357 -445
rect 1758 -605 1918 -445
rect 2319 -605 2479 -445
rect -2730 -955 -2570 -795
rect -2169 -955 -2009 -795
rect -1608 -955 -1448 -795
rect -1047 -955 -887 -795
rect -486 -955 -326 -795
rect 75 -955 235 -795
rect 636 -955 796 -795
rect 1197 -955 1357 -795
rect 1758 -955 1918 -795
rect 2319 -955 2479 -795
rect -2730 -1305 -2570 -1145
rect -2169 -1305 -2009 -1145
rect -1608 -1305 -1448 -1145
rect -1047 -1305 -887 -1145
rect -486 -1305 -326 -1145
rect 75 -1305 235 -1145
rect 636 -1305 796 -1145
rect 1197 -1305 1357 -1145
rect 1758 -1305 1918 -1145
rect 2319 -1305 2479 -1145
rect -2730 -1655 -2570 -1495
rect -2169 -1655 -2009 -1495
rect -1608 -1655 -1448 -1495
rect -1047 -1655 -887 -1495
rect -486 -1655 -326 -1495
rect 75 -1655 235 -1495
rect 636 -1655 796 -1495
rect 1197 -1655 1357 -1495
rect 1758 -1655 1918 -1495
rect 2319 -1655 2479 -1495
<< metal5 >>
rect -2730 1667 -2410 1750
rect -2169 1667 -1849 1750
rect -1608 1667 -1288 1750
rect -1047 1667 -727 1750
rect -486 1667 -166 1750
rect 75 1667 395 1750
rect 636 1667 956 1750
rect 1197 1667 1517 1750
rect 1758 1667 2078 1750
rect 2319 1667 2639 1750
rect -2742 1655 -2410 1667
rect -2742 1495 -2730 1655
rect -2570 1495 -2410 1655
rect -2742 1483 -2410 1495
rect -2181 1655 -1849 1667
rect -2181 1495 -2169 1655
rect -2009 1495 -1849 1655
rect -2181 1483 -1849 1495
rect -1620 1655 -1288 1667
rect -1620 1495 -1608 1655
rect -1448 1495 -1288 1655
rect -1620 1483 -1288 1495
rect -1059 1655 -727 1667
rect -1059 1495 -1047 1655
rect -887 1495 -727 1655
rect -1059 1483 -727 1495
rect -498 1655 -166 1667
rect -498 1495 -486 1655
rect -326 1495 -166 1655
rect -498 1483 -166 1495
rect 63 1655 395 1667
rect 63 1495 75 1655
rect 235 1495 395 1655
rect 63 1483 395 1495
rect 624 1655 956 1667
rect 624 1495 636 1655
rect 796 1495 956 1655
rect 624 1483 956 1495
rect 1185 1655 1517 1667
rect 1185 1495 1197 1655
rect 1357 1495 1517 1655
rect 1185 1483 1517 1495
rect 1746 1655 2078 1667
rect 1746 1495 1758 1655
rect 1918 1495 2078 1655
rect 1746 1483 2078 1495
rect 2307 1655 2639 1667
rect 2307 1495 2319 1655
rect 2479 1495 2639 1655
rect 2307 1483 2639 1495
rect -2730 1317 -2410 1483
rect -2169 1317 -1849 1483
rect -1608 1317 -1288 1483
rect -1047 1317 -727 1483
rect -486 1317 -166 1483
rect 75 1317 395 1483
rect 636 1317 956 1483
rect 1197 1317 1517 1483
rect 1758 1317 2078 1483
rect 2319 1317 2639 1483
rect -2742 1305 -2410 1317
rect -2742 1145 -2730 1305
rect -2570 1145 -2410 1305
rect -2742 1133 -2410 1145
rect -2181 1305 -1849 1317
rect -2181 1145 -2169 1305
rect -2009 1145 -1849 1305
rect -2181 1133 -1849 1145
rect -1620 1305 -1288 1317
rect -1620 1145 -1608 1305
rect -1448 1145 -1288 1305
rect -1620 1133 -1288 1145
rect -1059 1305 -727 1317
rect -1059 1145 -1047 1305
rect -887 1145 -727 1305
rect -1059 1133 -727 1145
rect -498 1305 -166 1317
rect -498 1145 -486 1305
rect -326 1145 -166 1305
rect -498 1133 -166 1145
rect 63 1305 395 1317
rect 63 1145 75 1305
rect 235 1145 395 1305
rect 63 1133 395 1145
rect 624 1305 956 1317
rect 624 1145 636 1305
rect 796 1145 956 1305
rect 624 1133 956 1145
rect 1185 1305 1517 1317
rect 1185 1145 1197 1305
rect 1357 1145 1517 1305
rect 1185 1133 1517 1145
rect 1746 1305 2078 1317
rect 1746 1145 1758 1305
rect 1918 1145 2078 1305
rect 1746 1133 2078 1145
rect 2307 1305 2639 1317
rect 2307 1145 2319 1305
rect 2479 1145 2639 1305
rect 2307 1133 2639 1145
rect -2730 967 -2410 1133
rect -2169 967 -1849 1133
rect -1608 967 -1288 1133
rect -1047 967 -727 1133
rect -486 967 -166 1133
rect 75 967 395 1133
rect 636 967 956 1133
rect 1197 967 1517 1133
rect 1758 967 2078 1133
rect 2319 967 2639 1133
rect -2742 955 -2410 967
rect -2742 795 -2730 955
rect -2570 795 -2410 955
rect -2742 783 -2410 795
rect -2181 955 -1849 967
rect -2181 795 -2169 955
rect -2009 795 -1849 955
rect -2181 783 -1849 795
rect -1620 955 -1288 967
rect -1620 795 -1608 955
rect -1448 795 -1288 955
rect -1620 783 -1288 795
rect -1059 955 -727 967
rect -1059 795 -1047 955
rect -887 795 -727 955
rect -1059 783 -727 795
rect -498 955 -166 967
rect -498 795 -486 955
rect -326 795 -166 955
rect -498 783 -166 795
rect 63 955 395 967
rect 63 795 75 955
rect 235 795 395 955
rect 63 783 395 795
rect 624 955 956 967
rect 624 795 636 955
rect 796 795 956 955
rect 624 783 956 795
rect 1185 955 1517 967
rect 1185 795 1197 955
rect 1357 795 1517 955
rect 1185 783 1517 795
rect 1746 955 2078 967
rect 1746 795 1758 955
rect 1918 795 2078 955
rect 1746 783 2078 795
rect 2307 955 2639 967
rect 2307 795 2319 955
rect 2479 795 2639 955
rect 2307 783 2639 795
rect -2730 617 -2410 783
rect -2169 617 -1849 783
rect -1608 617 -1288 783
rect -1047 617 -727 783
rect -486 617 -166 783
rect 75 617 395 783
rect 636 617 956 783
rect 1197 617 1517 783
rect 1758 617 2078 783
rect 2319 617 2639 783
rect -2742 605 -2410 617
rect -2742 445 -2730 605
rect -2570 445 -2410 605
rect -2742 433 -2410 445
rect -2181 605 -1849 617
rect -2181 445 -2169 605
rect -2009 445 -1849 605
rect -2181 433 -1849 445
rect -1620 605 -1288 617
rect -1620 445 -1608 605
rect -1448 445 -1288 605
rect -1620 433 -1288 445
rect -1059 605 -727 617
rect -1059 445 -1047 605
rect -887 445 -727 605
rect -1059 433 -727 445
rect -498 605 -166 617
rect -498 445 -486 605
rect -326 445 -166 605
rect -498 433 -166 445
rect 63 605 395 617
rect 63 445 75 605
rect 235 445 395 605
rect 63 433 395 445
rect 624 605 956 617
rect 624 445 636 605
rect 796 445 956 605
rect 624 433 956 445
rect 1185 605 1517 617
rect 1185 445 1197 605
rect 1357 445 1517 605
rect 1185 433 1517 445
rect 1746 605 2078 617
rect 1746 445 1758 605
rect 1918 445 2078 605
rect 1746 433 2078 445
rect 2307 605 2639 617
rect 2307 445 2319 605
rect 2479 445 2639 605
rect 2307 433 2639 445
rect -2730 267 -2410 433
rect -2169 267 -1849 433
rect -1608 267 -1288 433
rect -1047 267 -727 433
rect -486 267 -166 433
rect 75 267 395 433
rect 636 267 956 433
rect 1197 267 1517 433
rect 1758 267 2078 433
rect 2319 267 2639 433
rect -2742 255 -2410 267
rect -2742 95 -2730 255
rect -2570 95 -2410 255
rect -2742 83 -2410 95
rect -2181 255 -1849 267
rect -2181 95 -2169 255
rect -2009 95 -1849 255
rect -2181 83 -1849 95
rect -1620 255 -1288 267
rect -1620 95 -1608 255
rect -1448 95 -1288 255
rect -1620 83 -1288 95
rect -1059 255 -727 267
rect -1059 95 -1047 255
rect -887 95 -727 255
rect -1059 83 -727 95
rect -498 255 -166 267
rect -498 95 -486 255
rect -326 95 -166 255
rect -498 83 -166 95
rect 63 255 395 267
rect 63 95 75 255
rect 235 95 395 255
rect 63 83 395 95
rect 624 255 956 267
rect 624 95 636 255
rect 796 95 956 255
rect 624 83 956 95
rect 1185 255 1517 267
rect 1185 95 1197 255
rect 1357 95 1517 255
rect 1185 83 1517 95
rect 1746 255 2078 267
rect 1746 95 1758 255
rect 1918 95 2078 255
rect 1746 83 2078 95
rect 2307 255 2639 267
rect 2307 95 2319 255
rect 2479 95 2639 255
rect 2307 83 2639 95
rect -2730 -83 -2410 83
rect -2169 -83 -1849 83
rect -1608 -83 -1288 83
rect -1047 -83 -727 83
rect -486 -83 -166 83
rect 75 -83 395 83
rect 636 -83 956 83
rect 1197 -83 1517 83
rect 1758 -83 2078 83
rect 2319 -83 2639 83
rect -2742 -95 -2410 -83
rect -2742 -255 -2730 -95
rect -2570 -255 -2410 -95
rect -2742 -267 -2410 -255
rect -2181 -95 -1849 -83
rect -2181 -255 -2169 -95
rect -2009 -255 -1849 -95
rect -2181 -267 -1849 -255
rect -1620 -95 -1288 -83
rect -1620 -255 -1608 -95
rect -1448 -255 -1288 -95
rect -1620 -267 -1288 -255
rect -1059 -95 -727 -83
rect -1059 -255 -1047 -95
rect -887 -255 -727 -95
rect -1059 -267 -727 -255
rect -498 -95 -166 -83
rect -498 -255 -486 -95
rect -326 -255 -166 -95
rect -498 -267 -166 -255
rect 63 -95 395 -83
rect 63 -255 75 -95
rect 235 -255 395 -95
rect 63 -267 395 -255
rect 624 -95 956 -83
rect 624 -255 636 -95
rect 796 -255 956 -95
rect 624 -267 956 -255
rect 1185 -95 1517 -83
rect 1185 -255 1197 -95
rect 1357 -255 1517 -95
rect 1185 -267 1517 -255
rect 1746 -95 2078 -83
rect 1746 -255 1758 -95
rect 1918 -255 2078 -95
rect 1746 -267 2078 -255
rect 2307 -95 2639 -83
rect 2307 -255 2319 -95
rect 2479 -255 2639 -95
rect 2307 -267 2639 -255
rect -2730 -433 -2410 -267
rect -2169 -433 -1849 -267
rect -1608 -433 -1288 -267
rect -1047 -433 -727 -267
rect -486 -433 -166 -267
rect 75 -433 395 -267
rect 636 -433 956 -267
rect 1197 -433 1517 -267
rect 1758 -433 2078 -267
rect 2319 -433 2639 -267
rect -2742 -445 -2410 -433
rect -2742 -605 -2730 -445
rect -2570 -605 -2410 -445
rect -2742 -617 -2410 -605
rect -2181 -445 -1849 -433
rect -2181 -605 -2169 -445
rect -2009 -605 -1849 -445
rect -2181 -617 -1849 -605
rect -1620 -445 -1288 -433
rect -1620 -605 -1608 -445
rect -1448 -605 -1288 -445
rect -1620 -617 -1288 -605
rect -1059 -445 -727 -433
rect -1059 -605 -1047 -445
rect -887 -605 -727 -445
rect -1059 -617 -727 -605
rect -498 -445 -166 -433
rect -498 -605 -486 -445
rect -326 -605 -166 -445
rect -498 -617 -166 -605
rect 63 -445 395 -433
rect 63 -605 75 -445
rect 235 -605 395 -445
rect 63 -617 395 -605
rect 624 -445 956 -433
rect 624 -605 636 -445
rect 796 -605 956 -445
rect 624 -617 956 -605
rect 1185 -445 1517 -433
rect 1185 -605 1197 -445
rect 1357 -605 1517 -445
rect 1185 -617 1517 -605
rect 1746 -445 2078 -433
rect 1746 -605 1758 -445
rect 1918 -605 2078 -445
rect 1746 -617 2078 -605
rect 2307 -445 2639 -433
rect 2307 -605 2319 -445
rect 2479 -605 2639 -445
rect 2307 -617 2639 -605
rect -2730 -783 -2410 -617
rect -2169 -783 -1849 -617
rect -1608 -783 -1288 -617
rect -1047 -783 -727 -617
rect -486 -783 -166 -617
rect 75 -783 395 -617
rect 636 -783 956 -617
rect 1197 -783 1517 -617
rect 1758 -783 2078 -617
rect 2319 -783 2639 -617
rect -2742 -795 -2410 -783
rect -2742 -955 -2730 -795
rect -2570 -955 -2410 -795
rect -2742 -967 -2410 -955
rect -2181 -795 -1849 -783
rect -2181 -955 -2169 -795
rect -2009 -955 -1849 -795
rect -2181 -967 -1849 -955
rect -1620 -795 -1288 -783
rect -1620 -955 -1608 -795
rect -1448 -955 -1288 -795
rect -1620 -967 -1288 -955
rect -1059 -795 -727 -783
rect -1059 -955 -1047 -795
rect -887 -955 -727 -795
rect -1059 -967 -727 -955
rect -498 -795 -166 -783
rect -498 -955 -486 -795
rect -326 -955 -166 -795
rect -498 -967 -166 -955
rect 63 -795 395 -783
rect 63 -955 75 -795
rect 235 -955 395 -795
rect 63 -967 395 -955
rect 624 -795 956 -783
rect 624 -955 636 -795
rect 796 -955 956 -795
rect 624 -967 956 -955
rect 1185 -795 1517 -783
rect 1185 -955 1197 -795
rect 1357 -955 1517 -795
rect 1185 -967 1517 -955
rect 1746 -795 2078 -783
rect 1746 -955 1758 -795
rect 1918 -955 2078 -795
rect 1746 -967 2078 -955
rect 2307 -795 2639 -783
rect 2307 -955 2319 -795
rect 2479 -955 2639 -795
rect 2307 -967 2639 -955
rect -2730 -1133 -2410 -967
rect -2169 -1133 -1849 -967
rect -1608 -1133 -1288 -967
rect -1047 -1133 -727 -967
rect -486 -1133 -166 -967
rect 75 -1133 395 -967
rect 636 -1133 956 -967
rect 1197 -1133 1517 -967
rect 1758 -1133 2078 -967
rect 2319 -1133 2639 -967
rect -2742 -1145 -2410 -1133
rect -2742 -1305 -2730 -1145
rect -2570 -1305 -2410 -1145
rect -2742 -1317 -2410 -1305
rect -2181 -1145 -1849 -1133
rect -2181 -1305 -2169 -1145
rect -2009 -1305 -1849 -1145
rect -2181 -1317 -1849 -1305
rect -1620 -1145 -1288 -1133
rect -1620 -1305 -1608 -1145
rect -1448 -1305 -1288 -1145
rect -1620 -1317 -1288 -1305
rect -1059 -1145 -727 -1133
rect -1059 -1305 -1047 -1145
rect -887 -1305 -727 -1145
rect -1059 -1317 -727 -1305
rect -498 -1145 -166 -1133
rect -498 -1305 -486 -1145
rect -326 -1305 -166 -1145
rect -498 -1317 -166 -1305
rect 63 -1145 395 -1133
rect 63 -1305 75 -1145
rect 235 -1305 395 -1145
rect 63 -1317 395 -1305
rect 624 -1145 956 -1133
rect 624 -1305 636 -1145
rect 796 -1305 956 -1145
rect 624 -1317 956 -1305
rect 1185 -1145 1517 -1133
rect 1185 -1305 1197 -1145
rect 1357 -1305 1517 -1145
rect 1185 -1317 1517 -1305
rect 1746 -1145 2078 -1133
rect 1746 -1305 1758 -1145
rect 1918 -1305 2078 -1145
rect 1746 -1317 2078 -1305
rect 2307 -1145 2639 -1133
rect 2307 -1305 2319 -1145
rect 2479 -1305 2639 -1145
rect 2307 -1317 2639 -1305
rect -2730 -1483 -2410 -1317
rect -2169 -1483 -1849 -1317
rect -1608 -1483 -1288 -1317
rect -1047 -1483 -727 -1317
rect -486 -1483 -166 -1317
rect 75 -1483 395 -1317
rect 636 -1483 956 -1317
rect 1197 -1483 1517 -1317
rect 1758 -1483 2078 -1317
rect 2319 -1483 2639 -1317
rect -2742 -1495 -2410 -1483
rect -2742 -1655 -2730 -1495
rect -2570 -1655 -2410 -1495
rect -2742 -1667 -2410 -1655
rect -2181 -1495 -1849 -1483
rect -2181 -1655 -2169 -1495
rect -2009 -1655 -1849 -1495
rect -2181 -1667 -1849 -1655
rect -1620 -1495 -1288 -1483
rect -1620 -1655 -1608 -1495
rect -1448 -1655 -1288 -1495
rect -1620 -1667 -1288 -1655
rect -1059 -1495 -727 -1483
rect -1059 -1655 -1047 -1495
rect -887 -1655 -727 -1495
rect -1059 -1667 -727 -1655
rect -498 -1495 -166 -1483
rect -498 -1655 -486 -1495
rect -326 -1655 -166 -1495
rect -498 -1667 -166 -1655
rect 63 -1495 395 -1483
rect 63 -1655 75 -1495
rect 235 -1655 395 -1495
rect 63 -1667 395 -1655
rect 624 -1495 956 -1483
rect 624 -1655 636 -1495
rect 796 -1655 956 -1495
rect 624 -1667 956 -1655
rect 1185 -1495 1517 -1483
rect 1185 -1655 1197 -1495
rect 1357 -1655 1517 -1495
rect 1185 -1667 1517 -1655
rect 1746 -1495 2078 -1483
rect 1746 -1655 1758 -1495
rect 1918 -1655 2078 -1495
rect 1746 -1667 2078 -1655
rect 2307 -1495 2639 -1483
rect 2307 -1655 2319 -1495
rect 2479 -1655 2639 -1495
rect 2307 -1667 2639 -1655
rect -2730 -1750 -2410 -1667
rect -2169 -1750 -1849 -1667
rect -1608 -1750 -1288 -1667
rect -1047 -1750 -727 -1667
rect -486 -1750 -166 -1667
rect 75 -1750 395 -1667
rect 636 -1750 956 -1667
rect 1197 -1750 1517 -1667
rect 1758 -1750 2078 -1667
rect 2319 -1750 2639 -1667
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX 2249 1425 2549 1725
string parameters w 2.00 l 2.00 val 5.36 carea 1.00 cperi 0.17 nx 10 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>
