magic
tech sky130A
magscale 1 2
timestamp 1620848404
<< nwell >>
rect -850 2420 -50 5162
rect 3398 2420 4198 5162
<< psubdiff >>
rect -750 1720 -550 1820
rect -750 120 -700 1720
rect -600 120 -550 1720
rect -750 20 -550 120
rect 3902 1720 4102 1820
rect 3902 120 3952 1720
rect 4052 120 4102 1720
rect 3902 20 4102 120
<< nsubdiff >>
rect -750 4962 -550 5062
rect -750 2620 -700 4962
rect -600 2620 -550 4962
rect -750 2520 -550 2620
rect 3898 4962 4098 5062
rect 3898 2620 3948 4962
rect 4048 2620 4098 4962
rect 3898 2520 4098 2620
<< psubdiffcont >>
rect -700 120 -600 1720
rect 3952 120 4052 1720
<< nsubdiffcont >>
rect -700 2620 -600 4962
rect 3948 2620 4048 4962
<< locali >>
rect -716 4962 -584 4978
rect -716 2620 -700 4962
rect -600 2620 -584 4962
rect -716 2608 -584 2620
rect 3932 4962 4064 4978
rect 3932 2620 3948 4962
rect 4048 2620 4064 4962
rect 3932 2608 4064 2620
rect -716 1720 -584 1736
rect -716 120 -700 1720
rect -600 120 -584 1720
rect -716 104 -584 120
rect 3936 1720 4068 1736
rect 3936 120 3952 1720
rect 4052 120 4068 1720
rect 3936 104 4068 120
<< viali >>
rect -700 2620 -600 4962
rect 3948 2620 4048 4962
<< metal1 >>
rect -716 5314 -584 5324
rect -716 5210 -690 5314
rect -638 5210 -584 5314
rect -716 4962 -584 5210
rect 432 5314 504 5324
rect 432 5210 442 5314
rect 494 5210 504 5314
rect 432 5200 504 5210
rect 1004 5314 1076 5324
rect 1004 5210 1014 5314
rect 1066 5210 1076 5314
rect 1004 5200 1076 5210
rect 1576 5314 1648 5324
rect 1576 5210 1586 5314
rect 1638 5210 1648 5314
rect 1576 5200 1648 5210
rect 2148 5314 2220 5324
rect 2148 5210 2158 5314
rect 2210 5210 2220 5314
rect 2148 5200 2220 5210
rect 2720 5314 2792 5324
rect 2720 5210 2730 5314
rect 2782 5210 2792 5314
rect 2720 5200 2792 5210
rect 3292 5314 3360 5324
rect 3292 5210 3302 5314
rect 3354 5210 3360 5314
rect 3292 5200 3360 5210
rect 3932 5314 4064 5324
rect 3932 5210 3958 5314
rect 4010 5210 4064 5314
rect -716 2620 -700 4962
rect -600 2620 -584 4962
rect -716 2608 -584 2620
rect 456 2536 490 5200
rect 1028 2536 1062 5200
rect -2 2478 32 2536
rect 1600 2532 1634 5200
rect 2172 2532 2206 5200
rect 2744 2532 2778 5200
rect 3316 2532 3350 5200
rect 3932 4962 4064 5210
rect 3932 2620 3948 4962
rect 4048 2620 4064 4962
rect 3932 2608 4064 2620
rect 134 2480 354 2490
rect 134 2478 140 2480
rect -2 2438 140 2478
rect -2 1896 32 2438
rect 134 2422 140 2438
rect 348 2478 354 2480
rect 348 2442 444 2478
rect 348 2422 354 2442
rect 134 2420 354 2422
rect 570 2392 604 2532
rect 706 2484 926 2490
rect 706 2426 712 2484
rect 920 2426 926 2484
rect 706 2420 926 2426
rect 1142 2474 1176 2532
rect 1278 2480 1498 2486
rect 1278 2474 1284 2480
rect 1142 2438 1284 2474
rect 556 2386 620 2392
rect 556 2132 562 2386
rect 614 2132 620 2386
rect 556 2126 620 2132
rect 432 2086 504 2096
rect 432 1982 442 2086
rect 494 1982 504 2086
rect 432 1972 504 1982
rect 458 120 492 1972
rect 570 1896 604 2126
rect 1004 2086 1076 2096
rect 1004 1982 1014 2086
rect 1066 1982 1076 2086
rect 1004 1972 1076 1982
rect 1030 120 1064 1972
rect 1142 1896 1176 2438
rect 1278 2422 1284 2438
rect 1492 2474 1498 2480
rect 1492 2438 1588 2474
rect 1492 2422 1498 2438
rect 1278 2416 1498 2422
rect 1714 2392 1748 2532
rect 1850 2480 2070 2486
rect 1850 2422 1856 2480
rect 2064 2422 2070 2480
rect 1850 2416 2070 2422
rect 2286 2474 2320 2532
rect 2422 2480 2642 2486
rect 2422 2474 2428 2480
rect 2286 2438 2428 2474
rect 1700 2386 1764 2392
rect 1700 2132 1706 2386
rect 1758 2132 1764 2386
rect 1700 2126 1764 2132
rect 1576 2086 1648 2096
rect 1576 1982 1586 2086
rect 1638 1982 1648 2086
rect 1576 1972 1648 1982
rect 1602 120 1636 1972
rect 1714 1896 1748 2126
rect 2148 2086 2220 2096
rect 2148 1982 2158 2086
rect 2210 1982 2220 2086
rect 2148 1972 2220 1982
rect 2174 120 2208 1972
rect 2286 1896 2320 2438
rect 2422 2422 2428 2438
rect 2636 2474 2642 2480
rect 2636 2438 2732 2474
rect 2636 2422 2642 2438
rect 2422 2416 2642 2422
rect 2858 2392 2892 2532
rect 2994 2480 3214 2486
rect 2994 2422 3000 2480
rect 3208 2422 3214 2480
rect 2994 2416 3214 2422
rect 2844 2386 2908 2392
rect 2844 2132 2850 2386
rect 2902 2132 2908 2386
rect 2844 2126 2908 2132
rect 2720 2086 2792 2096
rect 2720 1982 2730 2086
rect 2782 1982 2792 2086
rect 2720 1972 2792 1982
rect 2746 120 2780 1972
rect 2858 1896 2892 2126
rect 3292 2086 3364 2096
rect 3292 1982 3302 2086
rect 3354 1982 3364 2086
rect 3292 1972 3364 1982
rect 3318 120 3352 1972
rect 154 -30 338 70
rect 154 -84 174 -30
rect 318 -84 338 -30
rect 154 -104 338 -84
rect 726 -170 910 56
rect 1298 -30 1482 30
rect 1298 -84 1318 -30
rect 1462 -84 1482 -30
rect 1298 -104 1482 -84
rect 726 -224 746 -170
rect 890 -224 910 -170
rect 726 -244 910 -224
rect 1870 -170 2054 56
rect 2442 -30 2626 30
rect 2442 -84 2462 -30
rect 2606 -84 2626 -30
rect 2442 -104 2626 -84
rect 1870 -224 1890 -170
rect 2034 -224 2054 -170
rect 1870 -244 2054 -224
rect 3014 -170 3198 56
rect 3014 -224 3034 -170
rect 3178 -224 3198 -170
rect 3014 -244 3198 -224
<< via1 >>
rect -690 5210 -638 5314
rect 442 5210 494 5314
rect 1014 5210 1066 5314
rect 1586 5210 1638 5314
rect 2158 5210 2210 5314
rect 2730 5210 2782 5314
rect 3302 5210 3354 5314
rect 3958 5210 4010 5314
rect 140 2422 348 2480
rect 712 2426 920 2484
rect 562 2132 614 2386
rect 442 1982 494 2086
rect 1014 1982 1066 2086
rect 1284 2422 1492 2480
rect 1856 2422 2064 2480
rect 1706 2132 1758 2386
rect 1586 1982 1638 2086
rect 2158 1982 2210 2086
rect 2428 2422 2636 2480
rect 3000 2422 3208 2480
rect 2850 2132 2902 2386
rect 2730 1982 2782 2086
rect 3302 1982 3354 2086
rect 174 -84 318 -30
rect 1318 -84 1462 -30
rect 746 -224 890 -170
rect 2462 -84 2606 -30
rect 1890 -224 2034 -170
rect 3034 -224 3178 -170
<< metal2 >>
rect -716 5314 4064 5324
rect -716 5210 -690 5314
rect -638 5210 442 5314
rect 494 5210 1014 5314
rect 1066 5210 1586 5314
rect 1638 5210 2158 5314
rect 2210 5210 2730 5314
rect 2782 5210 3302 5314
rect 3354 5210 3958 5314
rect 4010 5210 4064 5314
rect -716 5200 4064 5210
rect 134 2486 1180 2490
rect 134 2484 3214 2486
rect 134 2480 712 2484
rect 134 2422 140 2480
rect 348 2426 712 2480
rect 920 2480 3214 2484
rect 920 2426 1284 2480
rect 348 2422 1284 2426
rect 1492 2422 1856 2480
rect 2064 2422 2428 2480
rect 2636 2422 3000 2480
rect 3208 2422 3214 2480
rect 134 2420 3214 2422
rect 556 2386 3480 2392
rect 556 2132 562 2386
rect 614 2132 1706 2386
rect 1758 2132 2850 2386
rect 2902 2132 3480 2386
rect 556 2126 3480 2132
rect 432 2096 842 2098
rect 432 2086 3364 2096
rect 432 1982 442 2086
rect 494 1982 1014 2086
rect 1066 1982 1586 2086
rect 1638 1982 2158 2086
rect 2210 1982 2730 2086
rect 2782 1982 3302 2086
rect 3354 1982 3364 2086
rect 432 1972 3364 1982
rect 154 -30 2626 -24
rect 154 -84 174 -30
rect 318 -84 1318 -30
rect 1462 -84 2462 -30
rect 2606 -84 2626 -30
rect 154 -104 2626 -84
rect 726 -170 3198 -164
rect 726 -224 746 -170
rect 890 -224 1890 -170
rect 2034 -224 3034 -170
rect 3178 -224 3198 -170
rect 726 -244 3198 -224
use sky130_fd_pr__nfet_01v8_lvt_75T4HJ  sky130_fd_pr__nfet_01v8_lvt_75T4HJ_0
timestamp 1620840674
transform 1 0 1676 0 1 977
box -1688 -957 1688 957
use sky130_fd_pr__pfet_01v8_lvt_K54UQX  sky130_fd_pr__pfet_01v8_lvt_K54UQX_0
timestamp 1620836830
transform 1 0 1674 0 1 3774
box -1724 -1354 1724 1388
<< labels >>
flabel metal1 -2 2286 32 2378 1 FreeSans 800 0 0 0 vg
flabel metal2 1750 5200 1766 5324 1 FreeSans 800 0 0 0 VDD!
port 0 n
flabel metal2 2404 1972 2420 2096 1 FreeSans 800 0 0 0 Vq
port 5 n
flabel metal2 2346 -244 2362 -164 1 FreeSans 800 0 0 0 Va
port 2 n
flabel metal2 1574 -104 1590 -24 1 FreeSans 800 0 0 0 Vb
port 3 n
flabel metal2 3080 2126 3174 2392 1 FreeSans 800 0 0 0 Vgate
port 1 n
flabel psubdiffcont -700 120 -600 1720 1 FreeSans 800 0 0 0 GND!
port 4 n
flabel psubdiff 3902 20 4102 120 1 FreeSans 800 0 0 0 GND!
<< end >>
