magic
tech sky130A
magscale 1 2
timestamp 1621192096
<< psubdiff >>
rect 430 670 1470 694
rect 430 594 454 670
rect 1446 594 1470 670
rect 430 570 1470 594
rect -498 516 -50 540
rect -498 -60 -474 516
rect -74 -60 -50 516
rect 1952 516 2400 540
rect -498 -84 -50 -60
rect 1952 -60 1976 516
rect 2376 -60 2400 516
rect 1952 -84 2400 -60
<< psubdiffcont >>
rect 454 594 1446 670
rect -474 -60 -74 516
rect 1976 -60 2376 516
<< poly >>
rect 1438 404 1762 438
<< locali >>
rect 438 670 1462 686
rect 438 594 454 670
rect 1446 594 1462 670
rect 438 554 1462 594
rect -490 516 -58 532
rect -490 -60 -474 516
rect -74 -60 -58 516
rect 438 502 466 554
rect 518 502 1382 554
rect 1434 502 1462 554
rect 438 490 1462 502
rect 1960 516 2392 532
rect 464 404 522 438
rect 922 404 980 438
rect 1380 404 1438 438
rect -490 -76 -58 -60
rect 1960 -60 1976 516
rect 2376 -60 2392 516
rect 1960 -76 2392 -60
<< viali >>
rect 466 502 518 554
rect 1382 502 1434 554
<< metal1 >>
rect 454 554 530 566
rect 454 502 466 554
rect 518 502 530 554
rect 454 490 530 502
rect 1370 554 1446 566
rect 1370 502 1382 554
rect 1434 502 1446 554
rect 1370 490 1446 502
rect 148 438 380 450
rect 12 404 380 438
rect 12 366 56 404
rect 148 386 380 404
rect 12 -164 58 366
rect 470 -22 516 490
rect 2 -170 66 -164
rect 2 -222 8 -170
rect 60 -222 66 -170
rect 2 -228 66 -222
rect 928 -370 974 366
rect 1386 -22 1432 490
rect 1512 438 1744 450
rect 1512 404 1890 438
rect 1512 386 1744 404
rect 1844 -158 1890 404
rect 1836 -164 1900 -158
rect 1836 -216 1842 -164
rect 1894 -216 1900 -164
rect 1836 -222 1900 -216
rect 920 -376 984 -370
rect 920 -428 926 -376
rect 978 -428 984 -376
rect 920 -434 984 -428
<< via1 >>
rect 8 -222 60 -170
rect 1842 -216 1894 -164
rect 926 -428 978 -376
<< metal2 >>
rect 2 -164 1900 -158
rect 2 -170 1842 -164
rect 2 -222 8 -170
rect 60 -216 1842 -170
rect 1894 -216 1900 -164
rect 60 -222 1900 -216
rect 2 -228 1900 -222
rect 60 -376 1842 -368
rect 60 -428 926 -376
rect 978 -428 1842 -376
rect 60 -438 1842 -428
use sky130_fd_pr__nfet_01v8_lvt_NHDRDL  sky130_fd_pr__nfet_01v8_lvt_NHDRDL_0
timestamp 1620928018
transform 1 0 951 0 1 197
box -945 -257 945 257
<< labels >>
flabel metal2 60 -438 1842 -368 1 FreeSans 800 0 0 0 Vq
port 2 n
flabel metal2 60 -228 1842 -158 1 FreeSans 800 0 0 0 Vx
port 1 n
flabel locali 920 532 1002 560 1 FreeSans 800 0 0 0 GND!
port 3 n
<< end >>
