magic
tech sky130A
magscale 1 2
timestamp 1622081478
<< metal4 >>
rect -3179 2998 3179 3100
rect -3179 2762 2923 2998
rect 3159 2762 3179 2998
rect -3179 2678 3179 2762
rect -3179 2442 2923 2678
rect 3159 2442 3179 2678
rect -3179 2358 3179 2442
rect -3179 2122 2923 2358
rect 3159 2122 3179 2358
rect -3179 2038 3179 2122
rect -3179 1802 2923 2038
rect 3159 1802 3179 2038
rect -3179 1718 3179 1802
rect -3179 1482 2923 1718
rect 3159 1482 3179 1718
rect -3179 1398 3179 1482
rect -3179 1162 2923 1398
rect 3159 1162 3179 1398
rect -3179 1078 3179 1162
rect -3179 842 2923 1078
rect 3159 842 3179 1078
rect -3179 758 3179 842
rect -3179 522 2923 758
rect 3159 522 3179 758
rect -3179 438 3179 522
rect -3179 202 2923 438
rect 3159 202 3179 438
rect -3179 118 3179 202
rect -3179 -118 2923 118
rect 3159 -118 3179 118
rect -3179 -202 3179 -118
rect -3179 -438 2923 -202
rect 3159 -438 3179 -202
rect -3179 -522 3179 -438
rect -3179 -758 2923 -522
rect 3159 -758 3179 -522
rect -3179 -842 3179 -758
rect -3179 -1078 2923 -842
rect 3159 -1078 3179 -842
rect -3179 -1162 3179 -1078
rect -3179 -1398 2923 -1162
rect 3159 -1398 3179 -1162
rect -3179 -1482 3179 -1398
rect -3179 -1718 2923 -1482
rect 3159 -1718 3179 -1482
rect -3179 -1802 3179 -1718
rect -3179 -2038 2923 -1802
rect 3159 -2038 3179 -1802
rect -3179 -2122 3179 -2038
rect -3179 -2358 2923 -2122
rect 3159 -2358 3179 -2122
rect -3179 -2442 3179 -2358
rect -3179 -2678 2923 -2442
rect 3159 -2678 3179 -2442
rect -3179 -2762 3179 -2678
rect -3179 -2998 2923 -2762
rect 3159 -2998 3179 -2762
rect -3179 -3100 3179 -2998
<< via4 >>
rect 2923 2762 3159 2998
rect 2923 2442 3159 2678
rect 2923 2122 3159 2358
rect 2923 1802 3159 2038
rect 2923 1482 3159 1718
rect 2923 1162 3159 1398
rect 2923 842 3159 1078
rect 2923 522 3159 758
rect 2923 202 3159 438
rect 2923 -118 3159 118
rect 2923 -438 3159 -202
rect 2923 -758 3159 -522
rect 2923 -1078 3159 -842
rect 2923 -1398 3159 -1162
rect 2923 -1718 3159 -1482
rect 2923 -2038 3159 -1802
rect 2923 -2358 3159 -2122
rect 2923 -2678 3159 -2442
rect 2923 -2998 3159 -2762
<< mimcap2 >>
rect -3079 2838 2921 3000
rect -3079 -2838 -2893 2838
rect 2143 -2838 2921 2838
rect -3079 -3000 2921 -2838
<< mimcap2contact >>
rect -2893 -2838 2143 2838
<< metal5 >>
rect 2881 2998 3201 3101
rect -3063 2838 2313 2984
rect -3063 -2838 -2893 2838
rect 2143 -2838 2313 2838
rect -3063 -2984 2313 -2838
rect 2881 2762 2923 2998
rect 3159 2762 3201 2998
rect 2881 2678 3201 2762
rect 2881 2442 2923 2678
rect 3159 2442 3201 2678
rect 2881 2358 3201 2442
rect 2881 2122 2923 2358
rect 3159 2122 3201 2358
rect 2881 2038 3201 2122
rect 2881 1802 2923 2038
rect 3159 1802 3201 2038
rect 2881 1718 3201 1802
rect 2881 1482 2923 1718
rect 3159 1482 3201 1718
rect 2881 1398 3201 1482
rect 2881 1162 2923 1398
rect 3159 1162 3201 1398
rect 2881 1078 3201 1162
rect 2881 842 2923 1078
rect 3159 842 3201 1078
rect 2881 758 3201 842
rect 2881 522 2923 758
rect 3159 522 3201 758
rect 2881 438 3201 522
rect 2881 202 2923 438
rect 3159 202 3201 438
rect 2881 118 3201 202
rect 2881 -118 2923 118
rect 3159 -118 3201 118
rect 2881 -202 3201 -118
rect 2881 -438 2923 -202
rect 3159 -438 3201 -202
rect 2881 -522 3201 -438
rect 2881 -758 2923 -522
rect 3159 -758 3201 -522
rect 2881 -842 3201 -758
rect 2881 -1078 2923 -842
rect 3159 -1078 3201 -842
rect 2881 -1162 3201 -1078
rect 2881 -1398 2923 -1162
rect 3159 -1398 3201 -1162
rect 2881 -1482 3201 -1398
rect 2881 -1718 2923 -1482
rect 3159 -1718 3201 -1482
rect 2881 -1802 3201 -1718
rect 2881 -2038 2923 -1802
rect 3159 -2038 3201 -1802
rect 2881 -2122 3201 -2038
rect 2881 -2358 2923 -2122
rect 3159 -2358 3201 -2122
rect 2881 -2442 3201 -2358
rect 2881 -2678 2923 -2442
rect 3159 -2678 3201 -2442
rect 2881 -2762 3201 -2678
rect 2881 -2998 2923 -2762
rect 3159 -2998 3201 -2762
rect 2881 -3101 3201 -2998
<< properties >>
string FIXED_BBOX -3179 -3100 3021 3100
<< end >>
