magic
tech sky130A
magscale 1 2
timestamp 1620324069
<< nwell >>
rect -2813 -4400 2813 4400
<< pmoslvt >>
rect -2719 -4300 -2319 4300
rect -2261 -4300 -1861 4300
rect -1803 -4300 -1403 4300
rect -1345 -4300 -945 4300
rect -887 -4300 -487 4300
rect -429 -4300 -29 4300
rect 29 -4300 429 4300
rect 487 -4300 887 4300
rect 945 -4300 1345 4300
rect 1403 -4300 1803 4300
rect 1861 -4300 2261 4300
rect 2319 -4300 2719 4300
<< pdiff >>
rect -2777 4288 -2719 4300
rect -2777 -4288 -2765 4288
rect -2731 -4288 -2719 4288
rect -2777 -4300 -2719 -4288
rect -2319 4288 -2261 4300
rect -2319 -4288 -2307 4288
rect -2273 -4288 -2261 4288
rect -2319 -4300 -2261 -4288
rect -1861 4288 -1803 4300
rect -1861 -4288 -1849 4288
rect -1815 -4288 -1803 4288
rect -1861 -4300 -1803 -4288
rect -1403 4288 -1345 4300
rect -1403 -4288 -1391 4288
rect -1357 -4288 -1345 4288
rect -1403 -4300 -1345 -4288
rect -945 4288 -887 4300
rect -945 -4288 -933 4288
rect -899 -4288 -887 4288
rect -945 -4300 -887 -4288
rect -487 4288 -429 4300
rect -487 -4288 -475 4288
rect -441 -4288 -429 4288
rect -487 -4300 -429 -4288
rect -29 4288 29 4300
rect -29 -4288 -17 4288
rect 17 -4288 29 4288
rect -29 -4300 29 -4288
rect 429 4288 487 4300
rect 429 -4288 441 4288
rect 475 -4288 487 4288
rect 429 -4300 487 -4288
rect 887 4288 945 4300
rect 887 -4288 899 4288
rect 933 -4288 945 4288
rect 887 -4300 945 -4288
rect 1345 4288 1403 4300
rect 1345 -4288 1357 4288
rect 1391 -4288 1403 4288
rect 1345 -4300 1403 -4288
rect 1803 4288 1861 4300
rect 1803 -4288 1815 4288
rect 1849 -4288 1861 4288
rect 1803 -4300 1861 -4288
rect 2261 4288 2319 4300
rect 2261 -4288 2273 4288
rect 2307 -4288 2319 4288
rect 2261 -4300 2319 -4288
rect 2719 4288 2777 4300
rect 2719 -4288 2731 4288
rect 2765 -4288 2777 4288
rect 2719 -4300 2777 -4288
<< pdiffc >>
rect -2765 -4288 -2731 4288
rect -2307 -4288 -2273 4288
rect -1849 -4288 -1815 4288
rect -1391 -4288 -1357 4288
rect -933 -4288 -899 4288
rect -475 -4288 -441 4288
rect -17 -4288 17 4288
rect 441 -4288 475 4288
rect 899 -4288 933 4288
rect 1357 -4288 1391 4288
rect 1815 -4288 1849 4288
rect 2273 -4288 2307 4288
rect 2731 -4288 2765 4288
<< poly >>
rect -2719 4381 -2319 4397
rect -2719 4347 -2703 4381
rect -2335 4347 -2319 4381
rect -2719 4300 -2319 4347
rect -2261 4381 -1861 4397
rect -2261 4347 -2245 4381
rect -1877 4347 -1861 4381
rect -2261 4300 -1861 4347
rect -1803 4381 -1403 4397
rect -1803 4347 -1787 4381
rect -1419 4347 -1403 4381
rect -1803 4300 -1403 4347
rect -1345 4381 -945 4397
rect -1345 4347 -1329 4381
rect -961 4347 -945 4381
rect -1345 4300 -945 4347
rect -887 4381 -487 4397
rect -887 4347 -871 4381
rect -503 4347 -487 4381
rect -887 4300 -487 4347
rect -429 4381 -29 4397
rect -429 4347 -413 4381
rect -45 4347 -29 4381
rect -429 4300 -29 4347
rect 29 4381 429 4397
rect 29 4347 45 4381
rect 413 4347 429 4381
rect 29 4300 429 4347
rect 487 4381 887 4397
rect 487 4347 503 4381
rect 871 4347 887 4381
rect 487 4300 887 4347
rect 945 4381 1345 4397
rect 945 4347 961 4381
rect 1329 4347 1345 4381
rect 945 4300 1345 4347
rect 1403 4381 1803 4397
rect 1403 4347 1419 4381
rect 1787 4347 1803 4381
rect 1403 4300 1803 4347
rect 1861 4381 2261 4397
rect 1861 4347 1877 4381
rect 2245 4347 2261 4381
rect 1861 4300 2261 4347
rect 2319 4381 2719 4397
rect 2319 4347 2335 4381
rect 2703 4347 2719 4381
rect 2319 4300 2719 4347
rect -2719 -4347 -2319 -4300
rect -2719 -4381 -2703 -4347
rect -2335 -4381 -2319 -4347
rect -2719 -4397 -2319 -4381
rect -2261 -4347 -1861 -4300
rect -2261 -4381 -2245 -4347
rect -1877 -4381 -1861 -4347
rect -2261 -4397 -1861 -4381
rect -1803 -4347 -1403 -4300
rect -1803 -4381 -1787 -4347
rect -1419 -4381 -1403 -4347
rect -1803 -4397 -1403 -4381
rect -1345 -4347 -945 -4300
rect -1345 -4381 -1329 -4347
rect -961 -4381 -945 -4347
rect -1345 -4397 -945 -4381
rect -887 -4347 -487 -4300
rect -887 -4381 -871 -4347
rect -503 -4381 -487 -4347
rect -887 -4397 -487 -4381
rect -429 -4347 -29 -4300
rect -429 -4381 -413 -4347
rect -45 -4381 -29 -4347
rect -429 -4397 -29 -4381
rect 29 -4347 429 -4300
rect 29 -4381 45 -4347
rect 413 -4381 429 -4347
rect 29 -4397 429 -4381
rect 487 -4347 887 -4300
rect 487 -4381 503 -4347
rect 871 -4381 887 -4347
rect 487 -4397 887 -4381
rect 945 -4347 1345 -4300
rect 945 -4381 961 -4347
rect 1329 -4381 1345 -4347
rect 945 -4397 1345 -4381
rect 1403 -4347 1803 -4300
rect 1403 -4381 1419 -4347
rect 1787 -4381 1803 -4347
rect 1403 -4397 1803 -4381
rect 1861 -4347 2261 -4300
rect 1861 -4381 1877 -4347
rect 2245 -4381 2261 -4347
rect 1861 -4397 2261 -4381
rect 2319 -4347 2719 -4300
rect 2319 -4381 2335 -4347
rect 2703 -4381 2719 -4347
rect 2319 -4397 2719 -4381
<< polycont >>
rect -2703 4347 -2335 4381
rect -2245 4347 -1877 4381
rect -1787 4347 -1419 4381
rect -1329 4347 -961 4381
rect -871 4347 -503 4381
rect -413 4347 -45 4381
rect 45 4347 413 4381
rect 503 4347 871 4381
rect 961 4347 1329 4381
rect 1419 4347 1787 4381
rect 1877 4347 2245 4381
rect 2335 4347 2703 4381
rect -2703 -4381 -2335 -4347
rect -2245 -4381 -1877 -4347
rect -1787 -4381 -1419 -4347
rect -1329 -4381 -961 -4347
rect -871 -4381 -503 -4347
rect -413 -4381 -45 -4347
rect 45 -4381 413 -4347
rect 503 -4381 871 -4347
rect 961 -4381 1329 -4347
rect 1419 -4381 1787 -4347
rect 1877 -4381 2245 -4347
rect 2335 -4381 2703 -4347
<< locali >>
rect -2719 4347 -2703 4381
rect -2335 4347 -2319 4381
rect -2261 4347 -2245 4381
rect -1877 4347 -1861 4381
rect -1803 4347 -1787 4381
rect -1419 4347 -1403 4381
rect -1345 4347 -1329 4381
rect -961 4347 -945 4381
rect -887 4347 -871 4381
rect -503 4347 -487 4381
rect -429 4347 -413 4381
rect -45 4347 -29 4381
rect 29 4347 45 4381
rect 413 4347 429 4381
rect 487 4347 503 4381
rect 871 4347 887 4381
rect 945 4347 961 4381
rect 1329 4347 1345 4381
rect 1403 4347 1419 4381
rect 1787 4347 1803 4381
rect 1861 4347 1877 4381
rect 2245 4347 2261 4381
rect 2319 4347 2335 4381
rect 2703 4347 2719 4381
rect -2765 4288 -2731 4304
rect -2765 -4304 -2731 -4288
rect -2307 4288 -2273 4304
rect -2307 -4304 -2273 -4288
rect -1849 4288 -1815 4304
rect -1849 -4304 -1815 -4288
rect -1391 4288 -1357 4304
rect -1391 -4304 -1357 -4288
rect -933 4288 -899 4304
rect -933 -4304 -899 -4288
rect -475 4288 -441 4304
rect -475 -4304 -441 -4288
rect -17 4288 17 4304
rect -17 -4304 17 -4288
rect 441 4288 475 4304
rect 441 -4304 475 -4288
rect 899 4288 933 4304
rect 899 -4304 933 -4288
rect 1357 4288 1391 4304
rect 1357 -4304 1391 -4288
rect 1815 4288 1849 4304
rect 1815 -4304 1849 -4288
rect 2273 4288 2307 4304
rect 2273 -4304 2307 -4288
rect 2731 4288 2765 4304
rect 2731 -4304 2765 -4288
rect -2719 -4381 -2703 -4347
rect -2335 -4381 -2319 -4347
rect -2261 -4381 -2245 -4347
rect -1877 -4381 -1861 -4347
rect -1803 -4381 -1787 -4347
rect -1419 -4381 -1403 -4347
rect -1345 -4381 -1329 -4347
rect -961 -4381 -945 -4347
rect -887 -4381 -871 -4347
rect -503 -4381 -487 -4347
rect -429 -4381 -413 -4347
rect -45 -4381 -29 -4347
rect 29 -4381 45 -4347
rect 413 -4381 429 -4347
rect 487 -4381 503 -4347
rect 871 -4381 887 -4347
rect 945 -4381 961 -4347
rect 1329 -4381 1345 -4347
rect 1403 -4381 1419 -4347
rect 1787 -4381 1803 -4347
rect 1861 -4381 1877 -4347
rect 2245 -4381 2261 -4347
rect 2319 -4381 2335 -4347
rect 2703 -4381 2719 -4347
<< viali >>
rect -2703 4347 -2335 4381
rect -2245 4347 -1877 4381
rect -1787 4347 -1419 4381
rect -1329 4347 -961 4381
rect -871 4347 -503 4381
rect -413 4347 -45 4381
rect 45 4347 413 4381
rect 503 4347 871 4381
rect 961 4347 1329 4381
rect 1419 4347 1787 4381
rect 1877 4347 2245 4381
rect 2335 4347 2703 4381
rect -2765 -4288 -2731 4288
rect -2307 -4288 -2273 4288
rect -1849 -4288 -1815 4288
rect -1391 -4288 -1357 4288
rect -933 -4288 -899 4288
rect -475 -4288 -441 4288
rect -17 -4288 17 4288
rect 441 -4288 475 4288
rect 899 -4288 933 4288
rect 1357 -4288 1391 4288
rect 1815 -4288 1849 4288
rect 2273 -4288 2307 4288
rect 2731 -4288 2765 4288
rect -2703 -4381 -2335 -4347
rect -2245 -4381 -1877 -4347
rect -1787 -4381 -1419 -4347
rect -1329 -4381 -961 -4347
rect -871 -4381 -503 -4347
rect -413 -4381 -45 -4347
rect 45 -4381 413 -4347
rect 503 -4381 871 -4347
rect 961 -4381 1329 -4347
rect 1419 -4381 1787 -4347
rect 1877 -4381 2245 -4347
rect 2335 -4381 2703 -4347
<< metal1 >>
rect -2715 4381 -2323 4387
rect -2715 4347 -2703 4381
rect -2335 4347 -2323 4381
rect -2715 4341 -2323 4347
rect -2257 4381 -1865 4387
rect -2257 4347 -2245 4381
rect -1877 4347 -1865 4381
rect -2257 4341 -1865 4347
rect -1799 4381 -1407 4387
rect -1799 4347 -1787 4381
rect -1419 4347 -1407 4381
rect -1799 4341 -1407 4347
rect -1341 4381 -949 4387
rect -1341 4347 -1329 4381
rect -961 4347 -949 4381
rect -1341 4341 -949 4347
rect -883 4381 -491 4387
rect -883 4347 -871 4381
rect -503 4347 -491 4381
rect -883 4341 -491 4347
rect -425 4381 -33 4387
rect -425 4347 -413 4381
rect -45 4347 -33 4381
rect -425 4341 -33 4347
rect 33 4381 425 4387
rect 33 4347 45 4381
rect 413 4347 425 4381
rect 33 4341 425 4347
rect 491 4381 883 4387
rect 491 4347 503 4381
rect 871 4347 883 4381
rect 491 4341 883 4347
rect 949 4381 1341 4387
rect 949 4347 961 4381
rect 1329 4347 1341 4381
rect 949 4341 1341 4347
rect 1407 4381 1799 4387
rect 1407 4347 1419 4381
rect 1787 4347 1799 4381
rect 1407 4341 1799 4347
rect 1865 4381 2257 4387
rect 1865 4347 1877 4381
rect 2245 4347 2257 4381
rect 1865 4341 2257 4347
rect 2323 4381 2715 4387
rect 2323 4347 2335 4381
rect 2703 4347 2715 4381
rect 2323 4341 2715 4347
rect -2771 4288 -2725 4300
rect -2771 -4288 -2765 4288
rect -2731 -4288 -2725 4288
rect -2771 -4300 -2725 -4288
rect -2313 4288 -2267 4300
rect -2313 -4288 -2307 4288
rect -2273 -4288 -2267 4288
rect -2313 -4300 -2267 -4288
rect -1855 4288 -1809 4300
rect -1855 -4288 -1849 4288
rect -1815 -4288 -1809 4288
rect -1855 -4300 -1809 -4288
rect -1397 4288 -1351 4300
rect -1397 -4288 -1391 4288
rect -1357 -4288 -1351 4288
rect -1397 -4300 -1351 -4288
rect -939 4288 -893 4300
rect -939 -4288 -933 4288
rect -899 -4288 -893 4288
rect -939 -4300 -893 -4288
rect -481 4288 -435 4300
rect -481 -4288 -475 4288
rect -441 -4288 -435 4288
rect -481 -4300 -435 -4288
rect -23 4288 23 4300
rect -23 -4288 -17 4288
rect 17 -4288 23 4288
rect -23 -4300 23 -4288
rect 435 4288 481 4300
rect 435 -4288 441 4288
rect 475 -4288 481 4288
rect 435 -4300 481 -4288
rect 893 4288 939 4300
rect 893 -4288 899 4288
rect 933 -4288 939 4288
rect 893 -4300 939 -4288
rect 1351 4288 1397 4300
rect 1351 -4288 1357 4288
rect 1391 -4288 1397 4288
rect 1351 -4300 1397 -4288
rect 1809 4288 1855 4300
rect 1809 -4288 1815 4288
rect 1849 -4288 1855 4288
rect 1809 -4300 1855 -4288
rect 2267 4288 2313 4300
rect 2267 -4288 2273 4288
rect 2307 -4288 2313 4288
rect 2267 -4300 2313 -4288
rect 2725 4288 2771 4300
rect 2725 -4288 2731 4288
rect 2765 -4288 2771 4288
rect 2725 -4300 2771 -4288
rect -2715 -4347 -2323 -4341
rect -2715 -4381 -2703 -4347
rect -2335 -4381 -2323 -4347
rect -2715 -4387 -2323 -4381
rect -2257 -4347 -1865 -4341
rect -2257 -4381 -2245 -4347
rect -1877 -4381 -1865 -4347
rect -2257 -4387 -1865 -4381
rect -1799 -4347 -1407 -4341
rect -1799 -4381 -1787 -4347
rect -1419 -4381 -1407 -4347
rect -1799 -4387 -1407 -4381
rect -1341 -4347 -949 -4341
rect -1341 -4381 -1329 -4347
rect -961 -4381 -949 -4347
rect -1341 -4387 -949 -4381
rect -883 -4347 -491 -4341
rect -883 -4381 -871 -4347
rect -503 -4381 -491 -4347
rect -883 -4387 -491 -4381
rect -425 -4347 -33 -4341
rect -425 -4381 -413 -4347
rect -45 -4381 -33 -4347
rect -425 -4387 -33 -4381
rect 33 -4347 425 -4341
rect 33 -4381 45 -4347
rect 413 -4381 425 -4347
rect 33 -4387 425 -4381
rect 491 -4347 883 -4341
rect 491 -4381 503 -4347
rect 871 -4381 883 -4347
rect 491 -4387 883 -4381
rect 949 -4347 1341 -4341
rect 949 -4381 961 -4347
rect 1329 -4381 1341 -4347
rect 949 -4387 1341 -4381
rect 1407 -4347 1799 -4341
rect 1407 -4381 1419 -4347
rect 1787 -4381 1799 -4347
rect 1407 -4387 1799 -4381
rect 1865 -4347 2257 -4341
rect 1865 -4381 1877 -4347
rect 2245 -4381 2257 -4347
rect 1865 -4387 2257 -4381
rect 2323 -4347 2715 -4341
rect 2323 -4381 2335 -4347
rect 2703 -4381 2715 -4347
rect 2323 -4387 2715 -4381
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 43 l 2 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
