magic
tech sky130A
magscale 1 2
timestamp 1621285914
<< nwell >>
rect -9600 9500 7778 9502
rect -19400 1000 -9872 4342
rect -9600 1602 8666 9500
rect -9600 1600 -3680 1602
rect -2890 1600 1820 1602
rect 2610 1600 8666 1602
<< pwell >>
rect 12444 12133 18884 12234
rect 12444 11047 12545 12133
rect 13631 11047 13833 12133
rect 14919 11047 15121 12133
rect 16207 11047 16409 12133
rect 17495 11047 17697 12133
rect 18783 11047 18884 12133
rect 12444 10845 18884 11047
rect 12444 9759 12545 10845
rect 13631 9759 13833 10845
rect 14919 9759 15121 10845
rect 16207 9759 16409 10845
rect 17495 9759 17697 10845
rect 18783 9759 18884 10845
rect 12444 9557 18884 9759
rect 12444 8471 12545 9557
rect 13631 8471 13833 9557
rect 14919 8471 15121 9557
rect 16207 8471 16409 9557
rect 17495 8471 17697 9557
rect 18783 8471 18884 9557
rect 12444 8269 18884 8471
rect 12444 7183 12545 8269
rect 13631 7183 13833 8269
rect 14919 7183 15121 8269
rect 16207 7183 16409 8269
rect 17495 7183 17697 8269
rect 18783 7183 18884 8269
rect 12444 6981 18884 7183
rect 12444 5895 12545 6981
rect 13631 5895 13833 6981
rect 14919 5895 15121 6981
rect 16207 5895 16409 6981
rect 17495 5895 17697 6981
rect 18783 5895 18884 6981
rect 12444 5693 18884 5895
rect 12444 4607 12545 5693
rect 13631 4607 13833 5693
rect 14919 4607 15121 5693
rect 16207 4607 16409 5693
rect 17495 4607 17697 5693
rect 18783 4607 18884 5693
rect 12444 4405 18884 4607
rect 12444 3319 12545 4405
rect 13631 3319 13833 4405
rect 14919 3319 15121 4405
rect 16207 3319 16409 4405
rect 17495 3319 17697 4405
rect 18783 3319 18884 4405
rect 12444 3117 18884 3319
rect 12444 2031 12545 3117
rect 13631 2031 13833 3117
rect 14919 2031 15121 3117
rect 16207 2031 16409 3117
rect 17495 2031 17697 3117
rect 18783 2031 18884 3117
rect 12444 1930 18884 2031
<< nbase >>
rect 12571 11073 13605 12107
rect 13859 11073 14893 12107
rect 15147 11073 16181 12107
rect 16435 11073 17469 12107
rect 17723 11073 18757 12107
rect 12571 9785 13605 10819
rect 13859 9785 14893 10819
rect 15147 9785 16181 10819
rect 16435 9785 17469 10819
rect 17723 9785 18757 10819
rect 12571 8497 13605 9531
rect 13859 8497 14893 9531
rect 15147 8497 16181 9531
rect 16435 8497 17469 9531
rect 17723 8497 18757 9531
rect 12571 7209 13605 8243
rect 13859 7209 14893 8243
rect 15147 7209 16181 8243
rect 16435 7209 17469 8243
rect 17723 7209 18757 8243
rect 12571 5921 13605 6955
rect 13859 5921 14893 6955
rect 15147 5921 16181 6955
rect 16435 5921 17469 6955
rect 17723 5921 18757 6955
rect 12571 4633 13605 5667
rect 13859 4633 14893 5667
rect 15147 4633 16181 5667
rect 16435 4633 17469 5667
rect 17723 4633 18757 5667
rect 12571 3345 13605 4379
rect 13859 3345 14893 4379
rect 15147 3345 16181 4379
rect 16435 3345 17469 4379
rect 17723 3345 18757 4379
rect 12571 2057 13605 3091
rect 13859 2057 14893 3091
rect 15147 2057 16181 3091
rect 16435 2057 17469 3091
rect 17723 2057 18757 3091
<< pmoslvt >>
rect -18562 1662 -18162 4242
rect -17990 1662 -17590 4242
rect -17418 1662 -17018 4242
rect -16846 1662 -16446 4242
rect -16274 1662 -15874 4242
rect -15702 1662 -15302 4242
rect -15130 1662 -14730 4242
rect -14558 1662 -14158 4242
rect -13986 1662 -13586 4242
rect -13414 1662 -13014 4242
rect -12842 1662 -12442 4242
rect -12270 1662 -11870 4242
rect -11698 1662 -11298 4242
rect -11126 1662 -10726 4242
rect -8754 1700 -8354 9440
rect -8296 1700 -7896 9440
rect -7838 1700 -7438 9440
rect -7380 1700 -6980 9440
rect -6922 1700 -6522 9440
rect -6464 1700 -6064 9440
rect -6006 1700 -5606 9440
rect -5548 1700 -5148 9440
rect -5090 1700 -4690 9440
rect -4632 1700 -4232 9440
rect -4174 1700 -3774 9440
rect -2796 1700 -2396 9440
rect -2338 1700 -1938 9440
rect -1880 1700 -1480 9440
rect -1422 1700 -1022 9440
rect -964 1700 -564 9440
rect -506 1700 -106 9440
rect -48 1700 352 9440
rect 410 1700 810 9440
rect 868 1700 1268 9440
rect 1326 1700 1726 9440
rect 2704 1700 3104 9440
rect 3162 1700 3562 9440
rect 3620 1700 4020 9440
rect 4078 1700 4478 9440
rect 4536 1700 4936 9440
rect 4994 1700 5394 9440
rect 5452 1700 5852 9440
rect 5910 1700 6310 9440
rect 6368 1700 6768 9440
rect 6826 1700 7226 9440
rect 7284 1700 7684 9440
<< nmoslvt >>
rect -17176 8406 -11776 8806
rect -21766 5132 -21366 5532
rect -21308 5132 -20908 5532
rect -20850 5132 -20450 5532
rect -20392 5132 -19992 5532
rect -19934 5132 -19534 5532
rect -19476 5132 -19076 5532
rect -16836 4854 -16436 6654
rect -16264 4854 -15864 6654
rect -15692 4854 -15292 6654
rect -15120 4854 -14720 6654
rect -14548 4854 -14148 6654
rect -13976 4854 -13576 6654
rect -13404 4854 -13004 6654
rect -12832 4854 -12432 6654
<< ndiff >>
rect -17176 8852 -11776 8864
rect -17176 8818 -17164 8852
rect -11788 8818 -11776 8852
rect -17176 8806 -11776 8818
rect -17176 8394 -11776 8406
rect -17176 8360 -17164 8394
rect -11788 8360 -11776 8394
rect -17176 8348 -11776 8360
rect -21824 5520 -21766 5532
rect -21824 5144 -21812 5520
rect -21778 5144 -21766 5520
rect -21824 5132 -21766 5144
rect -21366 5520 -21308 5532
rect -21366 5144 -21354 5520
rect -21320 5144 -21308 5520
rect -21366 5132 -21308 5144
rect -20908 5520 -20850 5532
rect -20908 5144 -20896 5520
rect -20862 5144 -20850 5520
rect -20908 5132 -20850 5144
rect -20450 5520 -20392 5532
rect -20450 5144 -20438 5520
rect -20404 5144 -20392 5520
rect -20450 5132 -20392 5144
rect -19992 5520 -19934 5532
rect -19992 5144 -19980 5520
rect -19946 5144 -19934 5520
rect -19992 5132 -19934 5144
rect -19534 5520 -19476 5532
rect -19534 5144 -19522 5520
rect -19488 5144 -19476 5520
rect -19534 5132 -19476 5144
rect -19076 5520 -19018 5532
rect -19076 5144 -19064 5520
rect -19030 5144 -19018 5520
rect -19076 5132 -19018 5144
rect -16894 6642 -16836 6654
rect -16894 4866 -16882 6642
rect -16848 4866 -16836 6642
rect -16894 4854 -16836 4866
rect -16436 6642 -16378 6654
rect -16436 4866 -16424 6642
rect -16390 4866 -16378 6642
rect -16436 4854 -16378 4866
rect -16322 6642 -16264 6654
rect -16322 4866 -16310 6642
rect -16276 4866 -16264 6642
rect -16322 4854 -16264 4866
rect -15864 6642 -15806 6654
rect -15864 4866 -15852 6642
rect -15818 4866 -15806 6642
rect -15864 4854 -15806 4866
rect -15750 6642 -15692 6654
rect -15750 4866 -15738 6642
rect -15704 4866 -15692 6642
rect -15750 4854 -15692 4866
rect -15292 6642 -15234 6654
rect -15292 4866 -15280 6642
rect -15246 4866 -15234 6642
rect -15292 4854 -15234 4866
rect -15178 6642 -15120 6654
rect -15178 4866 -15166 6642
rect -15132 4866 -15120 6642
rect -15178 4854 -15120 4866
rect -14720 6642 -14662 6654
rect -14720 4866 -14708 6642
rect -14674 4866 -14662 6642
rect -14720 4854 -14662 4866
rect -14606 6642 -14548 6654
rect -14606 4866 -14594 6642
rect -14560 4866 -14548 6642
rect -14606 4854 -14548 4866
rect -14148 6642 -14090 6654
rect -14148 4866 -14136 6642
rect -14102 4866 -14090 6642
rect -14148 4854 -14090 4866
rect -14034 6642 -13976 6654
rect -14034 4866 -14022 6642
rect -13988 4866 -13976 6642
rect -14034 4854 -13976 4866
rect -13576 6642 -13518 6654
rect -13576 4866 -13564 6642
rect -13530 4866 -13518 6642
rect -13576 4854 -13518 4866
rect -13462 6642 -13404 6654
rect -13462 4866 -13450 6642
rect -13416 4866 -13404 6642
rect -13462 4854 -13404 4866
rect -13004 6642 -12946 6654
rect -13004 4866 -12992 6642
rect -12958 4866 -12946 6642
rect -13004 4854 -12946 4866
rect -12890 6642 -12832 6654
rect -12890 4866 -12878 6642
rect -12844 4866 -12832 6642
rect -12890 4854 -12832 4866
rect -12432 6642 -12374 6654
rect -12432 4866 -12420 6642
rect -12386 4866 -12374 6642
rect -12432 4854 -12374 4866
<< pdiff >>
rect 12748 11876 13428 11930
rect 12748 11842 12800 11876
rect 12834 11842 12890 11876
rect 12924 11842 12980 11876
rect 13014 11842 13070 11876
rect 13104 11842 13160 11876
rect 13194 11842 13250 11876
rect 13284 11842 13340 11876
rect 13374 11842 13428 11876
rect 12748 11786 13428 11842
rect 12748 11752 12800 11786
rect 12834 11752 12890 11786
rect 12924 11752 12980 11786
rect 13014 11752 13070 11786
rect 13104 11752 13160 11786
rect 13194 11752 13250 11786
rect 13284 11752 13340 11786
rect 13374 11752 13428 11786
rect 12748 11696 13428 11752
rect 12748 11662 12800 11696
rect 12834 11662 12890 11696
rect 12924 11662 12980 11696
rect 13014 11662 13070 11696
rect 13104 11662 13160 11696
rect 13194 11662 13250 11696
rect 13284 11662 13340 11696
rect 13374 11662 13428 11696
rect 12748 11606 13428 11662
rect 12748 11572 12800 11606
rect 12834 11572 12890 11606
rect 12924 11572 12980 11606
rect 13014 11572 13070 11606
rect 13104 11572 13160 11606
rect 13194 11572 13250 11606
rect 13284 11572 13340 11606
rect 13374 11572 13428 11606
rect 12748 11516 13428 11572
rect 12748 11482 12800 11516
rect 12834 11482 12890 11516
rect 12924 11482 12980 11516
rect 13014 11482 13070 11516
rect 13104 11482 13160 11516
rect 13194 11482 13250 11516
rect 13284 11482 13340 11516
rect 13374 11482 13428 11516
rect 12748 11426 13428 11482
rect 12748 11392 12800 11426
rect 12834 11392 12890 11426
rect 12924 11392 12980 11426
rect 13014 11392 13070 11426
rect 13104 11392 13160 11426
rect 13194 11392 13250 11426
rect 13284 11392 13340 11426
rect 13374 11392 13428 11426
rect 12748 11336 13428 11392
rect 12748 11302 12800 11336
rect 12834 11302 12890 11336
rect 12924 11302 12980 11336
rect 13014 11302 13070 11336
rect 13104 11302 13160 11336
rect 13194 11302 13250 11336
rect 13284 11302 13340 11336
rect 13374 11302 13428 11336
rect 12748 11250 13428 11302
rect 14036 11876 14716 11930
rect 14036 11842 14088 11876
rect 14122 11842 14178 11876
rect 14212 11842 14268 11876
rect 14302 11842 14358 11876
rect 14392 11842 14448 11876
rect 14482 11842 14538 11876
rect 14572 11842 14628 11876
rect 14662 11842 14716 11876
rect 14036 11786 14716 11842
rect 14036 11752 14088 11786
rect 14122 11752 14178 11786
rect 14212 11752 14268 11786
rect 14302 11752 14358 11786
rect 14392 11752 14448 11786
rect 14482 11752 14538 11786
rect 14572 11752 14628 11786
rect 14662 11752 14716 11786
rect 14036 11696 14716 11752
rect 14036 11662 14088 11696
rect 14122 11662 14178 11696
rect 14212 11662 14268 11696
rect 14302 11662 14358 11696
rect 14392 11662 14448 11696
rect 14482 11662 14538 11696
rect 14572 11662 14628 11696
rect 14662 11662 14716 11696
rect 14036 11606 14716 11662
rect 14036 11572 14088 11606
rect 14122 11572 14178 11606
rect 14212 11572 14268 11606
rect 14302 11572 14358 11606
rect 14392 11572 14448 11606
rect 14482 11572 14538 11606
rect 14572 11572 14628 11606
rect 14662 11572 14716 11606
rect 14036 11516 14716 11572
rect 14036 11482 14088 11516
rect 14122 11482 14178 11516
rect 14212 11482 14268 11516
rect 14302 11482 14358 11516
rect 14392 11482 14448 11516
rect 14482 11482 14538 11516
rect 14572 11482 14628 11516
rect 14662 11482 14716 11516
rect 14036 11426 14716 11482
rect 14036 11392 14088 11426
rect 14122 11392 14178 11426
rect 14212 11392 14268 11426
rect 14302 11392 14358 11426
rect 14392 11392 14448 11426
rect 14482 11392 14538 11426
rect 14572 11392 14628 11426
rect 14662 11392 14716 11426
rect 14036 11336 14716 11392
rect 14036 11302 14088 11336
rect 14122 11302 14178 11336
rect 14212 11302 14268 11336
rect 14302 11302 14358 11336
rect 14392 11302 14448 11336
rect 14482 11302 14538 11336
rect 14572 11302 14628 11336
rect 14662 11302 14716 11336
rect 14036 11250 14716 11302
rect 15324 11876 16004 11930
rect 15324 11842 15376 11876
rect 15410 11842 15466 11876
rect 15500 11842 15556 11876
rect 15590 11842 15646 11876
rect 15680 11842 15736 11876
rect 15770 11842 15826 11876
rect 15860 11842 15916 11876
rect 15950 11842 16004 11876
rect 15324 11786 16004 11842
rect 15324 11752 15376 11786
rect 15410 11752 15466 11786
rect 15500 11752 15556 11786
rect 15590 11752 15646 11786
rect 15680 11752 15736 11786
rect 15770 11752 15826 11786
rect 15860 11752 15916 11786
rect 15950 11752 16004 11786
rect 15324 11696 16004 11752
rect 15324 11662 15376 11696
rect 15410 11662 15466 11696
rect 15500 11662 15556 11696
rect 15590 11662 15646 11696
rect 15680 11662 15736 11696
rect 15770 11662 15826 11696
rect 15860 11662 15916 11696
rect 15950 11662 16004 11696
rect 15324 11606 16004 11662
rect 15324 11572 15376 11606
rect 15410 11572 15466 11606
rect 15500 11572 15556 11606
rect 15590 11572 15646 11606
rect 15680 11572 15736 11606
rect 15770 11572 15826 11606
rect 15860 11572 15916 11606
rect 15950 11572 16004 11606
rect 15324 11516 16004 11572
rect 15324 11482 15376 11516
rect 15410 11482 15466 11516
rect 15500 11482 15556 11516
rect 15590 11482 15646 11516
rect 15680 11482 15736 11516
rect 15770 11482 15826 11516
rect 15860 11482 15916 11516
rect 15950 11482 16004 11516
rect 15324 11426 16004 11482
rect 15324 11392 15376 11426
rect 15410 11392 15466 11426
rect 15500 11392 15556 11426
rect 15590 11392 15646 11426
rect 15680 11392 15736 11426
rect 15770 11392 15826 11426
rect 15860 11392 15916 11426
rect 15950 11392 16004 11426
rect 15324 11336 16004 11392
rect 15324 11302 15376 11336
rect 15410 11302 15466 11336
rect 15500 11302 15556 11336
rect 15590 11302 15646 11336
rect 15680 11302 15736 11336
rect 15770 11302 15826 11336
rect 15860 11302 15916 11336
rect 15950 11302 16004 11336
rect 15324 11250 16004 11302
rect 16612 11876 17292 11930
rect 16612 11842 16664 11876
rect 16698 11842 16754 11876
rect 16788 11842 16844 11876
rect 16878 11842 16934 11876
rect 16968 11842 17024 11876
rect 17058 11842 17114 11876
rect 17148 11842 17204 11876
rect 17238 11842 17292 11876
rect 16612 11786 17292 11842
rect 16612 11752 16664 11786
rect 16698 11752 16754 11786
rect 16788 11752 16844 11786
rect 16878 11752 16934 11786
rect 16968 11752 17024 11786
rect 17058 11752 17114 11786
rect 17148 11752 17204 11786
rect 17238 11752 17292 11786
rect 16612 11696 17292 11752
rect 16612 11662 16664 11696
rect 16698 11662 16754 11696
rect 16788 11662 16844 11696
rect 16878 11662 16934 11696
rect 16968 11662 17024 11696
rect 17058 11662 17114 11696
rect 17148 11662 17204 11696
rect 17238 11662 17292 11696
rect 16612 11606 17292 11662
rect 16612 11572 16664 11606
rect 16698 11572 16754 11606
rect 16788 11572 16844 11606
rect 16878 11572 16934 11606
rect 16968 11572 17024 11606
rect 17058 11572 17114 11606
rect 17148 11572 17204 11606
rect 17238 11572 17292 11606
rect 16612 11516 17292 11572
rect 16612 11482 16664 11516
rect 16698 11482 16754 11516
rect 16788 11482 16844 11516
rect 16878 11482 16934 11516
rect 16968 11482 17024 11516
rect 17058 11482 17114 11516
rect 17148 11482 17204 11516
rect 17238 11482 17292 11516
rect 16612 11426 17292 11482
rect 16612 11392 16664 11426
rect 16698 11392 16754 11426
rect 16788 11392 16844 11426
rect 16878 11392 16934 11426
rect 16968 11392 17024 11426
rect 17058 11392 17114 11426
rect 17148 11392 17204 11426
rect 17238 11392 17292 11426
rect 16612 11336 17292 11392
rect 16612 11302 16664 11336
rect 16698 11302 16754 11336
rect 16788 11302 16844 11336
rect 16878 11302 16934 11336
rect 16968 11302 17024 11336
rect 17058 11302 17114 11336
rect 17148 11302 17204 11336
rect 17238 11302 17292 11336
rect 16612 11250 17292 11302
rect 17900 11876 18580 11930
rect 17900 11842 17952 11876
rect 17986 11842 18042 11876
rect 18076 11842 18132 11876
rect 18166 11842 18222 11876
rect 18256 11842 18312 11876
rect 18346 11842 18402 11876
rect 18436 11842 18492 11876
rect 18526 11842 18580 11876
rect 17900 11786 18580 11842
rect 17900 11752 17952 11786
rect 17986 11752 18042 11786
rect 18076 11752 18132 11786
rect 18166 11752 18222 11786
rect 18256 11752 18312 11786
rect 18346 11752 18402 11786
rect 18436 11752 18492 11786
rect 18526 11752 18580 11786
rect 17900 11696 18580 11752
rect 17900 11662 17952 11696
rect 17986 11662 18042 11696
rect 18076 11662 18132 11696
rect 18166 11662 18222 11696
rect 18256 11662 18312 11696
rect 18346 11662 18402 11696
rect 18436 11662 18492 11696
rect 18526 11662 18580 11696
rect 17900 11606 18580 11662
rect 17900 11572 17952 11606
rect 17986 11572 18042 11606
rect 18076 11572 18132 11606
rect 18166 11572 18222 11606
rect 18256 11572 18312 11606
rect 18346 11572 18402 11606
rect 18436 11572 18492 11606
rect 18526 11572 18580 11606
rect 17900 11516 18580 11572
rect 17900 11482 17952 11516
rect 17986 11482 18042 11516
rect 18076 11482 18132 11516
rect 18166 11482 18222 11516
rect 18256 11482 18312 11516
rect 18346 11482 18402 11516
rect 18436 11482 18492 11516
rect 18526 11482 18580 11516
rect 17900 11426 18580 11482
rect 17900 11392 17952 11426
rect 17986 11392 18042 11426
rect 18076 11392 18132 11426
rect 18166 11392 18222 11426
rect 18256 11392 18312 11426
rect 18346 11392 18402 11426
rect 18436 11392 18492 11426
rect 18526 11392 18580 11426
rect 17900 11336 18580 11392
rect 17900 11302 17952 11336
rect 17986 11302 18042 11336
rect 18076 11302 18132 11336
rect 18166 11302 18222 11336
rect 18256 11302 18312 11336
rect 18346 11302 18402 11336
rect 18436 11302 18492 11336
rect 18526 11302 18580 11336
rect 17900 11250 18580 11302
rect 12748 10588 13428 10642
rect 12748 10554 12800 10588
rect 12834 10554 12890 10588
rect 12924 10554 12980 10588
rect 13014 10554 13070 10588
rect 13104 10554 13160 10588
rect 13194 10554 13250 10588
rect 13284 10554 13340 10588
rect 13374 10554 13428 10588
rect 12748 10498 13428 10554
rect 12748 10464 12800 10498
rect 12834 10464 12890 10498
rect 12924 10464 12980 10498
rect 13014 10464 13070 10498
rect 13104 10464 13160 10498
rect 13194 10464 13250 10498
rect 13284 10464 13340 10498
rect 13374 10464 13428 10498
rect 12748 10408 13428 10464
rect 12748 10374 12800 10408
rect 12834 10374 12890 10408
rect 12924 10374 12980 10408
rect 13014 10374 13070 10408
rect 13104 10374 13160 10408
rect 13194 10374 13250 10408
rect 13284 10374 13340 10408
rect 13374 10374 13428 10408
rect 12748 10318 13428 10374
rect 12748 10284 12800 10318
rect 12834 10284 12890 10318
rect 12924 10284 12980 10318
rect 13014 10284 13070 10318
rect 13104 10284 13160 10318
rect 13194 10284 13250 10318
rect 13284 10284 13340 10318
rect 13374 10284 13428 10318
rect 12748 10228 13428 10284
rect 12748 10194 12800 10228
rect 12834 10194 12890 10228
rect 12924 10194 12980 10228
rect 13014 10194 13070 10228
rect 13104 10194 13160 10228
rect 13194 10194 13250 10228
rect 13284 10194 13340 10228
rect 13374 10194 13428 10228
rect 12748 10138 13428 10194
rect 12748 10104 12800 10138
rect 12834 10104 12890 10138
rect 12924 10104 12980 10138
rect 13014 10104 13070 10138
rect 13104 10104 13160 10138
rect 13194 10104 13250 10138
rect 13284 10104 13340 10138
rect 13374 10104 13428 10138
rect 12748 10048 13428 10104
rect 12748 10014 12800 10048
rect 12834 10014 12890 10048
rect 12924 10014 12980 10048
rect 13014 10014 13070 10048
rect 13104 10014 13160 10048
rect 13194 10014 13250 10048
rect 13284 10014 13340 10048
rect 13374 10014 13428 10048
rect 12748 9962 13428 10014
rect 14036 10588 14716 10642
rect 14036 10554 14088 10588
rect 14122 10554 14178 10588
rect 14212 10554 14268 10588
rect 14302 10554 14358 10588
rect 14392 10554 14448 10588
rect 14482 10554 14538 10588
rect 14572 10554 14628 10588
rect 14662 10554 14716 10588
rect 14036 10498 14716 10554
rect 14036 10464 14088 10498
rect 14122 10464 14178 10498
rect 14212 10464 14268 10498
rect 14302 10464 14358 10498
rect 14392 10464 14448 10498
rect 14482 10464 14538 10498
rect 14572 10464 14628 10498
rect 14662 10464 14716 10498
rect 14036 10408 14716 10464
rect 14036 10374 14088 10408
rect 14122 10374 14178 10408
rect 14212 10374 14268 10408
rect 14302 10374 14358 10408
rect 14392 10374 14448 10408
rect 14482 10374 14538 10408
rect 14572 10374 14628 10408
rect 14662 10374 14716 10408
rect 14036 10318 14716 10374
rect 14036 10284 14088 10318
rect 14122 10284 14178 10318
rect 14212 10284 14268 10318
rect 14302 10284 14358 10318
rect 14392 10284 14448 10318
rect 14482 10284 14538 10318
rect 14572 10284 14628 10318
rect 14662 10284 14716 10318
rect 14036 10228 14716 10284
rect 14036 10194 14088 10228
rect 14122 10194 14178 10228
rect 14212 10194 14268 10228
rect 14302 10194 14358 10228
rect 14392 10194 14448 10228
rect 14482 10194 14538 10228
rect 14572 10194 14628 10228
rect 14662 10194 14716 10228
rect 14036 10138 14716 10194
rect 14036 10104 14088 10138
rect 14122 10104 14178 10138
rect 14212 10104 14268 10138
rect 14302 10104 14358 10138
rect 14392 10104 14448 10138
rect 14482 10104 14538 10138
rect 14572 10104 14628 10138
rect 14662 10104 14716 10138
rect 14036 10048 14716 10104
rect 14036 10014 14088 10048
rect 14122 10014 14178 10048
rect 14212 10014 14268 10048
rect 14302 10014 14358 10048
rect 14392 10014 14448 10048
rect 14482 10014 14538 10048
rect 14572 10014 14628 10048
rect 14662 10014 14716 10048
rect 14036 9962 14716 10014
rect 15324 10588 16004 10642
rect 15324 10554 15376 10588
rect 15410 10554 15466 10588
rect 15500 10554 15556 10588
rect 15590 10554 15646 10588
rect 15680 10554 15736 10588
rect 15770 10554 15826 10588
rect 15860 10554 15916 10588
rect 15950 10554 16004 10588
rect 15324 10498 16004 10554
rect 15324 10464 15376 10498
rect 15410 10464 15466 10498
rect 15500 10464 15556 10498
rect 15590 10464 15646 10498
rect 15680 10464 15736 10498
rect 15770 10464 15826 10498
rect 15860 10464 15916 10498
rect 15950 10464 16004 10498
rect 15324 10408 16004 10464
rect 15324 10374 15376 10408
rect 15410 10374 15466 10408
rect 15500 10374 15556 10408
rect 15590 10374 15646 10408
rect 15680 10374 15736 10408
rect 15770 10374 15826 10408
rect 15860 10374 15916 10408
rect 15950 10374 16004 10408
rect 15324 10318 16004 10374
rect 15324 10284 15376 10318
rect 15410 10284 15466 10318
rect 15500 10284 15556 10318
rect 15590 10284 15646 10318
rect 15680 10284 15736 10318
rect 15770 10284 15826 10318
rect 15860 10284 15916 10318
rect 15950 10284 16004 10318
rect 15324 10228 16004 10284
rect 15324 10194 15376 10228
rect 15410 10194 15466 10228
rect 15500 10194 15556 10228
rect 15590 10194 15646 10228
rect 15680 10194 15736 10228
rect 15770 10194 15826 10228
rect 15860 10194 15916 10228
rect 15950 10194 16004 10228
rect 15324 10138 16004 10194
rect 15324 10104 15376 10138
rect 15410 10104 15466 10138
rect 15500 10104 15556 10138
rect 15590 10104 15646 10138
rect 15680 10104 15736 10138
rect 15770 10104 15826 10138
rect 15860 10104 15916 10138
rect 15950 10104 16004 10138
rect 15324 10048 16004 10104
rect 15324 10014 15376 10048
rect 15410 10014 15466 10048
rect 15500 10014 15556 10048
rect 15590 10014 15646 10048
rect 15680 10014 15736 10048
rect 15770 10014 15826 10048
rect 15860 10014 15916 10048
rect 15950 10014 16004 10048
rect 15324 9962 16004 10014
rect 16612 10588 17292 10642
rect 16612 10554 16664 10588
rect 16698 10554 16754 10588
rect 16788 10554 16844 10588
rect 16878 10554 16934 10588
rect 16968 10554 17024 10588
rect 17058 10554 17114 10588
rect 17148 10554 17204 10588
rect 17238 10554 17292 10588
rect 16612 10498 17292 10554
rect 16612 10464 16664 10498
rect 16698 10464 16754 10498
rect 16788 10464 16844 10498
rect 16878 10464 16934 10498
rect 16968 10464 17024 10498
rect 17058 10464 17114 10498
rect 17148 10464 17204 10498
rect 17238 10464 17292 10498
rect 16612 10408 17292 10464
rect 16612 10374 16664 10408
rect 16698 10374 16754 10408
rect 16788 10374 16844 10408
rect 16878 10374 16934 10408
rect 16968 10374 17024 10408
rect 17058 10374 17114 10408
rect 17148 10374 17204 10408
rect 17238 10374 17292 10408
rect 16612 10318 17292 10374
rect 16612 10284 16664 10318
rect 16698 10284 16754 10318
rect 16788 10284 16844 10318
rect 16878 10284 16934 10318
rect 16968 10284 17024 10318
rect 17058 10284 17114 10318
rect 17148 10284 17204 10318
rect 17238 10284 17292 10318
rect 16612 10228 17292 10284
rect 16612 10194 16664 10228
rect 16698 10194 16754 10228
rect 16788 10194 16844 10228
rect 16878 10194 16934 10228
rect 16968 10194 17024 10228
rect 17058 10194 17114 10228
rect 17148 10194 17204 10228
rect 17238 10194 17292 10228
rect 16612 10138 17292 10194
rect 16612 10104 16664 10138
rect 16698 10104 16754 10138
rect 16788 10104 16844 10138
rect 16878 10104 16934 10138
rect 16968 10104 17024 10138
rect 17058 10104 17114 10138
rect 17148 10104 17204 10138
rect 17238 10104 17292 10138
rect 16612 10048 17292 10104
rect 16612 10014 16664 10048
rect 16698 10014 16754 10048
rect 16788 10014 16844 10048
rect 16878 10014 16934 10048
rect 16968 10014 17024 10048
rect 17058 10014 17114 10048
rect 17148 10014 17204 10048
rect 17238 10014 17292 10048
rect 16612 9962 17292 10014
rect 17900 10588 18580 10642
rect 17900 10554 17952 10588
rect 17986 10554 18042 10588
rect 18076 10554 18132 10588
rect 18166 10554 18222 10588
rect 18256 10554 18312 10588
rect 18346 10554 18402 10588
rect 18436 10554 18492 10588
rect 18526 10554 18580 10588
rect 17900 10498 18580 10554
rect 17900 10464 17952 10498
rect 17986 10464 18042 10498
rect 18076 10464 18132 10498
rect 18166 10464 18222 10498
rect 18256 10464 18312 10498
rect 18346 10464 18402 10498
rect 18436 10464 18492 10498
rect 18526 10464 18580 10498
rect 17900 10408 18580 10464
rect 17900 10374 17952 10408
rect 17986 10374 18042 10408
rect 18076 10374 18132 10408
rect 18166 10374 18222 10408
rect 18256 10374 18312 10408
rect 18346 10374 18402 10408
rect 18436 10374 18492 10408
rect 18526 10374 18580 10408
rect 17900 10318 18580 10374
rect 17900 10284 17952 10318
rect 17986 10284 18042 10318
rect 18076 10284 18132 10318
rect 18166 10284 18222 10318
rect 18256 10284 18312 10318
rect 18346 10284 18402 10318
rect 18436 10284 18492 10318
rect 18526 10284 18580 10318
rect 17900 10228 18580 10284
rect 17900 10194 17952 10228
rect 17986 10194 18042 10228
rect 18076 10194 18132 10228
rect 18166 10194 18222 10228
rect 18256 10194 18312 10228
rect 18346 10194 18402 10228
rect 18436 10194 18492 10228
rect 18526 10194 18580 10228
rect 17900 10138 18580 10194
rect 17900 10104 17952 10138
rect 17986 10104 18042 10138
rect 18076 10104 18132 10138
rect 18166 10104 18222 10138
rect 18256 10104 18312 10138
rect 18346 10104 18402 10138
rect 18436 10104 18492 10138
rect 18526 10104 18580 10138
rect 17900 10048 18580 10104
rect 17900 10014 17952 10048
rect 17986 10014 18042 10048
rect 18076 10014 18132 10048
rect 18166 10014 18222 10048
rect 18256 10014 18312 10048
rect 18346 10014 18402 10048
rect 18436 10014 18492 10048
rect 18526 10014 18580 10048
rect 17900 9962 18580 10014
rect -8812 9428 -8754 9440
rect -18620 4230 -18562 4242
rect -18620 1674 -18608 4230
rect -18574 1674 -18562 4230
rect -18620 1662 -18562 1674
rect -18162 4230 -18104 4242
rect -18162 1674 -18150 4230
rect -18116 1674 -18104 4230
rect -18162 1662 -18104 1674
rect -18048 4230 -17990 4242
rect -18048 1674 -18036 4230
rect -18002 1674 -17990 4230
rect -18048 1662 -17990 1674
rect -17590 4230 -17532 4242
rect -17590 1674 -17578 4230
rect -17544 1674 -17532 4230
rect -17590 1662 -17532 1674
rect -17476 4230 -17418 4242
rect -17476 1674 -17464 4230
rect -17430 1674 -17418 4230
rect -17476 1662 -17418 1674
rect -17018 4230 -16960 4242
rect -17018 1674 -17006 4230
rect -16972 1674 -16960 4230
rect -17018 1662 -16960 1674
rect -16904 4230 -16846 4242
rect -16904 1674 -16892 4230
rect -16858 1674 -16846 4230
rect -16904 1662 -16846 1674
rect -16446 4230 -16388 4242
rect -16446 1674 -16434 4230
rect -16400 1674 -16388 4230
rect -16446 1662 -16388 1674
rect -16332 4230 -16274 4242
rect -16332 1674 -16320 4230
rect -16286 1674 -16274 4230
rect -16332 1662 -16274 1674
rect -15874 4230 -15816 4242
rect -15874 1674 -15862 4230
rect -15828 1674 -15816 4230
rect -15874 1662 -15816 1674
rect -15760 4230 -15702 4242
rect -15760 1674 -15748 4230
rect -15714 1674 -15702 4230
rect -15760 1662 -15702 1674
rect -15302 4230 -15244 4242
rect -15302 1674 -15290 4230
rect -15256 1674 -15244 4230
rect -15302 1662 -15244 1674
rect -15188 4230 -15130 4242
rect -15188 1674 -15176 4230
rect -15142 1674 -15130 4230
rect -15188 1662 -15130 1674
rect -14730 4230 -14672 4242
rect -14730 1674 -14718 4230
rect -14684 1674 -14672 4230
rect -14730 1662 -14672 1674
rect -14616 4230 -14558 4242
rect -14616 1674 -14604 4230
rect -14570 1674 -14558 4230
rect -14616 1662 -14558 1674
rect -14158 4230 -14100 4242
rect -14158 1674 -14146 4230
rect -14112 1674 -14100 4230
rect -14158 1662 -14100 1674
rect -14044 4230 -13986 4242
rect -14044 1674 -14032 4230
rect -13998 1674 -13986 4230
rect -14044 1662 -13986 1674
rect -13586 4230 -13528 4242
rect -13586 1674 -13574 4230
rect -13540 1674 -13528 4230
rect -13586 1662 -13528 1674
rect -13472 4230 -13414 4242
rect -13472 1674 -13460 4230
rect -13426 1674 -13414 4230
rect -13472 1662 -13414 1674
rect -13014 4230 -12956 4242
rect -13014 1674 -13002 4230
rect -12968 1674 -12956 4230
rect -13014 1662 -12956 1674
rect -12900 4230 -12842 4242
rect -12900 1674 -12888 4230
rect -12854 1674 -12842 4230
rect -12900 1662 -12842 1674
rect -12442 4230 -12384 4242
rect -12442 1674 -12430 4230
rect -12396 1674 -12384 4230
rect -12442 1662 -12384 1674
rect -12328 4230 -12270 4242
rect -12328 1674 -12316 4230
rect -12282 1674 -12270 4230
rect -12328 1662 -12270 1674
rect -11870 4230 -11812 4242
rect -11870 1674 -11858 4230
rect -11824 1674 -11812 4230
rect -11870 1662 -11812 1674
rect -11756 4230 -11698 4242
rect -11756 1674 -11744 4230
rect -11710 1674 -11698 4230
rect -11756 1662 -11698 1674
rect -11298 4230 -11240 4242
rect -11298 1674 -11286 4230
rect -11252 1674 -11240 4230
rect -11298 1662 -11240 1674
rect -11184 4230 -11126 4242
rect -11184 1674 -11172 4230
rect -11138 1674 -11126 4230
rect -11184 1662 -11126 1674
rect -10726 4230 -10668 4242
rect -10726 1674 -10714 4230
rect -10680 1674 -10668 4230
rect -8812 1712 -8800 9428
rect -8766 1712 -8754 9428
rect -8812 1700 -8754 1712
rect -8354 9428 -8296 9440
rect -8354 1712 -8342 9428
rect -8308 1712 -8296 9428
rect -8354 1700 -8296 1712
rect -7896 9428 -7838 9440
rect -7896 1712 -7884 9428
rect -7850 1712 -7838 9428
rect -7896 1700 -7838 1712
rect -7438 9428 -7380 9440
rect -7438 1712 -7426 9428
rect -7392 1712 -7380 9428
rect -7438 1700 -7380 1712
rect -6980 9428 -6922 9440
rect -6980 1712 -6968 9428
rect -6934 1712 -6922 9428
rect -6980 1700 -6922 1712
rect -6522 9428 -6464 9440
rect -6522 1712 -6510 9428
rect -6476 1712 -6464 9428
rect -6522 1700 -6464 1712
rect -6064 9428 -6006 9440
rect -6064 1712 -6052 9428
rect -6018 1712 -6006 9428
rect -6064 1700 -6006 1712
rect -5606 9428 -5548 9440
rect -5606 1712 -5594 9428
rect -5560 1712 -5548 9428
rect -5606 1700 -5548 1712
rect -5148 9428 -5090 9440
rect -5148 1712 -5136 9428
rect -5102 1712 -5090 9428
rect -5148 1700 -5090 1712
rect -4690 9428 -4632 9440
rect -4690 1712 -4678 9428
rect -4644 1712 -4632 9428
rect -4690 1700 -4632 1712
rect -4232 9428 -4174 9440
rect -4232 1712 -4220 9428
rect -4186 1712 -4174 9428
rect -4232 1700 -4174 1712
rect -3774 9428 -3716 9440
rect -3774 1712 -3762 9428
rect -3728 1712 -3716 9428
rect -2854 9428 -2796 9440
rect -3774 1700 -3716 1712
rect -2854 1712 -2842 9428
rect -2808 1712 -2796 9428
rect -2854 1700 -2796 1712
rect -2396 9428 -2338 9440
rect -2396 1712 -2384 9428
rect -2350 1712 -2338 9428
rect -2396 1700 -2338 1712
rect -1938 9428 -1880 9440
rect -1938 1712 -1926 9428
rect -1892 1712 -1880 9428
rect -1938 1700 -1880 1712
rect -1480 9428 -1422 9440
rect -1480 1712 -1468 9428
rect -1434 1712 -1422 9428
rect -1480 1700 -1422 1712
rect -1022 9428 -964 9440
rect -1022 1712 -1010 9428
rect -976 1712 -964 9428
rect -1022 1700 -964 1712
rect -564 9428 -506 9440
rect -564 1712 -552 9428
rect -518 1712 -506 9428
rect -564 1700 -506 1712
rect -106 9428 -48 9440
rect -106 1712 -94 9428
rect -60 1712 -48 9428
rect -106 1700 -48 1712
rect 352 9428 410 9440
rect 352 1712 364 9428
rect 398 1712 410 9428
rect 352 1700 410 1712
rect 810 9428 868 9440
rect 810 1712 822 9428
rect 856 1712 868 9428
rect 810 1700 868 1712
rect 1268 9428 1326 9440
rect 1268 1712 1280 9428
rect 1314 1712 1326 9428
rect 1268 1700 1326 1712
rect 1726 9428 1784 9440
rect 1726 1712 1738 9428
rect 1772 1712 1784 9428
rect 2646 9428 2704 9440
rect 1726 1700 1784 1712
rect 2646 1712 2658 9428
rect 2692 1712 2704 9428
rect 2646 1700 2704 1712
rect 3104 9428 3162 9440
rect 3104 1712 3116 9428
rect 3150 1712 3162 9428
rect 3104 1700 3162 1712
rect 3562 9428 3620 9440
rect 3562 1712 3574 9428
rect 3608 1712 3620 9428
rect 3562 1700 3620 1712
rect 4020 9428 4078 9440
rect 4020 1712 4032 9428
rect 4066 1712 4078 9428
rect 4020 1700 4078 1712
rect 4478 9428 4536 9440
rect 4478 1712 4490 9428
rect 4524 1712 4536 9428
rect 4478 1700 4536 1712
rect 4936 9428 4994 9440
rect 4936 1712 4948 9428
rect 4982 1712 4994 9428
rect 4936 1700 4994 1712
rect 5394 9428 5452 9440
rect 5394 1712 5406 9428
rect 5440 1712 5452 9428
rect 5394 1700 5452 1712
rect 5852 9428 5910 9440
rect 5852 1712 5864 9428
rect 5898 1712 5910 9428
rect 5852 1700 5910 1712
rect 6310 9428 6368 9440
rect 6310 1712 6322 9428
rect 6356 1712 6368 9428
rect 6310 1700 6368 1712
rect 6768 9428 6826 9440
rect 6768 1712 6780 9428
rect 6814 1712 6826 9428
rect 6768 1700 6826 1712
rect 7226 9428 7284 9440
rect 7226 1712 7238 9428
rect 7272 1712 7284 9428
rect 7226 1700 7284 1712
rect 7684 9428 7742 9440
rect 7684 1712 7696 9428
rect 7730 1712 7742 9428
rect 12748 9300 13428 9354
rect 12748 9266 12800 9300
rect 12834 9266 12890 9300
rect 12924 9266 12980 9300
rect 13014 9266 13070 9300
rect 13104 9266 13160 9300
rect 13194 9266 13250 9300
rect 13284 9266 13340 9300
rect 13374 9266 13428 9300
rect 12748 9210 13428 9266
rect 12748 9176 12800 9210
rect 12834 9176 12890 9210
rect 12924 9176 12980 9210
rect 13014 9176 13070 9210
rect 13104 9176 13160 9210
rect 13194 9176 13250 9210
rect 13284 9176 13340 9210
rect 13374 9176 13428 9210
rect 12748 9120 13428 9176
rect 12748 9086 12800 9120
rect 12834 9086 12890 9120
rect 12924 9086 12980 9120
rect 13014 9086 13070 9120
rect 13104 9086 13160 9120
rect 13194 9086 13250 9120
rect 13284 9086 13340 9120
rect 13374 9086 13428 9120
rect 12748 9030 13428 9086
rect 12748 8996 12800 9030
rect 12834 8996 12890 9030
rect 12924 8996 12980 9030
rect 13014 8996 13070 9030
rect 13104 8996 13160 9030
rect 13194 8996 13250 9030
rect 13284 8996 13340 9030
rect 13374 8996 13428 9030
rect 12748 8940 13428 8996
rect 12748 8906 12800 8940
rect 12834 8906 12890 8940
rect 12924 8906 12980 8940
rect 13014 8906 13070 8940
rect 13104 8906 13160 8940
rect 13194 8906 13250 8940
rect 13284 8906 13340 8940
rect 13374 8906 13428 8940
rect 12748 8850 13428 8906
rect 12748 8816 12800 8850
rect 12834 8816 12890 8850
rect 12924 8816 12980 8850
rect 13014 8816 13070 8850
rect 13104 8816 13160 8850
rect 13194 8816 13250 8850
rect 13284 8816 13340 8850
rect 13374 8816 13428 8850
rect 12748 8760 13428 8816
rect 12748 8726 12800 8760
rect 12834 8726 12890 8760
rect 12924 8726 12980 8760
rect 13014 8726 13070 8760
rect 13104 8726 13160 8760
rect 13194 8726 13250 8760
rect 13284 8726 13340 8760
rect 13374 8726 13428 8760
rect 12748 8674 13428 8726
rect 14036 9300 14716 9354
rect 14036 9266 14088 9300
rect 14122 9266 14178 9300
rect 14212 9266 14268 9300
rect 14302 9266 14358 9300
rect 14392 9266 14448 9300
rect 14482 9266 14538 9300
rect 14572 9266 14628 9300
rect 14662 9266 14716 9300
rect 14036 9210 14716 9266
rect 14036 9176 14088 9210
rect 14122 9176 14178 9210
rect 14212 9176 14268 9210
rect 14302 9176 14358 9210
rect 14392 9176 14448 9210
rect 14482 9176 14538 9210
rect 14572 9176 14628 9210
rect 14662 9176 14716 9210
rect 14036 9120 14716 9176
rect 14036 9086 14088 9120
rect 14122 9086 14178 9120
rect 14212 9086 14268 9120
rect 14302 9086 14358 9120
rect 14392 9086 14448 9120
rect 14482 9086 14538 9120
rect 14572 9086 14628 9120
rect 14662 9086 14716 9120
rect 14036 9030 14716 9086
rect 14036 8996 14088 9030
rect 14122 8996 14178 9030
rect 14212 8996 14268 9030
rect 14302 8996 14358 9030
rect 14392 8996 14448 9030
rect 14482 8996 14538 9030
rect 14572 8996 14628 9030
rect 14662 8996 14716 9030
rect 14036 8940 14716 8996
rect 14036 8906 14088 8940
rect 14122 8906 14178 8940
rect 14212 8906 14268 8940
rect 14302 8906 14358 8940
rect 14392 8906 14448 8940
rect 14482 8906 14538 8940
rect 14572 8906 14628 8940
rect 14662 8906 14716 8940
rect 14036 8850 14716 8906
rect 14036 8816 14088 8850
rect 14122 8816 14178 8850
rect 14212 8816 14268 8850
rect 14302 8816 14358 8850
rect 14392 8816 14448 8850
rect 14482 8816 14538 8850
rect 14572 8816 14628 8850
rect 14662 8816 14716 8850
rect 14036 8760 14716 8816
rect 14036 8726 14088 8760
rect 14122 8726 14178 8760
rect 14212 8726 14268 8760
rect 14302 8726 14358 8760
rect 14392 8726 14448 8760
rect 14482 8726 14538 8760
rect 14572 8726 14628 8760
rect 14662 8726 14716 8760
rect 14036 8674 14716 8726
rect 15324 9300 16004 9354
rect 15324 9266 15376 9300
rect 15410 9266 15466 9300
rect 15500 9266 15556 9300
rect 15590 9266 15646 9300
rect 15680 9266 15736 9300
rect 15770 9266 15826 9300
rect 15860 9266 15916 9300
rect 15950 9266 16004 9300
rect 15324 9210 16004 9266
rect 15324 9176 15376 9210
rect 15410 9176 15466 9210
rect 15500 9176 15556 9210
rect 15590 9176 15646 9210
rect 15680 9176 15736 9210
rect 15770 9176 15826 9210
rect 15860 9176 15916 9210
rect 15950 9176 16004 9210
rect 15324 9120 16004 9176
rect 15324 9086 15376 9120
rect 15410 9086 15466 9120
rect 15500 9086 15556 9120
rect 15590 9086 15646 9120
rect 15680 9086 15736 9120
rect 15770 9086 15826 9120
rect 15860 9086 15916 9120
rect 15950 9086 16004 9120
rect 15324 9030 16004 9086
rect 15324 8996 15376 9030
rect 15410 8996 15466 9030
rect 15500 8996 15556 9030
rect 15590 8996 15646 9030
rect 15680 8996 15736 9030
rect 15770 8996 15826 9030
rect 15860 8996 15916 9030
rect 15950 8996 16004 9030
rect 15324 8940 16004 8996
rect 15324 8906 15376 8940
rect 15410 8906 15466 8940
rect 15500 8906 15556 8940
rect 15590 8906 15646 8940
rect 15680 8906 15736 8940
rect 15770 8906 15826 8940
rect 15860 8906 15916 8940
rect 15950 8906 16004 8940
rect 15324 8850 16004 8906
rect 15324 8816 15376 8850
rect 15410 8816 15466 8850
rect 15500 8816 15556 8850
rect 15590 8816 15646 8850
rect 15680 8816 15736 8850
rect 15770 8816 15826 8850
rect 15860 8816 15916 8850
rect 15950 8816 16004 8850
rect 15324 8760 16004 8816
rect 15324 8726 15376 8760
rect 15410 8726 15466 8760
rect 15500 8726 15556 8760
rect 15590 8726 15646 8760
rect 15680 8726 15736 8760
rect 15770 8726 15826 8760
rect 15860 8726 15916 8760
rect 15950 8726 16004 8760
rect 15324 8674 16004 8726
rect 16612 9300 17292 9354
rect 16612 9266 16664 9300
rect 16698 9266 16754 9300
rect 16788 9266 16844 9300
rect 16878 9266 16934 9300
rect 16968 9266 17024 9300
rect 17058 9266 17114 9300
rect 17148 9266 17204 9300
rect 17238 9266 17292 9300
rect 16612 9210 17292 9266
rect 16612 9176 16664 9210
rect 16698 9176 16754 9210
rect 16788 9176 16844 9210
rect 16878 9176 16934 9210
rect 16968 9176 17024 9210
rect 17058 9176 17114 9210
rect 17148 9176 17204 9210
rect 17238 9176 17292 9210
rect 16612 9120 17292 9176
rect 16612 9086 16664 9120
rect 16698 9086 16754 9120
rect 16788 9086 16844 9120
rect 16878 9086 16934 9120
rect 16968 9086 17024 9120
rect 17058 9086 17114 9120
rect 17148 9086 17204 9120
rect 17238 9086 17292 9120
rect 16612 9030 17292 9086
rect 16612 8996 16664 9030
rect 16698 8996 16754 9030
rect 16788 8996 16844 9030
rect 16878 8996 16934 9030
rect 16968 8996 17024 9030
rect 17058 8996 17114 9030
rect 17148 8996 17204 9030
rect 17238 8996 17292 9030
rect 16612 8940 17292 8996
rect 16612 8906 16664 8940
rect 16698 8906 16754 8940
rect 16788 8906 16844 8940
rect 16878 8906 16934 8940
rect 16968 8906 17024 8940
rect 17058 8906 17114 8940
rect 17148 8906 17204 8940
rect 17238 8906 17292 8940
rect 16612 8850 17292 8906
rect 16612 8816 16664 8850
rect 16698 8816 16754 8850
rect 16788 8816 16844 8850
rect 16878 8816 16934 8850
rect 16968 8816 17024 8850
rect 17058 8816 17114 8850
rect 17148 8816 17204 8850
rect 17238 8816 17292 8850
rect 16612 8760 17292 8816
rect 16612 8726 16664 8760
rect 16698 8726 16754 8760
rect 16788 8726 16844 8760
rect 16878 8726 16934 8760
rect 16968 8726 17024 8760
rect 17058 8726 17114 8760
rect 17148 8726 17204 8760
rect 17238 8726 17292 8760
rect 16612 8674 17292 8726
rect 17900 9300 18580 9354
rect 17900 9266 17952 9300
rect 17986 9266 18042 9300
rect 18076 9266 18132 9300
rect 18166 9266 18222 9300
rect 18256 9266 18312 9300
rect 18346 9266 18402 9300
rect 18436 9266 18492 9300
rect 18526 9266 18580 9300
rect 17900 9210 18580 9266
rect 17900 9176 17952 9210
rect 17986 9176 18042 9210
rect 18076 9176 18132 9210
rect 18166 9176 18222 9210
rect 18256 9176 18312 9210
rect 18346 9176 18402 9210
rect 18436 9176 18492 9210
rect 18526 9176 18580 9210
rect 17900 9120 18580 9176
rect 17900 9086 17952 9120
rect 17986 9086 18042 9120
rect 18076 9086 18132 9120
rect 18166 9086 18222 9120
rect 18256 9086 18312 9120
rect 18346 9086 18402 9120
rect 18436 9086 18492 9120
rect 18526 9086 18580 9120
rect 17900 9030 18580 9086
rect 17900 8996 17952 9030
rect 17986 8996 18042 9030
rect 18076 8996 18132 9030
rect 18166 8996 18222 9030
rect 18256 8996 18312 9030
rect 18346 8996 18402 9030
rect 18436 8996 18492 9030
rect 18526 8996 18580 9030
rect 17900 8940 18580 8996
rect 17900 8906 17952 8940
rect 17986 8906 18042 8940
rect 18076 8906 18132 8940
rect 18166 8906 18222 8940
rect 18256 8906 18312 8940
rect 18346 8906 18402 8940
rect 18436 8906 18492 8940
rect 18526 8906 18580 8940
rect 17900 8850 18580 8906
rect 17900 8816 17952 8850
rect 17986 8816 18042 8850
rect 18076 8816 18132 8850
rect 18166 8816 18222 8850
rect 18256 8816 18312 8850
rect 18346 8816 18402 8850
rect 18436 8816 18492 8850
rect 18526 8816 18580 8850
rect 17900 8760 18580 8816
rect 17900 8726 17952 8760
rect 17986 8726 18042 8760
rect 18076 8726 18132 8760
rect 18166 8726 18222 8760
rect 18256 8726 18312 8760
rect 18346 8726 18402 8760
rect 18436 8726 18492 8760
rect 18526 8726 18580 8760
rect 17900 8674 18580 8726
rect 12748 8012 13428 8066
rect 12748 7978 12800 8012
rect 12834 7978 12890 8012
rect 12924 7978 12980 8012
rect 13014 7978 13070 8012
rect 13104 7978 13160 8012
rect 13194 7978 13250 8012
rect 13284 7978 13340 8012
rect 13374 7978 13428 8012
rect 12748 7922 13428 7978
rect 12748 7888 12800 7922
rect 12834 7888 12890 7922
rect 12924 7888 12980 7922
rect 13014 7888 13070 7922
rect 13104 7888 13160 7922
rect 13194 7888 13250 7922
rect 13284 7888 13340 7922
rect 13374 7888 13428 7922
rect 12748 7832 13428 7888
rect 12748 7798 12800 7832
rect 12834 7798 12890 7832
rect 12924 7798 12980 7832
rect 13014 7798 13070 7832
rect 13104 7798 13160 7832
rect 13194 7798 13250 7832
rect 13284 7798 13340 7832
rect 13374 7798 13428 7832
rect 12748 7742 13428 7798
rect 12748 7708 12800 7742
rect 12834 7708 12890 7742
rect 12924 7708 12980 7742
rect 13014 7708 13070 7742
rect 13104 7708 13160 7742
rect 13194 7708 13250 7742
rect 13284 7708 13340 7742
rect 13374 7708 13428 7742
rect 12748 7652 13428 7708
rect 12748 7618 12800 7652
rect 12834 7618 12890 7652
rect 12924 7618 12980 7652
rect 13014 7618 13070 7652
rect 13104 7618 13160 7652
rect 13194 7618 13250 7652
rect 13284 7618 13340 7652
rect 13374 7618 13428 7652
rect 12748 7562 13428 7618
rect 12748 7528 12800 7562
rect 12834 7528 12890 7562
rect 12924 7528 12980 7562
rect 13014 7528 13070 7562
rect 13104 7528 13160 7562
rect 13194 7528 13250 7562
rect 13284 7528 13340 7562
rect 13374 7528 13428 7562
rect 12748 7472 13428 7528
rect 12748 7438 12800 7472
rect 12834 7438 12890 7472
rect 12924 7438 12980 7472
rect 13014 7438 13070 7472
rect 13104 7438 13160 7472
rect 13194 7438 13250 7472
rect 13284 7438 13340 7472
rect 13374 7438 13428 7472
rect 12748 7386 13428 7438
rect 14036 8012 14716 8066
rect 14036 7978 14088 8012
rect 14122 7978 14178 8012
rect 14212 7978 14268 8012
rect 14302 7978 14358 8012
rect 14392 7978 14448 8012
rect 14482 7978 14538 8012
rect 14572 7978 14628 8012
rect 14662 7978 14716 8012
rect 14036 7922 14716 7978
rect 14036 7888 14088 7922
rect 14122 7888 14178 7922
rect 14212 7888 14268 7922
rect 14302 7888 14358 7922
rect 14392 7888 14448 7922
rect 14482 7888 14538 7922
rect 14572 7888 14628 7922
rect 14662 7888 14716 7922
rect 14036 7832 14716 7888
rect 14036 7798 14088 7832
rect 14122 7798 14178 7832
rect 14212 7798 14268 7832
rect 14302 7798 14358 7832
rect 14392 7798 14448 7832
rect 14482 7798 14538 7832
rect 14572 7798 14628 7832
rect 14662 7798 14716 7832
rect 14036 7742 14716 7798
rect 14036 7708 14088 7742
rect 14122 7708 14178 7742
rect 14212 7708 14268 7742
rect 14302 7708 14358 7742
rect 14392 7708 14448 7742
rect 14482 7708 14538 7742
rect 14572 7708 14628 7742
rect 14662 7708 14716 7742
rect 14036 7652 14716 7708
rect 14036 7618 14088 7652
rect 14122 7618 14178 7652
rect 14212 7618 14268 7652
rect 14302 7618 14358 7652
rect 14392 7618 14448 7652
rect 14482 7618 14538 7652
rect 14572 7618 14628 7652
rect 14662 7618 14716 7652
rect 14036 7562 14716 7618
rect 14036 7528 14088 7562
rect 14122 7528 14178 7562
rect 14212 7528 14268 7562
rect 14302 7528 14358 7562
rect 14392 7528 14448 7562
rect 14482 7528 14538 7562
rect 14572 7528 14628 7562
rect 14662 7528 14716 7562
rect 14036 7472 14716 7528
rect 14036 7438 14088 7472
rect 14122 7438 14178 7472
rect 14212 7438 14268 7472
rect 14302 7438 14358 7472
rect 14392 7438 14448 7472
rect 14482 7438 14538 7472
rect 14572 7438 14628 7472
rect 14662 7438 14716 7472
rect 14036 7386 14716 7438
rect 15324 8012 16004 8066
rect 15324 7978 15376 8012
rect 15410 7978 15466 8012
rect 15500 7978 15556 8012
rect 15590 7978 15646 8012
rect 15680 7978 15736 8012
rect 15770 7978 15826 8012
rect 15860 7978 15916 8012
rect 15950 7978 16004 8012
rect 15324 7922 16004 7978
rect 15324 7888 15376 7922
rect 15410 7888 15466 7922
rect 15500 7888 15556 7922
rect 15590 7888 15646 7922
rect 15680 7888 15736 7922
rect 15770 7888 15826 7922
rect 15860 7888 15916 7922
rect 15950 7888 16004 7922
rect 15324 7832 16004 7888
rect 15324 7798 15376 7832
rect 15410 7798 15466 7832
rect 15500 7798 15556 7832
rect 15590 7798 15646 7832
rect 15680 7798 15736 7832
rect 15770 7798 15826 7832
rect 15860 7798 15916 7832
rect 15950 7798 16004 7832
rect 15324 7742 16004 7798
rect 15324 7708 15376 7742
rect 15410 7708 15466 7742
rect 15500 7708 15556 7742
rect 15590 7708 15646 7742
rect 15680 7708 15736 7742
rect 15770 7708 15826 7742
rect 15860 7708 15916 7742
rect 15950 7708 16004 7742
rect 15324 7652 16004 7708
rect 15324 7618 15376 7652
rect 15410 7618 15466 7652
rect 15500 7618 15556 7652
rect 15590 7618 15646 7652
rect 15680 7618 15736 7652
rect 15770 7618 15826 7652
rect 15860 7618 15916 7652
rect 15950 7618 16004 7652
rect 15324 7562 16004 7618
rect 15324 7528 15376 7562
rect 15410 7528 15466 7562
rect 15500 7528 15556 7562
rect 15590 7528 15646 7562
rect 15680 7528 15736 7562
rect 15770 7528 15826 7562
rect 15860 7528 15916 7562
rect 15950 7528 16004 7562
rect 15324 7472 16004 7528
rect 15324 7438 15376 7472
rect 15410 7438 15466 7472
rect 15500 7438 15556 7472
rect 15590 7438 15646 7472
rect 15680 7438 15736 7472
rect 15770 7438 15826 7472
rect 15860 7438 15916 7472
rect 15950 7438 16004 7472
rect 15324 7386 16004 7438
rect 16612 8012 17292 8066
rect 16612 7978 16664 8012
rect 16698 7978 16754 8012
rect 16788 7978 16844 8012
rect 16878 7978 16934 8012
rect 16968 7978 17024 8012
rect 17058 7978 17114 8012
rect 17148 7978 17204 8012
rect 17238 7978 17292 8012
rect 16612 7922 17292 7978
rect 16612 7888 16664 7922
rect 16698 7888 16754 7922
rect 16788 7888 16844 7922
rect 16878 7888 16934 7922
rect 16968 7888 17024 7922
rect 17058 7888 17114 7922
rect 17148 7888 17204 7922
rect 17238 7888 17292 7922
rect 16612 7832 17292 7888
rect 16612 7798 16664 7832
rect 16698 7798 16754 7832
rect 16788 7798 16844 7832
rect 16878 7798 16934 7832
rect 16968 7798 17024 7832
rect 17058 7798 17114 7832
rect 17148 7798 17204 7832
rect 17238 7798 17292 7832
rect 16612 7742 17292 7798
rect 16612 7708 16664 7742
rect 16698 7708 16754 7742
rect 16788 7708 16844 7742
rect 16878 7708 16934 7742
rect 16968 7708 17024 7742
rect 17058 7708 17114 7742
rect 17148 7708 17204 7742
rect 17238 7708 17292 7742
rect 16612 7652 17292 7708
rect 16612 7618 16664 7652
rect 16698 7618 16754 7652
rect 16788 7618 16844 7652
rect 16878 7618 16934 7652
rect 16968 7618 17024 7652
rect 17058 7618 17114 7652
rect 17148 7618 17204 7652
rect 17238 7618 17292 7652
rect 16612 7562 17292 7618
rect 16612 7528 16664 7562
rect 16698 7528 16754 7562
rect 16788 7528 16844 7562
rect 16878 7528 16934 7562
rect 16968 7528 17024 7562
rect 17058 7528 17114 7562
rect 17148 7528 17204 7562
rect 17238 7528 17292 7562
rect 16612 7472 17292 7528
rect 16612 7438 16664 7472
rect 16698 7438 16754 7472
rect 16788 7438 16844 7472
rect 16878 7438 16934 7472
rect 16968 7438 17024 7472
rect 17058 7438 17114 7472
rect 17148 7438 17204 7472
rect 17238 7438 17292 7472
rect 16612 7386 17292 7438
rect 17900 8012 18580 8066
rect 17900 7978 17952 8012
rect 17986 7978 18042 8012
rect 18076 7978 18132 8012
rect 18166 7978 18222 8012
rect 18256 7978 18312 8012
rect 18346 7978 18402 8012
rect 18436 7978 18492 8012
rect 18526 7978 18580 8012
rect 17900 7922 18580 7978
rect 17900 7888 17952 7922
rect 17986 7888 18042 7922
rect 18076 7888 18132 7922
rect 18166 7888 18222 7922
rect 18256 7888 18312 7922
rect 18346 7888 18402 7922
rect 18436 7888 18492 7922
rect 18526 7888 18580 7922
rect 17900 7832 18580 7888
rect 17900 7798 17952 7832
rect 17986 7798 18042 7832
rect 18076 7798 18132 7832
rect 18166 7798 18222 7832
rect 18256 7798 18312 7832
rect 18346 7798 18402 7832
rect 18436 7798 18492 7832
rect 18526 7798 18580 7832
rect 17900 7742 18580 7798
rect 17900 7708 17952 7742
rect 17986 7708 18042 7742
rect 18076 7708 18132 7742
rect 18166 7708 18222 7742
rect 18256 7708 18312 7742
rect 18346 7708 18402 7742
rect 18436 7708 18492 7742
rect 18526 7708 18580 7742
rect 17900 7652 18580 7708
rect 17900 7618 17952 7652
rect 17986 7618 18042 7652
rect 18076 7618 18132 7652
rect 18166 7618 18222 7652
rect 18256 7618 18312 7652
rect 18346 7618 18402 7652
rect 18436 7618 18492 7652
rect 18526 7618 18580 7652
rect 17900 7562 18580 7618
rect 17900 7528 17952 7562
rect 17986 7528 18042 7562
rect 18076 7528 18132 7562
rect 18166 7528 18222 7562
rect 18256 7528 18312 7562
rect 18346 7528 18402 7562
rect 18436 7528 18492 7562
rect 18526 7528 18580 7562
rect 17900 7472 18580 7528
rect 17900 7438 17952 7472
rect 17986 7438 18042 7472
rect 18076 7438 18132 7472
rect 18166 7438 18222 7472
rect 18256 7438 18312 7472
rect 18346 7438 18402 7472
rect 18436 7438 18492 7472
rect 18526 7438 18580 7472
rect 17900 7386 18580 7438
rect 12748 6724 13428 6778
rect 12748 6690 12800 6724
rect 12834 6690 12890 6724
rect 12924 6690 12980 6724
rect 13014 6690 13070 6724
rect 13104 6690 13160 6724
rect 13194 6690 13250 6724
rect 13284 6690 13340 6724
rect 13374 6690 13428 6724
rect 12748 6634 13428 6690
rect 12748 6600 12800 6634
rect 12834 6600 12890 6634
rect 12924 6600 12980 6634
rect 13014 6600 13070 6634
rect 13104 6600 13160 6634
rect 13194 6600 13250 6634
rect 13284 6600 13340 6634
rect 13374 6600 13428 6634
rect 12748 6544 13428 6600
rect 12748 6510 12800 6544
rect 12834 6510 12890 6544
rect 12924 6510 12980 6544
rect 13014 6510 13070 6544
rect 13104 6510 13160 6544
rect 13194 6510 13250 6544
rect 13284 6510 13340 6544
rect 13374 6510 13428 6544
rect 12748 6454 13428 6510
rect 12748 6420 12800 6454
rect 12834 6420 12890 6454
rect 12924 6420 12980 6454
rect 13014 6420 13070 6454
rect 13104 6420 13160 6454
rect 13194 6420 13250 6454
rect 13284 6420 13340 6454
rect 13374 6420 13428 6454
rect 12748 6364 13428 6420
rect 12748 6330 12800 6364
rect 12834 6330 12890 6364
rect 12924 6330 12980 6364
rect 13014 6330 13070 6364
rect 13104 6330 13160 6364
rect 13194 6330 13250 6364
rect 13284 6330 13340 6364
rect 13374 6330 13428 6364
rect 12748 6274 13428 6330
rect 12748 6240 12800 6274
rect 12834 6240 12890 6274
rect 12924 6240 12980 6274
rect 13014 6240 13070 6274
rect 13104 6240 13160 6274
rect 13194 6240 13250 6274
rect 13284 6240 13340 6274
rect 13374 6240 13428 6274
rect 12748 6184 13428 6240
rect 12748 6150 12800 6184
rect 12834 6150 12890 6184
rect 12924 6150 12980 6184
rect 13014 6150 13070 6184
rect 13104 6150 13160 6184
rect 13194 6150 13250 6184
rect 13284 6150 13340 6184
rect 13374 6150 13428 6184
rect 12748 6098 13428 6150
rect 14036 6724 14716 6778
rect 14036 6690 14088 6724
rect 14122 6690 14178 6724
rect 14212 6690 14268 6724
rect 14302 6690 14358 6724
rect 14392 6690 14448 6724
rect 14482 6690 14538 6724
rect 14572 6690 14628 6724
rect 14662 6690 14716 6724
rect 14036 6634 14716 6690
rect 14036 6600 14088 6634
rect 14122 6600 14178 6634
rect 14212 6600 14268 6634
rect 14302 6600 14358 6634
rect 14392 6600 14448 6634
rect 14482 6600 14538 6634
rect 14572 6600 14628 6634
rect 14662 6600 14716 6634
rect 14036 6544 14716 6600
rect 14036 6510 14088 6544
rect 14122 6510 14178 6544
rect 14212 6510 14268 6544
rect 14302 6510 14358 6544
rect 14392 6510 14448 6544
rect 14482 6510 14538 6544
rect 14572 6510 14628 6544
rect 14662 6510 14716 6544
rect 14036 6454 14716 6510
rect 14036 6420 14088 6454
rect 14122 6420 14178 6454
rect 14212 6420 14268 6454
rect 14302 6420 14358 6454
rect 14392 6420 14448 6454
rect 14482 6420 14538 6454
rect 14572 6420 14628 6454
rect 14662 6420 14716 6454
rect 14036 6364 14716 6420
rect 14036 6330 14088 6364
rect 14122 6330 14178 6364
rect 14212 6330 14268 6364
rect 14302 6330 14358 6364
rect 14392 6330 14448 6364
rect 14482 6330 14538 6364
rect 14572 6330 14628 6364
rect 14662 6330 14716 6364
rect 14036 6274 14716 6330
rect 14036 6240 14088 6274
rect 14122 6240 14178 6274
rect 14212 6240 14268 6274
rect 14302 6240 14358 6274
rect 14392 6240 14448 6274
rect 14482 6240 14538 6274
rect 14572 6240 14628 6274
rect 14662 6240 14716 6274
rect 14036 6184 14716 6240
rect 14036 6150 14088 6184
rect 14122 6150 14178 6184
rect 14212 6150 14268 6184
rect 14302 6150 14358 6184
rect 14392 6150 14448 6184
rect 14482 6150 14538 6184
rect 14572 6150 14628 6184
rect 14662 6150 14716 6184
rect 14036 6098 14716 6150
rect 15324 6724 16004 6778
rect 15324 6690 15376 6724
rect 15410 6690 15466 6724
rect 15500 6690 15556 6724
rect 15590 6690 15646 6724
rect 15680 6690 15736 6724
rect 15770 6690 15826 6724
rect 15860 6690 15916 6724
rect 15950 6690 16004 6724
rect 15324 6634 16004 6690
rect 15324 6600 15376 6634
rect 15410 6600 15466 6634
rect 15500 6600 15556 6634
rect 15590 6600 15646 6634
rect 15680 6600 15736 6634
rect 15770 6600 15826 6634
rect 15860 6600 15916 6634
rect 15950 6600 16004 6634
rect 15324 6544 16004 6600
rect 15324 6510 15376 6544
rect 15410 6510 15466 6544
rect 15500 6510 15556 6544
rect 15590 6510 15646 6544
rect 15680 6510 15736 6544
rect 15770 6510 15826 6544
rect 15860 6510 15916 6544
rect 15950 6510 16004 6544
rect 15324 6454 16004 6510
rect 15324 6420 15376 6454
rect 15410 6420 15466 6454
rect 15500 6420 15556 6454
rect 15590 6420 15646 6454
rect 15680 6420 15736 6454
rect 15770 6420 15826 6454
rect 15860 6420 15916 6454
rect 15950 6420 16004 6454
rect 15324 6364 16004 6420
rect 15324 6330 15376 6364
rect 15410 6330 15466 6364
rect 15500 6330 15556 6364
rect 15590 6330 15646 6364
rect 15680 6330 15736 6364
rect 15770 6330 15826 6364
rect 15860 6330 15916 6364
rect 15950 6330 16004 6364
rect 15324 6274 16004 6330
rect 15324 6240 15376 6274
rect 15410 6240 15466 6274
rect 15500 6240 15556 6274
rect 15590 6240 15646 6274
rect 15680 6240 15736 6274
rect 15770 6240 15826 6274
rect 15860 6240 15916 6274
rect 15950 6240 16004 6274
rect 15324 6184 16004 6240
rect 15324 6150 15376 6184
rect 15410 6150 15466 6184
rect 15500 6150 15556 6184
rect 15590 6150 15646 6184
rect 15680 6150 15736 6184
rect 15770 6150 15826 6184
rect 15860 6150 15916 6184
rect 15950 6150 16004 6184
rect 15324 6098 16004 6150
rect 16612 6724 17292 6778
rect 16612 6690 16664 6724
rect 16698 6690 16754 6724
rect 16788 6690 16844 6724
rect 16878 6690 16934 6724
rect 16968 6690 17024 6724
rect 17058 6690 17114 6724
rect 17148 6690 17204 6724
rect 17238 6690 17292 6724
rect 16612 6634 17292 6690
rect 16612 6600 16664 6634
rect 16698 6600 16754 6634
rect 16788 6600 16844 6634
rect 16878 6600 16934 6634
rect 16968 6600 17024 6634
rect 17058 6600 17114 6634
rect 17148 6600 17204 6634
rect 17238 6600 17292 6634
rect 16612 6544 17292 6600
rect 16612 6510 16664 6544
rect 16698 6510 16754 6544
rect 16788 6510 16844 6544
rect 16878 6510 16934 6544
rect 16968 6510 17024 6544
rect 17058 6510 17114 6544
rect 17148 6510 17204 6544
rect 17238 6510 17292 6544
rect 16612 6454 17292 6510
rect 16612 6420 16664 6454
rect 16698 6420 16754 6454
rect 16788 6420 16844 6454
rect 16878 6420 16934 6454
rect 16968 6420 17024 6454
rect 17058 6420 17114 6454
rect 17148 6420 17204 6454
rect 17238 6420 17292 6454
rect 16612 6364 17292 6420
rect 16612 6330 16664 6364
rect 16698 6330 16754 6364
rect 16788 6330 16844 6364
rect 16878 6330 16934 6364
rect 16968 6330 17024 6364
rect 17058 6330 17114 6364
rect 17148 6330 17204 6364
rect 17238 6330 17292 6364
rect 16612 6274 17292 6330
rect 16612 6240 16664 6274
rect 16698 6240 16754 6274
rect 16788 6240 16844 6274
rect 16878 6240 16934 6274
rect 16968 6240 17024 6274
rect 17058 6240 17114 6274
rect 17148 6240 17204 6274
rect 17238 6240 17292 6274
rect 16612 6184 17292 6240
rect 16612 6150 16664 6184
rect 16698 6150 16754 6184
rect 16788 6150 16844 6184
rect 16878 6150 16934 6184
rect 16968 6150 17024 6184
rect 17058 6150 17114 6184
rect 17148 6150 17204 6184
rect 17238 6150 17292 6184
rect 16612 6098 17292 6150
rect 17900 6724 18580 6778
rect 17900 6690 17952 6724
rect 17986 6690 18042 6724
rect 18076 6690 18132 6724
rect 18166 6690 18222 6724
rect 18256 6690 18312 6724
rect 18346 6690 18402 6724
rect 18436 6690 18492 6724
rect 18526 6690 18580 6724
rect 17900 6634 18580 6690
rect 17900 6600 17952 6634
rect 17986 6600 18042 6634
rect 18076 6600 18132 6634
rect 18166 6600 18222 6634
rect 18256 6600 18312 6634
rect 18346 6600 18402 6634
rect 18436 6600 18492 6634
rect 18526 6600 18580 6634
rect 17900 6544 18580 6600
rect 17900 6510 17952 6544
rect 17986 6510 18042 6544
rect 18076 6510 18132 6544
rect 18166 6510 18222 6544
rect 18256 6510 18312 6544
rect 18346 6510 18402 6544
rect 18436 6510 18492 6544
rect 18526 6510 18580 6544
rect 17900 6454 18580 6510
rect 17900 6420 17952 6454
rect 17986 6420 18042 6454
rect 18076 6420 18132 6454
rect 18166 6420 18222 6454
rect 18256 6420 18312 6454
rect 18346 6420 18402 6454
rect 18436 6420 18492 6454
rect 18526 6420 18580 6454
rect 17900 6364 18580 6420
rect 17900 6330 17952 6364
rect 17986 6330 18042 6364
rect 18076 6330 18132 6364
rect 18166 6330 18222 6364
rect 18256 6330 18312 6364
rect 18346 6330 18402 6364
rect 18436 6330 18492 6364
rect 18526 6330 18580 6364
rect 17900 6274 18580 6330
rect 17900 6240 17952 6274
rect 17986 6240 18042 6274
rect 18076 6240 18132 6274
rect 18166 6240 18222 6274
rect 18256 6240 18312 6274
rect 18346 6240 18402 6274
rect 18436 6240 18492 6274
rect 18526 6240 18580 6274
rect 17900 6184 18580 6240
rect 17900 6150 17952 6184
rect 17986 6150 18042 6184
rect 18076 6150 18132 6184
rect 18166 6150 18222 6184
rect 18256 6150 18312 6184
rect 18346 6150 18402 6184
rect 18436 6150 18492 6184
rect 18526 6150 18580 6184
rect 17900 6098 18580 6150
rect 12748 5436 13428 5490
rect 12748 5402 12800 5436
rect 12834 5402 12890 5436
rect 12924 5402 12980 5436
rect 13014 5402 13070 5436
rect 13104 5402 13160 5436
rect 13194 5402 13250 5436
rect 13284 5402 13340 5436
rect 13374 5402 13428 5436
rect 12748 5346 13428 5402
rect 12748 5312 12800 5346
rect 12834 5312 12890 5346
rect 12924 5312 12980 5346
rect 13014 5312 13070 5346
rect 13104 5312 13160 5346
rect 13194 5312 13250 5346
rect 13284 5312 13340 5346
rect 13374 5312 13428 5346
rect 12748 5256 13428 5312
rect 12748 5222 12800 5256
rect 12834 5222 12890 5256
rect 12924 5222 12980 5256
rect 13014 5222 13070 5256
rect 13104 5222 13160 5256
rect 13194 5222 13250 5256
rect 13284 5222 13340 5256
rect 13374 5222 13428 5256
rect 12748 5166 13428 5222
rect 12748 5132 12800 5166
rect 12834 5132 12890 5166
rect 12924 5132 12980 5166
rect 13014 5132 13070 5166
rect 13104 5132 13160 5166
rect 13194 5132 13250 5166
rect 13284 5132 13340 5166
rect 13374 5132 13428 5166
rect 12748 5076 13428 5132
rect 12748 5042 12800 5076
rect 12834 5042 12890 5076
rect 12924 5042 12980 5076
rect 13014 5042 13070 5076
rect 13104 5042 13160 5076
rect 13194 5042 13250 5076
rect 13284 5042 13340 5076
rect 13374 5042 13428 5076
rect 12748 4986 13428 5042
rect 12748 4952 12800 4986
rect 12834 4952 12890 4986
rect 12924 4952 12980 4986
rect 13014 4952 13070 4986
rect 13104 4952 13160 4986
rect 13194 4952 13250 4986
rect 13284 4952 13340 4986
rect 13374 4952 13428 4986
rect 12748 4896 13428 4952
rect 12748 4862 12800 4896
rect 12834 4862 12890 4896
rect 12924 4862 12980 4896
rect 13014 4862 13070 4896
rect 13104 4862 13160 4896
rect 13194 4862 13250 4896
rect 13284 4862 13340 4896
rect 13374 4862 13428 4896
rect 12748 4810 13428 4862
rect 14036 5436 14716 5490
rect 14036 5402 14088 5436
rect 14122 5402 14178 5436
rect 14212 5402 14268 5436
rect 14302 5402 14358 5436
rect 14392 5402 14448 5436
rect 14482 5402 14538 5436
rect 14572 5402 14628 5436
rect 14662 5402 14716 5436
rect 14036 5346 14716 5402
rect 14036 5312 14088 5346
rect 14122 5312 14178 5346
rect 14212 5312 14268 5346
rect 14302 5312 14358 5346
rect 14392 5312 14448 5346
rect 14482 5312 14538 5346
rect 14572 5312 14628 5346
rect 14662 5312 14716 5346
rect 14036 5256 14716 5312
rect 14036 5222 14088 5256
rect 14122 5222 14178 5256
rect 14212 5222 14268 5256
rect 14302 5222 14358 5256
rect 14392 5222 14448 5256
rect 14482 5222 14538 5256
rect 14572 5222 14628 5256
rect 14662 5222 14716 5256
rect 14036 5166 14716 5222
rect 14036 5132 14088 5166
rect 14122 5132 14178 5166
rect 14212 5132 14268 5166
rect 14302 5132 14358 5166
rect 14392 5132 14448 5166
rect 14482 5132 14538 5166
rect 14572 5132 14628 5166
rect 14662 5132 14716 5166
rect 14036 5076 14716 5132
rect 14036 5042 14088 5076
rect 14122 5042 14178 5076
rect 14212 5042 14268 5076
rect 14302 5042 14358 5076
rect 14392 5042 14448 5076
rect 14482 5042 14538 5076
rect 14572 5042 14628 5076
rect 14662 5042 14716 5076
rect 14036 4986 14716 5042
rect 14036 4952 14088 4986
rect 14122 4952 14178 4986
rect 14212 4952 14268 4986
rect 14302 4952 14358 4986
rect 14392 4952 14448 4986
rect 14482 4952 14538 4986
rect 14572 4952 14628 4986
rect 14662 4952 14716 4986
rect 14036 4896 14716 4952
rect 14036 4862 14088 4896
rect 14122 4862 14178 4896
rect 14212 4862 14268 4896
rect 14302 4862 14358 4896
rect 14392 4862 14448 4896
rect 14482 4862 14538 4896
rect 14572 4862 14628 4896
rect 14662 4862 14716 4896
rect 14036 4810 14716 4862
rect 15324 5436 16004 5490
rect 15324 5402 15376 5436
rect 15410 5402 15466 5436
rect 15500 5402 15556 5436
rect 15590 5402 15646 5436
rect 15680 5402 15736 5436
rect 15770 5402 15826 5436
rect 15860 5402 15916 5436
rect 15950 5402 16004 5436
rect 15324 5346 16004 5402
rect 15324 5312 15376 5346
rect 15410 5312 15466 5346
rect 15500 5312 15556 5346
rect 15590 5312 15646 5346
rect 15680 5312 15736 5346
rect 15770 5312 15826 5346
rect 15860 5312 15916 5346
rect 15950 5312 16004 5346
rect 15324 5256 16004 5312
rect 15324 5222 15376 5256
rect 15410 5222 15466 5256
rect 15500 5222 15556 5256
rect 15590 5222 15646 5256
rect 15680 5222 15736 5256
rect 15770 5222 15826 5256
rect 15860 5222 15916 5256
rect 15950 5222 16004 5256
rect 15324 5166 16004 5222
rect 15324 5132 15376 5166
rect 15410 5132 15466 5166
rect 15500 5132 15556 5166
rect 15590 5132 15646 5166
rect 15680 5132 15736 5166
rect 15770 5132 15826 5166
rect 15860 5132 15916 5166
rect 15950 5132 16004 5166
rect 15324 5076 16004 5132
rect 15324 5042 15376 5076
rect 15410 5042 15466 5076
rect 15500 5042 15556 5076
rect 15590 5042 15646 5076
rect 15680 5042 15736 5076
rect 15770 5042 15826 5076
rect 15860 5042 15916 5076
rect 15950 5042 16004 5076
rect 15324 4986 16004 5042
rect 15324 4952 15376 4986
rect 15410 4952 15466 4986
rect 15500 4952 15556 4986
rect 15590 4952 15646 4986
rect 15680 4952 15736 4986
rect 15770 4952 15826 4986
rect 15860 4952 15916 4986
rect 15950 4952 16004 4986
rect 15324 4896 16004 4952
rect 15324 4862 15376 4896
rect 15410 4862 15466 4896
rect 15500 4862 15556 4896
rect 15590 4862 15646 4896
rect 15680 4862 15736 4896
rect 15770 4862 15826 4896
rect 15860 4862 15916 4896
rect 15950 4862 16004 4896
rect 15324 4810 16004 4862
rect 16612 5436 17292 5490
rect 16612 5402 16664 5436
rect 16698 5402 16754 5436
rect 16788 5402 16844 5436
rect 16878 5402 16934 5436
rect 16968 5402 17024 5436
rect 17058 5402 17114 5436
rect 17148 5402 17204 5436
rect 17238 5402 17292 5436
rect 16612 5346 17292 5402
rect 16612 5312 16664 5346
rect 16698 5312 16754 5346
rect 16788 5312 16844 5346
rect 16878 5312 16934 5346
rect 16968 5312 17024 5346
rect 17058 5312 17114 5346
rect 17148 5312 17204 5346
rect 17238 5312 17292 5346
rect 16612 5256 17292 5312
rect 16612 5222 16664 5256
rect 16698 5222 16754 5256
rect 16788 5222 16844 5256
rect 16878 5222 16934 5256
rect 16968 5222 17024 5256
rect 17058 5222 17114 5256
rect 17148 5222 17204 5256
rect 17238 5222 17292 5256
rect 16612 5166 17292 5222
rect 16612 5132 16664 5166
rect 16698 5132 16754 5166
rect 16788 5132 16844 5166
rect 16878 5132 16934 5166
rect 16968 5132 17024 5166
rect 17058 5132 17114 5166
rect 17148 5132 17204 5166
rect 17238 5132 17292 5166
rect 16612 5076 17292 5132
rect 16612 5042 16664 5076
rect 16698 5042 16754 5076
rect 16788 5042 16844 5076
rect 16878 5042 16934 5076
rect 16968 5042 17024 5076
rect 17058 5042 17114 5076
rect 17148 5042 17204 5076
rect 17238 5042 17292 5076
rect 16612 4986 17292 5042
rect 16612 4952 16664 4986
rect 16698 4952 16754 4986
rect 16788 4952 16844 4986
rect 16878 4952 16934 4986
rect 16968 4952 17024 4986
rect 17058 4952 17114 4986
rect 17148 4952 17204 4986
rect 17238 4952 17292 4986
rect 16612 4896 17292 4952
rect 16612 4862 16664 4896
rect 16698 4862 16754 4896
rect 16788 4862 16844 4896
rect 16878 4862 16934 4896
rect 16968 4862 17024 4896
rect 17058 4862 17114 4896
rect 17148 4862 17204 4896
rect 17238 4862 17292 4896
rect 16612 4810 17292 4862
rect 17900 5436 18580 5490
rect 17900 5402 17952 5436
rect 17986 5402 18042 5436
rect 18076 5402 18132 5436
rect 18166 5402 18222 5436
rect 18256 5402 18312 5436
rect 18346 5402 18402 5436
rect 18436 5402 18492 5436
rect 18526 5402 18580 5436
rect 17900 5346 18580 5402
rect 17900 5312 17952 5346
rect 17986 5312 18042 5346
rect 18076 5312 18132 5346
rect 18166 5312 18222 5346
rect 18256 5312 18312 5346
rect 18346 5312 18402 5346
rect 18436 5312 18492 5346
rect 18526 5312 18580 5346
rect 17900 5256 18580 5312
rect 17900 5222 17952 5256
rect 17986 5222 18042 5256
rect 18076 5222 18132 5256
rect 18166 5222 18222 5256
rect 18256 5222 18312 5256
rect 18346 5222 18402 5256
rect 18436 5222 18492 5256
rect 18526 5222 18580 5256
rect 17900 5166 18580 5222
rect 17900 5132 17952 5166
rect 17986 5132 18042 5166
rect 18076 5132 18132 5166
rect 18166 5132 18222 5166
rect 18256 5132 18312 5166
rect 18346 5132 18402 5166
rect 18436 5132 18492 5166
rect 18526 5132 18580 5166
rect 17900 5076 18580 5132
rect 17900 5042 17952 5076
rect 17986 5042 18042 5076
rect 18076 5042 18132 5076
rect 18166 5042 18222 5076
rect 18256 5042 18312 5076
rect 18346 5042 18402 5076
rect 18436 5042 18492 5076
rect 18526 5042 18580 5076
rect 17900 4986 18580 5042
rect 17900 4952 17952 4986
rect 17986 4952 18042 4986
rect 18076 4952 18132 4986
rect 18166 4952 18222 4986
rect 18256 4952 18312 4986
rect 18346 4952 18402 4986
rect 18436 4952 18492 4986
rect 18526 4952 18580 4986
rect 17900 4896 18580 4952
rect 17900 4862 17952 4896
rect 17986 4862 18042 4896
rect 18076 4862 18132 4896
rect 18166 4862 18222 4896
rect 18256 4862 18312 4896
rect 18346 4862 18402 4896
rect 18436 4862 18492 4896
rect 18526 4862 18580 4896
rect 17900 4810 18580 4862
rect 12748 4148 13428 4202
rect 12748 4114 12800 4148
rect 12834 4114 12890 4148
rect 12924 4114 12980 4148
rect 13014 4114 13070 4148
rect 13104 4114 13160 4148
rect 13194 4114 13250 4148
rect 13284 4114 13340 4148
rect 13374 4114 13428 4148
rect 12748 4058 13428 4114
rect 12748 4024 12800 4058
rect 12834 4024 12890 4058
rect 12924 4024 12980 4058
rect 13014 4024 13070 4058
rect 13104 4024 13160 4058
rect 13194 4024 13250 4058
rect 13284 4024 13340 4058
rect 13374 4024 13428 4058
rect 12748 3968 13428 4024
rect 12748 3934 12800 3968
rect 12834 3934 12890 3968
rect 12924 3934 12980 3968
rect 13014 3934 13070 3968
rect 13104 3934 13160 3968
rect 13194 3934 13250 3968
rect 13284 3934 13340 3968
rect 13374 3934 13428 3968
rect 12748 3878 13428 3934
rect 12748 3844 12800 3878
rect 12834 3844 12890 3878
rect 12924 3844 12980 3878
rect 13014 3844 13070 3878
rect 13104 3844 13160 3878
rect 13194 3844 13250 3878
rect 13284 3844 13340 3878
rect 13374 3844 13428 3878
rect 12748 3788 13428 3844
rect 12748 3754 12800 3788
rect 12834 3754 12890 3788
rect 12924 3754 12980 3788
rect 13014 3754 13070 3788
rect 13104 3754 13160 3788
rect 13194 3754 13250 3788
rect 13284 3754 13340 3788
rect 13374 3754 13428 3788
rect 12748 3698 13428 3754
rect 12748 3664 12800 3698
rect 12834 3664 12890 3698
rect 12924 3664 12980 3698
rect 13014 3664 13070 3698
rect 13104 3664 13160 3698
rect 13194 3664 13250 3698
rect 13284 3664 13340 3698
rect 13374 3664 13428 3698
rect 12748 3608 13428 3664
rect 12748 3574 12800 3608
rect 12834 3574 12890 3608
rect 12924 3574 12980 3608
rect 13014 3574 13070 3608
rect 13104 3574 13160 3608
rect 13194 3574 13250 3608
rect 13284 3574 13340 3608
rect 13374 3574 13428 3608
rect 12748 3522 13428 3574
rect 14036 4148 14716 4202
rect 14036 4114 14088 4148
rect 14122 4114 14178 4148
rect 14212 4114 14268 4148
rect 14302 4114 14358 4148
rect 14392 4114 14448 4148
rect 14482 4114 14538 4148
rect 14572 4114 14628 4148
rect 14662 4114 14716 4148
rect 14036 4058 14716 4114
rect 14036 4024 14088 4058
rect 14122 4024 14178 4058
rect 14212 4024 14268 4058
rect 14302 4024 14358 4058
rect 14392 4024 14448 4058
rect 14482 4024 14538 4058
rect 14572 4024 14628 4058
rect 14662 4024 14716 4058
rect 14036 3968 14716 4024
rect 14036 3934 14088 3968
rect 14122 3934 14178 3968
rect 14212 3934 14268 3968
rect 14302 3934 14358 3968
rect 14392 3934 14448 3968
rect 14482 3934 14538 3968
rect 14572 3934 14628 3968
rect 14662 3934 14716 3968
rect 14036 3878 14716 3934
rect 14036 3844 14088 3878
rect 14122 3844 14178 3878
rect 14212 3844 14268 3878
rect 14302 3844 14358 3878
rect 14392 3844 14448 3878
rect 14482 3844 14538 3878
rect 14572 3844 14628 3878
rect 14662 3844 14716 3878
rect 14036 3788 14716 3844
rect 14036 3754 14088 3788
rect 14122 3754 14178 3788
rect 14212 3754 14268 3788
rect 14302 3754 14358 3788
rect 14392 3754 14448 3788
rect 14482 3754 14538 3788
rect 14572 3754 14628 3788
rect 14662 3754 14716 3788
rect 14036 3698 14716 3754
rect 14036 3664 14088 3698
rect 14122 3664 14178 3698
rect 14212 3664 14268 3698
rect 14302 3664 14358 3698
rect 14392 3664 14448 3698
rect 14482 3664 14538 3698
rect 14572 3664 14628 3698
rect 14662 3664 14716 3698
rect 14036 3608 14716 3664
rect 14036 3574 14088 3608
rect 14122 3574 14178 3608
rect 14212 3574 14268 3608
rect 14302 3574 14358 3608
rect 14392 3574 14448 3608
rect 14482 3574 14538 3608
rect 14572 3574 14628 3608
rect 14662 3574 14716 3608
rect 14036 3522 14716 3574
rect 15324 4148 16004 4202
rect 15324 4114 15376 4148
rect 15410 4114 15466 4148
rect 15500 4114 15556 4148
rect 15590 4114 15646 4148
rect 15680 4114 15736 4148
rect 15770 4114 15826 4148
rect 15860 4114 15916 4148
rect 15950 4114 16004 4148
rect 15324 4058 16004 4114
rect 15324 4024 15376 4058
rect 15410 4024 15466 4058
rect 15500 4024 15556 4058
rect 15590 4024 15646 4058
rect 15680 4024 15736 4058
rect 15770 4024 15826 4058
rect 15860 4024 15916 4058
rect 15950 4024 16004 4058
rect 15324 3968 16004 4024
rect 15324 3934 15376 3968
rect 15410 3934 15466 3968
rect 15500 3934 15556 3968
rect 15590 3934 15646 3968
rect 15680 3934 15736 3968
rect 15770 3934 15826 3968
rect 15860 3934 15916 3968
rect 15950 3934 16004 3968
rect 15324 3878 16004 3934
rect 15324 3844 15376 3878
rect 15410 3844 15466 3878
rect 15500 3844 15556 3878
rect 15590 3844 15646 3878
rect 15680 3844 15736 3878
rect 15770 3844 15826 3878
rect 15860 3844 15916 3878
rect 15950 3844 16004 3878
rect 15324 3788 16004 3844
rect 15324 3754 15376 3788
rect 15410 3754 15466 3788
rect 15500 3754 15556 3788
rect 15590 3754 15646 3788
rect 15680 3754 15736 3788
rect 15770 3754 15826 3788
rect 15860 3754 15916 3788
rect 15950 3754 16004 3788
rect 15324 3698 16004 3754
rect 15324 3664 15376 3698
rect 15410 3664 15466 3698
rect 15500 3664 15556 3698
rect 15590 3664 15646 3698
rect 15680 3664 15736 3698
rect 15770 3664 15826 3698
rect 15860 3664 15916 3698
rect 15950 3664 16004 3698
rect 15324 3608 16004 3664
rect 15324 3574 15376 3608
rect 15410 3574 15466 3608
rect 15500 3574 15556 3608
rect 15590 3574 15646 3608
rect 15680 3574 15736 3608
rect 15770 3574 15826 3608
rect 15860 3574 15916 3608
rect 15950 3574 16004 3608
rect 15324 3522 16004 3574
rect 16612 4148 17292 4202
rect 16612 4114 16664 4148
rect 16698 4114 16754 4148
rect 16788 4114 16844 4148
rect 16878 4114 16934 4148
rect 16968 4114 17024 4148
rect 17058 4114 17114 4148
rect 17148 4114 17204 4148
rect 17238 4114 17292 4148
rect 16612 4058 17292 4114
rect 16612 4024 16664 4058
rect 16698 4024 16754 4058
rect 16788 4024 16844 4058
rect 16878 4024 16934 4058
rect 16968 4024 17024 4058
rect 17058 4024 17114 4058
rect 17148 4024 17204 4058
rect 17238 4024 17292 4058
rect 16612 3968 17292 4024
rect 16612 3934 16664 3968
rect 16698 3934 16754 3968
rect 16788 3934 16844 3968
rect 16878 3934 16934 3968
rect 16968 3934 17024 3968
rect 17058 3934 17114 3968
rect 17148 3934 17204 3968
rect 17238 3934 17292 3968
rect 16612 3878 17292 3934
rect 16612 3844 16664 3878
rect 16698 3844 16754 3878
rect 16788 3844 16844 3878
rect 16878 3844 16934 3878
rect 16968 3844 17024 3878
rect 17058 3844 17114 3878
rect 17148 3844 17204 3878
rect 17238 3844 17292 3878
rect 16612 3788 17292 3844
rect 16612 3754 16664 3788
rect 16698 3754 16754 3788
rect 16788 3754 16844 3788
rect 16878 3754 16934 3788
rect 16968 3754 17024 3788
rect 17058 3754 17114 3788
rect 17148 3754 17204 3788
rect 17238 3754 17292 3788
rect 16612 3698 17292 3754
rect 16612 3664 16664 3698
rect 16698 3664 16754 3698
rect 16788 3664 16844 3698
rect 16878 3664 16934 3698
rect 16968 3664 17024 3698
rect 17058 3664 17114 3698
rect 17148 3664 17204 3698
rect 17238 3664 17292 3698
rect 16612 3608 17292 3664
rect 16612 3574 16664 3608
rect 16698 3574 16754 3608
rect 16788 3574 16844 3608
rect 16878 3574 16934 3608
rect 16968 3574 17024 3608
rect 17058 3574 17114 3608
rect 17148 3574 17204 3608
rect 17238 3574 17292 3608
rect 16612 3522 17292 3574
rect 17900 4148 18580 4202
rect 17900 4114 17952 4148
rect 17986 4114 18042 4148
rect 18076 4114 18132 4148
rect 18166 4114 18222 4148
rect 18256 4114 18312 4148
rect 18346 4114 18402 4148
rect 18436 4114 18492 4148
rect 18526 4114 18580 4148
rect 17900 4058 18580 4114
rect 17900 4024 17952 4058
rect 17986 4024 18042 4058
rect 18076 4024 18132 4058
rect 18166 4024 18222 4058
rect 18256 4024 18312 4058
rect 18346 4024 18402 4058
rect 18436 4024 18492 4058
rect 18526 4024 18580 4058
rect 17900 3968 18580 4024
rect 17900 3934 17952 3968
rect 17986 3934 18042 3968
rect 18076 3934 18132 3968
rect 18166 3934 18222 3968
rect 18256 3934 18312 3968
rect 18346 3934 18402 3968
rect 18436 3934 18492 3968
rect 18526 3934 18580 3968
rect 17900 3878 18580 3934
rect 17900 3844 17952 3878
rect 17986 3844 18042 3878
rect 18076 3844 18132 3878
rect 18166 3844 18222 3878
rect 18256 3844 18312 3878
rect 18346 3844 18402 3878
rect 18436 3844 18492 3878
rect 18526 3844 18580 3878
rect 17900 3788 18580 3844
rect 17900 3754 17952 3788
rect 17986 3754 18042 3788
rect 18076 3754 18132 3788
rect 18166 3754 18222 3788
rect 18256 3754 18312 3788
rect 18346 3754 18402 3788
rect 18436 3754 18492 3788
rect 18526 3754 18580 3788
rect 17900 3698 18580 3754
rect 17900 3664 17952 3698
rect 17986 3664 18042 3698
rect 18076 3664 18132 3698
rect 18166 3664 18222 3698
rect 18256 3664 18312 3698
rect 18346 3664 18402 3698
rect 18436 3664 18492 3698
rect 18526 3664 18580 3698
rect 17900 3608 18580 3664
rect 17900 3574 17952 3608
rect 17986 3574 18042 3608
rect 18076 3574 18132 3608
rect 18166 3574 18222 3608
rect 18256 3574 18312 3608
rect 18346 3574 18402 3608
rect 18436 3574 18492 3608
rect 18526 3574 18580 3608
rect 17900 3522 18580 3574
rect 12748 2860 13428 2914
rect 12748 2826 12800 2860
rect 12834 2826 12890 2860
rect 12924 2826 12980 2860
rect 13014 2826 13070 2860
rect 13104 2826 13160 2860
rect 13194 2826 13250 2860
rect 13284 2826 13340 2860
rect 13374 2826 13428 2860
rect 12748 2770 13428 2826
rect 12748 2736 12800 2770
rect 12834 2736 12890 2770
rect 12924 2736 12980 2770
rect 13014 2736 13070 2770
rect 13104 2736 13160 2770
rect 13194 2736 13250 2770
rect 13284 2736 13340 2770
rect 13374 2736 13428 2770
rect 12748 2680 13428 2736
rect 12748 2646 12800 2680
rect 12834 2646 12890 2680
rect 12924 2646 12980 2680
rect 13014 2646 13070 2680
rect 13104 2646 13160 2680
rect 13194 2646 13250 2680
rect 13284 2646 13340 2680
rect 13374 2646 13428 2680
rect 12748 2590 13428 2646
rect 12748 2556 12800 2590
rect 12834 2556 12890 2590
rect 12924 2556 12980 2590
rect 13014 2556 13070 2590
rect 13104 2556 13160 2590
rect 13194 2556 13250 2590
rect 13284 2556 13340 2590
rect 13374 2556 13428 2590
rect 12748 2500 13428 2556
rect 12748 2466 12800 2500
rect 12834 2466 12890 2500
rect 12924 2466 12980 2500
rect 13014 2466 13070 2500
rect 13104 2466 13160 2500
rect 13194 2466 13250 2500
rect 13284 2466 13340 2500
rect 13374 2466 13428 2500
rect 12748 2410 13428 2466
rect 12748 2376 12800 2410
rect 12834 2376 12890 2410
rect 12924 2376 12980 2410
rect 13014 2376 13070 2410
rect 13104 2376 13160 2410
rect 13194 2376 13250 2410
rect 13284 2376 13340 2410
rect 13374 2376 13428 2410
rect 12748 2320 13428 2376
rect 12748 2286 12800 2320
rect 12834 2286 12890 2320
rect 12924 2286 12980 2320
rect 13014 2286 13070 2320
rect 13104 2286 13160 2320
rect 13194 2286 13250 2320
rect 13284 2286 13340 2320
rect 13374 2286 13428 2320
rect 12748 2234 13428 2286
rect 14036 2860 14716 2914
rect 14036 2826 14088 2860
rect 14122 2826 14178 2860
rect 14212 2826 14268 2860
rect 14302 2826 14358 2860
rect 14392 2826 14448 2860
rect 14482 2826 14538 2860
rect 14572 2826 14628 2860
rect 14662 2826 14716 2860
rect 14036 2770 14716 2826
rect 14036 2736 14088 2770
rect 14122 2736 14178 2770
rect 14212 2736 14268 2770
rect 14302 2736 14358 2770
rect 14392 2736 14448 2770
rect 14482 2736 14538 2770
rect 14572 2736 14628 2770
rect 14662 2736 14716 2770
rect 14036 2680 14716 2736
rect 14036 2646 14088 2680
rect 14122 2646 14178 2680
rect 14212 2646 14268 2680
rect 14302 2646 14358 2680
rect 14392 2646 14448 2680
rect 14482 2646 14538 2680
rect 14572 2646 14628 2680
rect 14662 2646 14716 2680
rect 14036 2590 14716 2646
rect 14036 2556 14088 2590
rect 14122 2556 14178 2590
rect 14212 2556 14268 2590
rect 14302 2556 14358 2590
rect 14392 2556 14448 2590
rect 14482 2556 14538 2590
rect 14572 2556 14628 2590
rect 14662 2556 14716 2590
rect 14036 2500 14716 2556
rect 14036 2466 14088 2500
rect 14122 2466 14178 2500
rect 14212 2466 14268 2500
rect 14302 2466 14358 2500
rect 14392 2466 14448 2500
rect 14482 2466 14538 2500
rect 14572 2466 14628 2500
rect 14662 2466 14716 2500
rect 14036 2410 14716 2466
rect 14036 2376 14088 2410
rect 14122 2376 14178 2410
rect 14212 2376 14268 2410
rect 14302 2376 14358 2410
rect 14392 2376 14448 2410
rect 14482 2376 14538 2410
rect 14572 2376 14628 2410
rect 14662 2376 14716 2410
rect 14036 2320 14716 2376
rect 14036 2286 14088 2320
rect 14122 2286 14178 2320
rect 14212 2286 14268 2320
rect 14302 2286 14358 2320
rect 14392 2286 14448 2320
rect 14482 2286 14538 2320
rect 14572 2286 14628 2320
rect 14662 2286 14716 2320
rect 14036 2234 14716 2286
rect 15324 2860 16004 2914
rect 15324 2826 15376 2860
rect 15410 2826 15466 2860
rect 15500 2826 15556 2860
rect 15590 2826 15646 2860
rect 15680 2826 15736 2860
rect 15770 2826 15826 2860
rect 15860 2826 15916 2860
rect 15950 2826 16004 2860
rect 15324 2770 16004 2826
rect 15324 2736 15376 2770
rect 15410 2736 15466 2770
rect 15500 2736 15556 2770
rect 15590 2736 15646 2770
rect 15680 2736 15736 2770
rect 15770 2736 15826 2770
rect 15860 2736 15916 2770
rect 15950 2736 16004 2770
rect 15324 2680 16004 2736
rect 15324 2646 15376 2680
rect 15410 2646 15466 2680
rect 15500 2646 15556 2680
rect 15590 2646 15646 2680
rect 15680 2646 15736 2680
rect 15770 2646 15826 2680
rect 15860 2646 15916 2680
rect 15950 2646 16004 2680
rect 15324 2590 16004 2646
rect 15324 2556 15376 2590
rect 15410 2556 15466 2590
rect 15500 2556 15556 2590
rect 15590 2556 15646 2590
rect 15680 2556 15736 2590
rect 15770 2556 15826 2590
rect 15860 2556 15916 2590
rect 15950 2556 16004 2590
rect 15324 2500 16004 2556
rect 15324 2466 15376 2500
rect 15410 2466 15466 2500
rect 15500 2466 15556 2500
rect 15590 2466 15646 2500
rect 15680 2466 15736 2500
rect 15770 2466 15826 2500
rect 15860 2466 15916 2500
rect 15950 2466 16004 2500
rect 15324 2410 16004 2466
rect 15324 2376 15376 2410
rect 15410 2376 15466 2410
rect 15500 2376 15556 2410
rect 15590 2376 15646 2410
rect 15680 2376 15736 2410
rect 15770 2376 15826 2410
rect 15860 2376 15916 2410
rect 15950 2376 16004 2410
rect 15324 2320 16004 2376
rect 15324 2286 15376 2320
rect 15410 2286 15466 2320
rect 15500 2286 15556 2320
rect 15590 2286 15646 2320
rect 15680 2286 15736 2320
rect 15770 2286 15826 2320
rect 15860 2286 15916 2320
rect 15950 2286 16004 2320
rect 15324 2234 16004 2286
rect 16612 2860 17292 2914
rect 16612 2826 16664 2860
rect 16698 2826 16754 2860
rect 16788 2826 16844 2860
rect 16878 2826 16934 2860
rect 16968 2826 17024 2860
rect 17058 2826 17114 2860
rect 17148 2826 17204 2860
rect 17238 2826 17292 2860
rect 16612 2770 17292 2826
rect 16612 2736 16664 2770
rect 16698 2736 16754 2770
rect 16788 2736 16844 2770
rect 16878 2736 16934 2770
rect 16968 2736 17024 2770
rect 17058 2736 17114 2770
rect 17148 2736 17204 2770
rect 17238 2736 17292 2770
rect 16612 2680 17292 2736
rect 16612 2646 16664 2680
rect 16698 2646 16754 2680
rect 16788 2646 16844 2680
rect 16878 2646 16934 2680
rect 16968 2646 17024 2680
rect 17058 2646 17114 2680
rect 17148 2646 17204 2680
rect 17238 2646 17292 2680
rect 16612 2590 17292 2646
rect 16612 2556 16664 2590
rect 16698 2556 16754 2590
rect 16788 2556 16844 2590
rect 16878 2556 16934 2590
rect 16968 2556 17024 2590
rect 17058 2556 17114 2590
rect 17148 2556 17204 2590
rect 17238 2556 17292 2590
rect 16612 2500 17292 2556
rect 16612 2466 16664 2500
rect 16698 2466 16754 2500
rect 16788 2466 16844 2500
rect 16878 2466 16934 2500
rect 16968 2466 17024 2500
rect 17058 2466 17114 2500
rect 17148 2466 17204 2500
rect 17238 2466 17292 2500
rect 16612 2410 17292 2466
rect 16612 2376 16664 2410
rect 16698 2376 16754 2410
rect 16788 2376 16844 2410
rect 16878 2376 16934 2410
rect 16968 2376 17024 2410
rect 17058 2376 17114 2410
rect 17148 2376 17204 2410
rect 17238 2376 17292 2410
rect 16612 2320 17292 2376
rect 16612 2286 16664 2320
rect 16698 2286 16754 2320
rect 16788 2286 16844 2320
rect 16878 2286 16934 2320
rect 16968 2286 17024 2320
rect 17058 2286 17114 2320
rect 17148 2286 17204 2320
rect 17238 2286 17292 2320
rect 16612 2234 17292 2286
rect 17900 2860 18580 2914
rect 17900 2826 17952 2860
rect 17986 2826 18042 2860
rect 18076 2826 18132 2860
rect 18166 2826 18222 2860
rect 18256 2826 18312 2860
rect 18346 2826 18402 2860
rect 18436 2826 18492 2860
rect 18526 2826 18580 2860
rect 17900 2770 18580 2826
rect 17900 2736 17952 2770
rect 17986 2736 18042 2770
rect 18076 2736 18132 2770
rect 18166 2736 18222 2770
rect 18256 2736 18312 2770
rect 18346 2736 18402 2770
rect 18436 2736 18492 2770
rect 18526 2736 18580 2770
rect 17900 2680 18580 2736
rect 17900 2646 17952 2680
rect 17986 2646 18042 2680
rect 18076 2646 18132 2680
rect 18166 2646 18222 2680
rect 18256 2646 18312 2680
rect 18346 2646 18402 2680
rect 18436 2646 18492 2680
rect 18526 2646 18580 2680
rect 17900 2590 18580 2646
rect 17900 2556 17952 2590
rect 17986 2556 18042 2590
rect 18076 2556 18132 2590
rect 18166 2556 18222 2590
rect 18256 2556 18312 2590
rect 18346 2556 18402 2590
rect 18436 2556 18492 2590
rect 18526 2556 18580 2590
rect 17900 2500 18580 2556
rect 17900 2466 17952 2500
rect 17986 2466 18042 2500
rect 18076 2466 18132 2500
rect 18166 2466 18222 2500
rect 18256 2466 18312 2500
rect 18346 2466 18402 2500
rect 18436 2466 18492 2500
rect 18526 2466 18580 2500
rect 17900 2410 18580 2466
rect 17900 2376 17952 2410
rect 17986 2376 18042 2410
rect 18076 2376 18132 2410
rect 18166 2376 18222 2410
rect 18256 2376 18312 2410
rect 18346 2376 18402 2410
rect 18436 2376 18492 2410
rect 18526 2376 18580 2410
rect 17900 2320 18580 2376
rect 17900 2286 17952 2320
rect 17986 2286 18042 2320
rect 18076 2286 18132 2320
rect 18166 2286 18222 2320
rect 18256 2286 18312 2320
rect 18346 2286 18402 2320
rect 18436 2286 18492 2320
rect 18526 2286 18580 2320
rect 17900 2234 18580 2286
rect 7684 1700 7742 1712
rect -10726 1662 -10668 1674
<< ndiffc >>
rect -17164 8818 -11788 8852
rect -17164 8360 -11788 8394
rect -21812 5144 -21778 5520
rect -21354 5144 -21320 5520
rect -20896 5144 -20862 5520
rect -20438 5144 -20404 5520
rect -19980 5144 -19946 5520
rect -19522 5144 -19488 5520
rect -19064 5144 -19030 5520
rect -16882 4866 -16848 6642
rect -16424 4866 -16390 6642
rect -16310 4866 -16276 6642
rect -15852 4866 -15818 6642
rect -15738 4866 -15704 6642
rect -15280 4866 -15246 6642
rect -15166 4866 -15132 6642
rect -14708 4866 -14674 6642
rect -14594 4866 -14560 6642
rect -14136 4866 -14102 6642
rect -14022 4866 -13988 6642
rect -13564 4866 -13530 6642
rect -13450 4866 -13416 6642
rect -12992 4866 -12958 6642
rect -12878 4866 -12844 6642
rect -12420 4866 -12386 6642
<< pdiffc >>
rect 12800 11842 12834 11876
rect 12890 11842 12924 11876
rect 12980 11842 13014 11876
rect 13070 11842 13104 11876
rect 13160 11842 13194 11876
rect 13250 11842 13284 11876
rect 13340 11842 13374 11876
rect 12800 11752 12834 11786
rect 12890 11752 12924 11786
rect 12980 11752 13014 11786
rect 13070 11752 13104 11786
rect 13160 11752 13194 11786
rect 13250 11752 13284 11786
rect 13340 11752 13374 11786
rect 12800 11662 12834 11696
rect 12890 11662 12924 11696
rect 12980 11662 13014 11696
rect 13070 11662 13104 11696
rect 13160 11662 13194 11696
rect 13250 11662 13284 11696
rect 13340 11662 13374 11696
rect 12800 11572 12834 11606
rect 12890 11572 12924 11606
rect 12980 11572 13014 11606
rect 13070 11572 13104 11606
rect 13160 11572 13194 11606
rect 13250 11572 13284 11606
rect 13340 11572 13374 11606
rect 12800 11482 12834 11516
rect 12890 11482 12924 11516
rect 12980 11482 13014 11516
rect 13070 11482 13104 11516
rect 13160 11482 13194 11516
rect 13250 11482 13284 11516
rect 13340 11482 13374 11516
rect 12800 11392 12834 11426
rect 12890 11392 12924 11426
rect 12980 11392 13014 11426
rect 13070 11392 13104 11426
rect 13160 11392 13194 11426
rect 13250 11392 13284 11426
rect 13340 11392 13374 11426
rect 12800 11302 12834 11336
rect 12890 11302 12924 11336
rect 12980 11302 13014 11336
rect 13070 11302 13104 11336
rect 13160 11302 13194 11336
rect 13250 11302 13284 11336
rect 13340 11302 13374 11336
rect 14088 11842 14122 11876
rect 14178 11842 14212 11876
rect 14268 11842 14302 11876
rect 14358 11842 14392 11876
rect 14448 11842 14482 11876
rect 14538 11842 14572 11876
rect 14628 11842 14662 11876
rect 14088 11752 14122 11786
rect 14178 11752 14212 11786
rect 14268 11752 14302 11786
rect 14358 11752 14392 11786
rect 14448 11752 14482 11786
rect 14538 11752 14572 11786
rect 14628 11752 14662 11786
rect 14088 11662 14122 11696
rect 14178 11662 14212 11696
rect 14268 11662 14302 11696
rect 14358 11662 14392 11696
rect 14448 11662 14482 11696
rect 14538 11662 14572 11696
rect 14628 11662 14662 11696
rect 14088 11572 14122 11606
rect 14178 11572 14212 11606
rect 14268 11572 14302 11606
rect 14358 11572 14392 11606
rect 14448 11572 14482 11606
rect 14538 11572 14572 11606
rect 14628 11572 14662 11606
rect 14088 11482 14122 11516
rect 14178 11482 14212 11516
rect 14268 11482 14302 11516
rect 14358 11482 14392 11516
rect 14448 11482 14482 11516
rect 14538 11482 14572 11516
rect 14628 11482 14662 11516
rect 14088 11392 14122 11426
rect 14178 11392 14212 11426
rect 14268 11392 14302 11426
rect 14358 11392 14392 11426
rect 14448 11392 14482 11426
rect 14538 11392 14572 11426
rect 14628 11392 14662 11426
rect 14088 11302 14122 11336
rect 14178 11302 14212 11336
rect 14268 11302 14302 11336
rect 14358 11302 14392 11336
rect 14448 11302 14482 11336
rect 14538 11302 14572 11336
rect 14628 11302 14662 11336
rect 15376 11842 15410 11876
rect 15466 11842 15500 11876
rect 15556 11842 15590 11876
rect 15646 11842 15680 11876
rect 15736 11842 15770 11876
rect 15826 11842 15860 11876
rect 15916 11842 15950 11876
rect 15376 11752 15410 11786
rect 15466 11752 15500 11786
rect 15556 11752 15590 11786
rect 15646 11752 15680 11786
rect 15736 11752 15770 11786
rect 15826 11752 15860 11786
rect 15916 11752 15950 11786
rect 15376 11662 15410 11696
rect 15466 11662 15500 11696
rect 15556 11662 15590 11696
rect 15646 11662 15680 11696
rect 15736 11662 15770 11696
rect 15826 11662 15860 11696
rect 15916 11662 15950 11696
rect 15376 11572 15410 11606
rect 15466 11572 15500 11606
rect 15556 11572 15590 11606
rect 15646 11572 15680 11606
rect 15736 11572 15770 11606
rect 15826 11572 15860 11606
rect 15916 11572 15950 11606
rect 15376 11482 15410 11516
rect 15466 11482 15500 11516
rect 15556 11482 15590 11516
rect 15646 11482 15680 11516
rect 15736 11482 15770 11516
rect 15826 11482 15860 11516
rect 15916 11482 15950 11516
rect 15376 11392 15410 11426
rect 15466 11392 15500 11426
rect 15556 11392 15590 11426
rect 15646 11392 15680 11426
rect 15736 11392 15770 11426
rect 15826 11392 15860 11426
rect 15916 11392 15950 11426
rect 15376 11302 15410 11336
rect 15466 11302 15500 11336
rect 15556 11302 15590 11336
rect 15646 11302 15680 11336
rect 15736 11302 15770 11336
rect 15826 11302 15860 11336
rect 15916 11302 15950 11336
rect 16664 11842 16698 11876
rect 16754 11842 16788 11876
rect 16844 11842 16878 11876
rect 16934 11842 16968 11876
rect 17024 11842 17058 11876
rect 17114 11842 17148 11876
rect 17204 11842 17238 11876
rect 16664 11752 16698 11786
rect 16754 11752 16788 11786
rect 16844 11752 16878 11786
rect 16934 11752 16968 11786
rect 17024 11752 17058 11786
rect 17114 11752 17148 11786
rect 17204 11752 17238 11786
rect 16664 11662 16698 11696
rect 16754 11662 16788 11696
rect 16844 11662 16878 11696
rect 16934 11662 16968 11696
rect 17024 11662 17058 11696
rect 17114 11662 17148 11696
rect 17204 11662 17238 11696
rect 16664 11572 16698 11606
rect 16754 11572 16788 11606
rect 16844 11572 16878 11606
rect 16934 11572 16968 11606
rect 17024 11572 17058 11606
rect 17114 11572 17148 11606
rect 17204 11572 17238 11606
rect 16664 11482 16698 11516
rect 16754 11482 16788 11516
rect 16844 11482 16878 11516
rect 16934 11482 16968 11516
rect 17024 11482 17058 11516
rect 17114 11482 17148 11516
rect 17204 11482 17238 11516
rect 16664 11392 16698 11426
rect 16754 11392 16788 11426
rect 16844 11392 16878 11426
rect 16934 11392 16968 11426
rect 17024 11392 17058 11426
rect 17114 11392 17148 11426
rect 17204 11392 17238 11426
rect 16664 11302 16698 11336
rect 16754 11302 16788 11336
rect 16844 11302 16878 11336
rect 16934 11302 16968 11336
rect 17024 11302 17058 11336
rect 17114 11302 17148 11336
rect 17204 11302 17238 11336
rect 17952 11842 17986 11876
rect 18042 11842 18076 11876
rect 18132 11842 18166 11876
rect 18222 11842 18256 11876
rect 18312 11842 18346 11876
rect 18402 11842 18436 11876
rect 18492 11842 18526 11876
rect 17952 11752 17986 11786
rect 18042 11752 18076 11786
rect 18132 11752 18166 11786
rect 18222 11752 18256 11786
rect 18312 11752 18346 11786
rect 18402 11752 18436 11786
rect 18492 11752 18526 11786
rect 17952 11662 17986 11696
rect 18042 11662 18076 11696
rect 18132 11662 18166 11696
rect 18222 11662 18256 11696
rect 18312 11662 18346 11696
rect 18402 11662 18436 11696
rect 18492 11662 18526 11696
rect 17952 11572 17986 11606
rect 18042 11572 18076 11606
rect 18132 11572 18166 11606
rect 18222 11572 18256 11606
rect 18312 11572 18346 11606
rect 18402 11572 18436 11606
rect 18492 11572 18526 11606
rect 17952 11482 17986 11516
rect 18042 11482 18076 11516
rect 18132 11482 18166 11516
rect 18222 11482 18256 11516
rect 18312 11482 18346 11516
rect 18402 11482 18436 11516
rect 18492 11482 18526 11516
rect 17952 11392 17986 11426
rect 18042 11392 18076 11426
rect 18132 11392 18166 11426
rect 18222 11392 18256 11426
rect 18312 11392 18346 11426
rect 18402 11392 18436 11426
rect 18492 11392 18526 11426
rect 17952 11302 17986 11336
rect 18042 11302 18076 11336
rect 18132 11302 18166 11336
rect 18222 11302 18256 11336
rect 18312 11302 18346 11336
rect 18402 11302 18436 11336
rect 18492 11302 18526 11336
rect 12800 10554 12834 10588
rect 12890 10554 12924 10588
rect 12980 10554 13014 10588
rect 13070 10554 13104 10588
rect 13160 10554 13194 10588
rect 13250 10554 13284 10588
rect 13340 10554 13374 10588
rect 12800 10464 12834 10498
rect 12890 10464 12924 10498
rect 12980 10464 13014 10498
rect 13070 10464 13104 10498
rect 13160 10464 13194 10498
rect 13250 10464 13284 10498
rect 13340 10464 13374 10498
rect 12800 10374 12834 10408
rect 12890 10374 12924 10408
rect 12980 10374 13014 10408
rect 13070 10374 13104 10408
rect 13160 10374 13194 10408
rect 13250 10374 13284 10408
rect 13340 10374 13374 10408
rect 12800 10284 12834 10318
rect 12890 10284 12924 10318
rect 12980 10284 13014 10318
rect 13070 10284 13104 10318
rect 13160 10284 13194 10318
rect 13250 10284 13284 10318
rect 13340 10284 13374 10318
rect 12800 10194 12834 10228
rect 12890 10194 12924 10228
rect 12980 10194 13014 10228
rect 13070 10194 13104 10228
rect 13160 10194 13194 10228
rect 13250 10194 13284 10228
rect 13340 10194 13374 10228
rect 12800 10104 12834 10138
rect 12890 10104 12924 10138
rect 12980 10104 13014 10138
rect 13070 10104 13104 10138
rect 13160 10104 13194 10138
rect 13250 10104 13284 10138
rect 13340 10104 13374 10138
rect 12800 10014 12834 10048
rect 12890 10014 12924 10048
rect 12980 10014 13014 10048
rect 13070 10014 13104 10048
rect 13160 10014 13194 10048
rect 13250 10014 13284 10048
rect 13340 10014 13374 10048
rect 14088 10554 14122 10588
rect 14178 10554 14212 10588
rect 14268 10554 14302 10588
rect 14358 10554 14392 10588
rect 14448 10554 14482 10588
rect 14538 10554 14572 10588
rect 14628 10554 14662 10588
rect 14088 10464 14122 10498
rect 14178 10464 14212 10498
rect 14268 10464 14302 10498
rect 14358 10464 14392 10498
rect 14448 10464 14482 10498
rect 14538 10464 14572 10498
rect 14628 10464 14662 10498
rect 14088 10374 14122 10408
rect 14178 10374 14212 10408
rect 14268 10374 14302 10408
rect 14358 10374 14392 10408
rect 14448 10374 14482 10408
rect 14538 10374 14572 10408
rect 14628 10374 14662 10408
rect 14088 10284 14122 10318
rect 14178 10284 14212 10318
rect 14268 10284 14302 10318
rect 14358 10284 14392 10318
rect 14448 10284 14482 10318
rect 14538 10284 14572 10318
rect 14628 10284 14662 10318
rect 14088 10194 14122 10228
rect 14178 10194 14212 10228
rect 14268 10194 14302 10228
rect 14358 10194 14392 10228
rect 14448 10194 14482 10228
rect 14538 10194 14572 10228
rect 14628 10194 14662 10228
rect 14088 10104 14122 10138
rect 14178 10104 14212 10138
rect 14268 10104 14302 10138
rect 14358 10104 14392 10138
rect 14448 10104 14482 10138
rect 14538 10104 14572 10138
rect 14628 10104 14662 10138
rect 14088 10014 14122 10048
rect 14178 10014 14212 10048
rect 14268 10014 14302 10048
rect 14358 10014 14392 10048
rect 14448 10014 14482 10048
rect 14538 10014 14572 10048
rect 14628 10014 14662 10048
rect 15376 10554 15410 10588
rect 15466 10554 15500 10588
rect 15556 10554 15590 10588
rect 15646 10554 15680 10588
rect 15736 10554 15770 10588
rect 15826 10554 15860 10588
rect 15916 10554 15950 10588
rect 15376 10464 15410 10498
rect 15466 10464 15500 10498
rect 15556 10464 15590 10498
rect 15646 10464 15680 10498
rect 15736 10464 15770 10498
rect 15826 10464 15860 10498
rect 15916 10464 15950 10498
rect 15376 10374 15410 10408
rect 15466 10374 15500 10408
rect 15556 10374 15590 10408
rect 15646 10374 15680 10408
rect 15736 10374 15770 10408
rect 15826 10374 15860 10408
rect 15916 10374 15950 10408
rect 15376 10284 15410 10318
rect 15466 10284 15500 10318
rect 15556 10284 15590 10318
rect 15646 10284 15680 10318
rect 15736 10284 15770 10318
rect 15826 10284 15860 10318
rect 15916 10284 15950 10318
rect 15376 10194 15410 10228
rect 15466 10194 15500 10228
rect 15556 10194 15590 10228
rect 15646 10194 15680 10228
rect 15736 10194 15770 10228
rect 15826 10194 15860 10228
rect 15916 10194 15950 10228
rect 15376 10104 15410 10138
rect 15466 10104 15500 10138
rect 15556 10104 15590 10138
rect 15646 10104 15680 10138
rect 15736 10104 15770 10138
rect 15826 10104 15860 10138
rect 15916 10104 15950 10138
rect 15376 10014 15410 10048
rect 15466 10014 15500 10048
rect 15556 10014 15590 10048
rect 15646 10014 15680 10048
rect 15736 10014 15770 10048
rect 15826 10014 15860 10048
rect 15916 10014 15950 10048
rect 16664 10554 16698 10588
rect 16754 10554 16788 10588
rect 16844 10554 16878 10588
rect 16934 10554 16968 10588
rect 17024 10554 17058 10588
rect 17114 10554 17148 10588
rect 17204 10554 17238 10588
rect 16664 10464 16698 10498
rect 16754 10464 16788 10498
rect 16844 10464 16878 10498
rect 16934 10464 16968 10498
rect 17024 10464 17058 10498
rect 17114 10464 17148 10498
rect 17204 10464 17238 10498
rect 16664 10374 16698 10408
rect 16754 10374 16788 10408
rect 16844 10374 16878 10408
rect 16934 10374 16968 10408
rect 17024 10374 17058 10408
rect 17114 10374 17148 10408
rect 17204 10374 17238 10408
rect 16664 10284 16698 10318
rect 16754 10284 16788 10318
rect 16844 10284 16878 10318
rect 16934 10284 16968 10318
rect 17024 10284 17058 10318
rect 17114 10284 17148 10318
rect 17204 10284 17238 10318
rect 16664 10194 16698 10228
rect 16754 10194 16788 10228
rect 16844 10194 16878 10228
rect 16934 10194 16968 10228
rect 17024 10194 17058 10228
rect 17114 10194 17148 10228
rect 17204 10194 17238 10228
rect 16664 10104 16698 10138
rect 16754 10104 16788 10138
rect 16844 10104 16878 10138
rect 16934 10104 16968 10138
rect 17024 10104 17058 10138
rect 17114 10104 17148 10138
rect 17204 10104 17238 10138
rect 16664 10014 16698 10048
rect 16754 10014 16788 10048
rect 16844 10014 16878 10048
rect 16934 10014 16968 10048
rect 17024 10014 17058 10048
rect 17114 10014 17148 10048
rect 17204 10014 17238 10048
rect 17952 10554 17986 10588
rect 18042 10554 18076 10588
rect 18132 10554 18166 10588
rect 18222 10554 18256 10588
rect 18312 10554 18346 10588
rect 18402 10554 18436 10588
rect 18492 10554 18526 10588
rect 17952 10464 17986 10498
rect 18042 10464 18076 10498
rect 18132 10464 18166 10498
rect 18222 10464 18256 10498
rect 18312 10464 18346 10498
rect 18402 10464 18436 10498
rect 18492 10464 18526 10498
rect 17952 10374 17986 10408
rect 18042 10374 18076 10408
rect 18132 10374 18166 10408
rect 18222 10374 18256 10408
rect 18312 10374 18346 10408
rect 18402 10374 18436 10408
rect 18492 10374 18526 10408
rect 17952 10284 17986 10318
rect 18042 10284 18076 10318
rect 18132 10284 18166 10318
rect 18222 10284 18256 10318
rect 18312 10284 18346 10318
rect 18402 10284 18436 10318
rect 18492 10284 18526 10318
rect 17952 10194 17986 10228
rect 18042 10194 18076 10228
rect 18132 10194 18166 10228
rect 18222 10194 18256 10228
rect 18312 10194 18346 10228
rect 18402 10194 18436 10228
rect 18492 10194 18526 10228
rect 17952 10104 17986 10138
rect 18042 10104 18076 10138
rect 18132 10104 18166 10138
rect 18222 10104 18256 10138
rect 18312 10104 18346 10138
rect 18402 10104 18436 10138
rect 18492 10104 18526 10138
rect 17952 10014 17986 10048
rect 18042 10014 18076 10048
rect 18132 10014 18166 10048
rect 18222 10014 18256 10048
rect 18312 10014 18346 10048
rect 18402 10014 18436 10048
rect 18492 10014 18526 10048
rect -18608 1674 -18574 4230
rect -18150 1674 -18116 4230
rect -18036 1674 -18002 4230
rect -17578 1674 -17544 4230
rect -17464 1674 -17430 4230
rect -17006 1674 -16972 4230
rect -16892 1674 -16858 4230
rect -16434 1674 -16400 4230
rect -16320 1674 -16286 4230
rect -15862 1674 -15828 4230
rect -15748 1674 -15714 4230
rect -15290 1674 -15256 4230
rect -15176 1674 -15142 4230
rect -14718 1674 -14684 4230
rect -14604 1674 -14570 4230
rect -14146 1674 -14112 4230
rect -14032 1674 -13998 4230
rect -13574 1674 -13540 4230
rect -13460 1674 -13426 4230
rect -13002 1674 -12968 4230
rect -12888 1674 -12854 4230
rect -12430 1674 -12396 4230
rect -12316 1674 -12282 4230
rect -11858 1674 -11824 4230
rect -11744 1674 -11710 4230
rect -11286 1674 -11252 4230
rect -11172 1674 -11138 4230
rect -10714 1674 -10680 4230
rect -8800 1712 -8766 9428
rect -8342 1712 -8308 9428
rect -7884 1712 -7850 9428
rect -7426 1712 -7392 9428
rect -6968 1712 -6934 9428
rect -6510 1712 -6476 9428
rect -6052 1712 -6018 9428
rect -5594 1712 -5560 9428
rect -5136 1712 -5102 9428
rect -4678 1712 -4644 9428
rect -4220 1712 -4186 9428
rect -3762 1712 -3728 9428
rect -2842 1712 -2808 9428
rect -2384 1712 -2350 9428
rect -1926 1712 -1892 9428
rect -1468 1712 -1434 9428
rect -1010 1712 -976 9428
rect -552 1712 -518 9428
rect -94 1712 -60 9428
rect 364 1712 398 9428
rect 822 1712 856 9428
rect 1280 1712 1314 9428
rect 1738 1712 1772 9428
rect 2658 1712 2692 9428
rect 3116 1712 3150 9428
rect 3574 1712 3608 9428
rect 4032 1712 4066 9428
rect 4490 1712 4524 9428
rect 4948 1712 4982 9428
rect 5406 1712 5440 9428
rect 5864 1712 5898 9428
rect 6322 1712 6356 9428
rect 6780 1712 6814 9428
rect 7238 1712 7272 9428
rect 7696 1712 7730 9428
rect 12800 9266 12834 9300
rect 12890 9266 12924 9300
rect 12980 9266 13014 9300
rect 13070 9266 13104 9300
rect 13160 9266 13194 9300
rect 13250 9266 13284 9300
rect 13340 9266 13374 9300
rect 12800 9176 12834 9210
rect 12890 9176 12924 9210
rect 12980 9176 13014 9210
rect 13070 9176 13104 9210
rect 13160 9176 13194 9210
rect 13250 9176 13284 9210
rect 13340 9176 13374 9210
rect 12800 9086 12834 9120
rect 12890 9086 12924 9120
rect 12980 9086 13014 9120
rect 13070 9086 13104 9120
rect 13160 9086 13194 9120
rect 13250 9086 13284 9120
rect 13340 9086 13374 9120
rect 12800 8996 12834 9030
rect 12890 8996 12924 9030
rect 12980 8996 13014 9030
rect 13070 8996 13104 9030
rect 13160 8996 13194 9030
rect 13250 8996 13284 9030
rect 13340 8996 13374 9030
rect 12800 8906 12834 8940
rect 12890 8906 12924 8940
rect 12980 8906 13014 8940
rect 13070 8906 13104 8940
rect 13160 8906 13194 8940
rect 13250 8906 13284 8940
rect 13340 8906 13374 8940
rect 12800 8816 12834 8850
rect 12890 8816 12924 8850
rect 12980 8816 13014 8850
rect 13070 8816 13104 8850
rect 13160 8816 13194 8850
rect 13250 8816 13284 8850
rect 13340 8816 13374 8850
rect 12800 8726 12834 8760
rect 12890 8726 12924 8760
rect 12980 8726 13014 8760
rect 13070 8726 13104 8760
rect 13160 8726 13194 8760
rect 13250 8726 13284 8760
rect 13340 8726 13374 8760
rect 14088 9266 14122 9300
rect 14178 9266 14212 9300
rect 14268 9266 14302 9300
rect 14358 9266 14392 9300
rect 14448 9266 14482 9300
rect 14538 9266 14572 9300
rect 14628 9266 14662 9300
rect 14088 9176 14122 9210
rect 14178 9176 14212 9210
rect 14268 9176 14302 9210
rect 14358 9176 14392 9210
rect 14448 9176 14482 9210
rect 14538 9176 14572 9210
rect 14628 9176 14662 9210
rect 14088 9086 14122 9120
rect 14178 9086 14212 9120
rect 14268 9086 14302 9120
rect 14358 9086 14392 9120
rect 14448 9086 14482 9120
rect 14538 9086 14572 9120
rect 14628 9086 14662 9120
rect 14088 8996 14122 9030
rect 14178 8996 14212 9030
rect 14268 8996 14302 9030
rect 14358 8996 14392 9030
rect 14448 8996 14482 9030
rect 14538 8996 14572 9030
rect 14628 8996 14662 9030
rect 14088 8906 14122 8940
rect 14178 8906 14212 8940
rect 14268 8906 14302 8940
rect 14358 8906 14392 8940
rect 14448 8906 14482 8940
rect 14538 8906 14572 8940
rect 14628 8906 14662 8940
rect 14088 8816 14122 8850
rect 14178 8816 14212 8850
rect 14268 8816 14302 8850
rect 14358 8816 14392 8850
rect 14448 8816 14482 8850
rect 14538 8816 14572 8850
rect 14628 8816 14662 8850
rect 14088 8726 14122 8760
rect 14178 8726 14212 8760
rect 14268 8726 14302 8760
rect 14358 8726 14392 8760
rect 14448 8726 14482 8760
rect 14538 8726 14572 8760
rect 14628 8726 14662 8760
rect 15376 9266 15410 9300
rect 15466 9266 15500 9300
rect 15556 9266 15590 9300
rect 15646 9266 15680 9300
rect 15736 9266 15770 9300
rect 15826 9266 15860 9300
rect 15916 9266 15950 9300
rect 15376 9176 15410 9210
rect 15466 9176 15500 9210
rect 15556 9176 15590 9210
rect 15646 9176 15680 9210
rect 15736 9176 15770 9210
rect 15826 9176 15860 9210
rect 15916 9176 15950 9210
rect 15376 9086 15410 9120
rect 15466 9086 15500 9120
rect 15556 9086 15590 9120
rect 15646 9086 15680 9120
rect 15736 9086 15770 9120
rect 15826 9086 15860 9120
rect 15916 9086 15950 9120
rect 15376 8996 15410 9030
rect 15466 8996 15500 9030
rect 15556 8996 15590 9030
rect 15646 8996 15680 9030
rect 15736 8996 15770 9030
rect 15826 8996 15860 9030
rect 15916 8996 15950 9030
rect 15376 8906 15410 8940
rect 15466 8906 15500 8940
rect 15556 8906 15590 8940
rect 15646 8906 15680 8940
rect 15736 8906 15770 8940
rect 15826 8906 15860 8940
rect 15916 8906 15950 8940
rect 15376 8816 15410 8850
rect 15466 8816 15500 8850
rect 15556 8816 15590 8850
rect 15646 8816 15680 8850
rect 15736 8816 15770 8850
rect 15826 8816 15860 8850
rect 15916 8816 15950 8850
rect 15376 8726 15410 8760
rect 15466 8726 15500 8760
rect 15556 8726 15590 8760
rect 15646 8726 15680 8760
rect 15736 8726 15770 8760
rect 15826 8726 15860 8760
rect 15916 8726 15950 8760
rect 16664 9266 16698 9300
rect 16754 9266 16788 9300
rect 16844 9266 16878 9300
rect 16934 9266 16968 9300
rect 17024 9266 17058 9300
rect 17114 9266 17148 9300
rect 17204 9266 17238 9300
rect 16664 9176 16698 9210
rect 16754 9176 16788 9210
rect 16844 9176 16878 9210
rect 16934 9176 16968 9210
rect 17024 9176 17058 9210
rect 17114 9176 17148 9210
rect 17204 9176 17238 9210
rect 16664 9086 16698 9120
rect 16754 9086 16788 9120
rect 16844 9086 16878 9120
rect 16934 9086 16968 9120
rect 17024 9086 17058 9120
rect 17114 9086 17148 9120
rect 17204 9086 17238 9120
rect 16664 8996 16698 9030
rect 16754 8996 16788 9030
rect 16844 8996 16878 9030
rect 16934 8996 16968 9030
rect 17024 8996 17058 9030
rect 17114 8996 17148 9030
rect 17204 8996 17238 9030
rect 16664 8906 16698 8940
rect 16754 8906 16788 8940
rect 16844 8906 16878 8940
rect 16934 8906 16968 8940
rect 17024 8906 17058 8940
rect 17114 8906 17148 8940
rect 17204 8906 17238 8940
rect 16664 8816 16698 8850
rect 16754 8816 16788 8850
rect 16844 8816 16878 8850
rect 16934 8816 16968 8850
rect 17024 8816 17058 8850
rect 17114 8816 17148 8850
rect 17204 8816 17238 8850
rect 16664 8726 16698 8760
rect 16754 8726 16788 8760
rect 16844 8726 16878 8760
rect 16934 8726 16968 8760
rect 17024 8726 17058 8760
rect 17114 8726 17148 8760
rect 17204 8726 17238 8760
rect 17952 9266 17986 9300
rect 18042 9266 18076 9300
rect 18132 9266 18166 9300
rect 18222 9266 18256 9300
rect 18312 9266 18346 9300
rect 18402 9266 18436 9300
rect 18492 9266 18526 9300
rect 17952 9176 17986 9210
rect 18042 9176 18076 9210
rect 18132 9176 18166 9210
rect 18222 9176 18256 9210
rect 18312 9176 18346 9210
rect 18402 9176 18436 9210
rect 18492 9176 18526 9210
rect 17952 9086 17986 9120
rect 18042 9086 18076 9120
rect 18132 9086 18166 9120
rect 18222 9086 18256 9120
rect 18312 9086 18346 9120
rect 18402 9086 18436 9120
rect 18492 9086 18526 9120
rect 17952 8996 17986 9030
rect 18042 8996 18076 9030
rect 18132 8996 18166 9030
rect 18222 8996 18256 9030
rect 18312 8996 18346 9030
rect 18402 8996 18436 9030
rect 18492 8996 18526 9030
rect 17952 8906 17986 8940
rect 18042 8906 18076 8940
rect 18132 8906 18166 8940
rect 18222 8906 18256 8940
rect 18312 8906 18346 8940
rect 18402 8906 18436 8940
rect 18492 8906 18526 8940
rect 17952 8816 17986 8850
rect 18042 8816 18076 8850
rect 18132 8816 18166 8850
rect 18222 8816 18256 8850
rect 18312 8816 18346 8850
rect 18402 8816 18436 8850
rect 18492 8816 18526 8850
rect 17952 8726 17986 8760
rect 18042 8726 18076 8760
rect 18132 8726 18166 8760
rect 18222 8726 18256 8760
rect 18312 8726 18346 8760
rect 18402 8726 18436 8760
rect 18492 8726 18526 8760
rect 12800 7978 12834 8012
rect 12890 7978 12924 8012
rect 12980 7978 13014 8012
rect 13070 7978 13104 8012
rect 13160 7978 13194 8012
rect 13250 7978 13284 8012
rect 13340 7978 13374 8012
rect 12800 7888 12834 7922
rect 12890 7888 12924 7922
rect 12980 7888 13014 7922
rect 13070 7888 13104 7922
rect 13160 7888 13194 7922
rect 13250 7888 13284 7922
rect 13340 7888 13374 7922
rect 12800 7798 12834 7832
rect 12890 7798 12924 7832
rect 12980 7798 13014 7832
rect 13070 7798 13104 7832
rect 13160 7798 13194 7832
rect 13250 7798 13284 7832
rect 13340 7798 13374 7832
rect 12800 7708 12834 7742
rect 12890 7708 12924 7742
rect 12980 7708 13014 7742
rect 13070 7708 13104 7742
rect 13160 7708 13194 7742
rect 13250 7708 13284 7742
rect 13340 7708 13374 7742
rect 12800 7618 12834 7652
rect 12890 7618 12924 7652
rect 12980 7618 13014 7652
rect 13070 7618 13104 7652
rect 13160 7618 13194 7652
rect 13250 7618 13284 7652
rect 13340 7618 13374 7652
rect 12800 7528 12834 7562
rect 12890 7528 12924 7562
rect 12980 7528 13014 7562
rect 13070 7528 13104 7562
rect 13160 7528 13194 7562
rect 13250 7528 13284 7562
rect 13340 7528 13374 7562
rect 12800 7438 12834 7472
rect 12890 7438 12924 7472
rect 12980 7438 13014 7472
rect 13070 7438 13104 7472
rect 13160 7438 13194 7472
rect 13250 7438 13284 7472
rect 13340 7438 13374 7472
rect 14088 7978 14122 8012
rect 14178 7978 14212 8012
rect 14268 7978 14302 8012
rect 14358 7978 14392 8012
rect 14448 7978 14482 8012
rect 14538 7978 14572 8012
rect 14628 7978 14662 8012
rect 14088 7888 14122 7922
rect 14178 7888 14212 7922
rect 14268 7888 14302 7922
rect 14358 7888 14392 7922
rect 14448 7888 14482 7922
rect 14538 7888 14572 7922
rect 14628 7888 14662 7922
rect 14088 7798 14122 7832
rect 14178 7798 14212 7832
rect 14268 7798 14302 7832
rect 14358 7798 14392 7832
rect 14448 7798 14482 7832
rect 14538 7798 14572 7832
rect 14628 7798 14662 7832
rect 14088 7708 14122 7742
rect 14178 7708 14212 7742
rect 14268 7708 14302 7742
rect 14358 7708 14392 7742
rect 14448 7708 14482 7742
rect 14538 7708 14572 7742
rect 14628 7708 14662 7742
rect 14088 7618 14122 7652
rect 14178 7618 14212 7652
rect 14268 7618 14302 7652
rect 14358 7618 14392 7652
rect 14448 7618 14482 7652
rect 14538 7618 14572 7652
rect 14628 7618 14662 7652
rect 14088 7528 14122 7562
rect 14178 7528 14212 7562
rect 14268 7528 14302 7562
rect 14358 7528 14392 7562
rect 14448 7528 14482 7562
rect 14538 7528 14572 7562
rect 14628 7528 14662 7562
rect 14088 7438 14122 7472
rect 14178 7438 14212 7472
rect 14268 7438 14302 7472
rect 14358 7438 14392 7472
rect 14448 7438 14482 7472
rect 14538 7438 14572 7472
rect 14628 7438 14662 7472
rect 15376 7978 15410 8012
rect 15466 7978 15500 8012
rect 15556 7978 15590 8012
rect 15646 7978 15680 8012
rect 15736 7978 15770 8012
rect 15826 7978 15860 8012
rect 15916 7978 15950 8012
rect 15376 7888 15410 7922
rect 15466 7888 15500 7922
rect 15556 7888 15590 7922
rect 15646 7888 15680 7922
rect 15736 7888 15770 7922
rect 15826 7888 15860 7922
rect 15916 7888 15950 7922
rect 15376 7798 15410 7832
rect 15466 7798 15500 7832
rect 15556 7798 15590 7832
rect 15646 7798 15680 7832
rect 15736 7798 15770 7832
rect 15826 7798 15860 7832
rect 15916 7798 15950 7832
rect 15376 7708 15410 7742
rect 15466 7708 15500 7742
rect 15556 7708 15590 7742
rect 15646 7708 15680 7742
rect 15736 7708 15770 7742
rect 15826 7708 15860 7742
rect 15916 7708 15950 7742
rect 15376 7618 15410 7652
rect 15466 7618 15500 7652
rect 15556 7618 15590 7652
rect 15646 7618 15680 7652
rect 15736 7618 15770 7652
rect 15826 7618 15860 7652
rect 15916 7618 15950 7652
rect 15376 7528 15410 7562
rect 15466 7528 15500 7562
rect 15556 7528 15590 7562
rect 15646 7528 15680 7562
rect 15736 7528 15770 7562
rect 15826 7528 15860 7562
rect 15916 7528 15950 7562
rect 15376 7438 15410 7472
rect 15466 7438 15500 7472
rect 15556 7438 15590 7472
rect 15646 7438 15680 7472
rect 15736 7438 15770 7472
rect 15826 7438 15860 7472
rect 15916 7438 15950 7472
rect 16664 7978 16698 8012
rect 16754 7978 16788 8012
rect 16844 7978 16878 8012
rect 16934 7978 16968 8012
rect 17024 7978 17058 8012
rect 17114 7978 17148 8012
rect 17204 7978 17238 8012
rect 16664 7888 16698 7922
rect 16754 7888 16788 7922
rect 16844 7888 16878 7922
rect 16934 7888 16968 7922
rect 17024 7888 17058 7922
rect 17114 7888 17148 7922
rect 17204 7888 17238 7922
rect 16664 7798 16698 7832
rect 16754 7798 16788 7832
rect 16844 7798 16878 7832
rect 16934 7798 16968 7832
rect 17024 7798 17058 7832
rect 17114 7798 17148 7832
rect 17204 7798 17238 7832
rect 16664 7708 16698 7742
rect 16754 7708 16788 7742
rect 16844 7708 16878 7742
rect 16934 7708 16968 7742
rect 17024 7708 17058 7742
rect 17114 7708 17148 7742
rect 17204 7708 17238 7742
rect 16664 7618 16698 7652
rect 16754 7618 16788 7652
rect 16844 7618 16878 7652
rect 16934 7618 16968 7652
rect 17024 7618 17058 7652
rect 17114 7618 17148 7652
rect 17204 7618 17238 7652
rect 16664 7528 16698 7562
rect 16754 7528 16788 7562
rect 16844 7528 16878 7562
rect 16934 7528 16968 7562
rect 17024 7528 17058 7562
rect 17114 7528 17148 7562
rect 17204 7528 17238 7562
rect 16664 7438 16698 7472
rect 16754 7438 16788 7472
rect 16844 7438 16878 7472
rect 16934 7438 16968 7472
rect 17024 7438 17058 7472
rect 17114 7438 17148 7472
rect 17204 7438 17238 7472
rect 17952 7978 17986 8012
rect 18042 7978 18076 8012
rect 18132 7978 18166 8012
rect 18222 7978 18256 8012
rect 18312 7978 18346 8012
rect 18402 7978 18436 8012
rect 18492 7978 18526 8012
rect 17952 7888 17986 7922
rect 18042 7888 18076 7922
rect 18132 7888 18166 7922
rect 18222 7888 18256 7922
rect 18312 7888 18346 7922
rect 18402 7888 18436 7922
rect 18492 7888 18526 7922
rect 17952 7798 17986 7832
rect 18042 7798 18076 7832
rect 18132 7798 18166 7832
rect 18222 7798 18256 7832
rect 18312 7798 18346 7832
rect 18402 7798 18436 7832
rect 18492 7798 18526 7832
rect 17952 7708 17986 7742
rect 18042 7708 18076 7742
rect 18132 7708 18166 7742
rect 18222 7708 18256 7742
rect 18312 7708 18346 7742
rect 18402 7708 18436 7742
rect 18492 7708 18526 7742
rect 17952 7618 17986 7652
rect 18042 7618 18076 7652
rect 18132 7618 18166 7652
rect 18222 7618 18256 7652
rect 18312 7618 18346 7652
rect 18402 7618 18436 7652
rect 18492 7618 18526 7652
rect 17952 7528 17986 7562
rect 18042 7528 18076 7562
rect 18132 7528 18166 7562
rect 18222 7528 18256 7562
rect 18312 7528 18346 7562
rect 18402 7528 18436 7562
rect 18492 7528 18526 7562
rect 17952 7438 17986 7472
rect 18042 7438 18076 7472
rect 18132 7438 18166 7472
rect 18222 7438 18256 7472
rect 18312 7438 18346 7472
rect 18402 7438 18436 7472
rect 18492 7438 18526 7472
rect 12800 6690 12834 6724
rect 12890 6690 12924 6724
rect 12980 6690 13014 6724
rect 13070 6690 13104 6724
rect 13160 6690 13194 6724
rect 13250 6690 13284 6724
rect 13340 6690 13374 6724
rect 12800 6600 12834 6634
rect 12890 6600 12924 6634
rect 12980 6600 13014 6634
rect 13070 6600 13104 6634
rect 13160 6600 13194 6634
rect 13250 6600 13284 6634
rect 13340 6600 13374 6634
rect 12800 6510 12834 6544
rect 12890 6510 12924 6544
rect 12980 6510 13014 6544
rect 13070 6510 13104 6544
rect 13160 6510 13194 6544
rect 13250 6510 13284 6544
rect 13340 6510 13374 6544
rect 12800 6420 12834 6454
rect 12890 6420 12924 6454
rect 12980 6420 13014 6454
rect 13070 6420 13104 6454
rect 13160 6420 13194 6454
rect 13250 6420 13284 6454
rect 13340 6420 13374 6454
rect 12800 6330 12834 6364
rect 12890 6330 12924 6364
rect 12980 6330 13014 6364
rect 13070 6330 13104 6364
rect 13160 6330 13194 6364
rect 13250 6330 13284 6364
rect 13340 6330 13374 6364
rect 12800 6240 12834 6274
rect 12890 6240 12924 6274
rect 12980 6240 13014 6274
rect 13070 6240 13104 6274
rect 13160 6240 13194 6274
rect 13250 6240 13284 6274
rect 13340 6240 13374 6274
rect 12800 6150 12834 6184
rect 12890 6150 12924 6184
rect 12980 6150 13014 6184
rect 13070 6150 13104 6184
rect 13160 6150 13194 6184
rect 13250 6150 13284 6184
rect 13340 6150 13374 6184
rect 14088 6690 14122 6724
rect 14178 6690 14212 6724
rect 14268 6690 14302 6724
rect 14358 6690 14392 6724
rect 14448 6690 14482 6724
rect 14538 6690 14572 6724
rect 14628 6690 14662 6724
rect 14088 6600 14122 6634
rect 14178 6600 14212 6634
rect 14268 6600 14302 6634
rect 14358 6600 14392 6634
rect 14448 6600 14482 6634
rect 14538 6600 14572 6634
rect 14628 6600 14662 6634
rect 14088 6510 14122 6544
rect 14178 6510 14212 6544
rect 14268 6510 14302 6544
rect 14358 6510 14392 6544
rect 14448 6510 14482 6544
rect 14538 6510 14572 6544
rect 14628 6510 14662 6544
rect 14088 6420 14122 6454
rect 14178 6420 14212 6454
rect 14268 6420 14302 6454
rect 14358 6420 14392 6454
rect 14448 6420 14482 6454
rect 14538 6420 14572 6454
rect 14628 6420 14662 6454
rect 14088 6330 14122 6364
rect 14178 6330 14212 6364
rect 14268 6330 14302 6364
rect 14358 6330 14392 6364
rect 14448 6330 14482 6364
rect 14538 6330 14572 6364
rect 14628 6330 14662 6364
rect 14088 6240 14122 6274
rect 14178 6240 14212 6274
rect 14268 6240 14302 6274
rect 14358 6240 14392 6274
rect 14448 6240 14482 6274
rect 14538 6240 14572 6274
rect 14628 6240 14662 6274
rect 14088 6150 14122 6184
rect 14178 6150 14212 6184
rect 14268 6150 14302 6184
rect 14358 6150 14392 6184
rect 14448 6150 14482 6184
rect 14538 6150 14572 6184
rect 14628 6150 14662 6184
rect 15376 6690 15410 6724
rect 15466 6690 15500 6724
rect 15556 6690 15590 6724
rect 15646 6690 15680 6724
rect 15736 6690 15770 6724
rect 15826 6690 15860 6724
rect 15916 6690 15950 6724
rect 15376 6600 15410 6634
rect 15466 6600 15500 6634
rect 15556 6600 15590 6634
rect 15646 6600 15680 6634
rect 15736 6600 15770 6634
rect 15826 6600 15860 6634
rect 15916 6600 15950 6634
rect 15376 6510 15410 6544
rect 15466 6510 15500 6544
rect 15556 6510 15590 6544
rect 15646 6510 15680 6544
rect 15736 6510 15770 6544
rect 15826 6510 15860 6544
rect 15916 6510 15950 6544
rect 15376 6420 15410 6454
rect 15466 6420 15500 6454
rect 15556 6420 15590 6454
rect 15646 6420 15680 6454
rect 15736 6420 15770 6454
rect 15826 6420 15860 6454
rect 15916 6420 15950 6454
rect 15376 6330 15410 6364
rect 15466 6330 15500 6364
rect 15556 6330 15590 6364
rect 15646 6330 15680 6364
rect 15736 6330 15770 6364
rect 15826 6330 15860 6364
rect 15916 6330 15950 6364
rect 15376 6240 15410 6274
rect 15466 6240 15500 6274
rect 15556 6240 15590 6274
rect 15646 6240 15680 6274
rect 15736 6240 15770 6274
rect 15826 6240 15860 6274
rect 15916 6240 15950 6274
rect 15376 6150 15410 6184
rect 15466 6150 15500 6184
rect 15556 6150 15590 6184
rect 15646 6150 15680 6184
rect 15736 6150 15770 6184
rect 15826 6150 15860 6184
rect 15916 6150 15950 6184
rect 16664 6690 16698 6724
rect 16754 6690 16788 6724
rect 16844 6690 16878 6724
rect 16934 6690 16968 6724
rect 17024 6690 17058 6724
rect 17114 6690 17148 6724
rect 17204 6690 17238 6724
rect 16664 6600 16698 6634
rect 16754 6600 16788 6634
rect 16844 6600 16878 6634
rect 16934 6600 16968 6634
rect 17024 6600 17058 6634
rect 17114 6600 17148 6634
rect 17204 6600 17238 6634
rect 16664 6510 16698 6544
rect 16754 6510 16788 6544
rect 16844 6510 16878 6544
rect 16934 6510 16968 6544
rect 17024 6510 17058 6544
rect 17114 6510 17148 6544
rect 17204 6510 17238 6544
rect 16664 6420 16698 6454
rect 16754 6420 16788 6454
rect 16844 6420 16878 6454
rect 16934 6420 16968 6454
rect 17024 6420 17058 6454
rect 17114 6420 17148 6454
rect 17204 6420 17238 6454
rect 16664 6330 16698 6364
rect 16754 6330 16788 6364
rect 16844 6330 16878 6364
rect 16934 6330 16968 6364
rect 17024 6330 17058 6364
rect 17114 6330 17148 6364
rect 17204 6330 17238 6364
rect 16664 6240 16698 6274
rect 16754 6240 16788 6274
rect 16844 6240 16878 6274
rect 16934 6240 16968 6274
rect 17024 6240 17058 6274
rect 17114 6240 17148 6274
rect 17204 6240 17238 6274
rect 16664 6150 16698 6184
rect 16754 6150 16788 6184
rect 16844 6150 16878 6184
rect 16934 6150 16968 6184
rect 17024 6150 17058 6184
rect 17114 6150 17148 6184
rect 17204 6150 17238 6184
rect 17952 6690 17986 6724
rect 18042 6690 18076 6724
rect 18132 6690 18166 6724
rect 18222 6690 18256 6724
rect 18312 6690 18346 6724
rect 18402 6690 18436 6724
rect 18492 6690 18526 6724
rect 17952 6600 17986 6634
rect 18042 6600 18076 6634
rect 18132 6600 18166 6634
rect 18222 6600 18256 6634
rect 18312 6600 18346 6634
rect 18402 6600 18436 6634
rect 18492 6600 18526 6634
rect 17952 6510 17986 6544
rect 18042 6510 18076 6544
rect 18132 6510 18166 6544
rect 18222 6510 18256 6544
rect 18312 6510 18346 6544
rect 18402 6510 18436 6544
rect 18492 6510 18526 6544
rect 17952 6420 17986 6454
rect 18042 6420 18076 6454
rect 18132 6420 18166 6454
rect 18222 6420 18256 6454
rect 18312 6420 18346 6454
rect 18402 6420 18436 6454
rect 18492 6420 18526 6454
rect 17952 6330 17986 6364
rect 18042 6330 18076 6364
rect 18132 6330 18166 6364
rect 18222 6330 18256 6364
rect 18312 6330 18346 6364
rect 18402 6330 18436 6364
rect 18492 6330 18526 6364
rect 17952 6240 17986 6274
rect 18042 6240 18076 6274
rect 18132 6240 18166 6274
rect 18222 6240 18256 6274
rect 18312 6240 18346 6274
rect 18402 6240 18436 6274
rect 18492 6240 18526 6274
rect 17952 6150 17986 6184
rect 18042 6150 18076 6184
rect 18132 6150 18166 6184
rect 18222 6150 18256 6184
rect 18312 6150 18346 6184
rect 18402 6150 18436 6184
rect 18492 6150 18526 6184
rect 12800 5402 12834 5436
rect 12890 5402 12924 5436
rect 12980 5402 13014 5436
rect 13070 5402 13104 5436
rect 13160 5402 13194 5436
rect 13250 5402 13284 5436
rect 13340 5402 13374 5436
rect 12800 5312 12834 5346
rect 12890 5312 12924 5346
rect 12980 5312 13014 5346
rect 13070 5312 13104 5346
rect 13160 5312 13194 5346
rect 13250 5312 13284 5346
rect 13340 5312 13374 5346
rect 12800 5222 12834 5256
rect 12890 5222 12924 5256
rect 12980 5222 13014 5256
rect 13070 5222 13104 5256
rect 13160 5222 13194 5256
rect 13250 5222 13284 5256
rect 13340 5222 13374 5256
rect 12800 5132 12834 5166
rect 12890 5132 12924 5166
rect 12980 5132 13014 5166
rect 13070 5132 13104 5166
rect 13160 5132 13194 5166
rect 13250 5132 13284 5166
rect 13340 5132 13374 5166
rect 12800 5042 12834 5076
rect 12890 5042 12924 5076
rect 12980 5042 13014 5076
rect 13070 5042 13104 5076
rect 13160 5042 13194 5076
rect 13250 5042 13284 5076
rect 13340 5042 13374 5076
rect 12800 4952 12834 4986
rect 12890 4952 12924 4986
rect 12980 4952 13014 4986
rect 13070 4952 13104 4986
rect 13160 4952 13194 4986
rect 13250 4952 13284 4986
rect 13340 4952 13374 4986
rect 12800 4862 12834 4896
rect 12890 4862 12924 4896
rect 12980 4862 13014 4896
rect 13070 4862 13104 4896
rect 13160 4862 13194 4896
rect 13250 4862 13284 4896
rect 13340 4862 13374 4896
rect 14088 5402 14122 5436
rect 14178 5402 14212 5436
rect 14268 5402 14302 5436
rect 14358 5402 14392 5436
rect 14448 5402 14482 5436
rect 14538 5402 14572 5436
rect 14628 5402 14662 5436
rect 14088 5312 14122 5346
rect 14178 5312 14212 5346
rect 14268 5312 14302 5346
rect 14358 5312 14392 5346
rect 14448 5312 14482 5346
rect 14538 5312 14572 5346
rect 14628 5312 14662 5346
rect 14088 5222 14122 5256
rect 14178 5222 14212 5256
rect 14268 5222 14302 5256
rect 14358 5222 14392 5256
rect 14448 5222 14482 5256
rect 14538 5222 14572 5256
rect 14628 5222 14662 5256
rect 14088 5132 14122 5166
rect 14178 5132 14212 5166
rect 14268 5132 14302 5166
rect 14358 5132 14392 5166
rect 14448 5132 14482 5166
rect 14538 5132 14572 5166
rect 14628 5132 14662 5166
rect 14088 5042 14122 5076
rect 14178 5042 14212 5076
rect 14268 5042 14302 5076
rect 14358 5042 14392 5076
rect 14448 5042 14482 5076
rect 14538 5042 14572 5076
rect 14628 5042 14662 5076
rect 14088 4952 14122 4986
rect 14178 4952 14212 4986
rect 14268 4952 14302 4986
rect 14358 4952 14392 4986
rect 14448 4952 14482 4986
rect 14538 4952 14572 4986
rect 14628 4952 14662 4986
rect 14088 4862 14122 4896
rect 14178 4862 14212 4896
rect 14268 4862 14302 4896
rect 14358 4862 14392 4896
rect 14448 4862 14482 4896
rect 14538 4862 14572 4896
rect 14628 4862 14662 4896
rect 15376 5402 15410 5436
rect 15466 5402 15500 5436
rect 15556 5402 15590 5436
rect 15646 5402 15680 5436
rect 15736 5402 15770 5436
rect 15826 5402 15860 5436
rect 15916 5402 15950 5436
rect 15376 5312 15410 5346
rect 15466 5312 15500 5346
rect 15556 5312 15590 5346
rect 15646 5312 15680 5346
rect 15736 5312 15770 5346
rect 15826 5312 15860 5346
rect 15916 5312 15950 5346
rect 15376 5222 15410 5256
rect 15466 5222 15500 5256
rect 15556 5222 15590 5256
rect 15646 5222 15680 5256
rect 15736 5222 15770 5256
rect 15826 5222 15860 5256
rect 15916 5222 15950 5256
rect 15376 5132 15410 5166
rect 15466 5132 15500 5166
rect 15556 5132 15590 5166
rect 15646 5132 15680 5166
rect 15736 5132 15770 5166
rect 15826 5132 15860 5166
rect 15916 5132 15950 5166
rect 15376 5042 15410 5076
rect 15466 5042 15500 5076
rect 15556 5042 15590 5076
rect 15646 5042 15680 5076
rect 15736 5042 15770 5076
rect 15826 5042 15860 5076
rect 15916 5042 15950 5076
rect 15376 4952 15410 4986
rect 15466 4952 15500 4986
rect 15556 4952 15590 4986
rect 15646 4952 15680 4986
rect 15736 4952 15770 4986
rect 15826 4952 15860 4986
rect 15916 4952 15950 4986
rect 15376 4862 15410 4896
rect 15466 4862 15500 4896
rect 15556 4862 15590 4896
rect 15646 4862 15680 4896
rect 15736 4862 15770 4896
rect 15826 4862 15860 4896
rect 15916 4862 15950 4896
rect 16664 5402 16698 5436
rect 16754 5402 16788 5436
rect 16844 5402 16878 5436
rect 16934 5402 16968 5436
rect 17024 5402 17058 5436
rect 17114 5402 17148 5436
rect 17204 5402 17238 5436
rect 16664 5312 16698 5346
rect 16754 5312 16788 5346
rect 16844 5312 16878 5346
rect 16934 5312 16968 5346
rect 17024 5312 17058 5346
rect 17114 5312 17148 5346
rect 17204 5312 17238 5346
rect 16664 5222 16698 5256
rect 16754 5222 16788 5256
rect 16844 5222 16878 5256
rect 16934 5222 16968 5256
rect 17024 5222 17058 5256
rect 17114 5222 17148 5256
rect 17204 5222 17238 5256
rect 16664 5132 16698 5166
rect 16754 5132 16788 5166
rect 16844 5132 16878 5166
rect 16934 5132 16968 5166
rect 17024 5132 17058 5166
rect 17114 5132 17148 5166
rect 17204 5132 17238 5166
rect 16664 5042 16698 5076
rect 16754 5042 16788 5076
rect 16844 5042 16878 5076
rect 16934 5042 16968 5076
rect 17024 5042 17058 5076
rect 17114 5042 17148 5076
rect 17204 5042 17238 5076
rect 16664 4952 16698 4986
rect 16754 4952 16788 4986
rect 16844 4952 16878 4986
rect 16934 4952 16968 4986
rect 17024 4952 17058 4986
rect 17114 4952 17148 4986
rect 17204 4952 17238 4986
rect 16664 4862 16698 4896
rect 16754 4862 16788 4896
rect 16844 4862 16878 4896
rect 16934 4862 16968 4896
rect 17024 4862 17058 4896
rect 17114 4862 17148 4896
rect 17204 4862 17238 4896
rect 17952 5402 17986 5436
rect 18042 5402 18076 5436
rect 18132 5402 18166 5436
rect 18222 5402 18256 5436
rect 18312 5402 18346 5436
rect 18402 5402 18436 5436
rect 18492 5402 18526 5436
rect 17952 5312 17986 5346
rect 18042 5312 18076 5346
rect 18132 5312 18166 5346
rect 18222 5312 18256 5346
rect 18312 5312 18346 5346
rect 18402 5312 18436 5346
rect 18492 5312 18526 5346
rect 17952 5222 17986 5256
rect 18042 5222 18076 5256
rect 18132 5222 18166 5256
rect 18222 5222 18256 5256
rect 18312 5222 18346 5256
rect 18402 5222 18436 5256
rect 18492 5222 18526 5256
rect 17952 5132 17986 5166
rect 18042 5132 18076 5166
rect 18132 5132 18166 5166
rect 18222 5132 18256 5166
rect 18312 5132 18346 5166
rect 18402 5132 18436 5166
rect 18492 5132 18526 5166
rect 17952 5042 17986 5076
rect 18042 5042 18076 5076
rect 18132 5042 18166 5076
rect 18222 5042 18256 5076
rect 18312 5042 18346 5076
rect 18402 5042 18436 5076
rect 18492 5042 18526 5076
rect 17952 4952 17986 4986
rect 18042 4952 18076 4986
rect 18132 4952 18166 4986
rect 18222 4952 18256 4986
rect 18312 4952 18346 4986
rect 18402 4952 18436 4986
rect 18492 4952 18526 4986
rect 17952 4862 17986 4896
rect 18042 4862 18076 4896
rect 18132 4862 18166 4896
rect 18222 4862 18256 4896
rect 18312 4862 18346 4896
rect 18402 4862 18436 4896
rect 18492 4862 18526 4896
rect 12800 4114 12834 4148
rect 12890 4114 12924 4148
rect 12980 4114 13014 4148
rect 13070 4114 13104 4148
rect 13160 4114 13194 4148
rect 13250 4114 13284 4148
rect 13340 4114 13374 4148
rect 12800 4024 12834 4058
rect 12890 4024 12924 4058
rect 12980 4024 13014 4058
rect 13070 4024 13104 4058
rect 13160 4024 13194 4058
rect 13250 4024 13284 4058
rect 13340 4024 13374 4058
rect 12800 3934 12834 3968
rect 12890 3934 12924 3968
rect 12980 3934 13014 3968
rect 13070 3934 13104 3968
rect 13160 3934 13194 3968
rect 13250 3934 13284 3968
rect 13340 3934 13374 3968
rect 12800 3844 12834 3878
rect 12890 3844 12924 3878
rect 12980 3844 13014 3878
rect 13070 3844 13104 3878
rect 13160 3844 13194 3878
rect 13250 3844 13284 3878
rect 13340 3844 13374 3878
rect 12800 3754 12834 3788
rect 12890 3754 12924 3788
rect 12980 3754 13014 3788
rect 13070 3754 13104 3788
rect 13160 3754 13194 3788
rect 13250 3754 13284 3788
rect 13340 3754 13374 3788
rect 12800 3664 12834 3698
rect 12890 3664 12924 3698
rect 12980 3664 13014 3698
rect 13070 3664 13104 3698
rect 13160 3664 13194 3698
rect 13250 3664 13284 3698
rect 13340 3664 13374 3698
rect 12800 3574 12834 3608
rect 12890 3574 12924 3608
rect 12980 3574 13014 3608
rect 13070 3574 13104 3608
rect 13160 3574 13194 3608
rect 13250 3574 13284 3608
rect 13340 3574 13374 3608
rect 14088 4114 14122 4148
rect 14178 4114 14212 4148
rect 14268 4114 14302 4148
rect 14358 4114 14392 4148
rect 14448 4114 14482 4148
rect 14538 4114 14572 4148
rect 14628 4114 14662 4148
rect 14088 4024 14122 4058
rect 14178 4024 14212 4058
rect 14268 4024 14302 4058
rect 14358 4024 14392 4058
rect 14448 4024 14482 4058
rect 14538 4024 14572 4058
rect 14628 4024 14662 4058
rect 14088 3934 14122 3968
rect 14178 3934 14212 3968
rect 14268 3934 14302 3968
rect 14358 3934 14392 3968
rect 14448 3934 14482 3968
rect 14538 3934 14572 3968
rect 14628 3934 14662 3968
rect 14088 3844 14122 3878
rect 14178 3844 14212 3878
rect 14268 3844 14302 3878
rect 14358 3844 14392 3878
rect 14448 3844 14482 3878
rect 14538 3844 14572 3878
rect 14628 3844 14662 3878
rect 14088 3754 14122 3788
rect 14178 3754 14212 3788
rect 14268 3754 14302 3788
rect 14358 3754 14392 3788
rect 14448 3754 14482 3788
rect 14538 3754 14572 3788
rect 14628 3754 14662 3788
rect 14088 3664 14122 3698
rect 14178 3664 14212 3698
rect 14268 3664 14302 3698
rect 14358 3664 14392 3698
rect 14448 3664 14482 3698
rect 14538 3664 14572 3698
rect 14628 3664 14662 3698
rect 14088 3574 14122 3608
rect 14178 3574 14212 3608
rect 14268 3574 14302 3608
rect 14358 3574 14392 3608
rect 14448 3574 14482 3608
rect 14538 3574 14572 3608
rect 14628 3574 14662 3608
rect 15376 4114 15410 4148
rect 15466 4114 15500 4148
rect 15556 4114 15590 4148
rect 15646 4114 15680 4148
rect 15736 4114 15770 4148
rect 15826 4114 15860 4148
rect 15916 4114 15950 4148
rect 15376 4024 15410 4058
rect 15466 4024 15500 4058
rect 15556 4024 15590 4058
rect 15646 4024 15680 4058
rect 15736 4024 15770 4058
rect 15826 4024 15860 4058
rect 15916 4024 15950 4058
rect 15376 3934 15410 3968
rect 15466 3934 15500 3968
rect 15556 3934 15590 3968
rect 15646 3934 15680 3968
rect 15736 3934 15770 3968
rect 15826 3934 15860 3968
rect 15916 3934 15950 3968
rect 15376 3844 15410 3878
rect 15466 3844 15500 3878
rect 15556 3844 15590 3878
rect 15646 3844 15680 3878
rect 15736 3844 15770 3878
rect 15826 3844 15860 3878
rect 15916 3844 15950 3878
rect 15376 3754 15410 3788
rect 15466 3754 15500 3788
rect 15556 3754 15590 3788
rect 15646 3754 15680 3788
rect 15736 3754 15770 3788
rect 15826 3754 15860 3788
rect 15916 3754 15950 3788
rect 15376 3664 15410 3698
rect 15466 3664 15500 3698
rect 15556 3664 15590 3698
rect 15646 3664 15680 3698
rect 15736 3664 15770 3698
rect 15826 3664 15860 3698
rect 15916 3664 15950 3698
rect 15376 3574 15410 3608
rect 15466 3574 15500 3608
rect 15556 3574 15590 3608
rect 15646 3574 15680 3608
rect 15736 3574 15770 3608
rect 15826 3574 15860 3608
rect 15916 3574 15950 3608
rect 16664 4114 16698 4148
rect 16754 4114 16788 4148
rect 16844 4114 16878 4148
rect 16934 4114 16968 4148
rect 17024 4114 17058 4148
rect 17114 4114 17148 4148
rect 17204 4114 17238 4148
rect 16664 4024 16698 4058
rect 16754 4024 16788 4058
rect 16844 4024 16878 4058
rect 16934 4024 16968 4058
rect 17024 4024 17058 4058
rect 17114 4024 17148 4058
rect 17204 4024 17238 4058
rect 16664 3934 16698 3968
rect 16754 3934 16788 3968
rect 16844 3934 16878 3968
rect 16934 3934 16968 3968
rect 17024 3934 17058 3968
rect 17114 3934 17148 3968
rect 17204 3934 17238 3968
rect 16664 3844 16698 3878
rect 16754 3844 16788 3878
rect 16844 3844 16878 3878
rect 16934 3844 16968 3878
rect 17024 3844 17058 3878
rect 17114 3844 17148 3878
rect 17204 3844 17238 3878
rect 16664 3754 16698 3788
rect 16754 3754 16788 3788
rect 16844 3754 16878 3788
rect 16934 3754 16968 3788
rect 17024 3754 17058 3788
rect 17114 3754 17148 3788
rect 17204 3754 17238 3788
rect 16664 3664 16698 3698
rect 16754 3664 16788 3698
rect 16844 3664 16878 3698
rect 16934 3664 16968 3698
rect 17024 3664 17058 3698
rect 17114 3664 17148 3698
rect 17204 3664 17238 3698
rect 16664 3574 16698 3608
rect 16754 3574 16788 3608
rect 16844 3574 16878 3608
rect 16934 3574 16968 3608
rect 17024 3574 17058 3608
rect 17114 3574 17148 3608
rect 17204 3574 17238 3608
rect 17952 4114 17986 4148
rect 18042 4114 18076 4148
rect 18132 4114 18166 4148
rect 18222 4114 18256 4148
rect 18312 4114 18346 4148
rect 18402 4114 18436 4148
rect 18492 4114 18526 4148
rect 17952 4024 17986 4058
rect 18042 4024 18076 4058
rect 18132 4024 18166 4058
rect 18222 4024 18256 4058
rect 18312 4024 18346 4058
rect 18402 4024 18436 4058
rect 18492 4024 18526 4058
rect 17952 3934 17986 3968
rect 18042 3934 18076 3968
rect 18132 3934 18166 3968
rect 18222 3934 18256 3968
rect 18312 3934 18346 3968
rect 18402 3934 18436 3968
rect 18492 3934 18526 3968
rect 17952 3844 17986 3878
rect 18042 3844 18076 3878
rect 18132 3844 18166 3878
rect 18222 3844 18256 3878
rect 18312 3844 18346 3878
rect 18402 3844 18436 3878
rect 18492 3844 18526 3878
rect 17952 3754 17986 3788
rect 18042 3754 18076 3788
rect 18132 3754 18166 3788
rect 18222 3754 18256 3788
rect 18312 3754 18346 3788
rect 18402 3754 18436 3788
rect 18492 3754 18526 3788
rect 17952 3664 17986 3698
rect 18042 3664 18076 3698
rect 18132 3664 18166 3698
rect 18222 3664 18256 3698
rect 18312 3664 18346 3698
rect 18402 3664 18436 3698
rect 18492 3664 18526 3698
rect 17952 3574 17986 3608
rect 18042 3574 18076 3608
rect 18132 3574 18166 3608
rect 18222 3574 18256 3608
rect 18312 3574 18346 3608
rect 18402 3574 18436 3608
rect 18492 3574 18526 3608
rect 12800 2826 12834 2860
rect 12890 2826 12924 2860
rect 12980 2826 13014 2860
rect 13070 2826 13104 2860
rect 13160 2826 13194 2860
rect 13250 2826 13284 2860
rect 13340 2826 13374 2860
rect 12800 2736 12834 2770
rect 12890 2736 12924 2770
rect 12980 2736 13014 2770
rect 13070 2736 13104 2770
rect 13160 2736 13194 2770
rect 13250 2736 13284 2770
rect 13340 2736 13374 2770
rect 12800 2646 12834 2680
rect 12890 2646 12924 2680
rect 12980 2646 13014 2680
rect 13070 2646 13104 2680
rect 13160 2646 13194 2680
rect 13250 2646 13284 2680
rect 13340 2646 13374 2680
rect 12800 2556 12834 2590
rect 12890 2556 12924 2590
rect 12980 2556 13014 2590
rect 13070 2556 13104 2590
rect 13160 2556 13194 2590
rect 13250 2556 13284 2590
rect 13340 2556 13374 2590
rect 12800 2466 12834 2500
rect 12890 2466 12924 2500
rect 12980 2466 13014 2500
rect 13070 2466 13104 2500
rect 13160 2466 13194 2500
rect 13250 2466 13284 2500
rect 13340 2466 13374 2500
rect 12800 2376 12834 2410
rect 12890 2376 12924 2410
rect 12980 2376 13014 2410
rect 13070 2376 13104 2410
rect 13160 2376 13194 2410
rect 13250 2376 13284 2410
rect 13340 2376 13374 2410
rect 12800 2286 12834 2320
rect 12890 2286 12924 2320
rect 12980 2286 13014 2320
rect 13070 2286 13104 2320
rect 13160 2286 13194 2320
rect 13250 2286 13284 2320
rect 13340 2286 13374 2320
rect 14088 2826 14122 2860
rect 14178 2826 14212 2860
rect 14268 2826 14302 2860
rect 14358 2826 14392 2860
rect 14448 2826 14482 2860
rect 14538 2826 14572 2860
rect 14628 2826 14662 2860
rect 14088 2736 14122 2770
rect 14178 2736 14212 2770
rect 14268 2736 14302 2770
rect 14358 2736 14392 2770
rect 14448 2736 14482 2770
rect 14538 2736 14572 2770
rect 14628 2736 14662 2770
rect 14088 2646 14122 2680
rect 14178 2646 14212 2680
rect 14268 2646 14302 2680
rect 14358 2646 14392 2680
rect 14448 2646 14482 2680
rect 14538 2646 14572 2680
rect 14628 2646 14662 2680
rect 14088 2556 14122 2590
rect 14178 2556 14212 2590
rect 14268 2556 14302 2590
rect 14358 2556 14392 2590
rect 14448 2556 14482 2590
rect 14538 2556 14572 2590
rect 14628 2556 14662 2590
rect 14088 2466 14122 2500
rect 14178 2466 14212 2500
rect 14268 2466 14302 2500
rect 14358 2466 14392 2500
rect 14448 2466 14482 2500
rect 14538 2466 14572 2500
rect 14628 2466 14662 2500
rect 14088 2376 14122 2410
rect 14178 2376 14212 2410
rect 14268 2376 14302 2410
rect 14358 2376 14392 2410
rect 14448 2376 14482 2410
rect 14538 2376 14572 2410
rect 14628 2376 14662 2410
rect 14088 2286 14122 2320
rect 14178 2286 14212 2320
rect 14268 2286 14302 2320
rect 14358 2286 14392 2320
rect 14448 2286 14482 2320
rect 14538 2286 14572 2320
rect 14628 2286 14662 2320
rect 15376 2826 15410 2860
rect 15466 2826 15500 2860
rect 15556 2826 15590 2860
rect 15646 2826 15680 2860
rect 15736 2826 15770 2860
rect 15826 2826 15860 2860
rect 15916 2826 15950 2860
rect 15376 2736 15410 2770
rect 15466 2736 15500 2770
rect 15556 2736 15590 2770
rect 15646 2736 15680 2770
rect 15736 2736 15770 2770
rect 15826 2736 15860 2770
rect 15916 2736 15950 2770
rect 15376 2646 15410 2680
rect 15466 2646 15500 2680
rect 15556 2646 15590 2680
rect 15646 2646 15680 2680
rect 15736 2646 15770 2680
rect 15826 2646 15860 2680
rect 15916 2646 15950 2680
rect 15376 2556 15410 2590
rect 15466 2556 15500 2590
rect 15556 2556 15590 2590
rect 15646 2556 15680 2590
rect 15736 2556 15770 2590
rect 15826 2556 15860 2590
rect 15916 2556 15950 2590
rect 15376 2466 15410 2500
rect 15466 2466 15500 2500
rect 15556 2466 15590 2500
rect 15646 2466 15680 2500
rect 15736 2466 15770 2500
rect 15826 2466 15860 2500
rect 15916 2466 15950 2500
rect 15376 2376 15410 2410
rect 15466 2376 15500 2410
rect 15556 2376 15590 2410
rect 15646 2376 15680 2410
rect 15736 2376 15770 2410
rect 15826 2376 15860 2410
rect 15916 2376 15950 2410
rect 15376 2286 15410 2320
rect 15466 2286 15500 2320
rect 15556 2286 15590 2320
rect 15646 2286 15680 2320
rect 15736 2286 15770 2320
rect 15826 2286 15860 2320
rect 15916 2286 15950 2320
rect 16664 2826 16698 2860
rect 16754 2826 16788 2860
rect 16844 2826 16878 2860
rect 16934 2826 16968 2860
rect 17024 2826 17058 2860
rect 17114 2826 17148 2860
rect 17204 2826 17238 2860
rect 16664 2736 16698 2770
rect 16754 2736 16788 2770
rect 16844 2736 16878 2770
rect 16934 2736 16968 2770
rect 17024 2736 17058 2770
rect 17114 2736 17148 2770
rect 17204 2736 17238 2770
rect 16664 2646 16698 2680
rect 16754 2646 16788 2680
rect 16844 2646 16878 2680
rect 16934 2646 16968 2680
rect 17024 2646 17058 2680
rect 17114 2646 17148 2680
rect 17204 2646 17238 2680
rect 16664 2556 16698 2590
rect 16754 2556 16788 2590
rect 16844 2556 16878 2590
rect 16934 2556 16968 2590
rect 17024 2556 17058 2590
rect 17114 2556 17148 2590
rect 17204 2556 17238 2590
rect 16664 2466 16698 2500
rect 16754 2466 16788 2500
rect 16844 2466 16878 2500
rect 16934 2466 16968 2500
rect 17024 2466 17058 2500
rect 17114 2466 17148 2500
rect 17204 2466 17238 2500
rect 16664 2376 16698 2410
rect 16754 2376 16788 2410
rect 16844 2376 16878 2410
rect 16934 2376 16968 2410
rect 17024 2376 17058 2410
rect 17114 2376 17148 2410
rect 17204 2376 17238 2410
rect 16664 2286 16698 2320
rect 16754 2286 16788 2320
rect 16844 2286 16878 2320
rect 16934 2286 16968 2320
rect 17024 2286 17058 2320
rect 17114 2286 17148 2320
rect 17204 2286 17238 2320
rect 17952 2826 17986 2860
rect 18042 2826 18076 2860
rect 18132 2826 18166 2860
rect 18222 2826 18256 2860
rect 18312 2826 18346 2860
rect 18402 2826 18436 2860
rect 18492 2826 18526 2860
rect 17952 2736 17986 2770
rect 18042 2736 18076 2770
rect 18132 2736 18166 2770
rect 18222 2736 18256 2770
rect 18312 2736 18346 2770
rect 18402 2736 18436 2770
rect 18492 2736 18526 2770
rect 17952 2646 17986 2680
rect 18042 2646 18076 2680
rect 18132 2646 18166 2680
rect 18222 2646 18256 2680
rect 18312 2646 18346 2680
rect 18402 2646 18436 2680
rect 18492 2646 18526 2680
rect 17952 2556 17986 2590
rect 18042 2556 18076 2590
rect 18132 2556 18166 2590
rect 18222 2556 18256 2590
rect 18312 2556 18346 2590
rect 18402 2556 18436 2590
rect 18492 2556 18526 2590
rect 17952 2466 17986 2500
rect 18042 2466 18076 2500
rect 18132 2466 18166 2500
rect 18222 2466 18256 2500
rect 18312 2466 18346 2500
rect 18402 2466 18436 2500
rect 18492 2466 18526 2500
rect 17952 2376 17986 2410
rect 18042 2376 18076 2410
rect 18132 2376 18166 2410
rect 18222 2376 18256 2410
rect 18312 2376 18346 2410
rect 18402 2376 18436 2410
rect 18492 2376 18526 2410
rect 17952 2286 17986 2320
rect 18042 2286 18076 2320
rect 18132 2286 18166 2320
rect 18222 2286 18256 2320
rect 18312 2286 18346 2320
rect 18402 2286 18436 2320
rect 18492 2286 18526 2320
<< psubdiff >>
rect -21540 25036 -10308 25060
rect -21540 24270 -21516 25036
rect -10332 24270 -10308 25036
rect -21540 24246 -10308 24270
rect -9780 21500 -9162 21524
rect -9780 15196 -9756 21500
rect -9186 15196 -9162 21500
rect -6536 21500 -5918 21524
rect -9780 15172 -9162 15196
rect -6536 15196 -6512 21500
rect -5942 15196 -5918 21500
rect -1576 21500 -958 21524
rect -6536 15172 -5918 15196
rect -1576 15196 -1552 21500
rect -982 15196 -958 21500
rect -1576 15172 -958 15196
rect 13112 21500 13730 21524
rect 13112 15196 13136 21500
rect 13706 15196 13730 21500
rect 13112 15172 13730 15196
rect 12444 12202 18884 12234
rect 12444 12168 12578 12202
rect 12612 12168 12668 12202
rect 12702 12168 12758 12202
rect 12792 12168 12848 12202
rect 12882 12168 12938 12202
rect 12972 12168 13028 12202
rect 13062 12168 13118 12202
rect 13152 12168 13208 12202
rect 13242 12168 13298 12202
rect 13332 12168 13388 12202
rect 13422 12168 13478 12202
rect 13512 12168 13568 12202
rect 13602 12168 13866 12202
rect 13900 12168 13956 12202
rect 13990 12168 14046 12202
rect 14080 12168 14136 12202
rect 14170 12168 14226 12202
rect 14260 12168 14316 12202
rect 14350 12168 14406 12202
rect 14440 12168 14496 12202
rect 14530 12168 14586 12202
rect 14620 12168 14676 12202
rect 14710 12168 14766 12202
rect 14800 12168 14856 12202
rect 14890 12168 15154 12202
rect 15188 12168 15244 12202
rect 15278 12168 15334 12202
rect 15368 12168 15424 12202
rect 15458 12168 15514 12202
rect 15548 12168 15604 12202
rect 15638 12168 15694 12202
rect 15728 12168 15784 12202
rect 15818 12168 15874 12202
rect 15908 12168 15964 12202
rect 15998 12168 16054 12202
rect 16088 12168 16144 12202
rect 16178 12168 16442 12202
rect 16476 12168 16532 12202
rect 16566 12168 16622 12202
rect 16656 12168 16712 12202
rect 16746 12168 16802 12202
rect 16836 12168 16892 12202
rect 16926 12168 16982 12202
rect 17016 12168 17072 12202
rect 17106 12168 17162 12202
rect 17196 12168 17252 12202
rect 17286 12168 17342 12202
rect 17376 12168 17432 12202
rect 17466 12168 17730 12202
rect 17764 12168 17820 12202
rect 17854 12168 17910 12202
rect 17944 12168 18000 12202
rect 18034 12168 18090 12202
rect 18124 12168 18180 12202
rect 18214 12168 18270 12202
rect 18304 12168 18360 12202
rect 18394 12168 18450 12202
rect 18484 12168 18540 12202
rect 18574 12168 18630 12202
rect 18664 12168 18720 12202
rect 18754 12168 18884 12202
rect 12444 12133 18884 12168
rect 12444 12118 12545 12133
rect 12444 12084 12477 12118
rect 12511 12084 12545 12118
rect 12444 12028 12545 12084
rect 13631 12118 13833 12133
rect 13631 12084 13664 12118
rect 13698 12084 13765 12118
rect 13799 12084 13833 12118
rect 12444 11994 12477 12028
rect 12511 11994 12545 12028
rect 12444 11938 12545 11994
rect 12444 11904 12477 11938
rect 12511 11904 12545 11938
rect 12444 11848 12545 11904
rect 12444 11814 12477 11848
rect 12511 11814 12545 11848
rect 12444 11758 12545 11814
rect 12444 11724 12477 11758
rect 12511 11724 12545 11758
rect 12444 11668 12545 11724
rect 12444 11634 12477 11668
rect 12511 11634 12545 11668
rect 12444 11578 12545 11634
rect 12444 11544 12477 11578
rect 12511 11544 12545 11578
rect 12444 11488 12545 11544
rect 12444 11454 12477 11488
rect 12511 11454 12545 11488
rect 12444 11398 12545 11454
rect 12444 11364 12477 11398
rect 12511 11364 12545 11398
rect 12444 11308 12545 11364
rect 12444 11274 12477 11308
rect 12511 11274 12545 11308
rect 12444 11218 12545 11274
rect 12444 11184 12477 11218
rect 12511 11184 12545 11218
rect 12444 11128 12545 11184
rect 12444 11094 12477 11128
rect 12511 11094 12545 11128
rect 13631 12028 13833 12084
rect 14919 12118 15121 12133
rect 14919 12084 14952 12118
rect 14986 12084 15053 12118
rect 15087 12084 15121 12118
rect 13631 11994 13664 12028
rect 13698 11994 13765 12028
rect 13799 11994 13833 12028
rect 13631 11938 13833 11994
rect 13631 11904 13664 11938
rect 13698 11904 13765 11938
rect 13799 11904 13833 11938
rect 13631 11848 13833 11904
rect 13631 11814 13664 11848
rect 13698 11814 13765 11848
rect 13799 11814 13833 11848
rect 13631 11758 13833 11814
rect 13631 11724 13664 11758
rect 13698 11724 13765 11758
rect 13799 11724 13833 11758
rect 13631 11668 13833 11724
rect 13631 11634 13664 11668
rect 13698 11634 13765 11668
rect 13799 11634 13833 11668
rect 13631 11578 13833 11634
rect 13631 11544 13664 11578
rect 13698 11544 13765 11578
rect 13799 11544 13833 11578
rect 13631 11488 13833 11544
rect 13631 11454 13664 11488
rect 13698 11454 13765 11488
rect 13799 11454 13833 11488
rect 13631 11398 13833 11454
rect 13631 11364 13664 11398
rect 13698 11364 13765 11398
rect 13799 11364 13833 11398
rect 13631 11308 13833 11364
rect 13631 11274 13664 11308
rect 13698 11274 13765 11308
rect 13799 11274 13833 11308
rect 13631 11218 13833 11274
rect 13631 11184 13664 11218
rect 13698 11184 13765 11218
rect 13799 11184 13833 11218
rect 13631 11128 13833 11184
rect 12444 11047 12545 11094
rect 13631 11094 13664 11128
rect 13698 11094 13765 11128
rect 13799 11094 13833 11128
rect 14919 12028 15121 12084
rect 16207 12118 16409 12133
rect 16207 12084 16240 12118
rect 16274 12084 16341 12118
rect 16375 12084 16409 12118
rect 14919 11994 14952 12028
rect 14986 11994 15053 12028
rect 15087 11994 15121 12028
rect 14919 11938 15121 11994
rect 14919 11904 14952 11938
rect 14986 11904 15053 11938
rect 15087 11904 15121 11938
rect 14919 11848 15121 11904
rect 14919 11814 14952 11848
rect 14986 11814 15053 11848
rect 15087 11814 15121 11848
rect 14919 11758 15121 11814
rect 14919 11724 14952 11758
rect 14986 11724 15053 11758
rect 15087 11724 15121 11758
rect 14919 11668 15121 11724
rect 14919 11634 14952 11668
rect 14986 11634 15053 11668
rect 15087 11634 15121 11668
rect 14919 11578 15121 11634
rect 14919 11544 14952 11578
rect 14986 11544 15053 11578
rect 15087 11544 15121 11578
rect 14919 11488 15121 11544
rect 14919 11454 14952 11488
rect 14986 11454 15053 11488
rect 15087 11454 15121 11488
rect 14919 11398 15121 11454
rect 14919 11364 14952 11398
rect 14986 11364 15053 11398
rect 15087 11364 15121 11398
rect 14919 11308 15121 11364
rect 14919 11274 14952 11308
rect 14986 11274 15053 11308
rect 15087 11274 15121 11308
rect 14919 11218 15121 11274
rect 14919 11184 14952 11218
rect 14986 11184 15053 11218
rect 15087 11184 15121 11218
rect 14919 11128 15121 11184
rect 13631 11047 13833 11094
rect 14919 11094 14952 11128
rect 14986 11094 15053 11128
rect 15087 11094 15121 11128
rect 16207 12028 16409 12084
rect 17495 12118 17697 12133
rect 17495 12084 17528 12118
rect 17562 12084 17629 12118
rect 17663 12084 17697 12118
rect 16207 11994 16240 12028
rect 16274 11994 16341 12028
rect 16375 11994 16409 12028
rect 16207 11938 16409 11994
rect 16207 11904 16240 11938
rect 16274 11904 16341 11938
rect 16375 11904 16409 11938
rect 16207 11848 16409 11904
rect 16207 11814 16240 11848
rect 16274 11814 16341 11848
rect 16375 11814 16409 11848
rect 16207 11758 16409 11814
rect 16207 11724 16240 11758
rect 16274 11724 16341 11758
rect 16375 11724 16409 11758
rect 16207 11668 16409 11724
rect 16207 11634 16240 11668
rect 16274 11634 16341 11668
rect 16375 11634 16409 11668
rect 16207 11578 16409 11634
rect 16207 11544 16240 11578
rect 16274 11544 16341 11578
rect 16375 11544 16409 11578
rect 16207 11488 16409 11544
rect 16207 11454 16240 11488
rect 16274 11454 16341 11488
rect 16375 11454 16409 11488
rect 16207 11398 16409 11454
rect 16207 11364 16240 11398
rect 16274 11364 16341 11398
rect 16375 11364 16409 11398
rect 16207 11308 16409 11364
rect 16207 11274 16240 11308
rect 16274 11274 16341 11308
rect 16375 11274 16409 11308
rect 16207 11218 16409 11274
rect 16207 11184 16240 11218
rect 16274 11184 16341 11218
rect 16375 11184 16409 11218
rect 16207 11128 16409 11184
rect 14919 11047 15121 11094
rect 16207 11094 16240 11128
rect 16274 11094 16341 11128
rect 16375 11094 16409 11128
rect 17495 12028 17697 12084
rect 18783 12118 18884 12133
rect 18783 12084 18816 12118
rect 18850 12084 18884 12118
rect 17495 11994 17528 12028
rect 17562 11994 17629 12028
rect 17663 11994 17697 12028
rect 17495 11938 17697 11994
rect 17495 11904 17528 11938
rect 17562 11904 17629 11938
rect 17663 11904 17697 11938
rect 17495 11848 17697 11904
rect 17495 11814 17528 11848
rect 17562 11814 17629 11848
rect 17663 11814 17697 11848
rect 17495 11758 17697 11814
rect 17495 11724 17528 11758
rect 17562 11724 17629 11758
rect 17663 11724 17697 11758
rect 17495 11668 17697 11724
rect 17495 11634 17528 11668
rect 17562 11634 17629 11668
rect 17663 11634 17697 11668
rect 17495 11578 17697 11634
rect 17495 11544 17528 11578
rect 17562 11544 17629 11578
rect 17663 11544 17697 11578
rect 17495 11488 17697 11544
rect 17495 11454 17528 11488
rect 17562 11454 17629 11488
rect 17663 11454 17697 11488
rect 17495 11398 17697 11454
rect 17495 11364 17528 11398
rect 17562 11364 17629 11398
rect 17663 11364 17697 11398
rect 17495 11308 17697 11364
rect 17495 11274 17528 11308
rect 17562 11274 17629 11308
rect 17663 11274 17697 11308
rect 17495 11218 17697 11274
rect 17495 11184 17528 11218
rect 17562 11184 17629 11218
rect 17663 11184 17697 11218
rect 17495 11128 17697 11184
rect 16207 11047 16409 11094
rect 17495 11094 17528 11128
rect 17562 11094 17629 11128
rect 17663 11094 17697 11128
rect 18783 12028 18884 12084
rect 18783 11994 18816 12028
rect 18850 11994 18884 12028
rect 18783 11938 18884 11994
rect 18783 11904 18816 11938
rect 18850 11904 18884 11938
rect 18783 11848 18884 11904
rect 18783 11814 18816 11848
rect 18850 11814 18884 11848
rect 18783 11758 18884 11814
rect 18783 11724 18816 11758
rect 18850 11724 18884 11758
rect 18783 11668 18884 11724
rect 18783 11634 18816 11668
rect 18850 11634 18884 11668
rect 18783 11578 18884 11634
rect 18783 11544 18816 11578
rect 18850 11544 18884 11578
rect 18783 11488 18884 11544
rect 18783 11454 18816 11488
rect 18850 11454 18884 11488
rect 18783 11398 18884 11454
rect 18783 11364 18816 11398
rect 18850 11364 18884 11398
rect 18783 11308 18884 11364
rect 18783 11274 18816 11308
rect 18850 11274 18884 11308
rect 18783 11218 18884 11274
rect 18783 11184 18816 11218
rect 18850 11184 18884 11218
rect 18783 11128 18884 11184
rect 17495 11047 17697 11094
rect 18783 11094 18816 11128
rect 18850 11094 18884 11128
rect 18783 11047 18884 11094
rect 12444 11038 18884 11047
rect 12444 11004 12477 11038
rect 12511 11015 13664 11038
rect 12511 11004 12578 11015
rect 12444 10981 12578 11004
rect 12612 10981 12668 11015
rect 12702 10981 12758 11015
rect 12792 10981 12848 11015
rect 12882 10981 12938 11015
rect 12972 10981 13028 11015
rect 13062 10981 13118 11015
rect 13152 10981 13208 11015
rect 13242 10981 13298 11015
rect 13332 10981 13388 11015
rect 13422 10981 13478 11015
rect 13512 10981 13568 11015
rect 13602 11004 13664 11015
rect 13698 11004 13765 11038
rect 13799 11015 14952 11038
rect 13799 11004 13866 11015
rect 13602 10981 13866 11004
rect 13900 10981 13956 11015
rect 13990 10981 14046 11015
rect 14080 10981 14136 11015
rect 14170 10981 14226 11015
rect 14260 10981 14316 11015
rect 14350 10981 14406 11015
rect 14440 10981 14496 11015
rect 14530 10981 14586 11015
rect 14620 10981 14676 11015
rect 14710 10981 14766 11015
rect 14800 10981 14856 11015
rect 14890 11004 14952 11015
rect 14986 11004 15053 11038
rect 15087 11015 16240 11038
rect 15087 11004 15154 11015
rect 14890 10981 15154 11004
rect 15188 10981 15244 11015
rect 15278 10981 15334 11015
rect 15368 10981 15424 11015
rect 15458 10981 15514 11015
rect 15548 10981 15604 11015
rect 15638 10981 15694 11015
rect 15728 10981 15784 11015
rect 15818 10981 15874 11015
rect 15908 10981 15964 11015
rect 15998 10981 16054 11015
rect 16088 10981 16144 11015
rect 16178 11004 16240 11015
rect 16274 11004 16341 11038
rect 16375 11015 17528 11038
rect 16375 11004 16442 11015
rect 16178 10981 16442 11004
rect 16476 10981 16532 11015
rect 16566 10981 16622 11015
rect 16656 10981 16712 11015
rect 16746 10981 16802 11015
rect 16836 10981 16892 11015
rect 16926 10981 16982 11015
rect 17016 10981 17072 11015
rect 17106 10981 17162 11015
rect 17196 10981 17252 11015
rect 17286 10981 17342 11015
rect 17376 10981 17432 11015
rect 17466 11004 17528 11015
rect 17562 11004 17629 11038
rect 17663 11015 18816 11038
rect 17663 11004 17730 11015
rect 17466 10981 17730 11004
rect 17764 10981 17820 11015
rect 17854 10981 17910 11015
rect 17944 10981 18000 11015
rect 18034 10981 18090 11015
rect 18124 10981 18180 11015
rect 18214 10981 18270 11015
rect 18304 10981 18360 11015
rect 18394 10981 18450 11015
rect 18484 10981 18540 11015
rect 18574 10981 18630 11015
rect 18664 10981 18720 11015
rect 18754 11004 18816 11015
rect 18850 11004 18884 11038
rect 18754 10981 18884 11004
rect 12444 10914 18884 10981
rect 12444 10880 12578 10914
rect 12612 10880 12668 10914
rect 12702 10880 12758 10914
rect 12792 10880 12848 10914
rect 12882 10880 12938 10914
rect 12972 10880 13028 10914
rect 13062 10880 13118 10914
rect 13152 10880 13208 10914
rect 13242 10880 13298 10914
rect 13332 10880 13388 10914
rect 13422 10880 13478 10914
rect 13512 10880 13568 10914
rect 13602 10880 13866 10914
rect 13900 10880 13956 10914
rect 13990 10880 14046 10914
rect 14080 10880 14136 10914
rect 14170 10880 14226 10914
rect 14260 10880 14316 10914
rect 14350 10880 14406 10914
rect 14440 10880 14496 10914
rect 14530 10880 14586 10914
rect 14620 10880 14676 10914
rect 14710 10880 14766 10914
rect 14800 10880 14856 10914
rect 14890 10880 15154 10914
rect 15188 10880 15244 10914
rect 15278 10880 15334 10914
rect 15368 10880 15424 10914
rect 15458 10880 15514 10914
rect 15548 10880 15604 10914
rect 15638 10880 15694 10914
rect 15728 10880 15784 10914
rect 15818 10880 15874 10914
rect 15908 10880 15964 10914
rect 15998 10880 16054 10914
rect 16088 10880 16144 10914
rect 16178 10880 16442 10914
rect 16476 10880 16532 10914
rect 16566 10880 16622 10914
rect 16656 10880 16712 10914
rect 16746 10880 16802 10914
rect 16836 10880 16892 10914
rect 16926 10880 16982 10914
rect 17016 10880 17072 10914
rect 17106 10880 17162 10914
rect 17196 10880 17252 10914
rect 17286 10880 17342 10914
rect 17376 10880 17432 10914
rect 17466 10880 17730 10914
rect 17764 10880 17820 10914
rect 17854 10880 17910 10914
rect 17944 10880 18000 10914
rect 18034 10880 18090 10914
rect 18124 10880 18180 10914
rect 18214 10880 18270 10914
rect 18304 10880 18360 10914
rect 18394 10880 18450 10914
rect 18484 10880 18540 10914
rect 18574 10880 18630 10914
rect 18664 10880 18720 10914
rect 18754 10880 18884 10914
rect 12444 10845 18884 10880
rect 12444 10830 12545 10845
rect 12444 10796 12477 10830
rect 12511 10796 12545 10830
rect 12444 10740 12545 10796
rect 13631 10830 13833 10845
rect 13631 10796 13664 10830
rect 13698 10796 13765 10830
rect 13799 10796 13833 10830
rect 12444 10706 12477 10740
rect 12511 10706 12545 10740
rect 12444 10650 12545 10706
rect 12444 10616 12477 10650
rect 12511 10616 12545 10650
rect 12444 10560 12545 10616
rect 12444 10526 12477 10560
rect 12511 10526 12545 10560
rect 12444 10470 12545 10526
rect 12444 10436 12477 10470
rect 12511 10436 12545 10470
rect 12444 10380 12545 10436
rect 12444 10346 12477 10380
rect 12511 10346 12545 10380
rect 12444 10290 12545 10346
rect 12444 10256 12477 10290
rect 12511 10256 12545 10290
rect 12444 10200 12545 10256
rect 12444 10166 12477 10200
rect 12511 10166 12545 10200
rect 12444 10110 12545 10166
rect 12444 10076 12477 10110
rect 12511 10076 12545 10110
rect 12444 10020 12545 10076
rect 12444 9986 12477 10020
rect 12511 9986 12545 10020
rect 12444 9930 12545 9986
rect 12444 9896 12477 9930
rect 12511 9896 12545 9930
rect 12444 9840 12545 9896
rect 12444 9806 12477 9840
rect 12511 9806 12545 9840
rect 13631 10740 13833 10796
rect 14919 10830 15121 10845
rect 14919 10796 14952 10830
rect 14986 10796 15053 10830
rect 15087 10796 15121 10830
rect 13631 10706 13664 10740
rect 13698 10706 13765 10740
rect 13799 10706 13833 10740
rect 13631 10650 13833 10706
rect 13631 10616 13664 10650
rect 13698 10616 13765 10650
rect 13799 10616 13833 10650
rect 13631 10560 13833 10616
rect 13631 10526 13664 10560
rect 13698 10526 13765 10560
rect 13799 10526 13833 10560
rect 13631 10470 13833 10526
rect 13631 10436 13664 10470
rect 13698 10436 13765 10470
rect 13799 10436 13833 10470
rect 13631 10380 13833 10436
rect 13631 10346 13664 10380
rect 13698 10346 13765 10380
rect 13799 10346 13833 10380
rect 13631 10290 13833 10346
rect 13631 10256 13664 10290
rect 13698 10256 13765 10290
rect 13799 10256 13833 10290
rect 13631 10200 13833 10256
rect 13631 10166 13664 10200
rect 13698 10166 13765 10200
rect 13799 10166 13833 10200
rect 13631 10110 13833 10166
rect 13631 10076 13664 10110
rect 13698 10076 13765 10110
rect 13799 10076 13833 10110
rect 13631 10020 13833 10076
rect 13631 9986 13664 10020
rect 13698 9986 13765 10020
rect 13799 9986 13833 10020
rect 13631 9930 13833 9986
rect 13631 9896 13664 9930
rect 13698 9896 13765 9930
rect 13799 9896 13833 9930
rect 13631 9840 13833 9896
rect 12444 9759 12545 9806
rect 13631 9806 13664 9840
rect 13698 9806 13765 9840
rect 13799 9806 13833 9840
rect 14919 10740 15121 10796
rect 16207 10830 16409 10845
rect 16207 10796 16240 10830
rect 16274 10796 16341 10830
rect 16375 10796 16409 10830
rect 14919 10706 14952 10740
rect 14986 10706 15053 10740
rect 15087 10706 15121 10740
rect 14919 10650 15121 10706
rect 14919 10616 14952 10650
rect 14986 10616 15053 10650
rect 15087 10616 15121 10650
rect 14919 10560 15121 10616
rect 14919 10526 14952 10560
rect 14986 10526 15053 10560
rect 15087 10526 15121 10560
rect 14919 10470 15121 10526
rect 14919 10436 14952 10470
rect 14986 10436 15053 10470
rect 15087 10436 15121 10470
rect 14919 10380 15121 10436
rect 14919 10346 14952 10380
rect 14986 10346 15053 10380
rect 15087 10346 15121 10380
rect 14919 10290 15121 10346
rect 14919 10256 14952 10290
rect 14986 10256 15053 10290
rect 15087 10256 15121 10290
rect 14919 10200 15121 10256
rect 14919 10166 14952 10200
rect 14986 10166 15053 10200
rect 15087 10166 15121 10200
rect 14919 10110 15121 10166
rect 14919 10076 14952 10110
rect 14986 10076 15053 10110
rect 15087 10076 15121 10110
rect 14919 10020 15121 10076
rect 14919 9986 14952 10020
rect 14986 9986 15053 10020
rect 15087 9986 15121 10020
rect 14919 9930 15121 9986
rect 14919 9896 14952 9930
rect 14986 9896 15053 9930
rect 15087 9896 15121 9930
rect 14919 9840 15121 9896
rect 13631 9759 13833 9806
rect 14919 9806 14952 9840
rect 14986 9806 15053 9840
rect 15087 9806 15121 9840
rect 16207 10740 16409 10796
rect 17495 10830 17697 10845
rect 17495 10796 17528 10830
rect 17562 10796 17629 10830
rect 17663 10796 17697 10830
rect 16207 10706 16240 10740
rect 16274 10706 16341 10740
rect 16375 10706 16409 10740
rect 16207 10650 16409 10706
rect 16207 10616 16240 10650
rect 16274 10616 16341 10650
rect 16375 10616 16409 10650
rect 16207 10560 16409 10616
rect 16207 10526 16240 10560
rect 16274 10526 16341 10560
rect 16375 10526 16409 10560
rect 16207 10470 16409 10526
rect 16207 10436 16240 10470
rect 16274 10436 16341 10470
rect 16375 10436 16409 10470
rect 16207 10380 16409 10436
rect 16207 10346 16240 10380
rect 16274 10346 16341 10380
rect 16375 10346 16409 10380
rect 16207 10290 16409 10346
rect 16207 10256 16240 10290
rect 16274 10256 16341 10290
rect 16375 10256 16409 10290
rect 16207 10200 16409 10256
rect 16207 10166 16240 10200
rect 16274 10166 16341 10200
rect 16375 10166 16409 10200
rect 16207 10110 16409 10166
rect 16207 10076 16240 10110
rect 16274 10076 16341 10110
rect 16375 10076 16409 10110
rect 16207 10020 16409 10076
rect 16207 9986 16240 10020
rect 16274 9986 16341 10020
rect 16375 9986 16409 10020
rect 16207 9930 16409 9986
rect 16207 9896 16240 9930
rect 16274 9896 16341 9930
rect 16375 9896 16409 9930
rect 16207 9840 16409 9896
rect 14919 9759 15121 9806
rect 16207 9806 16240 9840
rect 16274 9806 16341 9840
rect 16375 9806 16409 9840
rect 17495 10740 17697 10796
rect 18783 10830 18884 10845
rect 18783 10796 18816 10830
rect 18850 10796 18884 10830
rect 17495 10706 17528 10740
rect 17562 10706 17629 10740
rect 17663 10706 17697 10740
rect 17495 10650 17697 10706
rect 17495 10616 17528 10650
rect 17562 10616 17629 10650
rect 17663 10616 17697 10650
rect 17495 10560 17697 10616
rect 17495 10526 17528 10560
rect 17562 10526 17629 10560
rect 17663 10526 17697 10560
rect 17495 10470 17697 10526
rect 17495 10436 17528 10470
rect 17562 10436 17629 10470
rect 17663 10436 17697 10470
rect 17495 10380 17697 10436
rect 17495 10346 17528 10380
rect 17562 10346 17629 10380
rect 17663 10346 17697 10380
rect 17495 10290 17697 10346
rect 17495 10256 17528 10290
rect 17562 10256 17629 10290
rect 17663 10256 17697 10290
rect 17495 10200 17697 10256
rect 17495 10166 17528 10200
rect 17562 10166 17629 10200
rect 17663 10166 17697 10200
rect 17495 10110 17697 10166
rect 17495 10076 17528 10110
rect 17562 10076 17629 10110
rect 17663 10076 17697 10110
rect 17495 10020 17697 10076
rect 17495 9986 17528 10020
rect 17562 9986 17629 10020
rect 17663 9986 17697 10020
rect 17495 9930 17697 9986
rect 17495 9896 17528 9930
rect 17562 9896 17629 9930
rect 17663 9896 17697 9930
rect 17495 9840 17697 9896
rect 16207 9759 16409 9806
rect 17495 9806 17528 9840
rect 17562 9806 17629 9840
rect 17663 9806 17697 9840
rect 18783 10740 18884 10796
rect 18783 10706 18816 10740
rect 18850 10706 18884 10740
rect 18783 10650 18884 10706
rect 18783 10616 18816 10650
rect 18850 10616 18884 10650
rect 18783 10560 18884 10616
rect 18783 10526 18816 10560
rect 18850 10526 18884 10560
rect 18783 10470 18884 10526
rect 18783 10436 18816 10470
rect 18850 10436 18884 10470
rect 18783 10380 18884 10436
rect 18783 10346 18816 10380
rect 18850 10346 18884 10380
rect 18783 10290 18884 10346
rect 18783 10256 18816 10290
rect 18850 10256 18884 10290
rect 18783 10200 18884 10256
rect 18783 10166 18816 10200
rect 18850 10166 18884 10200
rect 18783 10110 18884 10166
rect 18783 10076 18816 10110
rect 18850 10076 18884 10110
rect 18783 10020 18884 10076
rect 18783 9986 18816 10020
rect 18850 9986 18884 10020
rect 18783 9930 18884 9986
rect 18783 9896 18816 9930
rect 18850 9896 18884 9930
rect 18783 9840 18884 9896
rect 17495 9759 17697 9806
rect 18783 9806 18816 9840
rect 18850 9806 18884 9840
rect 18783 9759 18884 9806
rect 12444 9750 18884 9759
rect 12444 9716 12477 9750
rect 12511 9727 13664 9750
rect 12511 9716 12578 9727
rect 12444 9693 12578 9716
rect 12612 9693 12668 9727
rect 12702 9693 12758 9727
rect 12792 9693 12848 9727
rect 12882 9693 12938 9727
rect 12972 9693 13028 9727
rect 13062 9693 13118 9727
rect 13152 9693 13208 9727
rect 13242 9693 13298 9727
rect 13332 9693 13388 9727
rect 13422 9693 13478 9727
rect 13512 9693 13568 9727
rect 13602 9716 13664 9727
rect 13698 9716 13765 9750
rect 13799 9727 14952 9750
rect 13799 9716 13866 9727
rect 13602 9693 13866 9716
rect 13900 9693 13956 9727
rect 13990 9693 14046 9727
rect 14080 9693 14136 9727
rect 14170 9693 14226 9727
rect 14260 9693 14316 9727
rect 14350 9693 14406 9727
rect 14440 9693 14496 9727
rect 14530 9693 14586 9727
rect 14620 9693 14676 9727
rect 14710 9693 14766 9727
rect 14800 9693 14856 9727
rect 14890 9716 14952 9727
rect 14986 9716 15053 9750
rect 15087 9727 16240 9750
rect 15087 9716 15154 9727
rect 14890 9693 15154 9716
rect 15188 9693 15244 9727
rect 15278 9693 15334 9727
rect 15368 9693 15424 9727
rect 15458 9693 15514 9727
rect 15548 9693 15604 9727
rect 15638 9693 15694 9727
rect 15728 9693 15784 9727
rect 15818 9693 15874 9727
rect 15908 9693 15964 9727
rect 15998 9693 16054 9727
rect 16088 9693 16144 9727
rect 16178 9716 16240 9727
rect 16274 9716 16341 9750
rect 16375 9727 17528 9750
rect 16375 9716 16442 9727
rect 16178 9693 16442 9716
rect 16476 9693 16532 9727
rect 16566 9693 16622 9727
rect 16656 9693 16712 9727
rect 16746 9693 16802 9727
rect 16836 9693 16892 9727
rect 16926 9693 16982 9727
rect 17016 9693 17072 9727
rect 17106 9693 17162 9727
rect 17196 9693 17252 9727
rect 17286 9693 17342 9727
rect 17376 9693 17432 9727
rect 17466 9716 17528 9727
rect 17562 9716 17629 9750
rect 17663 9727 18816 9750
rect 17663 9716 17730 9727
rect 17466 9693 17730 9716
rect 17764 9693 17820 9727
rect 17854 9693 17910 9727
rect 17944 9693 18000 9727
rect 18034 9693 18090 9727
rect 18124 9693 18180 9727
rect 18214 9693 18270 9727
rect 18304 9693 18360 9727
rect 18394 9693 18450 9727
rect 18484 9693 18540 9727
rect 18574 9693 18630 9727
rect 18664 9693 18720 9727
rect 18754 9716 18816 9727
rect 18850 9716 18884 9750
rect 18754 9693 18884 9716
rect 12444 9626 18884 9693
rect 12444 9592 12578 9626
rect 12612 9592 12668 9626
rect 12702 9592 12758 9626
rect 12792 9592 12848 9626
rect 12882 9592 12938 9626
rect 12972 9592 13028 9626
rect 13062 9592 13118 9626
rect 13152 9592 13208 9626
rect 13242 9592 13298 9626
rect 13332 9592 13388 9626
rect 13422 9592 13478 9626
rect 13512 9592 13568 9626
rect 13602 9592 13866 9626
rect 13900 9592 13956 9626
rect 13990 9592 14046 9626
rect 14080 9592 14136 9626
rect 14170 9592 14226 9626
rect 14260 9592 14316 9626
rect 14350 9592 14406 9626
rect 14440 9592 14496 9626
rect 14530 9592 14586 9626
rect 14620 9592 14676 9626
rect 14710 9592 14766 9626
rect 14800 9592 14856 9626
rect 14890 9592 15154 9626
rect 15188 9592 15244 9626
rect 15278 9592 15334 9626
rect 15368 9592 15424 9626
rect 15458 9592 15514 9626
rect 15548 9592 15604 9626
rect 15638 9592 15694 9626
rect 15728 9592 15784 9626
rect 15818 9592 15874 9626
rect 15908 9592 15964 9626
rect 15998 9592 16054 9626
rect 16088 9592 16144 9626
rect 16178 9592 16442 9626
rect 16476 9592 16532 9626
rect 16566 9592 16622 9626
rect 16656 9592 16712 9626
rect 16746 9592 16802 9626
rect 16836 9592 16892 9626
rect 16926 9592 16982 9626
rect 17016 9592 17072 9626
rect 17106 9592 17162 9626
rect 17196 9592 17252 9626
rect 17286 9592 17342 9626
rect 17376 9592 17432 9626
rect 17466 9592 17730 9626
rect 17764 9592 17820 9626
rect 17854 9592 17910 9626
rect 17944 9592 18000 9626
rect 18034 9592 18090 9626
rect 18124 9592 18180 9626
rect 18214 9592 18270 9626
rect 18304 9592 18360 9626
rect 18394 9592 18450 9626
rect 18484 9592 18540 9626
rect 18574 9592 18630 9626
rect 18664 9592 18720 9626
rect 18754 9592 18884 9626
rect 12444 9557 18884 9592
rect 12444 9542 12545 9557
rect 12444 9508 12477 9542
rect 12511 9508 12545 9542
rect 12444 9452 12545 9508
rect 13631 9542 13833 9557
rect 13631 9508 13664 9542
rect 13698 9508 13765 9542
rect 13799 9508 13833 9542
rect -17906 9382 -11406 9406
rect -17906 9050 -17882 9382
rect -11430 9050 -11406 9382
rect -17906 9026 -11406 9050
rect -17484 6642 -17284 6742
rect -22332 5836 -18512 5860
rect -22332 5760 -20918 5836
rect -19926 5760 -18512 5836
rect -22332 5736 -18512 5760
rect -22328 5682 -21880 5736
rect -22328 5106 -22304 5682
rect -21904 5106 -21880 5682
rect -18962 5682 -18514 5736
rect -18962 5106 -18938 5682
rect -18538 5106 -18514 5682
rect -22328 5082 -21880 5106
rect -18962 5082 -18514 5106
rect -17484 5042 -17434 6642
rect -17334 5042 -17284 6642
rect -17484 4942 -17284 5042
rect -11984 6642 -11784 6742
rect -11984 5042 -11934 6642
rect -11834 5042 -11784 6642
rect -11984 4942 -11784 5042
rect 12444 9418 12477 9452
rect 12511 9418 12545 9452
rect 12444 9362 12545 9418
rect 12444 9328 12477 9362
rect 12511 9328 12545 9362
rect 12444 9272 12545 9328
rect 12444 9238 12477 9272
rect 12511 9238 12545 9272
rect 12444 9182 12545 9238
rect 12444 9148 12477 9182
rect 12511 9148 12545 9182
rect 12444 9092 12545 9148
rect 12444 9058 12477 9092
rect 12511 9058 12545 9092
rect 12444 9002 12545 9058
rect 12444 8968 12477 9002
rect 12511 8968 12545 9002
rect 12444 8912 12545 8968
rect 12444 8878 12477 8912
rect 12511 8878 12545 8912
rect 12444 8822 12545 8878
rect 12444 8788 12477 8822
rect 12511 8788 12545 8822
rect 12444 8732 12545 8788
rect 12444 8698 12477 8732
rect 12511 8698 12545 8732
rect 12444 8642 12545 8698
rect 12444 8608 12477 8642
rect 12511 8608 12545 8642
rect 12444 8552 12545 8608
rect 12444 8518 12477 8552
rect 12511 8518 12545 8552
rect 13631 9452 13833 9508
rect 14919 9542 15121 9557
rect 14919 9508 14952 9542
rect 14986 9508 15053 9542
rect 15087 9508 15121 9542
rect 13631 9418 13664 9452
rect 13698 9418 13765 9452
rect 13799 9418 13833 9452
rect 13631 9362 13833 9418
rect 13631 9328 13664 9362
rect 13698 9328 13765 9362
rect 13799 9328 13833 9362
rect 13631 9272 13833 9328
rect 13631 9238 13664 9272
rect 13698 9238 13765 9272
rect 13799 9238 13833 9272
rect 13631 9182 13833 9238
rect 13631 9148 13664 9182
rect 13698 9148 13765 9182
rect 13799 9148 13833 9182
rect 13631 9092 13833 9148
rect 13631 9058 13664 9092
rect 13698 9058 13765 9092
rect 13799 9058 13833 9092
rect 13631 9002 13833 9058
rect 13631 8968 13664 9002
rect 13698 8968 13765 9002
rect 13799 8968 13833 9002
rect 13631 8912 13833 8968
rect 13631 8878 13664 8912
rect 13698 8878 13765 8912
rect 13799 8878 13833 8912
rect 13631 8822 13833 8878
rect 13631 8788 13664 8822
rect 13698 8788 13765 8822
rect 13799 8788 13833 8822
rect 13631 8732 13833 8788
rect 13631 8698 13664 8732
rect 13698 8698 13765 8732
rect 13799 8698 13833 8732
rect 13631 8642 13833 8698
rect 13631 8608 13664 8642
rect 13698 8608 13765 8642
rect 13799 8608 13833 8642
rect 13631 8552 13833 8608
rect 12444 8471 12545 8518
rect 13631 8518 13664 8552
rect 13698 8518 13765 8552
rect 13799 8518 13833 8552
rect 14919 9452 15121 9508
rect 16207 9542 16409 9557
rect 16207 9508 16240 9542
rect 16274 9508 16341 9542
rect 16375 9508 16409 9542
rect 14919 9418 14952 9452
rect 14986 9418 15053 9452
rect 15087 9418 15121 9452
rect 14919 9362 15121 9418
rect 14919 9328 14952 9362
rect 14986 9328 15053 9362
rect 15087 9328 15121 9362
rect 14919 9272 15121 9328
rect 14919 9238 14952 9272
rect 14986 9238 15053 9272
rect 15087 9238 15121 9272
rect 14919 9182 15121 9238
rect 14919 9148 14952 9182
rect 14986 9148 15053 9182
rect 15087 9148 15121 9182
rect 14919 9092 15121 9148
rect 14919 9058 14952 9092
rect 14986 9058 15053 9092
rect 15087 9058 15121 9092
rect 14919 9002 15121 9058
rect 14919 8968 14952 9002
rect 14986 8968 15053 9002
rect 15087 8968 15121 9002
rect 14919 8912 15121 8968
rect 14919 8878 14952 8912
rect 14986 8878 15053 8912
rect 15087 8878 15121 8912
rect 14919 8822 15121 8878
rect 14919 8788 14952 8822
rect 14986 8788 15053 8822
rect 15087 8788 15121 8822
rect 14919 8732 15121 8788
rect 14919 8698 14952 8732
rect 14986 8698 15053 8732
rect 15087 8698 15121 8732
rect 14919 8642 15121 8698
rect 14919 8608 14952 8642
rect 14986 8608 15053 8642
rect 15087 8608 15121 8642
rect 14919 8552 15121 8608
rect 13631 8471 13833 8518
rect 14919 8518 14952 8552
rect 14986 8518 15053 8552
rect 15087 8518 15121 8552
rect 16207 9452 16409 9508
rect 17495 9542 17697 9557
rect 17495 9508 17528 9542
rect 17562 9508 17629 9542
rect 17663 9508 17697 9542
rect 16207 9418 16240 9452
rect 16274 9418 16341 9452
rect 16375 9418 16409 9452
rect 16207 9362 16409 9418
rect 16207 9328 16240 9362
rect 16274 9328 16341 9362
rect 16375 9328 16409 9362
rect 16207 9272 16409 9328
rect 16207 9238 16240 9272
rect 16274 9238 16341 9272
rect 16375 9238 16409 9272
rect 16207 9182 16409 9238
rect 16207 9148 16240 9182
rect 16274 9148 16341 9182
rect 16375 9148 16409 9182
rect 16207 9092 16409 9148
rect 16207 9058 16240 9092
rect 16274 9058 16341 9092
rect 16375 9058 16409 9092
rect 16207 9002 16409 9058
rect 16207 8968 16240 9002
rect 16274 8968 16341 9002
rect 16375 8968 16409 9002
rect 16207 8912 16409 8968
rect 16207 8878 16240 8912
rect 16274 8878 16341 8912
rect 16375 8878 16409 8912
rect 16207 8822 16409 8878
rect 16207 8788 16240 8822
rect 16274 8788 16341 8822
rect 16375 8788 16409 8822
rect 16207 8732 16409 8788
rect 16207 8698 16240 8732
rect 16274 8698 16341 8732
rect 16375 8698 16409 8732
rect 16207 8642 16409 8698
rect 16207 8608 16240 8642
rect 16274 8608 16341 8642
rect 16375 8608 16409 8642
rect 16207 8552 16409 8608
rect 14919 8471 15121 8518
rect 16207 8518 16240 8552
rect 16274 8518 16341 8552
rect 16375 8518 16409 8552
rect 17495 9452 17697 9508
rect 18783 9542 18884 9557
rect 18783 9508 18816 9542
rect 18850 9508 18884 9542
rect 17495 9418 17528 9452
rect 17562 9418 17629 9452
rect 17663 9418 17697 9452
rect 17495 9362 17697 9418
rect 17495 9328 17528 9362
rect 17562 9328 17629 9362
rect 17663 9328 17697 9362
rect 17495 9272 17697 9328
rect 17495 9238 17528 9272
rect 17562 9238 17629 9272
rect 17663 9238 17697 9272
rect 17495 9182 17697 9238
rect 17495 9148 17528 9182
rect 17562 9148 17629 9182
rect 17663 9148 17697 9182
rect 17495 9092 17697 9148
rect 17495 9058 17528 9092
rect 17562 9058 17629 9092
rect 17663 9058 17697 9092
rect 17495 9002 17697 9058
rect 17495 8968 17528 9002
rect 17562 8968 17629 9002
rect 17663 8968 17697 9002
rect 17495 8912 17697 8968
rect 17495 8878 17528 8912
rect 17562 8878 17629 8912
rect 17663 8878 17697 8912
rect 17495 8822 17697 8878
rect 17495 8788 17528 8822
rect 17562 8788 17629 8822
rect 17663 8788 17697 8822
rect 17495 8732 17697 8788
rect 17495 8698 17528 8732
rect 17562 8698 17629 8732
rect 17663 8698 17697 8732
rect 17495 8642 17697 8698
rect 17495 8608 17528 8642
rect 17562 8608 17629 8642
rect 17663 8608 17697 8642
rect 17495 8552 17697 8608
rect 16207 8471 16409 8518
rect 17495 8518 17528 8552
rect 17562 8518 17629 8552
rect 17663 8518 17697 8552
rect 18783 9452 18884 9508
rect 18783 9418 18816 9452
rect 18850 9418 18884 9452
rect 18783 9362 18884 9418
rect 18783 9328 18816 9362
rect 18850 9328 18884 9362
rect 18783 9272 18884 9328
rect 18783 9238 18816 9272
rect 18850 9238 18884 9272
rect 18783 9182 18884 9238
rect 18783 9148 18816 9182
rect 18850 9148 18884 9182
rect 18783 9092 18884 9148
rect 18783 9058 18816 9092
rect 18850 9058 18884 9092
rect 18783 9002 18884 9058
rect 18783 8968 18816 9002
rect 18850 8968 18884 9002
rect 18783 8912 18884 8968
rect 18783 8878 18816 8912
rect 18850 8878 18884 8912
rect 18783 8822 18884 8878
rect 18783 8788 18816 8822
rect 18850 8788 18884 8822
rect 18783 8732 18884 8788
rect 18783 8698 18816 8732
rect 18850 8698 18884 8732
rect 18783 8642 18884 8698
rect 18783 8608 18816 8642
rect 18850 8608 18884 8642
rect 18783 8552 18884 8608
rect 17495 8471 17697 8518
rect 18783 8518 18816 8552
rect 18850 8518 18884 8552
rect 18783 8471 18884 8518
rect 12444 8462 18884 8471
rect 12444 8428 12477 8462
rect 12511 8439 13664 8462
rect 12511 8428 12578 8439
rect 12444 8405 12578 8428
rect 12612 8405 12668 8439
rect 12702 8405 12758 8439
rect 12792 8405 12848 8439
rect 12882 8405 12938 8439
rect 12972 8405 13028 8439
rect 13062 8405 13118 8439
rect 13152 8405 13208 8439
rect 13242 8405 13298 8439
rect 13332 8405 13388 8439
rect 13422 8405 13478 8439
rect 13512 8405 13568 8439
rect 13602 8428 13664 8439
rect 13698 8428 13765 8462
rect 13799 8439 14952 8462
rect 13799 8428 13866 8439
rect 13602 8405 13866 8428
rect 13900 8405 13956 8439
rect 13990 8405 14046 8439
rect 14080 8405 14136 8439
rect 14170 8405 14226 8439
rect 14260 8405 14316 8439
rect 14350 8405 14406 8439
rect 14440 8405 14496 8439
rect 14530 8405 14586 8439
rect 14620 8405 14676 8439
rect 14710 8405 14766 8439
rect 14800 8405 14856 8439
rect 14890 8428 14952 8439
rect 14986 8428 15053 8462
rect 15087 8439 16240 8462
rect 15087 8428 15154 8439
rect 14890 8405 15154 8428
rect 15188 8405 15244 8439
rect 15278 8405 15334 8439
rect 15368 8405 15424 8439
rect 15458 8405 15514 8439
rect 15548 8405 15604 8439
rect 15638 8405 15694 8439
rect 15728 8405 15784 8439
rect 15818 8405 15874 8439
rect 15908 8405 15964 8439
rect 15998 8405 16054 8439
rect 16088 8405 16144 8439
rect 16178 8428 16240 8439
rect 16274 8428 16341 8462
rect 16375 8439 17528 8462
rect 16375 8428 16442 8439
rect 16178 8405 16442 8428
rect 16476 8405 16532 8439
rect 16566 8405 16622 8439
rect 16656 8405 16712 8439
rect 16746 8405 16802 8439
rect 16836 8405 16892 8439
rect 16926 8405 16982 8439
rect 17016 8405 17072 8439
rect 17106 8405 17162 8439
rect 17196 8405 17252 8439
rect 17286 8405 17342 8439
rect 17376 8405 17432 8439
rect 17466 8428 17528 8439
rect 17562 8428 17629 8462
rect 17663 8439 18816 8462
rect 17663 8428 17730 8439
rect 17466 8405 17730 8428
rect 17764 8405 17820 8439
rect 17854 8405 17910 8439
rect 17944 8405 18000 8439
rect 18034 8405 18090 8439
rect 18124 8405 18180 8439
rect 18214 8405 18270 8439
rect 18304 8405 18360 8439
rect 18394 8405 18450 8439
rect 18484 8405 18540 8439
rect 18574 8405 18630 8439
rect 18664 8405 18720 8439
rect 18754 8428 18816 8439
rect 18850 8428 18884 8462
rect 18754 8405 18884 8428
rect 12444 8338 18884 8405
rect 12444 8304 12578 8338
rect 12612 8304 12668 8338
rect 12702 8304 12758 8338
rect 12792 8304 12848 8338
rect 12882 8304 12938 8338
rect 12972 8304 13028 8338
rect 13062 8304 13118 8338
rect 13152 8304 13208 8338
rect 13242 8304 13298 8338
rect 13332 8304 13388 8338
rect 13422 8304 13478 8338
rect 13512 8304 13568 8338
rect 13602 8304 13866 8338
rect 13900 8304 13956 8338
rect 13990 8304 14046 8338
rect 14080 8304 14136 8338
rect 14170 8304 14226 8338
rect 14260 8304 14316 8338
rect 14350 8304 14406 8338
rect 14440 8304 14496 8338
rect 14530 8304 14586 8338
rect 14620 8304 14676 8338
rect 14710 8304 14766 8338
rect 14800 8304 14856 8338
rect 14890 8304 15154 8338
rect 15188 8304 15244 8338
rect 15278 8304 15334 8338
rect 15368 8304 15424 8338
rect 15458 8304 15514 8338
rect 15548 8304 15604 8338
rect 15638 8304 15694 8338
rect 15728 8304 15784 8338
rect 15818 8304 15874 8338
rect 15908 8304 15964 8338
rect 15998 8304 16054 8338
rect 16088 8304 16144 8338
rect 16178 8304 16442 8338
rect 16476 8304 16532 8338
rect 16566 8304 16622 8338
rect 16656 8304 16712 8338
rect 16746 8304 16802 8338
rect 16836 8304 16892 8338
rect 16926 8304 16982 8338
rect 17016 8304 17072 8338
rect 17106 8304 17162 8338
rect 17196 8304 17252 8338
rect 17286 8304 17342 8338
rect 17376 8304 17432 8338
rect 17466 8304 17730 8338
rect 17764 8304 17820 8338
rect 17854 8304 17910 8338
rect 17944 8304 18000 8338
rect 18034 8304 18090 8338
rect 18124 8304 18180 8338
rect 18214 8304 18270 8338
rect 18304 8304 18360 8338
rect 18394 8304 18450 8338
rect 18484 8304 18540 8338
rect 18574 8304 18630 8338
rect 18664 8304 18720 8338
rect 18754 8304 18884 8338
rect 12444 8269 18884 8304
rect 12444 8254 12545 8269
rect 12444 8220 12477 8254
rect 12511 8220 12545 8254
rect 12444 8164 12545 8220
rect 13631 8254 13833 8269
rect 13631 8220 13664 8254
rect 13698 8220 13765 8254
rect 13799 8220 13833 8254
rect 12444 8130 12477 8164
rect 12511 8130 12545 8164
rect 12444 8074 12545 8130
rect 12444 8040 12477 8074
rect 12511 8040 12545 8074
rect 12444 7984 12545 8040
rect 12444 7950 12477 7984
rect 12511 7950 12545 7984
rect 12444 7894 12545 7950
rect 12444 7860 12477 7894
rect 12511 7860 12545 7894
rect 12444 7804 12545 7860
rect 12444 7770 12477 7804
rect 12511 7770 12545 7804
rect 12444 7714 12545 7770
rect 12444 7680 12477 7714
rect 12511 7680 12545 7714
rect 12444 7624 12545 7680
rect 12444 7590 12477 7624
rect 12511 7590 12545 7624
rect 12444 7534 12545 7590
rect 12444 7500 12477 7534
rect 12511 7500 12545 7534
rect 12444 7444 12545 7500
rect 12444 7410 12477 7444
rect 12511 7410 12545 7444
rect 12444 7354 12545 7410
rect 12444 7320 12477 7354
rect 12511 7320 12545 7354
rect 12444 7264 12545 7320
rect 12444 7230 12477 7264
rect 12511 7230 12545 7264
rect 13631 8164 13833 8220
rect 14919 8254 15121 8269
rect 14919 8220 14952 8254
rect 14986 8220 15053 8254
rect 15087 8220 15121 8254
rect 13631 8130 13664 8164
rect 13698 8130 13765 8164
rect 13799 8130 13833 8164
rect 13631 8074 13833 8130
rect 13631 8040 13664 8074
rect 13698 8040 13765 8074
rect 13799 8040 13833 8074
rect 13631 7984 13833 8040
rect 13631 7950 13664 7984
rect 13698 7950 13765 7984
rect 13799 7950 13833 7984
rect 13631 7894 13833 7950
rect 13631 7860 13664 7894
rect 13698 7860 13765 7894
rect 13799 7860 13833 7894
rect 13631 7804 13833 7860
rect 13631 7770 13664 7804
rect 13698 7770 13765 7804
rect 13799 7770 13833 7804
rect 13631 7714 13833 7770
rect 13631 7680 13664 7714
rect 13698 7680 13765 7714
rect 13799 7680 13833 7714
rect 13631 7624 13833 7680
rect 13631 7590 13664 7624
rect 13698 7590 13765 7624
rect 13799 7590 13833 7624
rect 13631 7534 13833 7590
rect 13631 7500 13664 7534
rect 13698 7500 13765 7534
rect 13799 7500 13833 7534
rect 13631 7444 13833 7500
rect 13631 7410 13664 7444
rect 13698 7410 13765 7444
rect 13799 7410 13833 7444
rect 13631 7354 13833 7410
rect 13631 7320 13664 7354
rect 13698 7320 13765 7354
rect 13799 7320 13833 7354
rect 13631 7264 13833 7320
rect 12444 7183 12545 7230
rect 13631 7230 13664 7264
rect 13698 7230 13765 7264
rect 13799 7230 13833 7264
rect 14919 8164 15121 8220
rect 16207 8254 16409 8269
rect 16207 8220 16240 8254
rect 16274 8220 16341 8254
rect 16375 8220 16409 8254
rect 14919 8130 14952 8164
rect 14986 8130 15053 8164
rect 15087 8130 15121 8164
rect 14919 8074 15121 8130
rect 14919 8040 14952 8074
rect 14986 8040 15053 8074
rect 15087 8040 15121 8074
rect 14919 7984 15121 8040
rect 14919 7950 14952 7984
rect 14986 7950 15053 7984
rect 15087 7950 15121 7984
rect 14919 7894 15121 7950
rect 14919 7860 14952 7894
rect 14986 7860 15053 7894
rect 15087 7860 15121 7894
rect 14919 7804 15121 7860
rect 14919 7770 14952 7804
rect 14986 7770 15053 7804
rect 15087 7770 15121 7804
rect 14919 7714 15121 7770
rect 14919 7680 14952 7714
rect 14986 7680 15053 7714
rect 15087 7680 15121 7714
rect 14919 7624 15121 7680
rect 14919 7590 14952 7624
rect 14986 7590 15053 7624
rect 15087 7590 15121 7624
rect 14919 7534 15121 7590
rect 14919 7500 14952 7534
rect 14986 7500 15053 7534
rect 15087 7500 15121 7534
rect 14919 7444 15121 7500
rect 14919 7410 14952 7444
rect 14986 7410 15053 7444
rect 15087 7410 15121 7444
rect 14919 7354 15121 7410
rect 14919 7320 14952 7354
rect 14986 7320 15053 7354
rect 15087 7320 15121 7354
rect 14919 7264 15121 7320
rect 13631 7183 13833 7230
rect 14919 7230 14952 7264
rect 14986 7230 15053 7264
rect 15087 7230 15121 7264
rect 16207 8164 16409 8220
rect 17495 8254 17697 8269
rect 17495 8220 17528 8254
rect 17562 8220 17629 8254
rect 17663 8220 17697 8254
rect 16207 8130 16240 8164
rect 16274 8130 16341 8164
rect 16375 8130 16409 8164
rect 16207 8074 16409 8130
rect 16207 8040 16240 8074
rect 16274 8040 16341 8074
rect 16375 8040 16409 8074
rect 16207 7984 16409 8040
rect 16207 7950 16240 7984
rect 16274 7950 16341 7984
rect 16375 7950 16409 7984
rect 16207 7894 16409 7950
rect 16207 7860 16240 7894
rect 16274 7860 16341 7894
rect 16375 7860 16409 7894
rect 16207 7804 16409 7860
rect 16207 7770 16240 7804
rect 16274 7770 16341 7804
rect 16375 7770 16409 7804
rect 16207 7714 16409 7770
rect 16207 7680 16240 7714
rect 16274 7680 16341 7714
rect 16375 7680 16409 7714
rect 16207 7624 16409 7680
rect 16207 7590 16240 7624
rect 16274 7590 16341 7624
rect 16375 7590 16409 7624
rect 16207 7534 16409 7590
rect 16207 7500 16240 7534
rect 16274 7500 16341 7534
rect 16375 7500 16409 7534
rect 16207 7444 16409 7500
rect 16207 7410 16240 7444
rect 16274 7410 16341 7444
rect 16375 7410 16409 7444
rect 16207 7354 16409 7410
rect 16207 7320 16240 7354
rect 16274 7320 16341 7354
rect 16375 7320 16409 7354
rect 16207 7264 16409 7320
rect 14919 7183 15121 7230
rect 16207 7230 16240 7264
rect 16274 7230 16341 7264
rect 16375 7230 16409 7264
rect 17495 8164 17697 8220
rect 18783 8254 18884 8269
rect 18783 8220 18816 8254
rect 18850 8220 18884 8254
rect 17495 8130 17528 8164
rect 17562 8130 17629 8164
rect 17663 8130 17697 8164
rect 17495 8074 17697 8130
rect 17495 8040 17528 8074
rect 17562 8040 17629 8074
rect 17663 8040 17697 8074
rect 17495 7984 17697 8040
rect 17495 7950 17528 7984
rect 17562 7950 17629 7984
rect 17663 7950 17697 7984
rect 17495 7894 17697 7950
rect 17495 7860 17528 7894
rect 17562 7860 17629 7894
rect 17663 7860 17697 7894
rect 17495 7804 17697 7860
rect 17495 7770 17528 7804
rect 17562 7770 17629 7804
rect 17663 7770 17697 7804
rect 17495 7714 17697 7770
rect 17495 7680 17528 7714
rect 17562 7680 17629 7714
rect 17663 7680 17697 7714
rect 17495 7624 17697 7680
rect 17495 7590 17528 7624
rect 17562 7590 17629 7624
rect 17663 7590 17697 7624
rect 17495 7534 17697 7590
rect 17495 7500 17528 7534
rect 17562 7500 17629 7534
rect 17663 7500 17697 7534
rect 17495 7444 17697 7500
rect 17495 7410 17528 7444
rect 17562 7410 17629 7444
rect 17663 7410 17697 7444
rect 17495 7354 17697 7410
rect 17495 7320 17528 7354
rect 17562 7320 17629 7354
rect 17663 7320 17697 7354
rect 17495 7264 17697 7320
rect 16207 7183 16409 7230
rect 17495 7230 17528 7264
rect 17562 7230 17629 7264
rect 17663 7230 17697 7264
rect 18783 8164 18884 8220
rect 18783 8130 18816 8164
rect 18850 8130 18884 8164
rect 18783 8074 18884 8130
rect 18783 8040 18816 8074
rect 18850 8040 18884 8074
rect 18783 7984 18884 8040
rect 18783 7950 18816 7984
rect 18850 7950 18884 7984
rect 18783 7894 18884 7950
rect 18783 7860 18816 7894
rect 18850 7860 18884 7894
rect 18783 7804 18884 7860
rect 18783 7770 18816 7804
rect 18850 7770 18884 7804
rect 18783 7714 18884 7770
rect 18783 7680 18816 7714
rect 18850 7680 18884 7714
rect 18783 7624 18884 7680
rect 18783 7590 18816 7624
rect 18850 7590 18884 7624
rect 18783 7534 18884 7590
rect 18783 7500 18816 7534
rect 18850 7500 18884 7534
rect 18783 7444 18884 7500
rect 18783 7410 18816 7444
rect 18850 7410 18884 7444
rect 18783 7354 18884 7410
rect 18783 7320 18816 7354
rect 18850 7320 18884 7354
rect 18783 7264 18884 7320
rect 17495 7183 17697 7230
rect 18783 7230 18816 7264
rect 18850 7230 18884 7264
rect 18783 7183 18884 7230
rect 12444 7174 18884 7183
rect 12444 7140 12477 7174
rect 12511 7151 13664 7174
rect 12511 7140 12578 7151
rect 12444 7117 12578 7140
rect 12612 7117 12668 7151
rect 12702 7117 12758 7151
rect 12792 7117 12848 7151
rect 12882 7117 12938 7151
rect 12972 7117 13028 7151
rect 13062 7117 13118 7151
rect 13152 7117 13208 7151
rect 13242 7117 13298 7151
rect 13332 7117 13388 7151
rect 13422 7117 13478 7151
rect 13512 7117 13568 7151
rect 13602 7140 13664 7151
rect 13698 7140 13765 7174
rect 13799 7151 14952 7174
rect 13799 7140 13866 7151
rect 13602 7117 13866 7140
rect 13900 7117 13956 7151
rect 13990 7117 14046 7151
rect 14080 7117 14136 7151
rect 14170 7117 14226 7151
rect 14260 7117 14316 7151
rect 14350 7117 14406 7151
rect 14440 7117 14496 7151
rect 14530 7117 14586 7151
rect 14620 7117 14676 7151
rect 14710 7117 14766 7151
rect 14800 7117 14856 7151
rect 14890 7140 14952 7151
rect 14986 7140 15053 7174
rect 15087 7151 16240 7174
rect 15087 7140 15154 7151
rect 14890 7117 15154 7140
rect 15188 7117 15244 7151
rect 15278 7117 15334 7151
rect 15368 7117 15424 7151
rect 15458 7117 15514 7151
rect 15548 7117 15604 7151
rect 15638 7117 15694 7151
rect 15728 7117 15784 7151
rect 15818 7117 15874 7151
rect 15908 7117 15964 7151
rect 15998 7117 16054 7151
rect 16088 7117 16144 7151
rect 16178 7140 16240 7151
rect 16274 7140 16341 7174
rect 16375 7151 17528 7174
rect 16375 7140 16442 7151
rect 16178 7117 16442 7140
rect 16476 7117 16532 7151
rect 16566 7117 16622 7151
rect 16656 7117 16712 7151
rect 16746 7117 16802 7151
rect 16836 7117 16892 7151
rect 16926 7117 16982 7151
rect 17016 7117 17072 7151
rect 17106 7117 17162 7151
rect 17196 7117 17252 7151
rect 17286 7117 17342 7151
rect 17376 7117 17432 7151
rect 17466 7140 17528 7151
rect 17562 7140 17629 7174
rect 17663 7151 18816 7174
rect 17663 7140 17730 7151
rect 17466 7117 17730 7140
rect 17764 7117 17820 7151
rect 17854 7117 17910 7151
rect 17944 7117 18000 7151
rect 18034 7117 18090 7151
rect 18124 7117 18180 7151
rect 18214 7117 18270 7151
rect 18304 7117 18360 7151
rect 18394 7117 18450 7151
rect 18484 7117 18540 7151
rect 18574 7117 18630 7151
rect 18664 7117 18720 7151
rect 18754 7140 18816 7151
rect 18850 7140 18884 7174
rect 18754 7117 18884 7140
rect 12444 7050 18884 7117
rect 12444 7016 12578 7050
rect 12612 7016 12668 7050
rect 12702 7016 12758 7050
rect 12792 7016 12848 7050
rect 12882 7016 12938 7050
rect 12972 7016 13028 7050
rect 13062 7016 13118 7050
rect 13152 7016 13208 7050
rect 13242 7016 13298 7050
rect 13332 7016 13388 7050
rect 13422 7016 13478 7050
rect 13512 7016 13568 7050
rect 13602 7016 13866 7050
rect 13900 7016 13956 7050
rect 13990 7016 14046 7050
rect 14080 7016 14136 7050
rect 14170 7016 14226 7050
rect 14260 7016 14316 7050
rect 14350 7016 14406 7050
rect 14440 7016 14496 7050
rect 14530 7016 14586 7050
rect 14620 7016 14676 7050
rect 14710 7016 14766 7050
rect 14800 7016 14856 7050
rect 14890 7016 15154 7050
rect 15188 7016 15244 7050
rect 15278 7016 15334 7050
rect 15368 7016 15424 7050
rect 15458 7016 15514 7050
rect 15548 7016 15604 7050
rect 15638 7016 15694 7050
rect 15728 7016 15784 7050
rect 15818 7016 15874 7050
rect 15908 7016 15964 7050
rect 15998 7016 16054 7050
rect 16088 7016 16144 7050
rect 16178 7016 16442 7050
rect 16476 7016 16532 7050
rect 16566 7016 16622 7050
rect 16656 7016 16712 7050
rect 16746 7016 16802 7050
rect 16836 7016 16892 7050
rect 16926 7016 16982 7050
rect 17016 7016 17072 7050
rect 17106 7016 17162 7050
rect 17196 7016 17252 7050
rect 17286 7016 17342 7050
rect 17376 7016 17432 7050
rect 17466 7016 17730 7050
rect 17764 7016 17820 7050
rect 17854 7016 17910 7050
rect 17944 7016 18000 7050
rect 18034 7016 18090 7050
rect 18124 7016 18180 7050
rect 18214 7016 18270 7050
rect 18304 7016 18360 7050
rect 18394 7016 18450 7050
rect 18484 7016 18540 7050
rect 18574 7016 18630 7050
rect 18664 7016 18720 7050
rect 18754 7016 18884 7050
rect 12444 6981 18884 7016
rect 12444 6966 12545 6981
rect 12444 6932 12477 6966
rect 12511 6932 12545 6966
rect 12444 6876 12545 6932
rect 13631 6966 13833 6981
rect 13631 6932 13664 6966
rect 13698 6932 13765 6966
rect 13799 6932 13833 6966
rect 12444 6842 12477 6876
rect 12511 6842 12545 6876
rect 12444 6786 12545 6842
rect 12444 6752 12477 6786
rect 12511 6752 12545 6786
rect 12444 6696 12545 6752
rect 12444 6662 12477 6696
rect 12511 6662 12545 6696
rect 12444 6606 12545 6662
rect 12444 6572 12477 6606
rect 12511 6572 12545 6606
rect 12444 6516 12545 6572
rect 12444 6482 12477 6516
rect 12511 6482 12545 6516
rect 12444 6426 12545 6482
rect 12444 6392 12477 6426
rect 12511 6392 12545 6426
rect 12444 6336 12545 6392
rect 12444 6302 12477 6336
rect 12511 6302 12545 6336
rect 12444 6246 12545 6302
rect 12444 6212 12477 6246
rect 12511 6212 12545 6246
rect 12444 6156 12545 6212
rect 12444 6122 12477 6156
rect 12511 6122 12545 6156
rect 12444 6066 12545 6122
rect 12444 6032 12477 6066
rect 12511 6032 12545 6066
rect 12444 5976 12545 6032
rect 12444 5942 12477 5976
rect 12511 5942 12545 5976
rect 13631 6876 13833 6932
rect 14919 6966 15121 6981
rect 14919 6932 14952 6966
rect 14986 6932 15053 6966
rect 15087 6932 15121 6966
rect 13631 6842 13664 6876
rect 13698 6842 13765 6876
rect 13799 6842 13833 6876
rect 13631 6786 13833 6842
rect 13631 6752 13664 6786
rect 13698 6752 13765 6786
rect 13799 6752 13833 6786
rect 13631 6696 13833 6752
rect 13631 6662 13664 6696
rect 13698 6662 13765 6696
rect 13799 6662 13833 6696
rect 13631 6606 13833 6662
rect 13631 6572 13664 6606
rect 13698 6572 13765 6606
rect 13799 6572 13833 6606
rect 13631 6516 13833 6572
rect 13631 6482 13664 6516
rect 13698 6482 13765 6516
rect 13799 6482 13833 6516
rect 13631 6426 13833 6482
rect 13631 6392 13664 6426
rect 13698 6392 13765 6426
rect 13799 6392 13833 6426
rect 13631 6336 13833 6392
rect 13631 6302 13664 6336
rect 13698 6302 13765 6336
rect 13799 6302 13833 6336
rect 13631 6246 13833 6302
rect 13631 6212 13664 6246
rect 13698 6212 13765 6246
rect 13799 6212 13833 6246
rect 13631 6156 13833 6212
rect 13631 6122 13664 6156
rect 13698 6122 13765 6156
rect 13799 6122 13833 6156
rect 13631 6066 13833 6122
rect 13631 6032 13664 6066
rect 13698 6032 13765 6066
rect 13799 6032 13833 6066
rect 13631 5976 13833 6032
rect 12444 5895 12545 5942
rect 13631 5942 13664 5976
rect 13698 5942 13765 5976
rect 13799 5942 13833 5976
rect 14919 6876 15121 6932
rect 16207 6966 16409 6981
rect 16207 6932 16240 6966
rect 16274 6932 16341 6966
rect 16375 6932 16409 6966
rect 14919 6842 14952 6876
rect 14986 6842 15053 6876
rect 15087 6842 15121 6876
rect 14919 6786 15121 6842
rect 14919 6752 14952 6786
rect 14986 6752 15053 6786
rect 15087 6752 15121 6786
rect 14919 6696 15121 6752
rect 14919 6662 14952 6696
rect 14986 6662 15053 6696
rect 15087 6662 15121 6696
rect 14919 6606 15121 6662
rect 14919 6572 14952 6606
rect 14986 6572 15053 6606
rect 15087 6572 15121 6606
rect 14919 6516 15121 6572
rect 14919 6482 14952 6516
rect 14986 6482 15053 6516
rect 15087 6482 15121 6516
rect 14919 6426 15121 6482
rect 14919 6392 14952 6426
rect 14986 6392 15053 6426
rect 15087 6392 15121 6426
rect 14919 6336 15121 6392
rect 14919 6302 14952 6336
rect 14986 6302 15053 6336
rect 15087 6302 15121 6336
rect 14919 6246 15121 6302
rect 14919 6212 14952 6246
rect 14986 6212 15053 6246
rect 15087 6212 15121 6246
rect 14919 6156 15121 6212
rect 14919 6122 14952 6156
rect 14986 6122 15053 6156
rect 15087 6122 15121 6156
rect 14919 6066 15121 6122
rect 14919 6032 14952 6066
rect 14986 6032 15053 6066
rect 15087 6032 15121 6066
rect 14919 5976 15121 6032
rect 13631 5895 13833 5942
rect 14919 5942 14952 5976
rect 14986 5942 15053 5976
rect 15087 5942 15121 5976
rect 16207 6876 16409 6932
rect 17495 6966 17697 6981
rect 17495 6932 17528 6966
rect 17562 6932 17629 6966
rect 17663 6932 17697 6966
rect 16207 6842 16240 6876
rect 16274 6842 16341 6876
rect 16375 6842 16409 6876
rect 16207 6786 16409 6842
rect 16207 6752 16240 6786
rect 16274 6752 16341 6786
rect 16375 6752 16409 6786
rect 16207 6696 16409 6752
rect 16207 6662 16240 6696
rect 16274 6662 16341 6696
rect 16375 6662 16409 6696
rect 16207 6606 16409 6662
rect 16207 6572 16240 6606
rect 16274 6572 16341 6606
rect 16375 6572 16409 6606
rect 16207 6516 16409 6572
rect 16207 6482 16240 6516
rect 16274 6482 16341 6516
rect 16375 6482 16409 6516
rect 16207 6426 16409 6482
rect 16207 6392 16240 6426
rect 16274 6392 16341 6426
rect 16375 6392 16409 6426
rect 16207 6336 16409 6392
rect 16207 6302 16240 6336
rect 16274 6302 16341 6336
rect 16375 6302 16409 6336
rect 16207 6246 16409 6302
rect 16207 6212 16240 6246
rect 16274 6212 16341 6246
rect 16375 6212 16409 6246
rect 16207 6156 16409 6212
rect 16207 6122 16240 6156
rect 16274 6122 16341 6156
rect 16375 6122 16409 6156
rect 16207 6066 16409 6122
rect 16207 6032 16240 6066
rect 16274 6032 16341 6066
rect 16375 6032 16409 6066
rect 16207 5976 16409 6032
rect 14919 5895 15121 5942
rect 16207 5942 16240 5976
rect 16274 5942 16341 5976
rect 16375 5942 16409 5976
rect 17495 6876 17697 6932
rect 18783 6966 18884 6981
rect 18783 6932 18816 6966
rect 18850 6932 18884 6966
rect 17495 6842 17528 6876
rect 17562 6842 17629 6876
rect 17663 6842 17697 6876
rect 17495 6786 17697 6842
rect 17495 6752 17528 6786
rect 17562 6752 17629 6786
rect 17663 6752 17697 6786
rect 17495 6696 17697 6752
rect 17495 6662 17528 6696
rect 17562 6662 17629 6696
rect 17663 6662 17697 6696
rect 17495 6606 17697 6662
rect 17495 6572 17528 6606
rect 17562 6572 17629 6606
rect 17663 6572 17697 6606
rect 17495 6516 17697 6572
rect 17495 6482 17528 6516
rect 17562 6482 17629 6516
rect 17663 6482 17697 6516
rect 17495 6426 17697 6482
rect 17495 6392 17528 6426
rect 17562 6392 17629 6426
rect 17663 6392 17697 6426
rect 17495 6336 17697 6392
rect 17495 6302 17528 6336
rect 17562 6302 17629 6336
rect 17663 6302 17697 6336
rect 17495 6246 17697 6302
rect 17495 6212 17528 6246
rect 17562 6212 17629 6246
rect 17663 6212 17697 6246
rect 17495 6156 17697 6212
rect 17495 6122 17528 6156
rect 17562 6122 17629 6156
rect 17663 6122 17697 6156
rect 17495 6066 17697 6122
rect 17495 6032 17528 6066
rect 17562 6032 17629 6066
rect 17663 6032 17697 6066
rect 17495 5976 17697 6032
rect 16207 5895 16409 5942
rect 17495 5942 17528 5976
rect 17562 5942 17629 5976
rect 17663 5942 17697 5976
rect 18783 6876 18884 6932
rect 18783 6842 18816 6876
rect 18850 6842 18884 6876
rect 18783 6786 18884 6842
rect 18783 6752 18816 6786
rect 18850 6752 18884 6786
rect 18783 6696 18884 6752
rect 18783 6662 18816 6696
rect 18850 6662 18884 6696
rect 18783 6606 18884 6662
rect 18783 6572 18816 6606
rect 18850 6572 18884 6606
rect 18783 6516 18884 6572
rect 18783 6482 18816 6516
rect 18850 6482 18884 6516
rect 18783 6426 18884 6482
rect 18783 6392 18816 6426
rect 18850 6392 18884 6426
rect 18783 6336 18884 6392
rect 18783 6302 18816 6336
rect 18850 6302 18884 6336
rect 18783 6246 18884 6302
rect 18783 6212 18816 6246
rect 18850 6212 18884 6246
rect 18783 6156 18884 6212
rect 18783 6122 18816 6156
rect 18850 6122 18884 6156
rect 18783 6066 18884 6122
rect 18783 6032 18816 6066
rect 18850 6032 18884 6066
rect 18783 5976 18884 6032
rect 17495 5895 17697 5942
rect 18783 5942 18816 5976
rect 18850 5942 18884 5976
rect 18783 5895 18884 5942
rect 12444 5886 18884 5895
rect 12444 5852 12477 5886
rect 12511 5863 13664 5886
rect 12511 5852 12578 5863
rect 12444 5829 12578 5852
rect 12612 5829 12668 5863
rect 12702 5829 12758 5863
rect 12792 5829 12848 5863
rect 12882 5829 12938 5863
rect 12972 5829 13028 5863
rect 13062 5829 13118 5863
rect 13152 5829 13208 5863
rect 13242 5829 13298 5863
rect 13332 5829 13388 5863
rect 13422 5829 13478 5863
rect 13512 5829 13568 5863
rect 13602 5852 13664 5863
rect 13698 5852 13765 5886
rect 13799 5863 14952 5886
rect 13799 5852 13866 5863
rect 13602 5829 13866 5852
rect 13900 5829 13956 5863
rect 13990 5829 14046 5863
rect 14080 5829 14136 5863
rect 14170 5829 14226 5863
rect 14260 5829 14316 5863
rect 14350 5829 14406 5863
rect 14440 5829 14496 5863
rect 14530 5829 14586 5863
rect 14620 5829 14676 5863
rect 14710 5829 14766 5863
rect 14800 5829 14856 5863
rect 14890 5852 14952 5863
rect 14986 5852 15053 5886
rect 15087 5863 16240 5886
rect 15087 5852 15154 5863
rect 14890 5829 15154 5852
rect 15188 5829 15244 5863
rect 15278 5829 15334 5863
rect 15368 5829 15424 5863
rect 15458 5829 15514 5863
rect 15548 5829 15604 5863
rect 15638 5829 15694 5863
rect 15728 5829 15784 5863
rect 15818 5829 15874 5863
rect 15908 5829 15964 5863
rect 15998 5829 16054 5863
rect 16088 5829 16144 5863
rect 16178 5852 16240 5863
rect 16274 5852 16341 5886
rect 16375 5863 17528 5886
rect 16375 5852 16442 5863
rect 16178 5829 16442 5852
rect 16476 5829 16532 5863
rect 16566 5829 16622 5863
rect 16656 5829 16712 5863
rect 16746 5829 16802 5863
rect 16836 5829 16892 5863
rect 16926 5829 16982 5863
rect 17016 5829 17072 5863
rect 17106 5829 17162 5863
rect 17196 5829 17252 5863
rect 17286 5829 17342 5863
rect 17376 5829 17432 5863
rect 17466 5852 17528 5863
rect 17562 5852 17629 5886
rect 17663 5863 18816 5886
rect 17663 5852 17730 5863
rect 17466 5829 17730 5852
rect 17764 5829 17820 5863
rect 17854 5829 17910 5863
rect 17944 5829 18000 5863
rect 18034 5829 18090 5863
rect 18124 5829 18180 5863
rect 18214 5829 18270 5863
rect 18304 5829 18360 5863
rect 18394 5829 18450 5863
rect 18484 5829 18540 5863
rect 18574 5829 18630 5863
rect 18664 5829 18720 5863
rect 18754 5852 18816 5863
rect 18850 5852 18884 5886
rect 18754 5829 18884 5852
rect 12444 5762 18884 5829
rect 12444 5728 12578 5762
rect 12612 5728 12668 5762
rect 12702 5728 12758 5762
rect 12792 5728 12848 5762
rect 12882 5728 12938 5762
rect 12972 5728 13028 5762
rect 13062 5728 13118 5762
rect 13152 5728 13208 5762
rect 13242 5728 13298 5762
rect 13332 5728 13388 5762
rect 13422 5728 13478 5762
rect 13512 5728 13568 5762
rect 13602 5728 13866 5762
rect 13900 5728 13956 5762
rect 13990 5728 14046 5762
rect 14080 5728 14136 5762
rect 14170 5728 14226 5762
rect 14260 5728 14316 5762
rect 14350 5728 14406 5762
rect 14440 5728 14496 5762
rect 14530 5728 14586 5762
rect 14620 5728 14676 5762
rect 14710 5728 14766 5762
rect 14800 5728 14856 5762
rect 14890 5728 15154 5762
rect 15188 5728 15244 5762
rect 15278 5728 15334 5762
rect 15368 5728 15424 5762
rect 15458 5728 15514 5762
rect 15548 5728 15604 5762
rect 15638 5728 15694 5762
rect 15728 5728 15784 5762
rect 15818 5728 15874 5762
rect 15908 5728 15964 5762
rect 15998 5728 16054 5762
rect 16088 5728 16144 5762
rect 16178 5728 16442 5762
rect 16476 5728 16532 5762
rect 16566 5728 16622 5762
rect 16656 5728 16712 5762
rect 16746 5728 16802 5762
rect 16836 5728 16892 5762
rect 16926 5728 16982 5762
rect 17016 5728 17072 5762
rect 17106 5728 17162 5762
rect 17196 5728 17252 5762
rect 17286 5728 17342 5762
rect 17376 5728 17432 5762
rect 17466 5728 17730 5762
rect 17764 5728 17820 5762
rect 17854 5728 17910 5762
rect 17944 5728 18000 5762
rect 18034 5728 18090 5762
rect 18124 5728 18180 5762
rect 18214 5728 18270 5762
rect 18304 5728 18360 5762
rect 18394 5728 18450 5762
rect 18484 5728 18540 5762
rect 18574 5728 18630 5762
rect 18664 5728 18720 5762
rect 18754 5728 18884 5762
rect 12444 5693 18884 5728
rect 12444 5678 12545 5693
rect 12444 5644 12477 5678
rect 12511 5644 12545 5678
rect 12444 5588 12545 5644
rect 13631 5678 13833 5693
rect 13631 5644 13664 5678
rect 13698 5644 13765 5678
rect 13799 5644 13833 5678
rect 12444 5554 12477 5588
rect 12511 5554 12545 5588
rect 12444 5498 12545 5554
rect 12444 5464 12477 5498
rect 12511 5464 12545 5498
rect 12444 5408 12545 5464
rect 12444 5374 12477 5408
rect 12511 5374 12545 5408
rect 12444 5318 12545 5374
rect 12444 5284 12477 5318
rect 12511 5284 12545 5318
rect 12444 5228 12545 5284
rect 12444 5194 12477 5228
rect 12511 5194 12545 5228
rect 12444 5138 12545 5194
rect 12444 5104 12477 5138
rect 12511 5104 12545 5138
rect 12444 5048 12545 5104
rect 12444 5014 12477 5048
rect 12511 5014 12545 5048
rect 12444 4958 12545 5014
rect 12444 4924 12477 4958
rect 12511 4924 12545 4958
rect 12444 4868 12545 4924
rect 12444 4834 12477 4868
rect 12511 4834 12545 4868
rect 12444 4778 12545 4834
rect 12444 4744 12477 4778
rect 12511 4744 12545 4778
rect 12444 4688 12545 4744
rect 12444 4654 12477 4688
rect 12511 4654 12545 4688
rect 13631 5588 13833 5644
rect 14919 5678 15121 5693
rect 14919 5644 14952 5678
rect 14986 5644 15053 5678
rect 15087 5644 15121 5678
rect 13631 5554 13664 5588
rect 13698 5554 13765 5588
rect 13799 5554 13833 5588
rect 13631 5498 13833 5554
rect 13631 5464 13664 5498
rect 13698 5464 13765 5498
rect 13799 5464 13833 5498
rect 13631 5408 13833 5464
rect 13631 5374 13664 5408
rect 13698 5374 13765 5408
rect 13799 5374 13833 5408
rect 13631 5318 13833 5374
rect 13631 5284 13664 5318
rect 13698 5284 13765 5318
rect 13799 5284 13833 5318
rect 13631 5228 13833 5284
rect 13631 5194 13664 5228
rect 13698 5194 13765 5228
rect 13799 5194 13833 5228
rect 13631 5138 13833 5194
rect 13631 5104 13664 5138
rect 13698 5104 13765 5138
rect 13799 5104 13833 5138
rect 13631 5048 13833 5104
rect 13631 5014 13664 5048
rect 13698 5014 13765 5048
rect 13799 5014 13833 5048
rect 13631 4958 13833 5014
rect 13631 4924 13664 4958
rect 13698 4924 13765 4958
rect 13799 4924 13833 4958
rect 13631 4868 13833 4924
rect 13631 4834 13664 4868
rect 13698 4834 13765 4868
rect 13799 4834 13833 4868
rect 13631 4778 13833 4834
rect 13631 4744 13664 4778
rect 13698 4744 13765 4778
rect 13799 4744 13833 4778
rect 13631 4688 13833 4744
rect 12444 4607 12545 4654
rect 13631 4654 13664 4688
rect 13698 4654 13765 4688
rect 13799 4654 13833 4688
rect 14919 5588 15121 5644
rect 16207 5678 16409 5693
rect 16207 5644 16240 5678
rect 16274 5644 16341 5678
rect 16375 5644 16409 5678
rect 14919 5554 14952 5588
rect 14986 5554 15053 5588
rect 15087 5554 15121 5588
rect 14919 5498 15121 5554
rect 14919 5464 14952 5498
rect 14986 5464 15053 5498
rect 15087 5464 15121 5498
rect 14919 5408 15121 5464
rect 14919 5374 14952 5408
rect 14986 5374 15053 5408
rect 15087 5374 15121 5408
rect 14919 5318 15121 5374
rect 14919 5284 14952 5318
rect 14986 5284 15053 5318
rect 15087 5284 15121 5318
rect 14919 5228 15121 5284
rect 14919 5194 14952 5228
rect 14986 5194 15053 5228
rect 15087 5194 15121 5228
rect 14919 5138 15121 5194
rect 14919 5104 14952 5138
rect 14986 5104 15053 5138
rect 15087 5104 15121 5138
rect 14919 5048 15121 5104
rect 14919 5014 14952 5048
rect 14986 5014 15053 5048
rect 15087 5014 15121 5048
rect 14919 4958 15121 5014
rect 14919 4924 14952 4958
rect 14986 4924 15053 4958
rect 15087 4924 15121 4958
rect 14919 4868 15121 4924
rect 14919 4834 14952 4868
rect 14986 4834 15053 4868
rect 15087 4834 15121 4868
rect 14919 4778 15121 4834
rect 14919 4744 14952 4778
rect 14986 4744 15053 4778
rect 15087 4744 15121 4778
rect 14919 4688 15121 4744
rect 13631 4607 13833 4654
rect 14919 4654 14952 4688
rect 14986 4654 15053 4688
rect 15087 4654 15121 4688
rect 16207 5588 16409 5644
rect 17495 5678 17697 5693
rect 17495 5644 17528 5678
rect 17562 5644 17629 5678
rect 17663 5644 17697 5678
rect 16207 5554 16240 5588
rect 16274 5554 16341 5588
rect 16375 5554 16409 5588
rect 16207 5498 16409 5554
rect 16207 5464 16240 5498
rect 16274 5464 16341 5498
rect 16375 5464 16409 5498
rect 16207 5408 16409 5464
rect 16207 5374 16240 5408
rect 16274 5374 16341 5408
rect 16375 5374 16409 5408
rect 16207 5318 16409 5374
rect 16207 5284 16240 5318
rect 16274 5284 16341 5318
rect 16375 5284 16409 5318
rect 16207 5228 16409 5284
rect 16207 5194 16240 5228
rect 16274 5194 16341 5228
rect 16375 5194 16409 5228
rect 16207 5138 16409 5194
rect 16207 5104 16240 5138
rect 16274 5104 16341 5138
rect 16375 5104 16409 5138
rect 16207 5048 16409 5104
rect 16207 5014 16240 5048
rect 16274 5014 16341 5048
rect 16375 5014 16409 5048
rect 16207 4958 16409 5014
rect 16207 4924 16240 4958
rect 16274 4924 16341 4958
rect 16375 4924 16409 4958
rect 16207 4868 16409 4924
rect 16207 4834 16240 4868
rect 16274 4834 16341 4868
rect 16375 4834 16409 4868
rect 16207 4778 16409 4834
rect 16207 4744 16240 4778
rect 16274 4744 16341 4778
rect 16375 4744 16409 4778
rect 16207 4688 16409 4744
rect 14919 4607 15121 4654
rect 16207 4654 16240 4688
rect 16274 4654 16341 4688
rect 16375 4654 16409 4688
rect 17495 5588 17697 5644
rect 18783 5678 18884 5693
rect 18783 5644 18816 5678
rect 18850 5644 18884 5678
rect 17495 5554 17528 5588
rect 17562 5554 17629 5588
rect 17663 5554 17697 5588
rect 17495 5498 17697 5554
rect 17495 5464 17528 5498
rect 17562 5464 17629 5498
rect 17663 5464 17697 5498
rect 17495 5408 17697 5464
rect 17495 5374 17528 5408
rect 17562 5374 17629 5408
rect 17663 5374 17697 5408
rect 17495 5318 17697 5374
rect 17495 5284 17528 5318
rect 17562 5284 17629 5318
rect 17663 5284 17697 5318
rect 17495 5228 17697 5284
rect 17495 5194 17528 5228
rect 17562 5194 17629 5228
rect 17663 5194 17697 5228
rect 17495 5138 17697 5194
rect 17495 5104 17528 5138
rect 17562 5104 17629 5138
rect 17663 5104 17697 5138
rect 17495 5048 17697 5104
rect 17495 5014 17528 5048
rect 17562 5014 17629 5048
rect 17663 5014 17697 5048
rect 17495 4958 17697 5014
rect 17495 4924 17528 4958
rect 17562 4924 17629 4958
rect 17663 4924 17697 4958
rect 17495 4868 17697 4924
rect 17495 4834 17528 4868
rect 17562 4834 17629 4868
rect 17663 4834 17697 4868
rect 17495 4778 17697 4834
rect 17495 4744 17528 4778
rect 17562 4744 17629 4778
rect 17663 4744 17697 4778
rect 17495 4688 17697 4744
rect 16207 4607 16409 4654
rect 17495 4654 17528 4688
rect 17562 4654 17629 4688
rect 17663 4654 17697 4688
rect 18783 5588 18884 5644
rect 18783 5554 18816 5588
rect 18850 5554 18884 5588
rect 18783 5498 18884 5554
rect 18783 5464 18816 5498
rect 18850 5464 18884 5498
rect 18783 5408 18884 5464
rect 18783 5374 18816 5408
rect 18850 5374 18884 5408
rect 18783 5318 18884 5374
rect 18783 5284 18816 5318
rect 18850 5284 18884 5318
rect 18783 5228 18884 5284
rect 18783 5194 18816 5228
rect 18850 5194 18884 5228
rect 18783 5138 18884 5194
rect 18783 5104 18816 5138
rect 18850 5104 18884 5138
rect 18783 5048 18884 5104
rect 18783 5014 18816 5048
rect 18850 5014 18884 5048
rect 18783 4958 18884 5014
rect 18783 4924 18816 4958
rect 18850 4924 18884 4958
rect 18783 4868 18884 4924
rect 18783 4834 18816 4868
rect 18850 4834 18884 4868
rect 18783 4778 18884 4834
rect 18783 4744 18816 4778
rect 18850 4744 18884 4778
rect 18783 4688 18884 4744
rect 17495 4607 17697 4654
rect 18783 4654 18816 4688
rect 18850 4654 18884 4688
rect 18783 4607 18884 4654
rect 12444 4598 18884 4607
rect 12444 4564 12477 4598
rect 12511 4575 13664 4598
rect 12511 4564 12578 4575
rect 12444 4541 12578 4564
rect 12612 4541 12668 4575
rect 12702 4541 12758 4575
rect 12792 4541 12848 4575
rect 12882 4541 12938 4575
rect 12972 4541 13028 4575
rect 13062 4541 13118 4575
rect 13152 4541 13208 4575
rect 13242 4541 13298 4575
rect 13332 4541 13388 4575
rect 13422 4541 13478 4575
rect 13512 4541 13568 4575
rect 13602 4564 13664 4575
rect 13698 4564 13765 4598
rect 13799 4575 14952 4598
rect 13799 4564 13866 4575
rect 13602 4541 13866 4564
rect 13900 4541 13956 4575
rect 13990 4541 14046 4575
rect 14080 4541 14136 4575
rect 14170 4541 14226 4575
rect 14260 4541 14316 4575
rect 14350 4541 14406 4575
rect 14440 4541 14496 4575
rect 14530 4541 14586 4575
rect 14620 4541 14676 4575
rect 14710 4541 14766 4575
rect 14800 4541 14856 4575
rect 14890 4564 14952 4575
rect 14986 4564 15053 4598
rect 15087 4575 16240 4598
rect 15087 4564 15154 4575
rect 14890 4541 15154 4564
rect 15188 4541 15244 4575
rect 15278 4541 15334 4575
rect 15368 4541 15424 4575
rect 15458 4541 15514 4575
rect 15548 4541 15604 4575
rect 15638 4541 15694 4575
rect 15728 4541 15784 4575
rect 15818 4541 15874 4575
rect 15908 4541 15964 4575
rect 15998 4541 16054 4575
rect 16088 4541 16144 4575
rect 16178 4564 16240 4575
rect 16274 4564 16341 4598
rect 16375 4575 17528 4598
rect 16375 4564 16442 4575
rect 16178 4541 16442 4564
rect 16476 4541 16532 4575
rect 16566 4541 16622 4575
rect 16656 4541 16712 4575
rect 16746 4541 16802 4575
rect 16836 4541 16892 4575
rect 16926 4541 16982 4575
rect 17016 4541 17072 4575
rect 17106 4541 17162 4575
rect 17196 4541 17252 4575
rect 17286 4541 17342 4575
rect 17376 4541 17432 4575
rect 17466 4564 17528 4575
rect 17562 4564 17629 4598
rect 17663 4575 18816 4598
rect 17663 4564 17730 4575
rect 17466 4541 17730 4564
rect 17764 4541 17820 4575
rect 17854 4541 17910 4575
rect 17944 4541 18000 4575
rect 18034 4541 18090 4575
rect 18124 4541 18180 4575
rect 18214 4541 18270 4575
rect 18304 4541 18360 4575
rect 18394 4541 18450 4575
rect 18484 4541 18540 4575
rect 18574 4541 18630 4575
rect 18664 4541 18720 4575
rect 18754 4564 18816 4575
rect 18850 4564 18884 4598
rect 18754 4541 18884 4564
rect 12444 4474 18884 4541
rect 12444 4440 12578 4474
rect 12612 4440 12668 4474
rect 12702 4440 12758 4474
rect 12792 4440 12848 4474
rect 12882 4440 12938 4474
rect 12972 4440 13028 4474
rect 13062 4440 13118 4474
rect 13152 4440 13208 4474
rect 13242 4440 13298 4474
rect 13332 4440 13388 4474
rect 13422 4440 13478 4474
rect 13512 4440 13568 4474
rect 13602 4440 13866 4474
rect 13900 4440 13956 4474
rect 13990 4440 14046 4474
rect 14080 4440 14136 4474
rect 14170 4440 14226 4474
rect 14260 4440 14316 4474
rect 14350 4440 14406 4474
rect 14440 4440 14496 4474
rect 14530 4440 14586 4474
rect 14620 4440 14676 4474
rect 14710 4440 14766 4474
rect 14800 4440 14856 4474
rect 14890 4440 15154 4474
rect 15188 4440 15244 4474
rect 15278 4440 15334 4474
rect 15368 4440 15424 4474
rect 15458 4440 15514 4474
rect 15548 4440 15604 4474
rect 15638 4440 15694 4474
rect 15728 4440 15784 4474
rect 15818 4440 15874 4474
rect 15908 4440 15964 4474
rect 15998 4440 16054 4474
rect 16088 4440 16144 4474
rect 16178 4440 16442 4474
rect 16476 4440 16532 4474
rect 16566 4440 16622 4474
rect 16656 4440 16712 4474
rect 16746 4440 16802 4474
rect 16836 4440 16892 4474
rect 16926 4440 16982 4474
rect 17016 4440 17072 4474
rect 17106 4440 17162 4474
rect 17196 4440 17252 4474
rect 17286 4440 17342 4474
rect 17376 4440 17432 4474
rect 17466 4440 17730 4474
rect 17764 4440 17820 4474
rect 17854 4440 17910 4474
rect 17944 4440 18000 4474
rect 18034 4440 18090 4474
rect 18124 4440 18180 4474
rect 18214 4440 18270 4474
rect 18304 4440 18360 4474
rect 18394 4440 18450 4474
rect 18484 4440 18540 4474
rect 18574 4440 18630 4474
rect 18664 4440 18720 4474
rect 18754 4440 18884 4474
rect 12444 4405 18884 4440
rect 12444 4390 12545 4405
rect 12444 4356 12477 4390
rect 12511 4356 12545 4390
rect 12444 4300 12545 4356
rect 13631 4390 13833 4405
rect 13631 4356 13664 4390
rect 13698 4356 13765 4390
rect 13799 4356 13833 4390
rect 12444 4266 12477 4300
rect 12511 4266 12545 4300
rect 12444 4210 12545 4266
rect 12444 4176 12477 4210
rect 12511 4176 12545 4210
rect 12444 4120 12545 4176
rect 12444 4086 12477 4120
rect 12511 4086 12545 4120
rect 12444 4030 12545 4086
rect 12444 3996 12477 4030
rect 12511 3996 12545 4030
rect 12444 3940 12545 3996
rect 12444 3906 12477 3940
rect 12511 3906 12545 3940
rect 12444 3850 12545 3906
rect 12444 3816 12477 3850
rect 12511 3816 12545 3850
rect 12444 3760 12545 3816
rect 12444 3726 12477 3760
rect 12511 3726 12545 3760
rect 12444 3670 12545 3726
rect 12444 3636 12477 3670
rect 12511 3636 12545 3670
rect 12444 3580 12545 3636
rect 12444 3546 12477 3580
rect 12511 3546 12545 3580
rect 12444 3490 12545 3546
rect 12444 3456 12477 3490
rect 12511 3456 12545 3490
rect 12444 3400 12545 3456
rect 12444 3366 12477 3400
rect 12511 3366 12545 3400
rect 13631 4300 13833 4356
rect 14919 4390 15121 4405
rect 14919 4356 14952 4390
rect 14986 4356 15053 4390
rect 15087 4356 15121 4390
rect 13631 4266 13664 4300
rect 13698 4266 13765 4300
rect 13799 4266 13833 4300
rect 13631 4210 13833 4266
rect 13631 4176 13664 4210
rect 13698 4176 13765 4210
rect 13799 4176 13833 4210
rect 13631 4120 13833 4176
rect 13631 4086 13664 4120
rect 13698 4086 13765 4120
rect 13799 4086 13833 4120
rect 13631 4030 13833 4086
rect 13631 3996 13664 4030
rect 13698 3996 13765 4030
rect 13799 3996 13833 4030
rect 13631 3940 13833 3996
rect 13631 3906 13664 3940
rect 13698 3906 13765 3940
rect 13799 3906 13833 3940
rect 13631 3850 13833 3906
rect 13631 3816 13664 3850
rect 13698 3816 13765 3850
rect 13799 3816 13833 3850
rect 13631 3760 13833 3816
rect 13631 3726 13664 3760
rect 13698 3726 13765 3760
rect 13799 3726 13833 3760
rect 13631 3670 13833 3726
rect 13631 3636 13664 3670
rect 13698 3636 13765 3670
rect 13799 3636 13833 3670
rect 13631 3580 13833 3636
rect 13631 3546 13664 3580
rect 13698 3546 13765 3580
rect 13799 3546 13833 3580
rect 13631 3490 13833 3546
rect 13631 3456 13664 3490
rect 13698 3456 13765 3490
rect 13799 3456 13833 3490
rect 13631 3400 13833 3456
rect 12444 3319 12545 3366
rect 13631 3366 13664 3400
rect 13698 3366 13765 3400
rect 13799 3366 13833 3400
rect 14919 4300 15121 4356
rect 16207 4390 16409 4405
rect 16207 4356 16240 4390
rect 16274 4356 16341 4390
rect 16375 4356 16409 4390
rect 14919 4266 14952 4300
rect 14986 4266 15053 4300
rect 15087 4266 15121 4300
rect 14919 4210 15121 4266
rect 14919 4176 14952 4210
rect 14986 4176 15053 4210
rect 15087 4176 15121 4210
rect 14919 4120 15121 4176
rect 14919 4086 14952 4120
rect 14986 4086 15053 4120
rect 15087 4086 15121 4120
rect 14919 4030 15121 4086
rect 14919 3996 14952 4030
rect 14986 3996 15053 4030
rect 15087 3996 15121 4030
rect 14919 3940 15121 3996
rect 14919 3906 14952 3940
rect 14986 3906 15053 3940
rect 15087 3906 15121 3940
rect 14919 3850 15121 3906
rect 14919 3816 14952 3850
rect 14986 3816 15053 3850
rect 15087 3816 15121 3850
rect 14919 3760 15121 3816
rect 14919 3726 14952 3760
rect 14986 3726 15053 3760
rect 15087 3726 15121 3760
rect 14919 3670 15121 3726
rect 14919 3636 14952 3670
rect 14986 3636 15053 3670
rect 15087 3636 15121 3670
rect 14919 3580 15121 3636
rect 14919 3546 14952 3580
rect 14986 3546 15053 3580
rect 15087 3546 15121 3580
rect 14919 3490 15121 3546
rect 14919 3456 14952 3490
rect 14986 3456 15053 3490
rect 15087 3456 15121 3490
rect 14919 3400 15121 3456
rect 13631 3319 13833 3366
rect 14919 3366 14952 3400
rect 14986 3366 15053 3400
rect 15087 3366 15121 3400
rect 16207 4300 16409 4356
rect 17495 4390 17697 4405
rect 17495 4356 17528 4390
rect 17562 4356 17629 4390
rect 17663 4356 17697 4390
rect 16207 4266 16240 4300
rect 16274 4266 16341 4300
rect 16375 4266 16409 4300
rect 16207 4210 16409 4266
rect 16207 4176 16240 4210
rect 16274 4176 16341 4210
rect 16375 4176 16409 4210
rect 16207 4120 16409 4176
rect 16207 4086 16240 4120
rect 16274 4086 16341 4120
rect 16375 4086 16409 4120
rect 16207 4030 16409 4086
rect 16207 3996 16240 4030
rect 16274 3996 16341 4030
rect 16375 3996 16409 4030
rect 16207 3940 16409 3996
rect 16207 3906 16240 3940
rect 16274 3906 16341 3940
rect 16375 3906 16409 3940
rect 16207 3850 16409 3906
rect 16207 3816 16240 3850
rect 16274 3816 16341 3850
rect 16375 3816 16409 3850
rect 16207 3760 16409 3816
rect 16207 3726 16240 3760
rect 16274 3726 16341 3760
rect 16375 3726 16409 3760
rect 16207 3670 16409 3726
rect 16207 3636 16240 3670
rect 16274 3636 16341 3670
rect 16375 3636 16409 3670
rect 16207 3580 16409 3636
rect 16207 3546 16240 3580
rect 16274 3546 16341 3580
rect 16375 3546 16409 3580
rect 16207 3490 16409 3546
rect 16207 3456 16240 3490
rect 16274 3456 16341 3490
rect 16375 3456 16409 3490
rect 16207 3400 16409 3456
rect 14919 3319 15121 3366
rect 16207 3366 16240 3400
rect 16274 3366 16341 3400
rect 16375 3366 16409 3400
rect 17495 4300 17697 4356
rect 18783 4390 18884 4405
rect 18783 4356 18816 4390
rect 18850 4356 18884 4390
rect 17495 4266 17528 4300
rect 17562 4266 17629 4300
rect 17663 4266 17697 4300
rect 17495 4210 17697 4266
rect 17495 4176 17528 4210
rect 17562 4176 17629 4210
rect 17663 4176 17697 4210
rect 17495 4120 17697 4176
rect 17495 4086 17528 4120
rect 17562 4086 17629 4120
rect 17663 4086 17697 4120
rect 17495 4030 17697 4086
rect 17495 3996 17528 4030
rect 17562 3996 17629 4030
rect 17663 3996 17697 4030
rect 17495 3940 17697 3996
rect 17495 3906 17528 3940
rect 17562 3906 17629 3940
rect 17663 3906 17697 3940
rect 17495 3850 17697 3906
rect 17495 3816 17528 3850
rect 17562 3816 17629 3850
rect 17663 3816 17697 3850
rect 17495 3760 17697 3816
rect 17495 3726 17528 3760
rect 17562 3726 17629 3760
rect 17663 3726 17697 3760
rect 17495 3670 17697 3726
rect 17495 3636 17528 3670
rect 17562 3636 17629 3670
rect 17663 3636 17697 3670
rect 17495 3580 17697 3636
rect 17495 3546 17528 3580
rect 17562 3546 17629 3580
rect 17663 3546 17697 3580
rect 17495 3490 17697 3546
rect 17495 3456 17528 3490
rect 17562 3456 17629 3490
rect 17663 3456 17697 3490
rect 17495 3400 17697 3456
rect 16207 3319 16409 3366
rect 17495 3366 17528 3400
rect 17562 3366 17629 3400
rect 17663 3366 17697 3400
rect 18783 4300 18884 4356
rect 18783 4266 18816 4300
rect 18850 4266 18884 4300
rect 18783 4210 18884 4266
rect 18783 4176 18816 4210
rect 18850 4176 18884 4210
rect 18783 4120 18884 4176
rect 18783 4086 18816 4120
rect 18850 4086 18884 4120
rect 18783 4030 18884 4086
rect 18783 3996 18816 4030
rect 18850 3996 18884 4030
rect 18783 3940 18884 3996
rect 18783 3906 18816 3940
rect 18850 3906 18884 3940
rect 18783 3850 18884 3906
rect 18783 3816 18816 3850
rect 18850 3816 18884 3850
rect 18783 3760 18884 3816
rect 18783 3726 18816 3760
rect 18850 3726 18884 3760
rect 18783 3670 18884 3726
rect 18783 3636 18816 3670
rect 18850 3636 18884 3670
rect 18783 3580 18884 3636
rect 18783 3546 18816 3580
rect 18850 3546 18884 3580
rect 18783 3490 18884 3546
rect 18783 3456 18816 3490
rect 18850 3456 18884 3490
rect 18783 3400 18884 3456
rect 17495 3319 17697 3366
rect 18783 3366 18816 3400
rect 18850 3366 18884 3400
rect 18783 3319 18884 3366
rect 12444 3310 18884 3319
rect 12444 3276 12477 3310
rect 12511 3287 13664 3310
rect 12511 3276 12578 3287
rect 12444 3253 12578 3276
rect 12612 3253 12668 3287
rect 12702 3253 12758 3287
rect 12792 3253 12848 3287
rect 12882 3253 12938 3287
rect 12972 3253 13028 3287
rect 13062 3253 13118 3287
rect 13152 3253 13208 3287
rect 13242 3253 13298 3287
rect 13332 3253 13388 3287
rect 13422 3253 13478 3287
rect 13512 3253 13568 3287
rect 13602 3276 13664 3287
rect 13698 3276 13765 3310
rect 13799 3287 14952 3310
rect 13799 3276 13866 3287
rect 13602 3253 13866 3276
rect 13900 3253 13956 3287
rect 13990 3253 14046 3287
rect 14080 3253 14136 3287
rect 14170 3253 14226 3287
rect 14260 3253 14316 3287
rect 14350 3253 14406 3287
rect 14440 3253 14496 3287
rect 14530 3253 14586 3287
rect 14620 3253 14676 3287
rect 14710 3253 14766 3287
rect 14800 3253 14856 3287
rect 14890 3276 14952 3287
rect 14986 3276 15053 3310
rect 15087 3287 16240 3310
rect 15087 3276 15154 3287
rect 14890 3253 15154 3276
rect 15188 3253 15244 3287
rect 15278 3253 15334 3287
rect 15368 3253 15424 3287
rect 15458 3253 15514 3287
rect 15548 3253 15604 3287
rect 15638 3253 15694 3287
rect 15728 3253 15784 3287
rect 15818 3253 15874 3287
rect 15908 3253 15964 3287
rect 15998 3253 16054 3287
rect 16088 3253 16144 3287
rect 16178 3276 16240 3287
rect 16274 3276 16341 3310
rect 16375 3287 17528 3310
rect 16375 3276 16442 3287
rect 16178 3253 16442 3276
rect 16476 3253 16532 3287
rect 16566 3253 16622 3287
rect 16656 3253 16712 3287
rect 16746 3253 16802 3287
rect 16836 3253 16892 3287
rect 16926 3253 16982 3287
rect 17016 3253 17072 3287
rect 17106 3253 17162 3287
rect 17196 3253 17252 3287
rect 17286 3253 17342 3287
rect 17376 3253 17432 3287
rect 17466 3276 17528 3287
rect 17562 3276 17629 3310
rect 17663 3287 18816 3310
rect 17663 3276 17730 3287
rect 17466 3253 17730 3276
rect 17764 3253 17820 3287
rect 17854 3253 17910 3287
rect 17944 3253 18000 3287
rect 18034 3253 18090 3287
rect 18124 3253 18180 3287
rect 18214 3253 18270 3287
rect 18304 3253 18360 3287
rect 18394 3253 18450 3287
rect 18484 3253 18540 3287
rect 18574 3253 18630 3287
rect 18664 3253 18720 3287
rect 18754 3276 18816 3287
rect 18850 3276 18884 3310
rect 18754 3253 18884 3276
rect 12444 3186 18884 3253
rect 12444 3152 12578 3186
rect 12612 3152 12668 3186
rect 12702 3152 12758 3186
rect 12792 3152 12848 3186
rect 12882 3152 12938 3186
rect 12972 3152 13028 3186
rect 13062 3152 13118 3186
rect 13152 3152 13208 3186
rect 13242 3152 13298 3186
rect 13332 3152 13388 3186
rect 13422 3152 13478 3186
rect 13512 3152 13568 3186
rect 13602 3152 13866 3186
rect 13900 3152 13956 3186
rect 13990 3152 14046 3186
rect 14080 3152 14136 3186
rect 14170 3152 14226 3186
rect 14260 3152 14316 3186
rect 14350 3152 14406 3186
rect 14440 3152 14496 3186
rect 14530 3152 14586 3186
rect 14620 3152 14676 3186
rect 14710 3152 14766 3186
rect 14800 3152 14856 3186
rect 14890 3152 15154 3186
rect 15188 3152 15244 3186
rect 15278 3152 15334 3186
rect 15368 3152 15424 3186
rect 15458 3152 15514 3186
rect 15548 3152 15604 3186
rect 15638 3152 15694 3186
rect 15728 3152 15784 3186
rect 15818 3152 15874 3186
rect 15908 3152 15964 3186
rect 15998 3152 16054 3186
rect 16088 3152 16144 3186
rect 16178 3152 16442 3186
rect 16476 3152 16532 3186
rect 16566 3152 16622 3186
rect 16656 3152 16712 3186
rect 16746 3152 16802 3186
rect 16836 3152 16892 3186
rect 16926 3152 16982 3186
rect 17016 3152 17072 3186
rect 17106 3152 17162 3186
rect 17196 3152 17252 3186
rect 17286 3152 17342 3186
rect 17376 3152 17432 3186
rect 17466 3152 17730 3186
rect 17764 3152 17820 3186
rect 17854 3152 17910 3186
rect 17944 3152 18000 3186
rect 18034 3152 18090 3186
rect 18124 3152 18180 3186
rect 18214 3152 18270 3186
rect 18304 3152 18360 3186
rect 18394 3152 18450 3186
rect 18484 3152 18540 3186
rect 18574 3152 18630 3186
rect 18664 3152 18720 3186
rect 18754 3152 18884 3186
rect 12444 3117 18884 3152
rect 12444 3102 12545 3117
rect 12444 3068 12477 3102
rect 12511 3068 12545 3102
rect 12444 3012 12545 3068
rect 13631 3102 13833 3117
rect 13631 3068 13664 3102
rect 13698 3068 13765 3102
rect 13799 3068 13833 3102
rect 12444 2978 12477 3012
rect 12511 2978 12545 3012
rect 12444 2922 12545 2978
rect 12444 2888 12477 2922
rect 12511 2888 12545 2922
rect 12444 2832 12545 2888
rect 12444 2798 12477 2832
rect 12511 2798 12545 2832
rect 12444 2742 12545 2798
rect 12444 2708 12477 2742
rect 12511 2708 12545 2742
rect 12444 2652 12545 2708
rect 12444 2618 12477 2652
rect 12511 2618 12545 2652
rect 12444 2562 12545 2618
rect 12444 2528 12477 2562
rect 12511 2528 12545 2562
rect 12444 2472 12545 2528
rect 12444 2438 12477 2472
rect 12511 2438 12545 2472
rect 12444 2382 12545 2438
rect 12444 2348 12477 2382
rect 12511 2348 12545 2382
rect 12444 2292 12545 2348
rect 12444 2258 12477 2292
rect 12511 2258 12545 2292
rect 12444 2202 12545 2258
rect 12444 2168 12477 2202
rect 12511 2168 12545 2202
rect 12444 2112 12545 2168
rect 12444 2078 12477 2112
rect 12511 2078 12545 2112
rect 13631 3012 13833 3068
rect 14919 3102 15121 3117
rect 14919 3068 14952 3102
rect 14986 3068 15053 3102
rect 15087 3068 15121 3102
rect 13631 2978 13664 3012
rect 13698 2978 13765 3012
rect 13799 2978 13833 3012
rect 13631 2922 13833 2978
rect 13631 2888 13664 2922
rect 13698 2888 13765 2922
rect 13799 2888 13833 2922
rect 13631 2832 13833 2888
rect 13631 2798 13664 2832
rect 13698 2798 13765 2832
rect 13799 2798 13833 2832
rect 13631 2742 13833 2798
rect 13631 2708 13664 2742
rect 13698 2708 13765 2742
rect 13799 2708 13833 2742
rect 13631 2652 13833 2708
rect 13631 2618 13664 2652
rect 13698 2618 13765 2652
rect 13799 2618 13833 2652
rect 13631 2562 13833 2618
rect 13631 2528 13664 2562
rect 13698 2528 13765 2562
rect 13799 2528 13833 2562
rect 13631 2472 13833 2528
rect 13631 2438 13664 2472
rect 13698 2438 13765 2472
rect 13799 2438 13833 2472
rect 13631 2382 13833 2438
rect 13631 2348 13664 2382
rect 13698 2348 13765 2382
rect 13799 2348 13833 2382
rect 13631 2292 13833 2348
rect 13631 2258 13664 2292
rect 13698 2258 13765 2292
rect 13799 2258 13833 2292
rect 13631 2202 13833 2258
rect 13631 2168 13664 2202
rect 13698 2168 13765 2202
rect 13799 2168 13833 2202
rect 13631 2112 13833 2168
rect 12444 2031 12545 2078
rect 13631 2078 13664 2112
rect 13698 2078 13765 2112
rect 13799 2078 13833 2112
rect 14919 3012 15121 3068
rect 16207 3102 16409 3117
rect 16207 3068 16240 3102
rect 16274 3068 16341 3102
rect 16375 3068 16409 3102
rect 14919 2978 14952 3012
rect 14986 2978 15053 3012
rect 15087 2978 15121 3012
rect 14919 2922 15121 2978
rect 14919 2888 14952 2922
rect 14986 2888 15053 2922
rect 15087 2888 15121 2922
rect 14919 2832 15121 2888
rect 14919 2798 14952 2832
rect 14986 2798 15053 2832
rect 15087 2798 15121 2832
rect 14919 2742 15121 2798
rect 14919 2708 14952 2742
rect 14986 2708 15053 2742
rect 15087 2708 15121 2742
rect 14919 2652 15121 2708
rect 14919 2618 14952 2652
rect 14986 2618 15053 2652
rect 15087 2618 15121 2652
rect 14919 2562 15121 2618
rect 14919 2528 14952 2562
rect 14986 2528 15053 2562
rect 15087 2528 15121 2562
rect 14919 2472 15121 2528
rect 14919 2438 14952 2472
rect 14986 2438 15053 2472
rect 15087 2438 15121 2472
rect 14919 2382 15121 2438
rect 14919 2348 14952 2382
rect 14986 2348 15053 2382
rect 15087 2348 15121 2382
rect 14919 2292 15121 2348
rect 14919 2258 14952 2292
rect 14986 2258 15053 2292
rect 15087 2258 15121 2292
rect 14919 2202 15121 2258
rect 14919 2168 14952 2202
rect 14986 2168 15053 2202
rect 15087 2168 15121 2202
rect 14919 2112 15121 2168
rect 13631 2031 13833 2078
rect 14919 2078 14952 2112
rect 14986 2078 15053 2112
rect 15087 2078 15121 2112
rect 16207 3012 16409 3068
rect 17495 3102 17697 3117
rect 17495 3068 17528 3102
rect 17562 3068 17629 3102
rect 17663 3068 17697 3102
rect 16207 2978 16240 3012
rect 16274 2978 16341 3012
rect 16375 2978 16409 3012
rect 16207 2922 16409 2978
rect 16207 2888 16240 2922
rect 16274 2888 16341 2922
rect 16375 2888 16409 2922
rect 16207 2832 16409 2888
rect 16207 2798 16240 2832
rect 16274 2798 16341 2832
rect 16375 2798 16409 2832
rect 16207 2742 16409 2798
rect 16207 2708 16240 2742
rect 16274 2708 16341 2742
rect 16375 2708 16409 2742
rect 16207 2652 16409 2708
rect 16207 2618 16240 2652
rect 16274 2618 16341 2652
rect 16375 2618 16409 2652
rect 16207 2562 16409 2618
rect 16207 2528 16240 2562
rect 16274 2528 16341 2562
rect 16375 2528 16409 2562
rect 16207 2472 16409 2528
rect 16207 2438 16240 2472
rect 16274 2438 16341 2472
rect 16375 2438 16409 2472
rect 16207 2382 16409 2438
rect 16207 2348 16240 2382
rect 16274 2348 16341 2382
rect 16375 2348 16409 2382
rect 16207 2292 16409 2348
rect 16207 2258 16240 2292
rect 16274 2258 16341 2292
rect 16375 2258 16409 2292
rect 16207 2202 16409 2258
rect 16207 2168 16240 2202
rect 16274 2168 16341 2202
rect 16375 2168 16409 2202
rect 16207 2112 16409 2168
rect 14919 2031 15121 2078
rect 16207 2078 16240 2112
rect 16274 2078 16341 2112
rect 16375 2078 16409 2112
rect 17495 3012 17697 3068
rect 18783 3102 18884 3117
rect 18783 3068 18816 3102
rect 18850 3068 18884 3102
rect 17495 2978 17528 3012
rect 17562 2978 17629 3012
rect 17663 2978 17697 3012
rect 17495 2922 17697 2978
rect 17495 2888 17528 2922
rect 17562 2888 17629 2922
rect 17663 2888 17697 2922
rect 17495 2832 17697 2888
rect 17495 2798 17528 2832
rect 17562 2798 17629 2832
rect 17663 2798 17697 2832
rect 17495 2742 17697 2798
rect 17495 2708 17528 2742
rect 17562 2708 17629 2742
rect 17663 2708 17697 2742
rect 17495 2652 17697 2708
rect 17495 2618 17528 2652
rect 17562 2618 17629 2652
rect 17663 2618 17697 2652
rect 17495 2562 17697 2618
rect 17495 2528 17528 2562
rect 17562 2528 17629 2562
rect 17663 2528 17697 2562
rect 17495 2472 17697 2528
rect 17495 2438 17528 2472
rect 17562 2438 17629 2472
rect 17663 2438 17697 2472
rect 17495 2382 17697 2438
rect 17495 2348 17528 2382
rect 17562 2348 17629 2382
rect 17663 2348 17697 2382
rect 17495 2292 17697 2348
rect 17495 2258 17528 2292
rect 17562 2258 17629 2292
rect 17663 2258 17697 2292
rect 17495 2202 17697 2258
rect 17495 2168 17528 2202
rect 17562 2168 17629 2202
rect 17663 2168 17697 2202
rect 17495 2112 17697 2168
rect 16207 2031 16409 2078
rect 17495 2078 17528 2112
rect 17562 2078 17629 2112
rect 17663 2078 17697 2112
rect 18783 3012 18884 3068
rect 18783 2978 18816 3012
rect 18850 2978 18884 3012
rect 18783 2922 18884 2978
rect 18783 2888 18816 2922
rect 18850 2888 18884 2922
rect 18783 2832 18884 2888
rect 18783 2798 18816 2832
rect 18850 2798 18884 2832
rect 18783 2742 18884 2798
rect 18783 2708 18816 2742
rect 18850 2708 18884 2742
rect 18783 2652 18884 2708
rect 18783 2618 18816 2652
rect 18850 2618 18884 2652
rect 18783 2562 18884 2618
rect 18783 2528 18816 2562
rect 18850 2528 18884 2562
rect 18783 2472 18884 2528
rect 18783 2438 18816 2472
rect 18850 2438 18884 2472
rect 18783 2382 18884 2438
rect 18783 2348 18816 2382
rect 18850 2348 18884 2382
rect 18783 2292 18884 2348
rect 18783 2258 18816 2292
rect 18850 2258 18884 2292
rect 18783 2202 18884 2258
rect 18783 2168 18816 2202
rect 18850 2168 18884 2202
rect 18783 2112 18884 2168
rect 17495 2031 17697 2078
rect 18783 2078 18816 2112
rect 18850 2078 18884 2112
rect 18783 2031 18884 2078
rect 12444 2022 18884 2031
rect 12444 1988 12477 2022
rect 12511 1999 13664 2022
rect 12511 1988 12578 1999
rect 12444 1965 12578 1988
rect 12612 1965 12668 1999
rect 12702 1965 12758 1999
rect 12792 1965 12848 1999
rect 12882 1965 12938 1999
rect 12972 1965 13028 1999
rect 13062 1965 13118 1999
rect 13152 1965 13208 1999
rect 13242 1965 13298 1999
rect 13332 1965 13388 1999
rect 13422 1965 13478 1999
rect 13512 1965 13568 1999
rect 13602 1988 13664 1999
rect 13698 1988 13765 2022
rect 13799 1999 14952 2022
rect 13799 1988 13866 1999
rect 13602 1965 13866 1988
rect 13900 1965 13956 1999
rect 13990 1965 14046 1999
rect 14080 1965 14136 1999
rect 14170 1965 14226 1999
rect 14260 1965 14316 1999
rect 14350 1965 14406 1999
rect 14440 1965 14496 1999
rect 14530 1965 14586 1999
rect 14620 1965 14676 1999
rect 14710 1965 14766 1999
rect 14800 1965 14856 1999
rect 14890 1988 14952 1999
rect 14986 1988 15053 2022
rect 15087 1999 16240 2022
rect 15087 1988 15154 1999
rect 14890 1965 15154 1988
rect 15188 1965 15244 1999
rect 15278 1965 15334 1999
rect 15368 1965 15424 1999
rect 15458 1965 15514 1999
rect 15548 1965 15604 1999
rect 15638 1965 15694 1999
rect 15728 1965 15784 1999
rect 15818 1965 15874 1999
rect 15908 1965 15964 1999
rect 15998 1965 16054 1999
rect 16088 1965 16144 1999
rect 16178 1988 16240 1999
rect 16274 1988 16341 2022
rect 16375 1999 17528 2022
rect 16375 1988 16442 1999
rect 16178 1965 16442 1988
rect 16476 1965 16532 1999
rect 16566 1965 16622 1999
rect 16656 1965 16712 1999
rect 16746 1965 16802 1999
rect 16836 1965 16892 1999
rect 16926 1965 16982 1999
rect 17016 1965 17072 1999
rect 17106 1965 17162 1999
rect 17196 1965 17252 1999
rect 17286 1965 17342 1999
rect 17376 1965 17432 1999
rect 17466 1988 17528 1999
rect 17562 1988 17629 2022
rect 17663 1999 18816 2022
rect 17663 1988 17730 1999
rect 17466 1965 17730 1988
rect 17764 1965 17820 1999
rect 17854 1965 17910 1999
rect 17944 1965 18000 1999
rect 18034 1965 18090 1999
rect 18124 1965 18180 1999
rect 18214 1965 18270 1999
rect 18304 1965 18360 1999
rect 18394 1965 18450 1999
rect 18484 1965 18540 1999
rect 18574 1965 18630 1999
rect 18664 1965 18720 1999
rect 18754 1988 18816 1999
rect 18850 1988 18884 2022
rect 18754 1965 18884 1988
rect 12444 1930 18884 1965
<< nsubdiff >>
rect 12607 12052 13569 12071
rect 12607 12018 12718 12052
rect 12752 12018 12808 12052
rect 12842 12018 12898 12052
rect 12932 12018 12988 12052
rect 13022 12018 13078 12052
rect 13112 12018 13168 12052
rect 13202 12018 13258 12052
rect 13292 12018 13348 12052
rect 13382 12018 13438 12052
rect 13472 12018 13569 12052
rect 12607 11999 13569 12018
rect 12607 11958 12679 11999
rect 12607 11924 12626 11958
rect 12660 11924 12679 11958
rect 13497 11939 13569 11999
rect 12607 11868 12679 11924
rect 12607 11834 12626 11868
rect 12660 11834 12679 11868
rect 12607 11778 12679 11834
rect 12607 11744 12626 11778
rect 12660 11744 12679 11778
rect 12607 11688 12679 11744
rect 12607 11654 12626 11688
rect 12660 11654 12679 11688
rect 12607 11598 12679 11654
rect 12607 11564 12626 11598
rect 12660 11564 12679 11598
rect 12607 11508 12679 11564
rect 12607 11474 12626 11508
rect 12660 11474 12679 11508
rect 12607 11418 12679 11474
rect 12607 11384 12626 11418
rect 12660 11384 12679 11418
rect 12607 11328 12679 11384
rect 12607 11294 12626 11328
rect 12660 11294 12679 11328
rect 12607 11238 12679 11294
rect 13497 11905 13516 11939
rect 13550 11905 13569 11939
rect 13497 11849 13569 11905
rect 13497 11815 13516 11849
rect 13550 11815 13569 11849
rect 13497 11759 13569 11815
rect 13497 11725 13516 11759
rect 13550 11725 13569 11759
rect 13497 11669 13569 11725
rect 13497 11635 13516 11669
rect 13550 11635 13569 11669
rect 13497 11579 13569 11635
rect 13497 11545 13516 11579
rect 13550 11545 13569 11579
rect 13497 11489 13569 11545
rect 13497 11455 13516 11489
rect 13550 11455 13569 11489
rect 13497 11399 13569 11455
rect 13497 11365 13516 11399
rect 13550 11365 13569 11399
rect 13497 11309 13569 11365
rect 13497 11275 13516 11309
rect 13550 11275 13569 11309
rect 12607 11204 12626 11238
rect 12660 11204 12679 11238
rect 12607 11181 12679 11204
rect 13497 11219 13569 11275
rect 13497 11185 13516 11219
rect 13550 11185 13569 11219
rect 13497 11181 13569 11185
rect 12607 11162 13569 11181
rect 12607 11128 12684 11162
rect 12718 11128 12774 11162
rect 12808 11128 12864 11162
rect 12898 11128 12954 11162
rect 12988 11128 13044 11162
rect 13078 11128 13134 11162
rect 13168 11128 13224 11162
rect 13258 11128 13314 11162
rect 13348 11128 13404 11162
rect 13438 11128 13569 11162
rect 12607 11109 13569 11128
rect 13895 12052 14857 12071
rect 13895 12018 14006 12052
rect 14040 12018 14096 12052
rect 14130 12018 14186 12052
rect 14220 12018 14276 12052
rect 14310 12018 14366 12052
rect 14400 12018 14456 12052
rect 14490 12018 14546 12052
rect 14580 12018 14636 12052
rect 14670 12018 14726 12052
rect 14760 12018 14857 12052
rect 13895 11999 14857 12018
rect 13895 11958 13967 11999
rect 13895 11924 13914 11958
rect 13948 11924 13967 11958
rect 14785 11939 14857 11999
rect 13895 11868 13967 11924
rect 13895 11834 13914 11868
rect 13948 11834 13967 11868
rect 13895 11778 13967 11834
rect 13895 11744 13914 11778
rect 13948 11744 13967 11778
rect 13895 11688 13967 11744
rect 13895 11654 13914 11688
rect 13948 11654 13967 11688
rect 13895 11598 13967 11654
rect 13895 11564 13914 11598
rect 13948 11564 13967 11598
rect 13895 11508 13967 11564
rect 13895 11474 13914 11508
rect 13948 11474 13967 11508
rect 13895 11418 13967 11474
rect 13895 11384 13914 11418
rect 13948 11384 13967 11418
rect 13895 11328 13967 11384
rect 13895 11294 13914 11328
rect 13948 11294 13967 11328
rect 13895 11238 13967 11294
rect 14785 11905 14804 11939
rect 14838 11905 14857 11939
rect 14785 11849 14857 11905
rect 14785 11815 14804 11849
rect 14838 11815 14857 11849
rect 14785 11759 14857 11815
rect 14785 11725 14804 11759
rect 14838 11725 14857 11759
rect 14785 11669 14857 11725
rect 14785 11635 14804 11669
rect 14838 11635 14857 11669
rect 14785 11579 14857 11635
rect 14785 11545 14804 11579
rect 14838 11545 14857 11579
rect 14785 11489 14857 11545
rect 14785 11455 14804 11489
rect 14838 11455 14857 11489
rect 14785 11399 14857 11455
rect 14785 11365 14804 11399
rect 14838 11365 14857 11399
rect 14785 11309 14857 11365
rect 14785 11275 14804 11309
rect 14838 11275 14857 11309
rect 13895 11204 13914 11238
rect 13948 11204 13967 11238
rect 13895 11181 13967 11204
rect 14785 11219 14857 11275
rect 14785 11185 14804 11219
rect 14838 11185 14857 11219
rect 14785 11181 14857 11185
rect 13895 11162 14857 11181
rect 13895 11128 13972 11162
rect 14006 11128 14062 11162
rect 14096 11128 14152 11162
rect 14186 11128 14242 11162
rect 14276 11128 14332 11162
rect 14366 11128 14422 11162
rect 14456 11128 14512 11162
rect 14546 11128 14602 11162
rect 14636 11128 14692 11162
rect 14726 11128 14857 11162
rect 13895 11109 14857 11128
rect 15183 12052 16145 12071
rect 15183 12018 15294 12052
rect 15328 12018 15384 12052
rect 15418 12018 15474 12052
rect 15508 12018 15564 12052
rect 15598 12018 15654 12052
rect 15688 12018 15744 12052
rect 15778 12018 15834 12052
rect 15868 12018 15924 12052
rect 15958 12018 16014 12052
rect 16048 12018 16145 12052
rect 15183 11999 16145 12018
rect 15183 11958 15255 11999
rect 15183 11924 15202 11958
rect 15236 11924 15255 11958
rect 16073 11939 16145 11999
rect 15183 11868 15255 11924
rect 15183 11834 15202 11868
rect 15236 11834 15255 11868
rect 15183 11778 15255 11834
rect 15183 11744 15202 11778
rect 15236 11744 15255 11778
rect 15183 11688 15255 11744
rect 15183 11654 15202 11688
rect 15236 11654 15255 11688
rect 15183 11598 15255 11654
rect 15183 11564 15202 11598
rect 15236 11564 15255 11598
rect 15183 11508 15255 11564
rect 15183 11474 15202 11508
rect 15236 11474 15255 11508
rect 15183 11418 15255 11474
rect 15183 11384 15202 11418
rect 15236 11384 15255 11418
rect 15183 11328 15255 11384
rect 15183 11294 15202 11328
rect 15236 11294 15255 11328
rect 15183 11238 15255 11294
rect 16073 11905 16092 11939
rect 16126 11905 16145 11939
rect 16073 11849 16145 11905
rect 16073 11815 16092 11849
rect 16126 11815 16145 11849
rect 16073 11759 16145 11815
rect 16073 11725 16092 11759
rect 16126 11725 16145 11759
rect 16073 11669 16145 11725
rect 16073 11635 16092 11669
rect 16126 11635 16145 11669
rect 16073 11579 16145 11635
rect 16073 11545 16092 11579
rect 16126 11545 16145 11579
rect 16073 11489 16145 11545
rect 16073 11455 16092 11489
rect 16126 11455 16145 11489
rect 16073 11399 16145 11455
rect 16073 11365 16092 11399
rect 16126 11365 16145 11399
rect 16073 11309 16145 11365
rect 16073 11275 16092 11309
rect 16126 11275 16145 11309
rect 15183 11204 15202 11238
rect 15236 11204 15255 11238
rect 15183 11181 15255 11204
rect 16073 11219 16145 11275
rect 16073 11185 16092 11219
rect 16126 11185 16145 11219
rect 16073 11181 16145 11185
rect 15183 11162 16145 11181
rect 15183 11128 15260 11162
rect 15294 11128 15350 11162
rect 15384 11128 15440 11162
rect 15474 11128 15530 11162
rect 15564 11128 15620 11162
rect 15654 11128 15710 11162
rect 15744 11128 15800 11162
rect 15834 11128 15890 11162
rect 15924 11128 15980 11162
rect 16014 11128 16145 11162
rect 15183 11109 16145 11128
rect 16471 12052 17433 12071
rect 16471 12018 16582 12052
rect 16616 12018 16672 12052
rect 16706 12018 16762 12052
rect 16796 12018 16852 12052
rect 16886 12018 16942 12052
rect 16976 12018 17032 12052
rect 17066 12018 17122 12052
rect 17156 12018 17212 12052
rect 17246 12018 17302 12052
rect 17336 12018 17433 12052
rect 16471 11999 17433 12018
rect 16471 11958 16543 11999
rect 16471 11924 16490 11958
rect 16524 11924 16543 11958
rect 17361 11939 17433 11999
rect 16471 11868 16543 11924
rect 16471 11834 16490 11868
rect 16524 11834 16543 11868
rect 16471 11778 16543 11834
rect 16471 11744 16490 11778
rect 16524 11744 16543 11778
rect 16471 11688 16543 11744
rect 16471 11654 16490 11688
rect 16524 11654 16543 11688
rect 16471 11598 16543 11654
rect 16471 11564 16490 11598
rect 16524 11564 16543 11598
rect 16471 11508 16543 11564
rect 16471 11474 16490 11508
rect 16524 11474 16543 11508
rect 16471 11418 16543 11474
rect 16471 11384 16490 11418
rect 16524 11384 16543 11418
rect 16471 11328 16543 11384
rect 16471 11294 16490 11328
rect 16524 11294 16543 11328
rect 16471 11238 16543 11294
rect 17361 11905 17380 11939
rect 17414 11905 17433 11939
rect 17361 11849 17433 11905
rect 17361 11815 17380 11849
rect 17414 11815 17433 11849
rect 17361 11759 17433 11815
rect 17361 11725 17380 11759
rect 17414 11725 17433 11759
rect 17361 11669 17433 11725
rect 17361 11635 17380 11669
rect 17414 11635 17433 11669
rect 17361 11579 17433 11635
rect 17361 11545 17380 11579
rect 17414 11545 17433 11579
rect 17361 11489 17433 11545
rect 17361 11455 17380 11489
rect 17414 11455 17433 11489
rect 17361 11399 17433 11455
rect 17361 11365 17380 11399
rect 17414 11365 17433 11399
rect 17361 11309 17433 11365
rect 17361 11275 17380 11309
rect 17414 11275 17433 11309
rect 16471 11204 16490 11238
rect 16524 11204 16543 11238
rect 16471 11181 16543 11204
rect 17361 11219 17433 11275
rect 17361 11185 17380 11219
rect 17414 11185 17433 11219
rect 17361 11181 17433 11185
rect 16471 11162 17433 11181
rect 16471 11128 16548 11162
rect 16582 11128 16638 11162
rect 16672 11128 16728 11162
rect 16762 11128 16818 11162
rect 16852 11128 16908 11162
rect 16942 11128 16998 11162
rect 17032 11128 17088 11162
rect 17122 11128 17178 11162
rect 17212 11128 17268 11162
rect 17302 11128 17433 11162
rect 16471 11109 17433 11128
rect 17759 12052 18721 12071
rect 17759 12018 17870 12052
rect 17904 12018 17960 12052
rect 17994 12018 18050 12052
rect 18084 12018 18140 12052
rect 18174 12018 18230 12052
rect 18264 12018 18320 12052
rect 18354 12018 18410 12052
rect 18444 12018 18500 12052
rect 18534 12018 18590 12052
rect 18624 12018 18721 12052
rect 17759 11999 18721 12018
rect 17759 11958 17831 11999
rect 17759 11924 17778 11958
rect 17812 11924 17831 11958
rect 18649 11939 18721 11999
rect 17759 11868 17831 11924
rect 17759 11834 17778 11868
rect 17812 11834 17831 11868
rect 17759 11778 17831 11834
rect 17759 11744 17778 11778
rect 17812 11744 17831 11778
rect 17759 11688 17831 11744
rect 17759 11654 17778 11688
rect 17812 11654 17831 11688
rect 17759 11598 17831 11654
rect 17759 11564 17778 11598
rect 17812 11564 17831 11598
rect 17759 11508 17831 11564
rect 17759 11474 17778 11508
rect 17812 11474 17831 11508
rect 17759 11418 17831 11474
rect 17759 11384 17778 11418
rect 17812 11384 17831 11418
rect 17759 11328 17831 11384
rect 17759 11294 17778 11328
rect 17812 11294 17831 11328
rect 17759 11238 17831 11294
rect 18649 11905 18668 11939
rect 18702 11905 18721 11939
rect 18649 11849 18721 11905
rect 18649 11815 18668 11849
rect 18702 11815 18721 11849
rect 18649 11759 18721 11815
rect 18649 11725 18668 11759
rect 18702 11725 18721 11759
rect 18649 11669 18721 11725
rect 18649 11635 18668 11669
rect 18702 11635 18721 11669
rect 18649 11579 18721 11635
rect 18649 11545 18668 11579
rect 18702 11545 18721 11579
rect 18649 11489 18721 11545
rect 18649 11455 18668 11489
rect 18702 11455 18721 11489
rect 18649 11399 18721 11455
rect 18649 11365 18668 11399
rect 18702 11365 18721 11399
rect 18649 11309 18721 11365
rect 18649 11275 18668 11309
rect 18702 11275 18721 11309
rect 17759 11204 17778 11238
rect 17812 11204 17831 11238
rect 17759 11181 17831 11204
rect 18649 11219 18721 11275
rect 18649 11185 18668 11219
rect 18702 11185 18721 11219
rect 18649 11181 18721 11185
rect 17759 11162 18721 11181
rect 17759 11128 17836 11162
rect 17870 11128 17926 11162
rect 17960 11128 18016 11162
rect 18050 11128 18106 11162
rect 18140 11128 18196 11162
rect 18230 11128 18286 11162
rect 18320 11128 18376 11162
rect 18410 11128 18466 11162
rect 18500 11128 18556 11162
rect 18590 11128 18721 11162
rect 17759 11109 18721 11128
rect 12607 10764 13569 10783
rect 12607 10730 12718 10764
rect 12752 10730 12808 10764
rect 12842 10730 12898 10764
rect 12932 10730 12988 10764
rect 13022 10730 13078 10764
rect 13112 10730 13168 10764
rect 13202 10730 13258 10764
rect 13292 10730 13348 10764
rect 13382 10730 13438 10764
rect 13472 10730 13569 10764
rect 12607 10711 13569 10730
rect 12607 10670 12679 10711
rect 12607 10636 12626 10670
rect 12660 10636 12679 10670
rect 13497 10651 13569 10711
rect 12607 10580 12679 10636
rect 12607 10546 12626 10580
rect 12660 10546 12679 10580
rect 12607 10490 12679 10546
rect 12607 10456 12626 10490
rect 12660 10456 12679 10490
rect 12607 10400 12679 10456
rect 12607 10366 12626 10400
rect 12660 10366 12679 10400
rect 12607 10310 12679 10366
rect 12607 10276 12626 10310
rect 12660 10276 12679 10310
rect 12607 10220 12679 10276
rect 12607 10186 12626 10220
rect 12660 10186 12679 10220
rect 12607 10130 12679 10186
rect 12607 10096 12626 10130
rect 12660 10096 12679 10130
rect 12607 10040 12679 10096
rect 12607 10006 12626 10040
rect 12660 10006 12679 10040
rect 12607 9950 12679 10006
rect 13497 10617 13516 10651
rect 13550 10617 13569 10651
rect 13497 10561 13569 10617
rect 13497 10527 13516 10561
rect 13550 10527 13569 10561
rect 13497 10471 13569 10527
rect 13497 10437 13516 10471
rect 13550 10437 13569 10471
rect 13497 10381 13569 10437
rect 13497 10347 13516 10381
rect 13550 10347 13569 10381
rect 13497 10291 13569 10347
rect 13497 10257 13516 10291
rect 13550 10257 13569 10291
rect 13497 10201 13569 10257
rect 13497 10167 13516 10201
rect 13550 10167 13569 10201
rect 13497 10111 13569 10167
rect 13497 10077 13516 10111
rect 13550 10077 13569 10111
rect 13497 10021 13569 10077
rect 13497 9987 13516 10021
rect 13550 9987 13569 10021
rect 12607 9916 12626 9950
rect 12660 9916 12679 9950
rect 12607 9893 12679 9916
rect 13497 9931 13569 9987
rect 13497 9897 13516 9931
rect 13550 9897 13569 9931
rect 13497 9893 13569 9897
rect 12607 9874 13569 9893
rect 12607 9840 12684 9874
rect 12718 9840 12774 9874
rect 12808 9840 12864 9874
rect 12898 9840 12954 9874
rect 12988 9840 13044 9874
rect 13078 9840 13134 9874
rect 13168 9840 13224 9874
rect 13258 9840 13314 9874
rect 13348 9840 13404 9874
rect 13438 9840 13569 9874
rect 12607 9821 13569 9840
rect 13895 10764 14857 10783
rect 13895 10730 14006 10764
rect 14040 10730 14096 10764
rect 14130 10730 14186 10764
rect 14220 10730 14276 10764
rect 14310 10730 14366 10764
rect 14400 10730 14456 10764
rect 14490 10730 14546 10764
rect 14580 10730 14636 10764
rect 14670 10730 14726 10764
rect 14760 10730 14857 10764
rect 13895 10711 14857 10730
rect 13895 10670 13967 10711
rect 13895 10636 13914 10670
rect 13948 10636 13967 10670
rect 14785 10651 14857 10711
rect 13895 10580 13967 10636
rect 13895 10546 13914 10580
rect 13948 10546 13967 10580
rect 13895 10490 13967 10546
rect 13895 10456 13914 10490
rect 13948 10456 13967 10490
rect 13895 10400 13967 10456
rect 13895 10366 13914 10400
rect 13948 10366 13967 10400
rect 13895 10310 13967 10366
rect 13895 10276 13914 10310
rect 13948 10276 13967 10310
rect 13895 10220 13967 10276
rect 13895 10186 13914 10220
rect 13948 10186 13967 10220
rect 13895 10130 13967 10186
rect 13895 10096 13914 10130
rect 13948 10096 13967 10130
rect 13895 10040 13967 10096
rect 13895 10006 13914 10040
rect 13948 10006 13967 10040
rect 13895 9950 13967 10006
rect 14785 10617 14804 10651
rect 14838 10617 14857 10651
rect 14785 10561 14857 10617
rect 14785 10527 14804 10561
rect 14838 10527 14857 10561
rect 14785 10471 14857 10527
rect 14785 10437 14804 10471
rect 14838 10437 14857 10471
rect 14785 10381 14857 10437
rect 14785 10347 14804 10381
rect 14838 10347 14857 10381
rect 14785 10291 14857 10347
rect 14785 10257 14804 10291
rect 14838 10257 14857 10291
rect 14785 10201 14857 10257
rect 14785 10167 14804 10201
rect 14838 10167 14857 10201
rect 14785 10111 14857 10167
rect 14785 10077 14804 10111
rect 14838 10077 14857 10111
rect 14785 10021 14857 10077
rect 14785 9987 14804 10021
rect 14838 9987 14857 10021
rect 13895 9916 13914 9950
rect 13948 9916 13967 9950
rect 13895 9893 13967 9916
rect 14785 9931 14857 9987
rect 14785 9897 14804 9931
rect 14838 9897 14857 9931
rect 14785 9893 14857 9897
rect 13895 9874 14857 9893
rect 13895 9840 13972 9874
rect 14006 9840 14062 9874
rect 14096 9840 14152 9874
rect 14186 9840 14242 9874
rect 14276 9840 14332 9874
rect 14366 9840 14422 9874
rect 14456 9840 14512 9874
rect 14546 9840 14602 9874
rect 14636 9840 14692 9874
rect 14726 9840 14857 9874
rect 13895 9821 14857 9840
rect 15183 10764 16145 10783
rect 15183 10730 15294 10764
rect 15328 10730 15384 10764
rect 15418 10730 15474 10764
rect 15508 10730 15564 10764
rect 15598 10730 15654 10764
rect 15688 10730 15744 10764
rect 15778 10730 15834 10764
rect 15868 10730 15924 10764
rect 15958 10730 16014 10764
rect 16048 10730 16145 10764
rect 15183 10711 16145 10730
rect 15183 10670 15255 10711
rect 15183 10636 15202 10670
rect 15236 10636 15255 10670
rect 16073 10651 16145 10711
rect 15183 10580 15255 10636
rect 15183 10546 15202 10580
rect 15236 10546 15255 10580
rect 15183 10490 15255 10546
rect 15183 10456 15202 10490
rect 15236 10456 15255 10490
rect 15183 10400 15255 10456
rect 15183 10366 15202 10400
rect 15236 10366 15255 10400
rect 15183 10310 15255 10366
rect 15183 10276 15202 10310
rect 15236 10276 15255 10310
rect 15183 10220 15255 10276
rect 15183 10186 15202 10220
rect 15236 10186 15255 10220
rect 15183 10130 15255 10186
rect 15183 10096 15202 10130
rect 15236 10096 15255 10130
rect 15183 10040 15255 10096
rect 15183 10006 15202 10040
rect 15236 10006 15255 10040
rect 15183 9950 15255 10006
rect 16073 10617 16092 10651
rect 16126 10617 16145 10651
rect 16073 10561 16145 10617
rect 16073 10527 16092 10561
rect 16126 10527 16145 10561
rect 16073 10471 16145 10527
rect 16073 10437 16092 10471
rect 16126 10437 16145 10471
rect 16073 10381 16145 10437
rect 16073 10347 16092 10381
rect 16126 10347 16145 10381
rect 16073 10291 16145 10347
rect 16073 10257 16092 10291
rect 16126 10257 16145 10291
rect 16073 10201 16145 10257
rect 16073 10167 16092 10201
rect 16126 10167 16145 10201
rect 16073 10111 16145 10167
rect 16073 10077 16092 10111
rect 16126 10077 16145 10111
rect 16073 10021 16145 10077
rect 16073 9987 16092 10021
rect 16126 9987 16145 10021
rect 15183 9916 15202 9950
rect 15236 9916 15255 9950
rect 15183 9893 15255 9916
rect 16073 9931 16145 9987
rect 16073 9897 16092 9931
rect 16126 9897 16145 9931
rect 16073 9893 16145 9897
rect 15183 9874 16145 9893
rect 15183 9840 15260 9874
rect 15294 9840 15350 9874
rect 15384 9840 15440 9874
rect 15474 9840 15530 9874
rect 15564 9840 15620 9874
rect 15654 9840 15710 9874
rect 15744 9840 15800 9874
rect 15834 9840 15890 9874
rect 15924 9840 15980 9874
rect 16014 9840 16145 9874
rect 15183 9821 16145 9840
rect 16471 10764 17433 10783
rect 16471 10730 16582 10764
rect 16616 10730 16672 10764
rect 16706 10730 16762 10764
rect 16796 10730 16852 10764
rect 16886 10730 16942 10764
rect 16976 10730 17032 10764
rect 17066 10730 17122 10764
rect 17156 10730 17212 10764
rect 17246 10730 17302 10764
rect 17336 10730 17433 10764
rect 16471 10711 17433 10730
rect 16471 10670 16543 10711
rect 16471 10636 16490 10670
rect 16524 10636 16543 10670
rect 17361 10651 17433 10711
rect 16471 10580 16543 10636
rect 16471 10546 16490 10580
rect 16524 10546 16543 10580
rect 16471 10490 16543 10546
rect 16471 10456 16490 10490
rect 16524 10456 16543 10490
rect 16471 10400 16543 10456
rect 16471 10366 16490 10400
rect 16524 10366 16543 10400
rect 16471 10310 16543 10366
rect 16471 10276 16490 10310
rect 16524 10276 16543 10310
rect 16471 10220 16543 10276
rect 16471 10186 16490 10220
rect 16524 10186 16543 10220
rect 16471 10130 16543 10186
rect 16471 10096 16490 10130
rect 16524 10096 16543 10130
rect 16471 10040 16543 10096
rect 16471 10006 16490 10040
rect 16524 10006 16543 10040
rect 16471 9950 16543 10006
rect 17361 10617 17380 10651
rect 17414 10617 17433 10651
rect 17361 10561 17433 10617
rect 17361 10527 17380 10561
rect 17414 10527 17433 10561
rect 17361 10471 17433 10527
rect 17361 10437 17380 10471
rect 17414 10437 17433 10471
rect 17361 10381 17433 10437
rect 17361 10347 17380 10381
rect 17414 10347 17433 10381
rect 17361 10291 17433 10347
rect 17361 10257 17380 10291
rect 17414 10257 17433 10291
rect 17361 10201 17433 10257
rect 17361 10167 17380 10201
rect 17414 10167 17433 10201
rect 17361 10111 17433 10167
rect 17361 10077 17380 10111
rect 17414 10077 17433 10111
rect 17361 10021 17433 10077
rect 17361 9987 17380 10021
rect 17414 9987 17433 10021
rect 16471 9916 16490 9950
rect 16524 9916 16543 9950
rect 16471 9893 16543 9916
rect 17361 9931 17433 9987
rect 17361 9897 17380 9931
rect 17414 9897 17433 9931
rect 17361 9893 17433 9897
rect 16471 9874 17433 9893
rect 16471 9840 16548 9874
rect 16582 9840 16638 9874
rect 16672 9840 16728 9874
rect 16762 9840 16818 9874
rect 16852 9840 16908 9874
rect 16942 9840 16998 9874
rect 17032 9840 17088 9874
rect 17122 9840 17178 9874
rect 17212 9840 17268 9874
rect 17302 9840 17433 9874
rect 16471 9821 17433 9840
rect 17759 10764 18721 10783
rect 17759 10730 17870 10764
rect 17904 10730 17960 10764
rect 17994 10730 18050 10764
rect 18084 10730 18140 10764
rect 18174 10730 18230 10764
rect 18264 10730 18320 10764
rect 18354 10730 18410 10764
rect 18444 10730 18500 10764
rect 18534 10730 18590 10764
rect 18624 10730 18721 10764
rect 17759 10711 18721 10730
rect 17759 10670 17831 10711
rect 17759 10636 17778 10670
rect 17812 10636 17831 10670
rect 18649 10651 18721 10711
rect 17759 10580 17831 10636
rect 17759 10546 17778 10580
rect 17812 10546 17831 10580
rect 17759 10490 17831 10546
rect 17759 10456 17778 10490
rect 17812 10456 17831 10490
rect 17759 10400 17831 10456
rect 17759 10366 17778 10400
rect 17812 10366 17831 10400
rect 17759 10310 17831 10366
rect 17759 10276 17778 10310
rect 17812 10276 17831 10310
rect 17759 10220 17831 10276
rect 17759 10186 17778 10220
rect 17812 10186 17831 10220
rect 17759 10130 17831 10186
rect 17759 10096 17778 10130
rect 17812 10096 17831 10130
rect 17759 10040 17831 10096
rect 17759 10006 17778 10040
rect 17812 10006 17831 10040
rect 17759 9950 17831 10006
rect 18649 10617 18668 10651
rect 18702 10617 18721 10651
rect 18649 10561 18721 10617
rect 18649 10527 18668 10561
rect 18702 10527 18721 10561
rect 18649 10471 18721 10527
rect 18649 10437 18668 10471
rect 18702 10437 18721 10471
rect 18649 10381 18721 10437
rect 18649 10347 18668 10381
rect 18702 10347 18721 10381
rect 18649 10291 18721 10347
rect 18649 10257 18668 10291
rect 18702 10257 18721 10291
rect 18649 10201 18721 10257
rect 18649 10167 18668 10201
rect 18702 10167 18721 10201
rect 18649 10111 18721 10167
rect 18649 10077 18668 10111
rect 18702 10077 18721 10111
rect 18649 10021 18721 10077
rect 18649 9987 18668 10021
rect 18702 9987 18721 10021
rect 17759 9916 17778 9950
rect 17812 9916 17831 9950
rect 17759 9893 17831 9916
rect 18649 9931 18721 9987
rect 18649 9897 18668 9931
rect 18702 9897 18721 9931
rect 18649 9893 18721 9897
rect 17759 9874 18721 9893
rect 17759 9840 17836 9874
rect 17870 9840 17926 9874
rect 17960 9840 18016 9874
rect 18050 9840 18106 9874
rect 18140 9840 18196 9874
rect 18230 9840 18286 9874
rect 18320 9840 18376 9874
rect 18410 9840 18466 9874
rect 18500 9840 18556 9874
rect 18590 9840 18721 9874
rect 17759 9821 18721 9840
rect -9500 9102 -8900 9302
rect -19300 4142 -19100 4242
rect -19300 1800 -19250 4142
rect -19150 1800 -19100 4142
rect -19300 1700 -19100 1800
rect -10172 4142 -9972 4242
rect -10172 1800 -10122 4142
rect -10022 1800 -9972 4142
rect -9500 2102 -9300 9102
rect -9100 2102 -8900 9102
rect -9500 1902 -8900 2102
rect -10172 1700 -9972 1800
rect -3590 9102 -2990 9302
rect -3590 2102 -3390 9102
rect -3190 2102 -2990 9102
rect -3590 1902 -2990 2102
rect 1910 9102 2510 9302
rect 1910 2102 2110 9102
rect 2310 2102 2510 9102
rect 1910 1902 2510 2102
rect 7866 9100 8466 9300
rect 7866 2100 8066 9100
rect 8266 2100 8466 9100
rect 7866 1900 8466 2100
rect 12607 9476 13569 9495
rect 12607 9442 12718 9476
rect 12752 9442 12808 9476
rect 12842 9442 12898 9476
rect 12932 9442 12988 9476
rect 13022 9442 13078 9476
rect 13112 9442 13168 9476
rect 13202 9442 13258 9476
rect 13292 9442 13348 9476
rect 13382 9442 13438 9476
rect 13472 9442 13569 9476
rect 12607 9423 13569 9442
rect 12607 9382 12679 9423
rect 12607 9348 12626 9382
rect 12660 9348 12679 9382
rect 13497 9363 13569 9423
rect 12607 9292 12679 9348
rect 12607 9258 12626 9292
rect 12660 9258 12679 9292
rect 12607 9202 12679 9258
rect 12607 9168 12626 9202
rect 12660 9168 12679 9202
rect 12607 9112 12679 9168
rect 12607 9078 12626 9112
rect 12660 9078 12679 9112
rect 12607 9022 12679 9078
rect 12607 8988 12626 9022
rect 12660 8988 12679 9022
rect 12607 8932 12679 8988
rect 12607 8898 12626 8932
rect 12660 8898 12679 8932
rect 12607 8842 12679 8898
rect 12607 8808 12626 8842
rect 12660 8808 12679 8842
rect 12607 8752 12679 8808
rect 12607 8718 12626 8752
rect 12660 8718 12679 8752
rect 12607 8662 12679 8718
rect 13497 9329 13516 9363
rect 13550 9329 13569 9363
rect 13497 9273 13569 9329
rect 13497 9239 13516 9273
rect 13550 9239 13569 9273
rect 13497 9183 13569 9239
rect 13497 9149 13516 9183
rect 13550 9149 13569 9183
rect 13497 9093 13569 9149
rect 13497 9059 13516 9093
rect 13550 9059 13569 9093
rect 13497 9003 13569 9059
rect 13497 8969 13516 9003
rect 13550 8969 13569 9003
rect 13497 8913 13569 8969
rect 13497 8879 13516 8913
rect 13550 8879 13569 8913
rect 13497 8823 13569 8879
rect 13497 8789 13516 8823
rect 13550 8789 13569 8823
rect 13497 8733 13569 8789
rect 13497 8699 13516 8733
rect 13550 8699 13569 8733
rect 12607 8628 12626 8662
rect 12660 8628 12679 8662
rect 12607 8605 12679 8628
rect 13497 8643 13569 8699
rect 13497 8609 13516 8643
rect 13550 8609 13569 8643
rect 13497 8605 13569 8609
rect 12607 8586 13569 8605
rect 12607 8552 12684 8586
rect 12718 8552 12774 8586
rect 12808 8552 12864 8586
rect 12898 8552 12954 8586
rect 12988 8552 13044 8586
rect 13078 8552 13134 8586
rect 13168 8552 13224 8586
rect 13258 8552 13314 8586
rect 13348 8552 13404 8586
rect 13438 8552 13569 8586
rect 12607 8533 13569 8552
rect 13895 9476 14857 9495
rect 13895 9442 14006 9476
rect 14040 9442 14096 9476
rect 14130 9442 14186 9476
rect 14220 9442 14276 9476
rect 14310 9442 14366 9476
rect 14400 9442 14456 9476
rect 14490 9442 14546 9476
rect 14580 9442 14636 9476
rect 14670 9442 14726 9476
rect 14760 9442 14857 9476
rect 13895 9423 14857 9442
rect 13895 9382 13967 9423
rect 13895 9348 13914 9382
rect 13948 9348 13967 9382
rect 14785 9363 14857 9423
rect 13895 9292 13967 9348
rect 13895 9258 13914 9292
rect 13948 9258 13967 9292
rect 13895 9202 13967 9258
rect 13895 9168 13914 9202
rect 13948 9168 13967 9202
rect 13895 9112 13967 9168
rect 13895 9078 13914 9112
rect 13948 9078 13967 9112
rect 13895 9022 13967 9078
rect 13895 8988 13914 9022
rect 13948 8988 13967 9022
rect 13895 8932 13967 8988
rect 13895 8898 13914 8932
rect 13948 8898 13967 8932
rect 13895 8842 13967 8898
rect 13895 8808 13914 8842
rect 13948 8808 13967 8842
rect 13895 8752 13967 8808
rect 13895 8718 13914 8752
rect 13948 8718 13967 8752
rect 13895 8662 13967 8718
rect 14785 9329 14804 9363
rect 14838 9329 14857 9363
rect 14785 9273 14857 9329
rect 14785 9239 14804 9273
rect 14838 9239 14857 9273
rect 14785 9183 14857 9239
rect 14785 9149 14804 9183
rect 14838 9149 14857 9183
rect 14785 9093 14857 9149
rect 14785 9059 14804 9093
rect 14838 9059 14857 9093
rect 14785 9003 14857 9059
rect 14785 8969 14804 9003
rect 14838 8969 14857 9003
rect 14785 8913 14857 8969
rect 14785 8879 14804 8913
rect 14838 8879 14857 8913
rect 14785 8823 14857 8879
rect 14785 8789 14804 8823
rect 14838 8789 14857 8823
rect 14785 8733 14857 8789
rect 14785 8699 14804 8733
rect 14838 8699 14857 8733
rect 13895 8628 13914 8662
rect 13948 8628 13967 8662
rect 13895 8605 13967 8628
rect 14785 8643 14857 8699
rect 14785 8609 14804 8643
rect 14838 8609 14857 8643
rect 14785 8605 14857 8609
rect 13895 8586 14857 8605
rect 13895 8552 13972 8586
rect 14006 8552 14062 8586
rect 14096 8552 14152 8586
rect 14186 8552 14242 8586
rect 14276 8552 14332 8586
rect 14366 8552 14422 8586
rect 14456 8552 14512 8586
rect 14546 8552 14602 8586
rect 14636 8552 14692 8586
rect 14726 8552 14857 8586
rect 13895 8533 14857 8552
rect 15183 9476 16145 9495
rect 15183 9442 15294 9476
rect 15328 9442 15384 9476
rect 15418 9442 15474 9476
rect 15508 9442 15564 9476
rect 15598 9442 15654 9476
rect 15688 9442 15744 9476
rect 15778 9442 15834 9476
rect 15868 9442 15924 9476
rect 15958 9442 16014 9476
rect 16048 9442 16145 9476
rect 15183 9423 16145 9442
rect 15183 9382 15255 9423
rect 15183 9348 15202 9382
rect 15236 9348 15255 9382
rect 16073 9363 16145 9423
rect 15183 9292 15255 9348
rect 15183 9258 15202 9292
rect 15236 9258 15255 9292
rect 15183 9202 15255 9258
rect 15183 9168 15202 9202
rect 15236 9168 15255 9202
rect 15183 9112 15255 9168
rect 15183 9078 15202 9112
rect 15236 9078 15255 9112
rect 15183 9022 15255 9078
rect 15183 8988 15202 9022
rect 15236 8988 15255 9022
rect 15183 8932 15255 8988
rect 15183 8898 15202 8932
rect 15236 8898 15255 8932
rect 15183 8842 15255 8898
rect 15183 8808 15202 8842
rect 15236 8808 15255 8842
rect 15183 8752 15255 8808
rect 15183 8718 15202 8752
rect 15236 8718 15255 8752
rect 15183 8662 15255 8718
rect 16073 9329 16092 9363
rect 16126 9329 16145 9363
rect 16073 9273 16145 9329
rect 16073 9239 16092 9273
rect 16126 9239 16145 9273
rect 16073 9183 16145 9239
rect 16073 9149 16092 9183
rect 16126 9149 16145 9183
rect 16073 9093 16145 9149
rect 16073 9059 16092 9093
rect 16126 9059 16145 9093
rect 16073 9003 16145 9059
rect 16073 8969 16092 9003
rect 16126 8969 16145 9003
rect 16073 8913 16145 8969
rect 16073 8879 16092 8913
rect 16126 8879 16145 8913
rect 16073 8823 16145 8879
rect 16073 8789 16092 8823
rect 16126 8789 16145 8823
rect 16073 8733 16145 8789
rect 16073 8699 16092 8733
rect 16126 8699 16145 8733
rect 15183 8628 15202 8662
rect 15236 8628 15255 8662
rect 15183 8605 15255 8628
rect 16073 8643 16145 8699
rect 16073 8609 16092 8643
rect 16126 8609 16145 8643
rect 16073 8605 16145 8609
rect 15183 8586 16145 8605
rect 15183 8552 15260 8586
rect 15294 8552 15350 8586
rect 15384 8552 15440 8586
rect 15474 8552 15530 8586
rect 15564 8552 15620 8586
rect 15654 8552 15710 8586
rect 15744 8552 15800 8586
rect 15834 8552 15890 8586
rect 15924 8552 15980 8586
rect 16014 8552 16145 8586
rect 15183 8533 16145 8552
rect 16471 9476 17433 9495
rect 16471 9442 16582 9476
rect 16616 9442 16672 9476
rect 16706 9442 16762 9476
rect 16796 9442 16852 9476
rect 16886 9442 16942 9476
rect 16976 9442 17032 9476
rect 17066 9442 17122 9476
rect 17156 9442 17212 9476
rect 17246 9442 17302 9476
rect 17336 9442 17433 9476
rect 16471 9423 17433 9442
rect 16471 9382 16543 9423
rect 16471 9348 16490 9382
rect 16524 9348 16543 9382
rect 17361 9363 17433 9423
rect 16471 9292 16543 9348
rect 16471 9258 16490 9292
rect 16524 9258 16543 9292
rect 16471 9202 16543 9258
rect 16471 9168 16490 9202
rect 16524 9168 16543 9202
rect 16471 9112 16543 9168
rect 16471 9078 16490 9112
rect 16524 9078 16543 9112
rect 16471 9022 16543 9078
rect 16471 8988 16490 9022
rect 16524 8988 16543 9022
rect 16471 8932 16543 8988
rect 16471 8898 16490 8932
rect 16524 8898 16543 8932
rect 16471 8842 16543 8898
rect 16471 8808 16490 8842
rect 16524 8808 16543 8842
rect 16471 8752 16543 8808
rect 16471 8718 16490 8752
rect 16524 8718 16543 8752
rect 16471 8662 16543 8718
rect 17361 9329 17380 9363
rect 17414 9329 17433 9363
rect 17361 9273 17433 9329
rect 17361 9239 17380 9273
rect 17414 9239 17433 9273
rect 17361 9183 17433 9239
rect 17361 9149 17380 9183
rect 17414 9149 17433 9183
rect 17361 9093 17433 9149
rect 17361 9059 17380 9093
rect 17414 9059 17433 9093
rect 17361 9003 17433 9059
rect 17361 8969 17380 9003
rect 17414 8969 17433 9003
rect 17361 8913 17433 8969
rect 17361 8879 17380 8913
rect 17414 8879 17433 8913
rect 17361 8823 17433 8879
rect 17361 8789 17380 8823
rect 17414 8789 17433 8823
rect 17361 8733 17433 8789
rect 17361 8699 17380 8733
rect 17414 8699 17433 8733
rect 16471 8628 16490 8662
rect 16524 8628 16543 8662
rect 16471 8605 16543 8628
rect 17361 8643 17433 8699
rect 17361 8609 17380 8643
rect 17414 8609 17433 8643
rect 17361 8605 17433 8609
rect 16471 8586 17433 8605
rect 16471 8552 16548 8586
rect 16582 8552 16638 8586
rect 16672 8552 16728 8586
rect 16762 8552 16818 8586
rect 16852 8552 16908 8586
rect 16942 8552 16998 8586
rect 17032 8552 17088 8586
rect 17122 8552 17178 8586
rect 17212 8552 17268 8586
rect 17302 8552 17433 8586
rect 16471 8533 17433 8552
rect 17759 9476 18721 9495
rect 17759 9442 17870 9476
rect 17904 9442 17960 9476
rect 17994 9442 18050 9476
rect 18084 9442 18140 9476
rect 18174 9442 18230 9476
rect 18264 9442 18320 9476
rect 18354 9442 18410 9476
rect 18444 9442 18500 9476
rect 18534 9442 18590 9476
rect 18624 9442 18721 9476
rect 17759 9423 18721 9442
rect 17759 9382 17831 9423
rect 17759 9348 17778 9382
rect 17812 9348 17831 9382
rect 18649 9363 18721 9423
rect 17759 9292 17831 9348
rect 17759 9258 17778 9292
rect 17812 9258 17831 9292
rect 17759 9202 17831 9258
rect 17759 9168 17778 9202
rect 17812 9168 17831 9202
rect 17759 9112 17831 9168
rect 17759 9078 17778 9112
rect 17812 9078 17831 9112
rect 17759 9022 17831 9078
rect 17759 8988 17778 9022
rect 17812 8988 17831 9022
rect 17759 8932 17831 8988
rect 17759 8898 17778 8932
rect 17812 8898 17831 8932
rect 17759 8842 17831 8898
rect 17759 8808 17778 8842
rect 17812 8808 17831 8842
rect 17759 8752 17831 8808
rect 17759 8718 17778 8752
rect 17812 8718 17831 8752
rect 17759 8662 17831 8718
rect 18649 9329 18668 9363
rect 18702 9329 18721 9363
rect 18649 9273 18721 9329
rect 18649 9239 18668 9273
rect 18702 9239 18721 9273
rect 18649 9183 18721 9239
rect 18649 9149 18668 9183
rect 18702 9149 18721 9183
rect 18649 9093 18721 9149
rect 18649 9059 18668 9093
rect 18702 9059 18721 9093
rect 18649 9003 18721 9059
rect 18649 8969 18668 9003
rect 18702 8969 18721 9003
rect 18649 8913 18721 8969
rect 18649 8879 18668 8913
rect 18702 8879 18721 8913
rect 18649 8823 18721 8879
rect 18649 8789 18668 8823
rect 18702 8789 18721 8823
rect 18649 8733 18721 8789
rect 18649 8699 18668 8733
rect 18702 8699 18721 8733
rect 17759 8628 17778 8662
rect 17812 8628 17831 8662
rect 17759 8605 17831 8628
rect 18649 8643 18721 8699
rect 18649 8609 18668 8643
rect 18702 8609 18721 8643
rect 18649 8605 18721 8609
rect 17759 8586 18721 8605
rect 17759 8552 17836 8586
rect 17870 8552 17926 8586
rect 17960 8552 18016 8586
rect 18050 8552 18106 8586
rect 18140 8552 18196 8586
rect 18230 8552 18286 8586
rect 18320 8552 18376 8586
rect 18410 8552 18466 8586
rect 18500 8552 18556 8586
rect 18590 8552 18721 8586
rect 17759 8533 18721 8552
rect 12607 8188 13569 8207
rect 12607 8154 12718 8188
rect 12752 8154 12808 8188
rect 12842 8154 12898 8188
rect 12932 8154 12988 8188
rect 13022 8154 13078 8188
rect 13112 8154 13168 8188
rect 13202 8154 13258 8188
rect 13292 8154 13348 8188
rect 13382 8154 13438 8188
rect 13472 8154 13569 8188
rect 12607 8135 13569 8154
rect 12607 8094 12679 8135
rect 12607 8060 12626 8094
rect 12660 8060 12679 8094
rect 13497 8075 13569 8135
rect 12607 8004 12679 8060
rect 12607 7970 12626 8004
rect 12660 7970 12679 8004
rect 12607 7914 12679 7970
rect 12607 7880 12626 7914
rect 12660 7880 12679 7914
rect 12607 7824 12679 7880
rect 12607 7790 12626 7824
rect 12660 7790 12679 7824
rect 12607 7734 12679 7790
rect 12607 7700 12626 7734
rect 12660 7700 12679 7734
rect 12607 7644 12679 7700
rect 12607 7610 12626 7644
rect 12660 7610 12679 7644
rect 12607 7554 12679 7610
rect 12607 7520 12626 7554
rect 12660 7520 12679 7554
rect 12607 7464 12679 7520
rect 12607 7430 12626 7464
rect 12660 7430 12679 7464
rect 12607 7374 12679 7430
rect 13497 8041 13516 8075
rect 13550 8041 13569 8075
rect 13497 7985 13569 8041
rect 13497 7951 13516 7985
rect 13550 7951 13569 7985
rect 13497 7895 13569 7951
rect 13497 7861 13516 7895
rect 13550 7861 13569 7895
rect 13497 7805 13569 7861
rect 13497 7771 13516 7805
rect 13550 7771 13569 7805
rect 13497 7715 13569 7771
rect 13497 7681 13516 7715
rect 13550 7681 13569 7715
rect 13497 7625 13569 7681
rect 13497 7591 13516 7625
rect 13550 7591 13569 7625
rect 13497 7535 13569 7591
rect 13497 7501 13516 7535
rect 13550 7501 13569 7535
rect 13497 7445 13569 7501
rect 13497 7411 13516 7445
rect 13550 7411 13569 7445
rect 12607 7340 12626 7374
rect 12660 7340 12679 7374
rect 12607 7317 12679 7340
rect 13497 7355 13569 7411
rect 13497 7321 13516 7355
rect 13550 7321 13569 7355
rect 13497 7317 13569 7321
rect 12607 7298 13569 7317
rect 12607 7264 12684 7298
rect 12718 7264 12774 7298
rect 12808 7264 12864 7298
rect 12898 7264 12954 7298
rect 12988 7264 13044 7298
rect 13078 7264 13134 7298
rect 13168 7264 13224 7298
rect 13258 7264 13314 7298
rect 13348 7264 13404 7298
rect 13438 7264 13569 7298
rect 12607 7245 13569 7264
rect 13895 8188 14857 8207
rect 13895 8154 14006 8188
rect 14040 8154 14096 8188
rect 14130 8154 14186 8188
rect 14220 8154 14276 8188
rect 14310 8154 14366 8188
rect 14400 8154 14456 8188
rect 14490 8154 14546 8188
rect 14580 8154 14636 8188
rect 14670 8154 14726 8188
rect 14760 8154 14857 8188
rect 13895 8135 14857 8154
rect 13895 8094 13967 8135
rect 13895 8060 13914 8094
rect 13948 8060 13967 8094
rect 14785 8075 14857 8135
rect 13895 8004 13967 8060
rect 13895 7970 13914 8004
rect 13948 7970 13967 8004
rect 13895 7914 13967 7970
rect 13895 7880 13914 7914
rect 13948 7880 13967 7914
rect 13895 7824 13967 7880
rect 13895 7790 13914 7824
rect 13948 7790 13967 7824
rect 13895 7734 13967 7790
rect 13895 7700 13914 7734
rect 13948 7700 13967 7734
rect 13895 7644 13967 7700
rect 13895 7610 13914 7644
rect 13948 7610 13967 7644
rect 13895 7554 13967 7610
rect 13895 7520 13914 7554
rect 13948 7520 13967 7554
rect 13895 7464 13967 7520
rect 13895 7430 13914 7464
rect 13948 7430 13967 7464
rect 13895 7374 13967 7430
rect 14785 8041 14804 8075
rect 14838 8041 14857 8075
rect 14785 7985 14857 8041
rect 14785 7951 14804 7985
rect 14838 7951 14857 7985
rect 14785 7895 14857 7951
rect 14785 7861 14804 7895
rect 14838 7861 14857 7895
rect 14785 7805 14857 7861
rect 14785 7771 14804 7805
rect 14838 7771 14857 7805
rect 14785 7715 14857 7771
rect 14785 7681 14804 7715
rect 14838 7681 14857 7715
rect 14785 7625 14857 7681
rect 14785 7591 14804 7625
rect 14838 7591 14857 7625
rect 14785 7535 14857 7591
rect 14785 7501 14804 7535
rect 14838 7501 14857 7535
rect 14785 7445 14857 7501
rect 14785 7411 14804 7445
rect 14838 7411 14857 7445
rect 13895 7340 13914 7374
rect 13948 7340 13967 7374
rect 13895 7317 13967 7340
rect 14785 7355 14857 7411
rect 14785 7321 14804 7355
rect 14838 7321 14857 7355
rect 14785 7317 14857 7321
rect 13895 7298 14857 7317
rect 13895 7264 13972 7298
rect 14006 7264 14062 7298
rect 14096 7264 14152 7298
rect 14186 7264 14242 7298
rect 14276 7264 14332 7298
rect 14366 7264 14422 7298
rect 14456 7264 14512 7298
rect 14546 7264 14602 7298
rect 14636 7264 14692 7298
rect 14726 7264 14857 7298
rect 13895 7245 14857 7264
rect 15183 8188 16145 8207
rect 15183 8154 15294 8188
rect 15328 8154 15384 8188
rect 15418 8154 15474 8188
rect 15508 8154 15564 8188
rect 15598 8154 15654 8188
rect 15688 8154 15744 8188
rect 15778 8154 15834 8188
rect 15868 8154 15924 8188
rect 15958 8154 16014 8188
rect 16048 8154 16145 8188
rect 15183 8135 16145 8154
rect 15183 8094 15255 8135
rect 15183 8060 15202 8094
rect 15236 8060 15255 8094
rect 16073 8075 16145 8135
rect 15183 8004 15255 8060
rect 15183 7970 15202 8004
rect 15236 7970 15255 8004
rect 15183 7914 15255 7970
rect 15183 7880 15202 7914
rect 15236 7880 15255 7914
rect 15183 7824 15255 7880
rect 15183 7790 15202 7824
rect 15236 7790 15255 7824
rect 15183 7734 15255 7790
rect 15183 7700 15202 7734
rect 15236 7700 15255 7734
rect 15183 7644 15255 7700
rect 15183 7610 15202 7644
rect 15236 7610 15255 7644
rect 15183 7554 15255 7610
rect 15183 7520 15202 7554
rect 15236 7520 15255 7554
rect 15183 7464 15255 7520
rect 15183 7430 15202 7464
rect 15236 7430 15255 7464
rect 15183 7374 15255 7430
rect 16073 8041 16092 8075
rect 16126 8041 16145 8075
rect 16073 7985 16145 8041
rect 16073 7951 16092 7985
rect 16126 7951 16145 7985
rect 16073 7895 16145 7951
rect 16073 7861 16092 7895
rect 16126 7861 16145 7895
rect 16073 7805 16145 7861
rect 16073 7771 16092 7805
rect 16126 7771 16145 7805
rect 16073 7715 16145 7771
rect 16073 7681 16092 7715
rect 16126 7681 16145 7715
rect 16073 7625 16145 7681
rect 16073 7591 16092 7625
rect 16126 7591 16145 7625
rect 16073 7535 16145 7591
rect 16073 7501 16092 7535
rect 16126 7501 16145 7535
rect 16073 7445 16145 7501
rect 16073 7411 16092 7445
rect 16126 7411 16145 7445
rect 15183 7340 15202 7374
rect 15236 7340 15255 7374
rect 15183 7317 15255 7340
rect 16073 7355 16145 7411
rect 16073 7321 16092 7355
rect 16126 7321 16145 7355
rect 16073 7317 16145 7321
rect 15183 7298 16145 7317
rect 15183 7264 15260 7298
rect 15294 7264 15350 7298
rect 15384 7264 15440 7298
rect 15474 7264 15530 7298
rect 15564 7264 15620 7298
rect 15654 7264 15710 7298
rect 15744 7264 15800 7298
rect 15834 7264 15890 7298
rect 15924 7264 15980 7298
rect 16014 7264 16145 7298
rect 15183 7245 16145 7264
rect 16471 8188 17433 8207
rect 16471 8154 16582 8188
rect 16616 8154 16672 8188
rect 16706 8154 16762 8188
rect 16796 8154 16852 8188
rect 16886 8154 16942 8188
rect 16976 8154 17032 8188
rect 17066 8154 17122 8188
rect 17156 8154 17212 8188
rect 17246 8154 17302 8188
rect 17336 8154 17433 8188
rect 16471 8135 17433 8154
rect 16471 8094 16543 8135
rect 16471 8060 16490 8094
rect 16524 8060 16543 8094
rect 17361 8075 17433 8135
rect 16471 8004 16543 8060
rect 16471 7970 16490 8004
rect 16524 7970 16543 8004
rect 16471 7914 16543 7970
rect 16471 7880 16490 7914
rect 16524 7880 16543 7914
rect 16471 7824 16543 7880
rect 16471 7790 16490 7824
rect 16524 7790 16543 7824
rect 16471 7734 16543 7790
rect 16471 7700 16490 7734
rect 16524 7700 16543 7734
rect 16471 7644 16543 7700
rect 16471 7610 16490 7644
rect 16524 7610 16543 7644
rect 16471 7554 16543 7610
rect 16471 7520 16490 7554
rect 16524 7520 16543 7554
rect 16471 7464 16543 7520
rect 16471 7430 16490 7464
rect 16524 7430 16543 7464
rect 16471 7374 16543 7430
rect 17361 8041 17380 8075
rect 17414 8041 17433 8075
rect 17361 7985 17433 8041
rect 17361 7951 17380 7985
rect 17414 7951 17433 7985
rect 17361 7895 17433 7951
rect 17361 7861 17380 7895
rect 17414 7861 17433 7895
rect 17361 7805 17433 7861
rect 17361 7771 17380 7805
rect 17414 7771 17433 7805
rect 17361 7715 17433 7771
rect 17361 7681 17380 7715
rect 17414 7681 17433 7715
rect 17361 7625 17433 7681
rect 17361 7591 17380 7625
rect 17414 7591 17433 7625
rect 17361 7535 17433 7591
rect 17361 7501 17380 7535
rect 17414 7501 17433 7535
rect 17361 7445 17433 7501
rect 17361 7411 17380 7445
rect 17414 7411 17433 7445
rect 16471 7340 16490 7374
rect 16524 7340 16543 7374
rect 16471 7317 16543 7340
rect 17361 7355 17433 7411
rect 17361 7321 17380 7355
rect 17414 7321 17433 7355
rect 17361 7317 17433 7321
rect 16471 7298 17433 7317
rect 16471 7264 16548 7298
rect 16582 7264 16638 7298
rect 16672 7264 16728 7298
rect 16762 7264 16818 7298
rect 16852 7264 16908 7298
rect 16942 7264 16998 7298
rect 17032 7264 17088 7298
rect 17122 7264 17178 7298
rect 17212 7264 17268 7298
rect 17302 7264 17433 7298
rect 16471 7245 17433 7264
rect 17759 8188 18721 8207
rect 17759 8154 17870 8188
rect 17904 8154 17960 8188
rect 17994 8154 18050 8188
rect 18084 8154 18140 8188
rect 18174 8154 18230 8188
rect 18264 8154 18320 8188
rect 18354 8154 18410 8188
rect 18444 8154 18500 8188
rect 18534 8154 18590 8188
rect 18624 8154 18721 8188
rect 17759 8135 18721 8154
rect 17759 8094 17831 8135
rect 17759 8060 17778 8094
rect 17812 8060 17831 8094
rect 18649 8075 18721 8135
rect 17759 8004 17831 8060
rect 17759 7970 17778 8004
rect 17812 7970 17831 8004
rect 17759 7914 17831 7970
rect 17759 7880 17778 7914
rect 17812 7880 17831 7914
rect 17759 7824 17831 7880
rect 17759 7790 17778 7824
rect 17812 7790 17831 7824
rect 17759 7734 17831 7790
rect 17759 7700 17778 7734
rect 17812 7700 17831 7734
rect 17759 7644 17831 7700
rect 17759 7610 17778 7644
rect 17812 7610 17831 7644
rect 17759 7554 17831 7610
rect 17759 7520 17778 7554
rect 17812 7520 17831 7554
rect 17759 7464 17831 7520
rect 17759 7430 17778 7464
rect 17812 7430 17831 7464
rect 17759 7374 17831 7430
rect 18649 8041 18668 8075
rect 18702 8041 18721 8075
rect 18649 7985 18721 8041
rect 18649 7951 18668 7985
rect 18702 7951 18721 7985
rect 18649 7895 18721 7951
rect 18649 7861 18668 7895
rect 18702 7861 18721 7895
rect 18649 7805 18721 7861
rect 18649 7771 18668 7805
rect 18702 7771 18721 7805
rect 18649 7715 18721 7771
rect 18649 7681 18668 7715
rect 18702 7681 18721 7715
rect 18649 7625 18721 7681
rect 18649 7591 18668 7625
rect 18702 7591 18721 7625
rect 18649 7535 18721 7591
rect 18649 7501 18668 7535
rect 18702 7501 18721 7535
rect 18649 7445 18721 7501
rect 18649 7411 18668 7445
rect 18702 7411 18721 7445
rect 17759 7340 17778 7374
rect 17812 7340 17831 7374
rect 17759 7317 17831 7340
rect 18649 7355 18721 7411
rect 18649 7321 18668 7355
rect 18702 7321 18721 7355
rect 18649 7317 18721 7321
rect 17759 7298 18721 7317
rect 17759 7264 17836 7298
rect 17870 7264 17926 7298
rect 17960 7264 18016 7298
rect 18050 7264 18106 7298
rect 18140 7264 18196 7298
rect 18230 7264 18286 7298
rect 18320 7264 18376 7298
rect 18410 7264 18466 7298
rect 18500 7264 18556 7298
rect 18590 7264 18721 7298
rect 17759 7245 18721 7264
rect 12607 6900 13569 6919
rect 12607 6866 12718 6900
rect 12752 6866 12808 6900
rect 12842 6866 12898 6900
rect 12932 6866 12988 6900
rect 13022 6866 13078 6900
rect 13112 6866 13168 6900
rect 13202 6866 13258 6900
rect 13292 6866 13348 6900
rect 13382 6866 13438 6900
rect 13472 6866 13569 6900
rect 12607 6847 13569 6866
rect 12607 6806 12679 6847
rect 12607 6772 12626 6806
rect 12660 6772 12679 6806
rect 13497 6787 13569 6847
rect 12607 6716 12679 6772
rect 12607 6682 12626 6716
rect 12660 6682 12679 6716
rect 12607 6626 12679 6682
rect 12607 6592 12626 6626
rect 12660 6592 12679 6626
rect 12607 6536 12679 6592
rect 12607 6502 12626 6536
rect 12660 6502 12679 6536
rect 12607 6446 12679 6502
rect 12607 6412 12626 6446
rect 12660 6412 12679 6446
rect 12607 6356 12679 6412
rect 12607 6322 12626 6356
rect 12660 6322 12679 6356
rect 12607 6266 12679 6322
rect 12607 6232 12626 6266
rect 12660 6232 12679 6266
rect 12607 6176 12679 6232
rect 12607 6142 12626 6176
rect 12660 6142 12679 6176
rect 12607 6086 12679 6142
rect 13497 6753 13516 6787
rect 13550 6753 13569 6787
rect 13497 6697 13569 6753
rect 13497 6663 13516 6697
rect 13550 6663 13569 6697
rect 13497 6607 13569 6663
rect 13497 6573 13516 6607
rect 13550 6573 13569 6607
rect 13497 6517 13569 6573
rect 13497 6483 13516 6517
rect 13550 6483 13569 6517
rect 13497 6427 13569 6483
rect 13497 6393 13516 6427
rect 13550 6393 13569 6427
rect 13497 6337 13569 6393
rect 13497 6303 13516 6337
rect 13550 6303 13569 6337
rect 13497 6247 13569 6303
rect 13497 6213 13516 6247
rect 13550 6213 13569 6247
rect 13497 6157 13569 6213
rect 13497 6123 13516 6157
rect 13550 6123 13569 6157
rect 12607 6052 12626 6086
rect 12660 6052 12679 6086
rect 12607 6029 12679 6052
rect 13497 6067 13569 6123
rect 13497 6033 13516 6067
rect 13550 6033 13569 6067
rect 13497 6029 13569 6033
rect 12607 6010 13569 6029
rect 12607 5976 12684 6010
rect 12718 5976 12774 6010
rect 12808 5976 12864 6010
rect 12898 5976 12954 6010
rect 12988 5976 13044 6010
rect 13078 5976 13134 6010
rect 13168 5976 13224 6010
rect 13258 5976 13314 6010
rect 13348 5976 13404 6010
rect 13438 5976 13569 6010
rect 12607 5957 13569 5976
rect 13895 6900 14857 6919
rect 13895 6866 14006 6900
rect 14040 6866 14096 6900
rect 14130 6866 14186 6900
rect 14220 6866 14276 6900
rect 14310 6866 14366 6900
rect 14400 6866 14456 6900
rect 14490 6866 14546 6900
rect 14580 6866 14636 6900
rect 14670 6866 14726 6900
rect 14760 6866 14857 6900
rect 13895 6847 14857 6866
rect 13895 6806 13967 6847
rect 13895 6772 13914 6806
rect 13948 6772 13967 6806
rect 14785 6787 14857 6847
rect 13895 6716 13967 6772
rect 13895 6682 13914 6716
rect 13948 6682 13967 6716
rect 13895 6626 13967 6682
rect 13895 6592 13914 6626
rect 13948 6592 13967 6626
rect 13895 6536 13967 6592
rect 13895 6502 13914 6536
rect 13948 6502 13967 6536
rect 13895 6446 13967 6502
rect 13895 6412 13914 6446
rect 13948 6412 13967 6446
rect 13895 6356 13967 6412
rect 13895 6322 13914 6356
rect 13948 6322 13967 6356
rect 13895 6266 13967 6322
rect 13895 6232 13914 6266
rect 13948 6232 13967 6266
rect 13895 6176 13967 6232
rect 13895 6142 13914 6176
rect 13948 6142 13967 6176
rect 13895 6086 13967 6142
rect 14785 6753 14804 6787
rect 14838 6753 14857 6787
rect 14785 6697 14857 6753
rect 14785 6663 14804 6697
rect 14838 6663 14857 6697
rect 14785 6607 14857 6663
rect 14785 6573 14804 6607
rect 14838 6573 14857 6607
rect 14785 6517 14857 6573
rect 14785 6483 14804 6517
rect 14838 6483 14857 6517
rect 14785 6427 14857 6483
rect 14785 6393 14804 6427
rect 14838 6393 14857 6427
rect 14785 6337 14857 6393
rect 14785 6303 14804 6337
rect 14838 6303 14857 6337
rect 14785 6247 14857 6303
rect 14785 6213 14804 6247
rect 14838 6213 14857 6247
rect 14785 6157 14857 6213
rect 14785 6123 14804 6157
rect 14838 6123 14857 6157
rect 13895 6052 13914 6086
rect 13948 6052 13967 6086
rect 13895 6029 13967 6052
rect 14785 6067 14857 6123
rect 14785 6033 14804 6067
rect 14838 6033 14857 6067
rect 14785 6029 14857 6033
rect 13895 6010 14857 6029
rect 13895 5976 13972 6010
rect 14006 5976 14062 6010
rect 14096 5976 14152 6010
rect 14186 5976 14242 6010
rect 14276 5976 14332 6010
rect 14366 5976 14422 6010
rect 14456 5976 14512 6010
rect 14546 5976 14602 6010
rect 14636 5976 14692 6010
rect 14726 5976 14857 6010
rect 13895 5957 14857 5976
rect 15183 6900 16145 6919
rect 15183 6866 15294 6900
rect 15328 6866 15384 6900
rect 15418 6866 15474 6900
rect 15508 6866 15564 6900
rect 15598 6866 15654 6900
rect 15688 6866 15744 6900
rect 15778 6866 15834 6900
rect 15868 6866 15924 6900
rect 15958 6866 16014 6900
rect 16048 6866 16145 6900
rect 15183 6847 16145 6866
rect 15183 6806 15255 6847
rect 15183 6772 15202 6806
rect 15236 6772 15255 6806
rect 16073 6787 16145 6847
rect 15183 6716 15255 6772
rect 15183 6682 15202 6716
rect 15236 6682 15255 6716
rect 15183 6626 15255 6682
rect 15183 6592 15202 6626
rect 15236 6592 15255 6626
rect 15183 6536 15255 6592
rect 15183 6502 15202 6536
rect 15236 6502 15255 6536
rect 15183 6446 15255 6502
rect 15183 6412 15202 6446
rect 15236 6412 15255 6446
rect 15183 6356 15255 6412
rect 15183 6322 15202 6356
rect 15236 6322 15255 6356
rect 15183 6266 15255 6322
rect 15183 6232 15202 6266
rect 15236 6232 15255 6266
rect 15183 6176 15255 6232
rect 15183 6142 15202 6176
rect 15236 6142 15255 6176
rect 15183 6086 15255 6142
rect 16073 6753 16092 6787
rect 16126 6753 16145 6787
rect 16073 6697 16145 6753
rect 16073 6663 16092 6697
rect 16126 6663 16145 6697
rect 16073 6607 16145 6663
rect 16073 6573 16092 6607
rect 16126 6573 16145 6607
rect 16073 6517 16145 6573
rect 16073 6483 16092 6517
rect 16126 6483 16145 6517
rect 16073 6427 16145 6483
rect 16073 6393 16092 6427
rect 16126 6393 16145 6427
rect 16073 6337 16145 6393
rect 16073 6303 16092 6337
rect 16126 6303 16145 6337
rect 16073 6247 16145 6303
rect 16073 6213 16092 6247
rect 16126 6213 16145 6247
rect 16073 6157 16145 6213
rect 16073 6123 16092 6157
rect 16126 6123 16145 6157
rect 15183 6052 15202 6086
rect 15236 6052 15255 6086
rect 15183 6029 15255 6052
rect 16073 6067 16145 6123
rect 16073 6033 16092 6067
rect 16126 6033 16145 6067
rect 16073 6029 16145 6033
rect 15183 6010 16145 6029
rect 15183 5976 15260 6010
rect 15294 5976 15350 6010
rect 15384 5976 15440 6010
rect 15474 5976 15530 6010
rect 15564 5976 15620 6010
rect 15654 5976 15710 6010
rect 15744 5976 15800 6010
rect 15834 5976 15890 6010
rect 15924 5976 15980 6010
rect 16014 5976 16145 6010
rect 15183 5957 16145 5976
rect 16471 6900 17433 6919
rect 16471 6866 16582 6900
rect 16616 6866 16672 6900
rect 16706 6866 16762 6900
rect 16796 6866 16852 6900
rect 16886 6866 16942 6900
rect 16976 6866 17032 6900
rect 17066 6866 17122 6900
rect 17156 6866 17212 6900
rect 17246 6866 17302 6900
rect 17336 6866 17433 6900
rect 16471 6847 17433 6866
rect 16471 6806 16543 6847
rect 16471 6772 16490 6806
rect 16524 6772 16543 6806
rect 17361 6787 17433 6847
rect 16471 6716 16543 6772
rect 16471 6682 16490 6716
rect 16524 6682 16543 6716
rect 16471 6626 16543 6682
rect 16471 6592 16490 6626
rect 16524 6592 16543 6626
rect 16471 6536 16543 6592
rect 16471 6502 16490 6536
rect 16524 6502 16543 6536
rect 16471 6446 16543 6502
rect 16471 6412 16490 6446
rect 16524 6412 16543 6446
rect 16471 6356 16543 6412
rect 16471 6322 16490 6356
rect 16524 6322 16543 6356
rect 16471 6266 16543 6322
rect 16471 6232 16490 6266
rect 16524 6232 16543 6266
rect 16471 6176 16543 6232
rect 16471 6142 16490 6176
rect 16524 6142 16543 6176
rect 16471 6086 16543 6142
rect 17361 6753 17380 6787
rect 17414 6753 17433 6787
rect 17361 6697 17433 6753
rect 17361 6663 17380 6697
rect 17414 6663 17433 6697
rect 17361 6607 17433 6663
rect 17361 6573 17380 6607
rect 17414 6573 17433 6607
rect 17361 6517 17433 6573
rect 17361 6483 17380 6517
rect 17414 6483 17433 6517
rect 17361 6427 17433 6483
rect 17361 6393 17380 6427
rect 17414 6393 17433 6427
rect 17361 6337 17433 6393
rect 17361 6303 17380 6337
rect 17414 6303 17433 6337
rect 17361 6247 17433 6303
rect 17361 6213 17380 6247
rect 17414 6213 17433 6247
rect 17361 6157 17433 6213
rect 17361 6123 17380 6157
rect 17414 6123 17433 6157
rect 16471 6052 16490 6086
rect 16524 6052 16543 6086
rect 16471 6029 16543 6052
rect 17361 6067 17433 6123
rect 17361 6033 17380 6067
rect 17414 6033 17433 6067
rect 17361 6029 17433 6033
rect 16471 6010 17433 6029
rect 16471 5976 16548 6010
rect 16582 5976 16638 6010
rect 16672 5976 16728 6010
rect 16762 5976 16818 6010
rect 16852 5976 16908 6010
rect 16942 5976 16998 6010
rect 17032 5976 17088 6010
rect 17122 5976 17178 6010
rect 17212 5976 17268 6010
rect 17302 5976 17433 6010
rect 16471 5957 17433 5976
rect 17759 6900 18721 6919
rect 17759 6866 17870 6900
rect 17904 6866 17960 6900
rect 17994 6866 18050 6900
rect 18084 6866 18140 6900
rect 18174 6866 18230 6900
rect 18264 6866 18320 6900
rect 18354 6866 18410 6900
rect 18444 6866 18500 6900
rect 18534 6866 18590 6900
rect 18624 6866 18721 6900
rect 17759 6847 18721 6866
rect 17759 6806 17831 6847
rect 17759 6772 17778 6806
rect 17812 6772 17831 6806
rect 18649 6787 18721 6847
rect 17759 6716 17831 6772
rect 17759 6682 17778 6716
rect 17812 6682 17831 6716
rect 17759 6626 17831 6682
rect 17759 6592 17778 6626
rect 17812 6592 17831 6626
rect 17759 6536 17831 6592
rect 17759 6502 17778 6536
rect 17812 6502 17831 6536
rect 17759 6446 17831 6502
rect 17759 6412 17778 6446
rect 17812 6412 17831 6446
rect 17759 6356 17831 6412
rect 17759 6322 17778 6356
rect 17812 6322 17831 6356
rect 17759 6266 17831 6322
rect 17759 6232 17778 6266
rect 17812 6232 17831 6266
rect 17759 6176 17831 6232
rect 17759 6142 17778 6176
rect 17812 6142 17831 6176
rect 17759 6086 17831 6142
rect 18649 6753 18668 6787
rect 18702 6753 18721 6787
rect 18649 6697 18721 6753
rect 18649 6663 18668 6697
rect 18702 6663 18721 6697
rect 18649 6607 18721 6663
rect 18649 6573 18668 6607
rect 18702 6573 18721 6607
rect 18649 6517 18721 6573
rect 18649 6483 18668 6517
rect 18702 6483 18721 6517
rect 18649 6427 18721 6483
rect 18649 6393 18668 6427
rect 18702 6393 18721 6427
rect 18649 6337 18721 6393
rect 18649 6303 18668 6337
rect 18702 6303 18721 6337
rect 18649 6247 18721 6303
rect 18649 6213 18668 6247
rect 18702 6213 18721 6247
rect 18649 6157 18721 6213
rect 18649 6123 18668 6157
rect 18702 6123 18721 6157
rect 17759 6052 17778 6086
rect 17812 6052 17831 6086
rect 17759 6029 17831 6052
rect 18649 6067 18721 6123
rect 18649 6033 18668 6067
rect 18702 6033 18721 6067
rect 18649 6029 18721 6033
rect 17759 6010 18721 6029
rect 17759 5976 17836 6010
rect 17870 5976 17926 6010
rect 17960 5976 18016 6010
rect 18050 5976 18106 6010
rect 18140 5976 18196 6010
rect 18230 5976 18286 6010
rect 18320 5976 18376 6010
rect 18410 5976 18466 6010
rect 18500 5976 18556 6010
rect 18590 5976 18721 6010
rect 17759 5957 18721 5976
rect 12607 5612 13569 5631
rect 12607 5578 12718 5612
rect 12752 5578 12808 5612
rect 12842 5578 12898 5612
rect 12932 5578 12988 5612
rect 13022 5578 13078 5612
rect 13112 5578 13168 5612
rect 13202 5578 13258 5612
rect 13292 5578 13348 5612
rect 13382 5578 13438 5612
rect 13472 5578 13569 5612
rect 12607 5559 13569 5578
rect 12607 5518 12679 5559
rect 12607 5484 12626 5518
rect 12660 5484 12679 5518
rect 13497 5499 13569 5559
rect 12607 5428 12679 5484
rect 12607 5394 12626 5428
rect 12660 5394 12679 5428
rect 12607 5338 12679 5394
rect 12607 5304 12626 5338
rect 12660 5304 12679 5338
rect 12607 5248 12679 5304
rect 12607 5214 12626 5248
rect 12660 5214 12679 5248
rect 12607 5158 12679 5214
rect 12607 5124 12626 5158
rect 12660 5124 12679 5158
rect 12607 5068 12679 5124
rect 12607 5034 12626 5068
rect 12660 5034 12679 5068
rect 12607 4978 12679 5034
rect 12607 4944 12626 4978
rect 12660 4944 12679 4978
rect 12607 4888 12679 4944
rect 12607 4854 12626 4888
rect 12660 4854 12679 4888
rect 12607 4798 12679 4854
rect 13497 5465 13516 5499
rect 13550 5465 13569 5499
rect 13497 5409 13569 5465
rect 13497 5375 13516 5409
rect 13550 5375 13569 5409
rect 13497 5319 13569 5375
rect 13497 5285 13516 5319
rect 13550 5285 13569 5319
rect 13497 5229 13569 5285
rect 13497 5195 13516 5229
rect 13550 5195 13569 5229
rect 13497 5139 13569 5195
rect 13497 5105 13516 5139
rect 13550 5105 13569 5139
rect 13497 5049 13569 5105
rect 13497 5015 13516 5049
rect 13550 5015 13569 5049
rect 13497 4959 13569 5015
rect 13497 4925 13516 4959
rect 13550 4925 13569 4959
rect 13497 4869 13569 4925
rect 13497 4835 13516 4869
rect 13550 4835 13569 4869
rect 12607 4764 12626 4798
rect 12660 4764 12679 4798
rect 12607 4741 12679 4764
rect 13497 4779 13569 4835
rect 13497 4745 13516 4779
rect 13550 4745 13569 4779
rect 13497 4741 13569 4745
rect 12607 4722 13569 4741
rect 12607 4688 12684 4722
rect 12718 4688 12774 4722
rect 12808 4688 12864 4722
rect 12898 4688 12954 4722
rect 12988 4688 13044 4722
rect 13078 4688 13134 4722
rect 13168 4688 13224 4722
rect 13258 4688 13314 4722
rect 13348 4688 13404 4722
rect 13438 4688 13569 4722
rect 12607 4669 13569 4688
rect 13895 5612 14857 5631
rect 13895 5578 14006 5612
rect 14040 5578 14096 5612
rect 14130 5578 14186 5612
rect 14220 5578 14276 5612
rect 14310 5578 14366 5612
rect 14400 5578 14456 5612
rect 14490 5578 14546 5612
rect 14580 5578 14636 5612
rect 14670 5578 14726 5612
rect 14760 5578 14857 5612
rect 13895 5559 14857 5578
rect 13895 5518 13967 5559
rect 13895 5484 13914 5518
rect 13948 5484 13967 5518
rect 14785 5499 14857 5559
rect 13895 5428 13967 5484
rect 13895 5394 13914 5428
rect 13948 5394 13967 5428
rect 13895 5338 13967 5394
rect 13895 5304 13914 5338
rect 13948 5304 13967 5338
rect 13895 5248 13967 5304
rect 13895 5214 13914 5248
rect 13948 5214 13967 5248
rect 13895 5158 13967 5214
rect 13895 5124 13914 5158
rect 13948 5124 13967 5158
rect 13895 5068 13967 5124
rect 13895 5034 13914 5068
rect 13948 5034 13967 5068
rect 13895 4978 13967 5034
rect 13895 4944 13914 4978
rect 13948 4944 13967 4978
rect 13895 4888 13967 4944
rect 13895 4854 13914 4888
rect 13948 4854 13967 4888
rect 13895 4798 13967 4854
rect 14785 5465 14804 5499
rect 14838 5465 14857 5499
rect 14785 5409 14857 5465
rect 14785 5375 14804 5409
rect 14838 5375 14857 5409
rect 14785 5319 14857 5375
rect 14785 5285 14804 5319
rect 14838 5285 14857 5319
rect 14785 5229 14857 5285
rect 14785 5195 14804 5229
rect 14838 5195 14857 5229
rect 14785 5139 14857 5195
rect 14785 5105 14804 5139
rect 14838 5105 14857 5139
rect 14785 5049 14857 5105
rect 14785 5015 14804 5049
rect 14838 5015 14857 5049
rect 14785 4959 14857 5015
rect 14785 4925 14804 4959
rect 14838 4925 14857 4959
rect 14785 4869 14857 4925
rect 14785 4835 14804 4869
rect 14838 4835 14857 4869
rect 13895 4764 13914 4798
rect 13948 4764 13967 4798
rect 13895 4741 13967 4764
rect 14785 4779 14857 4835
rect 14785 4745 14804 4779
rect 14838 4745 14857 4779
rect 14785 4741 14857 4745
rect 13895 4722 14857 4741
rect 13895 4688 13972 4722
rect 14006 4688 14062 4722
rect 14096 4688 14152 4722
rect 14186 4688 14242 4722
rect 14276 4688 14332 4722
rect 14366 4688 14422 4722
rect 14456 4688 14512 4722
rect 14546 4688 14602 4722
rect 14636 4688 14692 4722
rect 14726 4688 14857 4722
rect 13895 4669 14857 4688
rect 15183 5612 16145 5631
rect 15183 5578 15294 5612
rect 15328 5578 15384 5612
rect 15418 5578 15474 5612
rect 15508 5578 15564 5612
rect 15598 5578 15654 5612
rect 15688 5578 15744 5612
rect 15778 5578 15834 5612
rect 15868 5578 15924 5612
rect 15958 5578 16014 5612
rect 16048 5578 16145 5612
rect 15183 5559 16145 5578
rect 15183 5518 15255 5559
rect 15183 5484 15202 5518
rect 15236 5484 15255 5518
rect 16073 5499 16145 5559
rect 15183 5428 15255 5484
rect 15183 5394 15202 5428
rect 15236 5394 15255 5428
rect 15183 5338 15255 5394
rect 15183 5304 15202 5338
rect 15236 5304 15255 5338
rect 15183 5248 15255 5304
rect 15183 5214 15202 5248
rect 15236 5214 15255 5248
rect 15183 5158 15255 5214
rect 15183 5124 15202 5158
rect 15236 5124 15255 5158
rect 15183 5068 15255 5124
rect 15183 5034 15202 5068
rect 15236 5034 15255 5068
rect 15183 4978 15255 5034
rect 15183 4944 15202 4978
rect 15236 4944 15255 4978
rect 15183 4888 15255 4944
rect 15183 4854 15202 4888
rect 15236 4854 15255 4888
rect 15183 4798 15255 4854
rect 16073 5465 16092 5499
rect 16126 5465 16145 5499
rect 16073 5409 16145 5465
rect 16073 5375 16092 5409
rect 16126 5375 16145 5409
rect 16073 5319 16145 5375
rect 16073 5285 16092 5319
rect 16126 5285 16145 5319
rect 16073 5229 16145 5285
rect 16073 5195 16092 5229
rect 16126 5195 16145 5229
rect 16073 5139 16145 5195
rect 16073 5105 16092 5139
rect 16126 5105 16145 5139
rect 16073 5049 16145 5105
rect 16073 5015 16092 5049
rect 16126 5015 16145 5049
rect 16073 4959 16145 5015
rect 16073 4925 16092 4959
rect 16126 4925 16145 4959
rect 16073 4869 16145 4925
rect 16073 4835 16092 4869
rect 16126 4835 16145 4869
rect 15183 4764 15202 4798
rect 15236 4764 15255 4798
rect 15183 4741 15255 4764
rect 16073 4779 16145 4835
rect 16073 4745 16092 4779
rect 16126 4745 16145 4779
rect 16073 4741 16145 4745
rect 15183 4722 16145 4741
rect 15183 4688 15260 4722
rect 15294 4688 15350 4722
rect 15384 4688 15440 4722
rect 15474 4688 15530 4722
rect 15564 4688 15620 4722
rect 15654 4688 15710 4722
rect 15744 4688 15800 4722
rect 15834 4688 15890 4722
rect 15924 4688 15980 4722
rect 16014 4688 16145 4722
rect 15183 4669 16145 4688
rect 16471 5612 17433 5631
rect 16471 5578 16582 5612
rect 16616 5578 16672 5612
rect 16706 5578 16762 5612
rect 16796 5578 16852 5612
rect 16886 5578 16942 5612
rect 16976 5578 17032 5612
rect 17066 5578 17122 5612
rect 17156 5578 17212 5612
rect 17246 5578 17302 5612
rect 17336 5578 17433 5612
rect 16471 5559 17433 5578
rect 16471 5518 16543 5559
rect 16471 5484 16490 5518
rect 16524 5484 16543 5518
rect 17361 5499 17433 5559
rect 16471 5428 16543 5484
rect 16471 5394 16490 5428
rect 16524 5394 16543 5428
rect 16471 5338 16543 5394
rect 16471 5304 16490 5338
rect 16524 5304 16543 5338
rect 16471 5248 16543 5304
rect 16471 5214 16490 5248
rect 16524 5214 16543 5248
rect 16471 5158 16543 5214
rect 16471 5124 16490 5158
rect 16524 5124 16543 5158
rect 16471 5068 16543 5124
rect 16471 5034 16490 5068
rect 16524 5034 16543 5068
rect 16471 4978 16543 5034
rect 16471 4944 16490 4978
rect 16524 4944 16543 4978
rect 16471 4888 16543 4944
rect 16471 4854 16490 4888
rect 16524 4854 16543 4888
rect 16471 4798 16543 4854
rect 17361 5465 17380 5499
rect 17414 5465 17433 5499
rect 17361 5409 17433 5465
rect 17361 5375 17380 5409
rect 17414 5375 17433 5409
rect 17361 5319 17433 5375
rect 17361 5285 17380 5319
rect 17414 5285 17433 5319
rect 17361 5229 17433 5285
rect 17361 5195 17380 5229
rect 17414 5195 17433 5229
rect 17361 5139 17433 5195
rect 17361 5105 17380 5139
rect 17414 5105 17433 5139
rect 17361 5049 17433 5105
rect 17361 5015 17380 5049
rect 17414 5015 17433 5049
rect 17361 4959 17433 5015
rect 17361 4925 17380 4959
rect 17414 4925 17433 4959
rect 17361 4869 17433 4925
rect 17361 4835 17380 4869
rect 17414 4835 17433 4869
rect 16471 4764 16490 4798
rect 16524 4764 16543 4798
rect 16471 4741 16543 4764
rect 17361 4779 17433 4835
rect 17361 4745 17380 4779
rect 17414 4745 17433 4779
rect 17361 4741 17433 4745
rect 16471 4722 17433 4741
rect 16471 4688 16548 4722
rect 16582 4688 16638 4722
rect 16672 4688 16728 4722
rect 16762 4688 16818 4722
rect 16852 4688 16908 4722
rect 16942 4688 16998 4722
rect 17032 4688 17088 4722
rect 17122 4688 17178 4722
rect 17212 4688 17268 4722
rect 17302 4688 17433 4722
rect 16471 4669 17433 4688
rect 17759 5612 18721 5631
rect 17759 5578 17870 5612
rect 17904 5578 17960 5612
rect 17994 5578 18050 5612
rect 18084 5578 18140 5612
rect 18174 5578 18230 5612
rect 18264 5578 18320 5612
rect 18354 5578 18410 5612
rect 18444 5578 18500 5612
rect 18534 5578 18590 5612
rect 18624 5578 18721 5612
rect 17759 5559 18721 5578
rect 17759 5518 17831 5559
rect 17759 5484 17778 5518
rect 17812 5484 17831 5518
rect 18649 5499 18721 5559
rect 17759 5428 17831 5484
rect 17759 5394 17778 5428
rect 17812 5394 17831 5428
rect 17759 5338 17831 5394
rect 17759 5304 17778 5338
rect 17812 5304 17831 5338
rect 17759 5248 17831 5304
rect 17759 5214 17778 5248
rect 17812 5214 17831 5248
rect 17759 5158 17831 5214
rect 17759 5124 17778 5158
rect 17812 5124 17831 5158
rect 17759 5068 17831 5124
rect 17759 5034 17778 5068
rect 17812 5034 17831 5068
rect 17759 4978 17831 5034
rect 17759 4944 17778 4978
rect 17812 4944 17831 4978
rect 17759 4888 17831 4944
rect 17759 4854 17778 4888
rect 17812 4854 17831 4888
rect 17759 4798 17831 4854
rect 18649 5465 18668 5499
rect 18702 5465 18721 5499
rect 18649 5409 18721 5465
rect 18649 5375 18668 5409
rect 18702 5375 18721 5409
rect 18649 5319 18721 5375
rect 18649 5285 18668 5319
rect 18702 5285 18721 5319
rect 18649 5229 18721 5285
rect 18649 5195 18668 5229
rect 18702 5195 18721 5229
rect 18649 5139 18721 5195
rect 18649 5105 18668 5139
rect 18702 5105 18721 5139
rect 18649 5049 18721 5105
rect 18649 5015 18668 5049
rect 18702 5015 18721 5049
rect 18649 4959 18721 5015
rect 18649 4925 18668 4959
rect 18702 4925 18721 4959
rect 18649 4869 18721 4925
rect 18649 4835 18668 4869
rect 18702 4835 18721 4869
rect 17759 4764 17778 4798
rect 17812 4764 17831 4798
rect 17759 4741 17831 4764
rect 18649 4779 18721 4835
rect 18649 4745 18668 4779
rect 18702 4745 18721 4779
rect 18649 4741 18721 4745
rect 17759 4722 18721 4741
rect 17759 4688 17836 4722
rect 17870 4688 17926 4722
rect 17960 4688 18016 4722
rect 18050 4688 18106 4722
rect 18140 4688 18196 4722
rect 18230 4688 18286 4722
rect 18320 4688 18376 4722
rect 18410 4688 18466 4722
rect 18500 4688 18556 4722
rect 18590 4688 18721 4722
rect 17759 4669 18721 4688
rect 12607 4324 13569 4343
rect 12607 4290 12718 4324
rect 12752 4290 12808 4324
rect 12842 4290 12898 4324
rect 12932 4290 12988 4324
rect 13022 4290 13078 4324
rect 13112 4290 13168 4324
rect 13202 4290 13258 4324
rect 13292 4290 13348 4324
rect 13382 4290 13438 4324
rect 13472 4290 13569 4324
rect 12607 4271 13569 4290
rect 12607 4230 12679 4271
rect 12607 4196 12626 4230
rect 12660 4196 12679 4230
rect 13497 4211 13569 4271
rect 12607 4140 12679 4196
rect 12607 4106 12626 4140
rect 12660 4106 12679 4140
rect 12607 4050 12679 4106
rect 12607 4016 12626 4050
rect 12660 4016 12679 4050
rect 12607 3960 12679 4016
rect 12607 3926 12626 3960
rect 12660 3926 12679 3960
rect 12607 3870 12679 3926
rect 12607 3836 12626 3870
rect 12660 3836 12679 3870
rect 12607 3780 12679 3836
rect 12607 3746 12626 3780
rect 12660 3746 12679 3780
rect 12607 3690 12679 3746
rect 12607 3656 12626 3690
rect 12660 3656 12679 3690
rect 12607 3600 12679 3656
rect 12607 3566 12626 3600
rect 12660 3566 12679 3600
rect 12607 3510 12679 3566
rect 13497 4177 13516 4211
rect 13550 4177 13569 4211
rect 13497 4121 13569 4177
rect 13497 4087 13516 4121
rect 13550 4087 13569 4121
rect 13497 4031 13569 4087
rect 13497 3997 13516 4031
rect 13550 3997 13569 4031
rect 13497 3941 13569 3997
rect 13497 3907 13516 3941
rect 13550 3907 13569 3941
rect 13497 3851 13569 3907
rect 13497 3817 13516 3851
rect 13550 3817 13569 3851
rect 13497 3761 13569 3817
rect 13497 3727 13516 3761
rect 13550 3727 13569 3761
rect 13497 3671 13569 3727
rect 13497 3637 13516 3671
rect 13550 3637 13569 3671
rect 13497 3581 13569 3637
rect 13497 3547 13516 3581
rect 13550 3547 13569 3581
rect 12607 3476 12626 3510
rect 12660 3476 12679 3510
rect 12607 3453 12679 3476
rect 13497 3491 13569 3547
rect 13497 3457 13516 3491
rect 13550 3457 13569 3491
rect 13497 3453 13569 3457
rect 12607 3434 13569 3453
rect 12607 3400 12684 3434
rect 12718 3400 12774 3434
rect 12808 3400 12864 3434
rect 12898 3400 12954 3434
rect 12988 3400 13044 3434
rect 13078 3400 13134 3434
rect 13168 3400 13224 3434
rect 13258 3400 13314 3434
rect 13348 3400 13404 3434
rect 13438 3400 13569 3434
rect 12607 3381 13569 3400
rect 13895 4324 14857 4343
rect 13895 4290 14006 4324
rect 14040 4290 14096 4324
rect 14130 4290 14186 4324
rect 14220 4290 14276 4324
rect 14310 4290 14366 4324
rect 14400 4290 14456 4324
rect 14490 4290 14546 4324
rect 14580 4290 14636 4324
rect 14670 4290 14726 4324
rect 14760 4290 14857 4324
rect 13895 4271 14857 4290
rect 13895 4230 13967 4271
rect 13895 4196 13914 4230
rect 13948 4196 13967 4230
rect 14785 4211 14857 4271
rect 13895 4140 13967 4196
rect 13895 4106 13914 4140
rect 13948 4106 13967 4140
rect 13895 4050 13967 4106
rect 13895 4016 13914 4050
rect 13948 4016 13967 4050
rect 13895 3960 13967 4016
rect 13895 3926 13914 3960
rect 13948 3926 13967 3960
rect 13895 3870 13967 3926
rect 13895 3836 13914 3870
rect 13948 3836 13967 3870
rect 13895 3780 13967 3836
rect 13895 3746 13914 3780
rect 13948 3746 13967 3780
rect 13895 3690 13967 3746
rect 13895 3656 13914 3690
rect 13948 3656 13967 3690
rect 13895 3600 13967 3656
rect 13895 3566 13914 3600
rect 13948 3566 13967 3600
rect 13895 3510 13967 3566
rect 14785 4177 14804 4211
rect 14838 4177 14857 4211
rect 14785 4121 14857 4177
rect 14785 4087 14804 4121
rect 14838 4087 14857 4121
rect 14785 4031 14857 4087
rect 14785 3997 14804 4031
rect 14838 3997 14857 4031
rect 14785 3941 14857 3997
rect 14785 3907 14804 3941
rect 14838 3907 14857 3941
rect 14785 3851 14857 3907
rect 14785 3817 14804 3851
rect 14838 3817 14857 3851
rect 14785 3761 14857 3817
rect 14785 3727 14804 3761
rect 14838 3727 14857 3761
rect 14785 3671 14857 3727
rect 14785 3637 14804 3671
rect 14838 3637 14857 3671
rect 14785 3581 14857 3637
rect 14785 3547 14804 3581
rect 14838 3547 14857 3581
rect 13895 3476 13914 3510
rect 13948 3476 13967 3510
rect 13895 3453 13967 3476
rect 14785 3491 14857 3547
rect 14785 3457 14804 3491
rect 14838 3457 14857 3491
rect 14785 3453 14857 3457
rect 13895 3434 14857 3453
rect 13895 3400 13972 3434
rect 14006 3400 14062 3434
rect 14096 3400 14152 3434
rect 14186 3400 14242 3434
rect 14276 3400 14332 3434
rect 14366 3400 14422 3434
rect 14456 3400 14512 3434
rect 14546 3400 14602 3434
rect 14636 3400 14692 3434
rect 14726 3400 14857 3434
rect 13895 3381 14857 3400
rect 15183 4324 16145 4343
rect 15183 4290 15294 4324
rect 15328 4290 15384 4324
rect 15418 4290 15474 4324
rect 15508 4290 15564 4324
rect 15598 4290 15654 4324
rect 15688 4290 15744 4324
rect 15778 4290 15834 4324
rect 15868 4290 15924 4324
rect 15958 4290 16014 4324
rect 16048 4290 16145 4324
rect 15183 4271 16145 4290
rect 15183 4230 15255 4271
rect 15183 4196 15202 4230
rect 15236 4196 15255 4230
rect 16073 4211 16145 4271
rect 15183 4140 15255 4196
rect 15183 4106 15202 4140
rect 15236 4106 15255 4140
rect 15183 4050 15255 4106
rect 15183 4016 15202 4050
rect 15236 4016 15255 4050
rect 15183 3960 15255 4016
rect 15183 3926 15202 3960
rect 15236 3926 15255 3960
rect 15183 3870 15255 3926
rect 15183 3836 15202 3870
rect 15236 3836 15255 3870
rect 15183 3780 15255 3836
rect 15183 3746 15202 3780
rect 15236 3746 15255 3780
rect 15183 3690 15255 3746
rect 15183 3656 15202 3690
rect 15236 3656 15255 3690
rect 15183 3600 15255 3656
rect 15183 3566 15202 3600
rect 15236 3566 15255 3600
rect 15183 3510 15255 3566
rect 16073 4177 16092 4211
rect 16126 4177 16145 4211
rect 16073 4121 16145 4177
rect 16073 4087 16092 4121
rect 16126 4087 16145 4121
rect 16073 4031 16145 4087
rect 16073 3997 16092 4031
rect 16126 3997 16145 4031
rect 16073 3941 16145 3997
rect 16073 3907 16092 3941
rect 16126 3907 16145 3941
rect 16073 3851 16145 3907
rect 16073 3817 16092 3851
rect 16126 3817 16145 3851
rect 16073 3761 16145 3817
rect 16073 3727 16092 3761
rect 16126 3727 16145 3761
rect 16073 3671 16145 3727
rect 16073 3637 16092 3671
rect 16126 3637 16145 3671
rect 16073 3581 16145 3637
rect 16073 3547 16092 3581
rect 16126 3547 16145 3581
rect 15183 3476 15202 3510
rect 15236 3476 15255 3510
rect 15183 3453 15255 3476
rect 16073 3491 16145 3547
rect 16073 3457 16092 3491
rect 16126 3457 16145 3491
rect 16073 3453 16145 3457
rect 15183 3434 16145 3453
rect 15183 3400 15260 3434
rect 15294 3400 15350 3434
rect 15384 3400 15440 3434
rect 15474 3400 15530 3434
rect 15564 3400 15620 3434
rect 15654 3400 15710 3434
rect 15744 3400 15800 3434
rect 15834 3400 15890 3434
rect 15924 3400 15980 3434
rect 16014 3400 16145 3434
rect 15183 3381 16145 3400
rect 16471 4324 17433 4343
rect 16471 4290 16582 4324
rect 16616 4290 16672 4324
rect 16706 4290 16762 4324
rect 16796 4290 16852 4324
rect 16886 4290 16942 4324
rect 16976 4290 17032 4324
rect 17066 4290 17122 4324
rect 17156 4290 17212 4324
rect 17246 4290 17302 4324
rect 17336 4290 17433 4324
rect 16471 4271 17433 4290
rect 16471 4230 16543 4271
rect 16471 4196 16490 4230
rect 16524 4196 16543 4230
rect 17361 4211 17433 4271
rect 16471 4140 16543 4196
rect 16471 4106 16490 4140
rect 16524 4106 16543 4140
rect 16471 4050 16543 4106
rect 16471 4016 16490 4050
rect 16524 4016 16543 4050
rect 16471 3960 16543 4016
rect 16471 3926 16490 3960
rect 16524 3926 16543 3960
rect 16471 3870 16543 3926
rect 16471 3836 16490 3870
rect 16524 3836 16543 3870
rect 16471 3780 16543 3836
rect 16471 3746 16490 3780
rect 16524 3746 16543 3780
rect 16471 3690 16543 3746
rect 16471 3656 16490 3690
rect 16524 3656 16543 3690
rect 16471 3600 16543 3656
rect 16471 3566 16490 3600
rect 16524 3566 16543 3600
rect 16471 3510 16543 3566
rect 17361 4177 17380 4211
rect 17414 4177 17433 4211
rect 17361 4121 17433 4177
rect 17361 4087 17380 4121
rect 17414 4087 17433 4121
rect 17361 4031 17433 4087
rect 17361 3997 17380 4031
rect 17414 3997 17433 4031
rect 17361 3941 17433 3997
rect 17361 3907 17380 3941
rect 17414 3907 17433 3941
rect 17361 3851 17433 3907
rect 17361 3817 17380 3851
rect 17414 3817 17433 3851
rect 17361 3761 17433 3817
rect 17361 3727 17380 3761
rect 17414 3727 17433 3761
rect 17361 3671 17433 3727
rect 17361 3637 17380 3671
rect 17414 3637 17433 3671
rect 17361 3581 17433 3637
rect 17361 3547 17380 3581
rect 17414 3547 17433 3581
rect 16471 3476 16490 3510
rect 16524 3476 16543 3510
rect 16471 3453 16543 3476
rect 17361 3491 17433 3547
rect 17361 3457 17380 3491
rect 17414 3457 17433 3491
rect 17361 3453 17433 3457
rect 16471 3434 17433 3453
rect 16471 3400 16548 3434
rect 16582 3400 16638 3434
rect 16672 3400 16728 3434
rect 16762 3400 16818 3434
rect 16852 3400 16908 3434
rect 16942 3400 16998 3434
rect 17032 3400 17088 3434
rect 17122 3400 17178 3434
rect 17212 3400 17268 3434
rect 17302 3400 17433 3434
rect 16471 3381 17433 3400
rect 17759 4324 18721 4343
rect 17759 4290 17870 4324
rect 17904 4290 17960 4324
rect 17994 4290 18050 4324
rect 18084 4290 18140 4324
rect 18174 4290 18230 4324
rect 18264 4290 18320 4324
rect 18354 4290 18410 4324
rect 18444 4290 18500 4324
rect 18534 4290 18590 4324
rect 18624 4290 18721 4324
rect 17759 4271 18721 4290
rect 17759 4230 17831 4271
rect 17759 4196 17778 4230
rect 17812 4196 17831 4230
rect 18649 4211 18721 4271
rect 17759 4140 17831 4196
rect 17759 4106 17778 4140
rect 17812 4106 17831 4140
rect 17759 4050 17831 4106
rect 17759 4016 17778 4050
rect 17812 4016 17831 4050
rect 17759 3960 17831 4016
rect 17759 3926 17778 3960
rect 17812 3926 17831 3960
rect 17759 3870 17831 3926
rect 17759 3836 17778 3870
rect 17812 3836 17831 3870
rect 17759 3780 17831 3836
rect 17759 3746 17778 3780
rect 17812 3746 17831 3780
rect 17759 3690 17831 3746
rect 17759 3656 17778 3690
rect 17812 3656 17831 3690
rect 17759 3600 17831 3656
rect 17759 3566 17778 3600
rect 17812 3566 17831 3600
rect 17759 3510 17831 3566
rect 18649 4177 18668 4211
rect 18702 4177 18721 4211
rect 18649 4121 18721 4177
rect 18649 4087 18668 4121
rect 18702 4087 18721 4121
rect 18649 4031 18721 4087
rect 18649 3997 18668 4031
rect 18702 3997 18721 4031
rect 18649 3941 18721 3997
rect 18649 3907 18668 3941
rect 18702 3907 18721 3941
rect 18649 3851 18721 3907
rect 18649 3817 18668 3851
rect 18702 3817 18721 3851
rect 18649 3761 18721 3817
rect 18649 3727 18668 3761
rect 18702 3727 18721 3761
rect 18649 3671 18721 3727
rect 18649 3637 18668 3671
rect 18702 3637 18721 3671
rect 18649 3581 18721 3637
rect 18649 3547 18668 3581
rect 18702 3547 18721 3581
rect 17759 3476 17778 3510
rect 17812 3476 17831 3510
rect 17759 3453 17831 3476
rect 18649 3491 18721 3547
rect 18649 3457 18668 3491
rect 18702 3457 18721 3491
rect 18649 3453 18721 3457
rect 17759 3434 18721 3453
rect 17759 3400 17836 3434
rect 17870 3400 17926 3434
rect 17960 3400 18016 3434
rect 18050 3400 18106 3434
rect 18140 3400 18196 3434
rect 18230 3400 18286 3434
rect 18320 3400 18376 3434
rect 18410 3400 18466 3434
rect 18500 3400 18556 3434
rect 18590 3400 18721 3434
rect 17759 3381 18721 3400
rect 12607 3036 13569 3055
rect 12607 3002 12718 3036
rect 12752 3002 12808 3036
rect 12842 3002 12898 3036
rect 12932 3002 12988 3036
rect 13022 3002 13078 3036
rect 13112 3002 13168 3036
rect 13202 3002 13258 3036
rect 13292 3002 13348 3036
rect 13382 3002 13438 3036
rect 13472 3002 13569 3036
rect 12607 2983 13569 3002
rect 12607 2942 12679 2983
rect 12607 2908 12626 2942
rect 12660 2908 12679 2942
rect 13497 2923 13569 2983
rect 12607 2852 12679 2908
rect 12607 2818 12626 2852
rect 12660 2818 12679 2852
rect 12607 2762 12679 2818
rect 12607 2728 12626 2762
rect 12660 2728 12679 2762
rect 12607 2672 12679 2728
rect 12607 2638 12626 2672
rect 12660 2638 12679 2672
rect 12607 2582 12679 2638
rect 12607 2548 12626 2582
rect 12660 2548 12679 2582
rect 12607 2492 12679 2548
rect 12607 2458 12626 2492
rect 12660 2458 12679 2492
rect 12607 2402 12679 2458
rect 12607 2368 12626 2402
rect 12660 2368 12679 2402
rect 12607 2312 12679 2368
rect 12607 2278 12626 2312
rect 12660 2278 12679 2312
rect 12607 2222 12679 2278
rect 13497 2889 13516 2923
rect 13550 2889 13569 2923
rect 13497 2833 13569 2889
rect 13497 2799 13516 2833
rect 13550 2799 13569 2833
rect 13497 2743 13569 2799
rect 13497 2709 13516 2743
rect 13550 2709 13569 2743
rect 13497 2653 13569 2709
rect 13497 2619 13516 2653
rect 13550 2619 13569 2653
rect 13497 2563 13569 2619
rect 13497 2529 13516 2563
rect 13550 2529 13569 2563
rect 13497 2473 13569 2529
rect 13497 2439 13516 2473
rect 13550 2439 13569 2473
rect 13497 2383 13569 2439
rect 13497 2349 13516 2383
rect 13550 2349 13569 2383
rect 13497 2293 13569 2349
rect 13497 2259 13516 2293
rect 13550 2259 13569 2293
rect 12607 2188 12626 2222
rect 12660 2188 12679 2222
rect 12607 2165 12679 2188
rect 13497 2203 13569 2259
rect 13497 2169 13516 2203
rect 13550 2169 13569 2203
rect 13497 2165 13569 2169
rect 12607 2146 13569 2165
rect 12607 2112 12684 2146
rect 12718 2112 12774 2146
rect 12808 2112 12864 2146
rect 12898 2112 12954 2146
rect 12988 2112 13044 2146
rect 13078 2112 13134 2146
rect 13168 2112 13224 2146
rect 13258 2112 13314 2146
rect 13348 2112 13404 2146
rect 13438 2112 13569 2146
rect 12607 2093 13569 2112
rect 13895 3036 14857 3055
rect 13895 3002 14006 3036
rect 14040 3002 14096 3036
rect 14130 3002 14186 3036
rect 14220 3002 14276 3036
rect 14310 3002 14366 3036
rect 14400 3002 14456 3036
rect 14490 3002 14546 3036
rect 14580 3002 14636 3036
rect 14670 3002 14726 3036
rect 14760 3002 14857 3036
rect 13895 2983 14857 3002
rect 13895 2942 13967 2983
rect 13895 2908 13914 2942
rect 13948 2908 13967 2942
rect 14785 2923 14857 2983
rect 13895 2852 13967 2908
rect 13895 2818 13914 2852
rect 13948 2818 13967 2852
rect 13895 2762 13967 2818
rect 13895 2728 13914 2762
rect 13948 2728 13967 2762
rect 13895 2672 13967 2728
rect 13895 2638 13914 2672
rect 13948 2638 13967 2672
rect 13895 2582 13967 2638
rect 13895 2548 13914 2582
rect 13948 2548 13967 2582
rect 13895 2492 13967 2548
rect 13895 2458 13914 2492
rect 13948 2458 13967 2492
rect 13895 2402 13967 2458
rect 13895 2368 13914 2402
rect 13948 2368 13967 2402
rect 13895 2312 13967 2368
rect 13895 2278 13914 2312
rect 13948 2278 13967 2312
rect 13895 2222 13967 2278
rect 14785 2889 14804 2923
rect 14838 2889 14857 2923
rect 14785 2833 14857 2889
rect 14785 2799 14804 2833
rect 14838 2799 14857 2833
rect 14785 2743 14857 2799
rect 14785 2709 14804 2743
rect 14838 2709 14857 2743
rect 14785 2653 14857 2709
rect 14785 2619 14804 2653
rect 14838 2619 14857 2653
rect 14785 2563 14857 2619
rect 14785 2529 14804 2563
rect 14838 2529 14857 2563
rect 14785 2473 14857 2529
rect 14785 2439 14804 2473
rect 14838 2439 14857 2473
rect 14785 2383 14857 2439
rect 14785 2349 14804 2383
rect 14838 2349 14857 2383
rect 14785 2293 14857 2349
rect 14785 2259 14804 2293
rect 14838 2259 14857 2293
rect 13895 2188 13914 2222
rect 13948 2188 13967 2222
rect 13895 2165 13967 2188
rect 14785 2203 14857 2259
rect 14785 2169 14804 2203
rect 14838 2169 14857 2203
rect 14785 2165 14857 2169
rect 13895 2146 14857 2165
rect 13895 2112 13972 2146
rect 14006 2112 14062 2146
rect 14096 2112 14152 2146
rect 14186 2112 14242 2146
rect 14276 2112 14332 2146
rect 14366 2112 14422 2146
rect 14456 2112 14512 2146
rect 14546 2112 14602 2146
rect 14636 2112 14692 2146
rect 14726 2112 14857 2146
rect 13895 2093 14857 2112
rect 15183 3036 16145 3055
rect 15183 3002 15294 3036
rect 15328 3002 15384 3036
rect 15418 3002 15474 3036
rect 15508 3002 15564 3036
rect 15598 3002 15654 3036
rect 15688 3002 15744 3036
rect 15778 3002 15834 3036
rect 15868 3002 15924 3036
rect 15958 3002 16014 3036
rect 16048 3002 16145 3036
rect 15183 2983 16145 3002
rect 15183 2942 15255 2983
rect 15183 2908 15202 2942
rect 15236 2908 15255 2942
rect 16073 2923 16145 2983
rect 15183 2852 15255 2908
rect 15183 2818 15202 2852
rect 15236 2818 15255 2852
rect 15183 2762 15255 2818
rect 15183 2728 15202 2762
rect 15236 2728 15255 2762
rect 15183 2672 15255 2728
rect 15183 2638 15202 2672
rect 15236 2638 15255 2672
rect 15183 2582 15255 2638
rect 15183 2548 15202 2582
rect 15236 2548 15255 2582
rect 15183 2492 15255 2548
rect 15183 2458 15202 2492
rect 15236 2458 15255 2492
rect 15183 2402 15255 2458
rect 15183 2368 15202 2402
rect 15236 2368 15255 2402
rect 15183 2312 15255 2368
rect 15183 2278 15202 2312
rect 15236 2278 15255 2312
rect 15183 2222 15255 2278
rect 16073 2889 16092 2923
rect 16126 2889 16145 2923
rect 16073 2833 16145 2889
rect 16073 2799 16092 2833
rect 16126 2799 16145 2833
rect 16073 2743 16145 2799
rect 16073 2709 16092 2743
rect 16126 2709 16145 2743
rect 16073 2653 16145 2709
rect 16073 2619 16092 2653
rect 16126 2619 16145 2653
rect 16073 2563 16145 2619
rect 16073 2529 16092 2563
rect 16126 2529 16145 2563
rect 16073 2473 16145 2529
rect 16073 2439 16092 2473
rect 16126 2439 16145 2473
rect 16073 2383 16145 2439
rect 16073 2349 16092 2383
rect 16126 2349 16145 2383
rect 16073 2293 16145 2349
rect 16073 2259 16092 2293
rect 16126 2259 16145 2293
rect 15183 2188 15202 2222
rect 15236 2188 15255 2222
rect 15183 2165 15255 2188
rect 16073 2203 16145 2259
rect 16073 2169 16092 2203
rect 16126 2169 16145 2203
rect 16073 2165 16145 2169
rect 15183 2146 16145 2165
rect 15183 2112 15260 2146
rect 15294 2112 15350 2146
rect 15384 2112 15440 2146
rect 15474 2112 15530 2146
rect 15564 2112 15620 2146
rect 15654 2112 15710 2146
rect 15744 2112 15800 2146
rect 15834 2112 15890 2146
rect 15924 2112 15980 2146
rect 16014 2112 16145 2146
rect 15183 2093 16145 2112
rect 16471 3036 17433 3055
rect 16471 3002 16582 3036
rect 16616 3002 16672 3036
rect 16706 3002 16762 3036
rect 16796 3002 16852 3036
rect 16886 3002 16942 3036
rect 16976 3002 17032 3036
rect 17066 3002 17122 3036
rect 17156 3002 17212 3036
rect 17246 3002 17302 3036
rect 17336 3002 17433 3036
rect 16471 2983 17433 3002
rect 16471 2942 16543 2983
rect 16471 2908 16490 2942
rect 16524 2908 16543 2942
rect 17361 2923 17433 2983
rect 16471 2852 16543 2908
rect 16471 2818 16490 2852
rect 16524 2818 16543 2852
rect 16471 2762 16543 2818
rect 16471 2728 16490 2762
rect 16524 2728 16543 2762
rect 16471 2672 16543 2728
rect 16471 2638 16490 2672
rect 16524 2638 16543 2672
rect 16471 2582 16543 2638
rect 16471 2548 16490 2582
rect 16524 2548 16543 2582
rect 16471 2492 16543 2548
rect 16471 2458 16490 2492
rect 16524 2458 16543 2492
rect 16471 2402 16543 2458
rect 16471 2368 16490 2402
rect 16524 2368 16543 2402
rect 16471 2312 16543 2368
rect 16471 2278 16490 2312
rect 16524 2278 16543 2312
rect 16471 2222 16543 2278
rect 17361 2889 17380 2923
rect 17414 2889 17433 2923
rect 17361 2833 17433 2889
rect 17361 2799 17380 2833
rect 17414 2799 17433 2833
rect 17361 2743 17433 2799
rect 17361 2709 17380 2743
rect 17414 2709 17433 2743
rect 17361 2653 17433 2709
rect 17361 2619 17380 2653
rect 17414 2619 17433 2653
rect 17361 2563 17433 2619
rect 17361 2529 17380 2563
rect 17414 2529 17433 2563
rect 17361 2473 17433 2529
rect 17361 2439 17380 2473
rect 17414 2439 17433 2473
rect 17361 2383 17433 2439
rect 17361 2349 17380 2383
rect 17414 2349 17433 2383
rect 17361 2293 17433 2349
rect 17361 2259 17380 2293
rect 17414 2259 17433 2293
rect 16471 2188 16490 2222
rect 16524 2188 16543 2222
rect 16471 2165 16543 2188
rect 17361 2203 17433 2259
rect 17361 2169 17380 2203
rect 17414 2169 17433 2203
rect 17361 2165 17433 2169
rect 16471 2146 17433 2165
rect 16471 2112 16548 2146
rect 16582 2112 16638 2146
rect 16672 2112 16728 2146
rect 16762 2112 16818 2146
rect 16852 2112 16908 2146
rect 16942 2112 16998 2146
rect 17032 2112 17088 2146
rect 17122 2112 17178 2146
rect 17212 2112 17268 2146
rect 17302 2112 17433 2146
rect 16471 2093 17433 2112
rect 17759 3036 18721 3055
rect 17759 3002 17870 3036
rect 17904 3002 17960 3036
rect 17994 3002 18050 3036
rect 18084 3002 18140 3036
rect 18174 3002 18230 3036
rect 18264 3002 18320 3036
rect 18354 3002 18410 3036
rect 18444 3002 18500 3036
rect 18534 3002 18590 3036
rect 18624 3002 18721 3036
rect 17759 2983 18721 3002
rect 17759 2942 17831 2983
rect 17759 2908 17778 2942
rect 17812 2908 17831 2942
rect 18649 2923 18721 2983
rect 17759 2852 17831 2908
rect 17759 2818 17778 2852
rect 17812 2818 17831 2852
rect 17759 2762 17831 2818
rect 17759 2728 17778 2762
rect 17812 2728 17831 2762
rect 17759 2672 17831 2728
rect 17759 2638 17778 2672
rect 17812 2638 17831 2672
rect 17759 2582 17831 2638
rect 17759 2548 17778 2582
rect 17812 2548 17831 2582
rect 17759 2492 17831 2548
rect 17759 2458 17778 2492
rect 17812 2458 17831 2492
rect 17759 2402 17831 2458
rect 17759 2368 17778 2402
rect 17812 2368 17831 2402
rect 17759 2312 17831 2368
rect 17759 2278 17778 2312
rect 17812 2278 17831 2312
rect 17759 2222 17831 2278
rect 18649 2889 18668 2923
rect 18702 2889 18721 2923
rect 18649 2833 18721 2889
rect 18649 2799 18668 2833
rect 18702 2799 18721 2833
rect 18649 2743 18721 2799
rect 18649 2709 18668 2743
rect 18702 2709 18721 2743
rect 18649 2653 18721 2709
rect 18649 2619 18668 2653
rect 18702 2619 18721 2653
rect 18649 2563 18721 2619
rect 18649 2529 18668 2563
rect 18702 2529 18721 2563
rect 18649 2473 18721 2529
rect 18649 2439 18668 2473
rect 18702 2439 18721 2473
rect 18649 2383 18721 2439
rect 18649 2349 18668 2383
rect 18702 2349 18721 2383
rect 18649 2293 18721 2349
rect 18649 2259 18668 2293
rect 18702 2259 18721 2293
rect 17759 2188 17778 2222
rect 17812 2188 17831 2222
rect 17759 2165 17831 2188
rect 18649 2203 18721 2259
rect 18649 2169 18668 2203
rect 18702 2169 18721 2203
rect 18649 2165 18721 2169
rect 17759 2146 18721 2165
rect 17759 2112 17836 2146
rect 17870 2112 17926 2146
rect 17960 2112 18016 2146
rect 18050 2112 18106 2146
rect 18140 2112 18196 2146
rect 18230 2112 18286 2146
rect 18320 2112 18376 2146
rect 18410 2112 18466 2146
rect 18500 2112 18556 2146
rect 18590 2112 18721 2146
rect 17759 2093 18721 2112
rect -15768 1296 -13226 1346
rect -15768 1196 -15668 1296
rect -13326 1196 -13226 1296
rect -15768 1146 -13226 1196
<< psubdiffcont >>
rect -21516 24270 -10332 25036
rect -9756 15196 -9186 21500
rect -6512 15196 -5942 21500
rect -1552 15196 -982 21500
rect 13136 15196 13706 21500
rect 12578 12168 12612 12202
rect 12668 12168 12702 12202
rect 12758 12168 12792 12202
rect 12848 12168 12882 12202
rect 12938 12168 12972 12202
rect 13028 12168 13062 12202
rect 13118 12168 13152 12202
rect 13208 12168 13242 12202
rect 13298 12168 13332 12202
rect 13388 12168 13422 12202
rect 13478 12168 13512 12202
rect 13568 12168 13602 12202
rect 13866 12168 13900 12202
rect 13956 12168 13990 12202
rect 14046 12168 14080 12202
rect 14136 12168 14170 12202
rect 14226 12168 14260 12202
rect 14316 12168 14350 12202
rect 14406 12168 14440 12202
rect 14496 12168 14530 12202
rect 14586 12168 14620 12202
rect 14676 12168 14710 12202
rect 14766 12168 14800 12202
rect 14856 12168 14890 12202
rect 15154 12168 15188 12202
rect 15244 12168 15278 12202
rect 15334 12168 15368 12202
rect 15424 12168 15458 12202
rect 15514 12168 15548 12202
rect 15604 12168 15638 12202
rect 15694 12168 15728 12202
rect 15784 12168 15818 12202
rect 15874 12168 15908 12202
rect 15964 12168 15998 12202
rect 16054 12168 16088 12202
rect 16144 12168 16178 12202
rect 16442 12168 16476 12202
rect 16532 12168 16566 12202
rect 16622 12168 16656 12202
rect 16712 12168 16746 12202
rect 16802 12168 16836 12202
rect 16892 12168 16926 12202
rect 16982 12168 17016 12202
rect 17072 12168 17106 12202
rect 17162 12168 17196 12202
rect 17252 12168 17286 12202
rect 17342 12168 17376 12202
rect 17432 12168 17466 12202
rect 17730 12168 17764 12202
rect 17820 12168 17854 12202
rect 17910 12168 17944 12202
rect 18000 12168 18034 12202
rect 18090 12168 18124 12202
rect 18180 12168 18214 12202
rect 18270 12168 18304 12202
rect 18360 12168 18394 12202
rect 18450 12168 18484 12202
rect 18540 12168 18574 12202
rect 18630 12168 18664 12202
rect 18720 12168 18754 12202
rect 12477 12084 12511 12118
rect 13664 12084 13698 12118
rect 13765 12084 13799 12118
rect 12477 11994 12511 12028
rect 12477 11904 12511 11938
rect 12477 11814 12511 11848
rect 12477 11724 12511 11758
rect 12477 11634 12511 11668
rect 12477 11544 12511 11578
rect 12477 11454 12511 11488
rect 12477 11364 12511 11398
rect 12477 11274 12511 11308
rect 12477 11184 12511 11218
rect 12477 11094 12511 11128
rect 14952 12084 14986 12118
rect 15053 12084 15087 12118
rect 13664 11994 13698 12028
rect 13765 11994 13799 12028
rect 13664 11904 13698 11938
rect 13765 11904 13799 11938
rect 13664 11814 13698 11848
rect 13765 11814 13799 11848
rect 13664 11724 13698 11758
rect 13765 11724 13799 11758
rect 13664 11634 13698 11668
rect 13765 11634 13799 11668
rect 13664 11544 13698 11578
rect 13765 11544 13799 11578
rect 13664 11454 13698 11488
rect 13765 11454 13799 11488
rect 13664 11364 13698 11398
rect 13765 11364 13799 11398
rect 13664 11274 13698 11308
rect 13765 11274 13799 11308
rect 13664 11184 13698 11218
rect 13765 11184 13799 11218
rect 13664 11094 13698 11128
rect 13765 11094 13799 11128
rect 16240 12084 16274 12118
rect 16341 12084 16375 12118
rect 14952 11994 14986 12028
rect 15053 11994 15087 12028
rect 14952 11904 14986 11938
rect 15053 11904 15087 11938
rect 14952 11814 14986 11848
rect 15053 11814 15087 11848
rect 14952 11724 14986 11758
rect 15053 11724 15087 11758
rect 14952 11634 14986 11668
rect 15053 11634 15087 11668
rect 14952 11544 14986 11578
rect 15053 11544 15087 11578
rect 14952 11454 14986 11488
rect 15053 11454 15087 11488
rect 14952 11364 14986 11398
rect 15053 11364 15087 11398
rect 14952 11274 14986 11308
rect 15053 11274 15087 11308
rect 14952 11184 14986 11218
rect 15053 11184 15087 11218
rect 14952 11094 14986 11128
rect 15053 11094 15087 11128
rect 17528 12084 17562 12118
rect 17629 12084 17663 12118
rect 16240 11994 16274 12028
rect 16341 11994 16375 12028
rect 16240 11904 16274 11938
rect 16341 11904 16375 11938
rect 16240 11814 16274 11848
rect 16341 11814 16375 11848
rect 16240 11724 16274 11758
rect 16341 11724 16375 11758
rect 16240 11634 16274 11668
rect 16341 11634 16375 11668
rect 16240 11544 16274 11578
rect 16341 11544 16375 11578
rect 16240 11454 16274 11488
rect 16341 11454 16375 11488
rect 16240 11364 16274 11398
rect 16341 11364 16375 11398
rect 16240 11274 16274 11308
rect 16341 11274 16375 11308
rect 16240 11184 16274 11218
rect 16341 11184 16375 11218
rect 16240 11094 16274 11128
rect 16341 11094 16375 11128
rect 18816 12084 18850 12118
rect 17528 11994 17562 12028
rect 17629 11994 17663 12028
rect 17528 11904 17562 11938
rect 17629 11904 17663 11938
rect 17528 11814 17562 11848
rect 17629 11814 17663 11848
rect 17528 11724 17562 11758
rect 17629 11724 17663 11758
rect 17528 11634 17562 11668
rect 17629 11634 17663 11668
rect 17528 11544 17562 11578
rect 17629 11544 17663 11578
rect 17528 11454 17562 11488
rect 17629 11454 17663 11488
rect 17528 11364 17562 11398
rect 17629 11364 17663 11398
rect 17528 11274 17562 11308
rect 17629 11274 17663 11308
rect 17528 11184 17562 11218
rect 17629 11184 17663 11218
rect 17528 11094 17562 11128
rect 17629 11094 17663 11128
rect 18816 11994 18850 12028
rect 18816 11904 18850 11938
rect 18816 11814 18850 11848
rect 18816 11724 18850 11758
rect 18816 11634 18850 11668
rect 18816 11544 18850 11578
rect 18816 11454 18850 11488
rect 18816 11364 18850 11398
rect 18816 11274 18850 11308
rect 18816 11184 18850 11218
rect 18816 11094 18850 11128
rect 12477 11004 12511 11038
rect 12578 10981 12612 11015
rect 12668 10981 12702 11015
rect 12758 10981 12792 11015
rect 12848 10981 12882 11015
rect 12938 10981 12972 11015
rect 13028 10981 13062 11015
rect 13118 10981 13152 11015
rect 13208 10981 13242 11015
rect 13298 10981 13332 11015
rect 13388 10981 13422 11015
rect 13478 10981 13512 11015
rect 13568 10981 13602 11015
rect 13664 11004 13698 11038
rect 13765 11004 13799 11038
rect 13866 10981 13900 11015
rect 13956 10981 13990 11015
rect 14046 10981 14080 11015
rect 14136 10981 14170 11015
rect 14226 10981 14260 11015
rect 14316 10981 14350 11015
rect 14406 10981 14440 11015
rect 14496 10981 14530 11015
rect 14586 10981 14620 11015
rect 14676 10981 14710 11015
rect 14766 10981 14800 11015
rect 14856 10981 14890 11015
rect 14952 11004 14986 11038
rect 15053 11004 15087 11038
rect 15154 10981 15188 11015
rect 15244 10981 15278 11015
rect 15334 10981 15368 11015
rect 15424 10981 15458 11015
rect 15514 10981 15548 11015
rect 15604 10981 15638 11015
rect 15694 10981 15728 11015
rect 15784 10981 15818 11015
rect 15874 10981 15908 11015
rect 15964 10981 15998 11015
rect 16054 10981 16088 11015
rect 16144 10981 16178 11015
rect 16240 11004 16274 11038
rect 16341 11004 16375 11038
rect 16442 10981 16476 11015
rect 16532 10981 16566 11015
rect 16622 10981 16656 11015
rect 16712 10981 16746 11015
rect 16802 10981 16836 11015
rect 16892 10981 16926 11015
rect 16982 10981 17016 11015
rect 17072 10981 17106 11015
rect 17162 10981 17196 11015
rect 17252 10981 17286 11015
rect 17342 10981 17376 11015
rect 17432 10981 17466 11015
rect 17528 11004 17562 11038
rect 17629 11004 17663 11038
rect 17730 10981 17764 11015
rect 17820 10981 17854 11015
rect 17910 10981 17944 11015
rect 18000 10981 18034 11015
rect 18090 10981 18124 11015
rect 18180 10981 18214 11015
rect 18270 10981 18304 11015
rect 18360 10981 18394 11015
rect 18450 10981 18484 11015
rect 18540 10981 18574 11015
rect 18630 10981 18664 11015
rect 18720 10981 18754 11015
rect 18816 11004 18850 11038
rect 12578 10880 12612 10914
rect 12668 10880 12702 10914
rect 12758 10880 12792 10914
rect 12848 10880 12882 10914
rect 12938 10880 12972 10914
rect 13028 10880 13062 10914
rect 13118 10880 13152 10914
rect 13208 10880 13242 10914
rect 13298 10880 13332 10914
rect 13388 10880 13422 10914
rect 13478 10880 13512 10914
rect 13568 10880 13602 10914
rect 13866 10880 13900 10914
rect 13956 10880 13990 10914
rect 14046 10880 14080 10914
rect 14136 10880 14170 10914
rect 14226 10880 14260 10914
rect 14316 10880 14350 10914
rect 14406 10880 14440 10914
rect 14496 10880 14530 10914
rect 14586 10880 14620 10914
rect 14676 10880 14710 10914
rect 14766 10880 14800 10914
rect 14856 10880 14890 10914
rect 15154 10880 15188 10914
rect 15244 10880 15278 10914
rect 15334 10880 15368 10914
rect 15424 10880 15458 10914
rect 15514 10880 15548 10914
rect 15604 10880 15638 10914
rect 15694 10880 15728 10914
rect 15784 10880 15818 10914
rect 15874 10880 15908 10914
rect 15964 10880 15998 10914
rect 16054 10880 16088 10914
rect 16144 10880 16178 10914
rect 16442 10880 16476 10914
rect 16532 10880 16566 10914
rect 16622 10880 16656 10914
rect 16712 10880 16746 10914
rect 16802 10880 16836 10914
rect 16892 10880 16926 10914
rect 16982 10880 17016 10914
rect 17072 10880 17106 10914
rect 17162 10880 17196 10914
rect 17252 10880 17286 10914
rect 17342 10880 17376 10914
rect 17432 10880 17466 10914
rect 17730 10880 17764 10914
rect 17820 10880 17854 10914
rect 17910 10880 17944 10914
rect 18000 10880 18034 10914
rect 18090 10880 18124 10914
rect 18180 10880 18214 10914
rect 18270 10880 18304 10914
rect 18360 10880 18394 10914
rect 18450 10880 18484 10914
rect 18540 10880 18574 10914
rect 18630 10880 18664 10914
rect 18720 10880 18754 10914
rect 12477 10796 12511 10830
rect 13664 10796 13698 10830
rect 13765 10796 13799 10830
rect 12477 10706 12511 10740
rect 12477 10616 12511 10650
rect 12477 10526 12511 10560
rect 12477 10436 12511 10470
rect 12477 10346 12511 10380
rect 12477 10256 12511 10290
rect 12477 10166 12511 10200
rect 12477 10076 12511 10110
rect 12477 9986 12511 10020
rect 12477 9896 12511 9930
rect 12477 9806 12511 9840
rect 14952 10796 14986 10830
rect 15053 10796 15087 10830
rect 13664 10706 13698 10740
rect 13765 10706 13799 10740
rect 13664 10616 13698 10650
rect 13765 10616 13799 10650
rect 13664 10526 13698 10560
rect 13765 10526 13799 10560
rect 13664 10436 13698 10470
rect 13765 10436 13799 10470
rect 13664 10346 13698 10380
rect 13765 10346 13799 10380
rect 13664 10256 13698 10290
rect 13765 10256 13799 10290
rect 13664 10166 13698 10200
rect 13765 10166 13799 10200
rect 13664 10076 13698 10110
rect 13765 10076 13799 10110
rect 13664 9986 13698 10020
rect 13765 9986 13799 10020
rect 13664 9896 13698 9930
rect 13765 9896 13799 9930
rect 13664 9806 13698 9840
rect 13765 9806 13799 9840
rect 16240 10796 16274 10830
rect 16341 10796 16375 10830
rect 14952 10706 14986 10740
rect 15053 10706 15087 10740
rect 14952 10616 14986 10650
rect 15053 10616 15087 10650
rect 14952 10526 14986 10560
rect 15053 10526 15087 10560
rect 14952 10436 14986 10470
rect 15053 10436 15087 10470
rect 14952 10346 14986 10380
rect 15053 10346 15087 10380
rect 14952 10256 14986 10290
rect 15053 10256 15087 10290
rect 14952 10166 14986 10200
rect 15053 10166 15087 10200
rect 14952 10076 14986 10110
rect 15053 10076 15087 10110
rect 14952 9986 14986 10020
rect 15053 9986 15087 10020
rect 14952 9896 14986 9930
rect 15053 9896 15087 9930
rect 14952 9806 14986 9840
rect 15053 9806 15087 9840
rect 17528 10796 17562 10830
rect 17629 10796 17663 10830
rect 16240 10706 16274 10740
rect 16341 10706 16375 10740
rect 16240 10616 16274 10650
rect 16341 10616 16375 10650
rect 16240 10526 16274 10560
rect 16341 10526 16375 10560
rect 16240 10436 16274 10470
rect 16341 10436 16375 10470
rect 16240 10346 16274 10380
rect 16341 10346 16375 10380
rect 16240 10256 16274 10290
rect 16341 10256 16375 10290
rect 16240 10166 16274 10200
rect 16341 10166 16375 10200
rect 16240 10076 16274 10110
rect 16341 10076 16375 10110
rect 16240 9986 16274 10020
rect 16341 9986 16375 10020
rect 16240 9896 16274 9930
rect 16341 9896 16375 9930
rect 16240 9806 16274 9840
rect 16341 9806 16375 9840
rect 18816 10796 18850 10830
rect 17528 10706 17562 10740
rect 17629 10706 17663 10740
rect 17528 10616 17562 10650
rect 17629 10616 17663 10650
rect 17528 10526 17562 10560
rect 17629 10526 17663 10560
rect 17528 10436 17562 10470
rect 17629 10436 17663 10470
rect 17528 10346 17562 10380
rect 17629 10346 17663 10380
rect 17528 10256 17562 10290
rect 17629 10256 17663 10290
rect 17528 10166 17562 10200
rect 17629 10166 17663 10200
rect 17528 10076 17562 10110
rect 17629 10076 17663 10110
rect 17528 9986 17562 10020
rect 17629 9986 17663 10020
rect 17528 9896 17562 9930
rect 17629 9896 17663 9930
rect 17528 9806 17562 9840
rect 17629 9806 17663 9840
rect 18816 10706 18850 10740
rect 18816 10616 18850 10650
rect 18816 10526 18850 10560
rect 18816 10436 18850 10470
rect 18816 10346 18850 10380
rect 18816 10256 18850 10290
rect 18816 10166 18850 10200
rect 18816 10076 18850 10110
rect 18816 9986 18850 10020
rect 18816 9896 18850 9930
rect 18816 9806 18850 9840
rect 12477 9716 12511 9750
rect 12578 9693 12612 9727
rect 12668 9693 12702 9727
rect 12758 9693 12792 9727
rect 12848 9693 12882 9727
rect 12938 9693 12972 9727
rect 13028 9693 13062 9727
rect 13118 9693 13152 9727
rect 13208 9693 13242 9727
rect 13298 9693 13332 9727
rect 13388 9693 13422 9727
rect 13478 9693 13512 9727
rect 13568 9693 13602 9727
rect 13664 9716 13698 9750
rect 13765 9716 13799 9750
rect 13866 9693 13900 9727
rect 13956 9693 13990 9727
rect 14046 9693 14080 9727
rect 14136 9693 14170 9727
rect 14226 9693 14260 9727
rect 14316 9693 14350 9727
rect 14406 9693 14440 9727
rect 14496 9693 14530 9727
rect 14586 9693 14620 9727
rect 14676 9693 14710 9727
rect 14766 9693 14800 9727
rect 14856 9693 14890 9727
rect 14952 9716 14986 9750
rect 15053 9716 15087 9750
rect 15154 9693 15188 9727
rect 15244 9693 15278 9727
rect 15334 9693 15368 9727
rect 15424 9693 15458 9727
rect 15514 9693 15548 9727
rect 15604 9693 15638 9727
rect 15694 9693 15728 9727
rect 15784 9693 15818 9727
rect 15874 9693 15908 9727
rect 15964 9693 15998 9727
rect 16054 9693 16088 9727
rect 16144 9693 16178 9727
rect 16240 9716 16274 9750
rect 16341 9716 16375 9750
rect 16442 9693 16476 9727
rect 16532 9693 16566 9727
rect 16622 9693 16656 9727
rect 16712 9693 16746 9727
rect 16802 9693 16836 9727
rect 16892 9693 16926 9727
rect 16982 9693 17016 9727
rect 17072 9693 17106 9727
rect 17162 9693 17196 9727
rect 17252 9693 17286 9727
rect 17342 9693 17376 9727
rect 17432 9693 17466 9727
rect 17528 9716 17562 9750
rect 17629 9716 17663 9750
rect 17730 9693 17764 9727
rect 17820 9693 17854 9727
rect 17910 9693 17944 9727
rect 18000 9693 18034 9727
rect 18090 9693 18124 9727
rect 18180 9693 18214 9727
rect 18270 9693 18304 9727
rect 18360 9693 18394 9727
rect 18450 9693 18484 9727
rect 18540 9693 18574 9727
rect 18630 9693 18664 9727
rect 18720 9693 18754 9727
rect 18816 9716 18850 9750
rect 12578 9592 12612 9626
rect 12668 9592 12702 9626
rect 12758 9592 12792 9626
rect 12848 9592 12882 9626
rect 12938 9592 12972 9626
rect 13028 9592 13062 9626
rect 13118 9592 13152 9626
rect 13208 9592 13242 9626
rect 13298 9592 13332 9626
rect 13388 9592 13422 9626
rect 13478 9592 13512 9626
rect 13568 9592 13602 9626
rect 13866 9592 13900 9626
rect 13956 9592 13990 9626
rect 14046 9592 14080 9626
rect 14136 9592 14170 9626
rect 14226 9592 14260 9626
rect 14316 9592 14350 9626
rect 14406 9592 14440 9626
rect 14496 9592 14530 9626
rect 14586 9592 14620 9626
rect 14676 9592 14710 9626
rect 14766 9592 14800 9626
rect 14856 9592 14890 9626
rect 15154 9592 15188 9626
rect 15244 9592 15278 9626
rect 15334 9592 15368 9626
rect 15424 9592 15458 9626
rect 15514 9592 15548 9626
rect 15604 9592 15638 9626
rect 15694 9592 15728 9626
rect 15784 9592 15818 9626
rect 15874 9592 15908 9626
rect 15964 9592 15998 9626
rect 16054 9592 16088 9626
rect 16144 9592 16178 9626
rect 16442 9592 16476 9626
rect 16532 9592 16566 9626
rect 16622 9592 16656 9626
rect 16712 9592 16746 9626
rect 16802 9592 16836 9626
rect 16892 9592 16926 9626
rect 16982 9592 17016 9626
rect 17072 9592 17106 9626
rect 17162 9592 17196 9626
rect 17252 9592 17286 9626
rect 17342 9592 17376 9626
rect 17432 9592 17466 9626
rect 17730 9592 17764 9626
rect 17820 9592 17854 9626
rect 17910 9592 17944 9626
rect 18000 9592 18034 9626
rect 18090 9592 18124 9626
rect 18180 9592 18214 9626
rect 18270 9592 18304 9626
rect 18360 9592 18394 9626
rect 18450 9592 18484 9626
rect 18540 9592 18574 9626
rect 18630 9592 18664 9626
rect 18720 9592 18754 9626
rect 12477 9508 12511 9542
rect 13664 9508 13698 9542
rect 13765 9508 13799 9542
rect -17882 9050 -11430 9382
rect -20918 5760 -19926 5836
rect -22304 5106 -21904 5682
rect -18938 5106 -18538 5682
rect -17434 5042 -17334 6642
rect -11934 5042 -11834 6642
rect 12477 9418 12511 9452
rect 12477 9328 12511 9362
rect 12477 9238 12511 9272
rect 12477 9148 12511 9182
rect 12477 9058 12511 9092
rect 12477 8968 12511 9002
rect 12477 8878 12511 8912
rect 12477 8788 12511 8822
rect 12477 8698 12511 8732
rect 12477 8608 12511 8642
rect 12477 8518 12511 8552
rect 14952 9508 14986 9542
rect 15053 9508 15087 9542
rect 13664 9418 13698 9452
rect 13765 9418 13799 9452
rect 13664 9328 13698 9362
rect 13765 9328 13799 9362
rect 13664 9238 13698 9272
rect 13765 9238 13799 9272
rect 13664 9148 13698 9182
rect 13765 9148 13799 9182
rect 13664 9058 13698 9092
rect 13765 9058 13799 9092
rect 13664 8968 13698 9002
rect 13765 8968 13799 9002
rect 13664 8878 13698 8912
rect 13765 8878 13799 8912
rect 13664 8788 13698 8822
rect 13765 8788 13799 8822
rect 13664 8698 13698 8732
rect 13765 8698 13799 8732
rect 13664 8608 13698 8642
rect 13765 8608 13799 8642
rect 13664 8518 13698 8552
rect 13765 8518 13799 8552
rect 16240 9508 16274 9542
rect 16341 9508 16375 9542
rect 14952 9418 14986 9452
rect 15053 9418 15087 9452
rect 14952 9328 14986 9362
rect 15053 9328 15087 9362
rect 14952 9238 14986 9272
rect 15053 9238 15087 9272
rect 14952 9148 14986 9182
rect 15053 9148 15087 9182
rect 14952 9058 14986 9092
rect 15053 9058 15087 9092
rect 14952 8968 14986 9002
rect 15053 8968 15087 9002
rect 14952 8878 14986 8912
rect 15053 8878 15087 8912
rect 14952 8788 14986 8822
rect 15053 8788 15087 8822
rect 14952 8698 14986 8732
rect 15053 8698 15087 8732
rect 14952 8608 14986 8642
rect 15053 8608 15087 8642
rect 14952 8518 14986 8552
rect 15053 8518 15087 8552
rect 17528 9508 17562 9542
rect 17629 9508 17663 9542
rect 16240 9418 16274 9452
rect 16341 9418 16375 9452
rect 16240 9328 16274 9362
rect 16341 9328 16375 9362
rect 16240 9238 16274 9272
rect 16341 9238 16375 9272
rect 16240 9148 16274 9182
rect 16341 9148 16375 9182
rect 16240 9058 16274 9092
rect 16341 9058 16375 9092
rect 16240 8968 16274 9002
rect 16341 8968 16375 9002
rect 16240 8878 16274 8912
rect 16341 8878 16375 8912
rect 16240 8788 16274 8822
rect 16341 8788 16375 8822
rect 16240 8698 16274 8732
rect 16341 8698 16375 8732
rect 16240 8608 16274 8642
rect 16341 8608 16375 8642
rect 16240 8518 16274 8552
rect 16341 8518 16375 8552
rect 18816 9508 18850 9542
rect 17528 9418 17562 9452
rect 17629 9418 17663 9452
rect 17528 9328 17562 9362
rect 17629 9328 17663 9362
rect 17528 9238 17562 9272
rect 17629 9238 17663 9272
rect 17528 9148 17562 9182
rect 17629 9148 17663 9182
rect 17528 9058 17562 9092
rect 17629 9058 17663 9092
rect 17528 8968 17562 9002
rect 17629 8968 17663 9002
rect 17528 8878 17562 8912
rect 17629 8878 17663 8912
rect 17528 8788 17562 8822
rect 17629 8788 17663 8822
rect 17528 8698 17562 8732
rect 17629 8698 17663 8732
rect 17528 8608 17562 8642
rect 17629 8608 17663 8642
rect 17528 8518 17562 8552
rect 17629 8518 17663 8552
rect 18816 9418 18850 9452
rect 18816 9328 18850 9362
rect 18816 9238 18850 9272
rect 18816 9148 18850 9182
rect 18816 9058 18850 9092
rect 18816 8968 18850 9002
rect 18816 8878 18850 8912
rect 18816 8788 18850 8822
rect 18816 8698 18850 8732
rect 18816 8608 18850 8642
rect 18816 8518 18850 8552
rect 12477 8428 12511 8462
rect 12578 8405 12612 8439
rect 12668 8405 12702 8439
rect 12758 8405 12792 8439
rect 12848 8405 12882 8439
rect 12938 8405 12972 8439
rect 13028 8405 13062 8439
rect 13118 8405 13152 8439
rect 13208 8405 13242 8439
rect 13298 8405 13332 8439
rect 13388 8405 13422 8439
rect 13478 8405 13512 8439
rect 13568 8405 13602 8439
rect 13664 8428 13698 8462
rect 13765 8428 13799 8462
rect 13866 8405 13900 8439
rect 13956 8405 13990 8439
rect 14046 8405 14080 8439
rect 14136 8405 14170 8439
rect 14226 8405 14260 8439
rect 14316 8405 14350 8439
rect 14406 8405 14440 8439
rect 14496 8405 14530 8439
rect 14586 8405 14620 8439
rect 14676 8405 14710 8439
rect 14766 8405 14800 8439
rect 14856 8405 14890 8439
rect 14952 8428 14986 8462
rect 15053 8428 15087 8462
rect 15154 8405 15188 8439
rect 15244 8405 15278 8439
rect 15334 8405 15368 8439
rect 15424 8405 15458 8439
rect 15514 8405 15548 8439
rect 15604 8405 15638 8439
rect 15694 8405 15728 8439
rect 15784 8405 15818 8439
rect 15874 8405 15908 8439
rect 15964 8405 15998 8439
rect 16054 8405 16088 8439
rect 16144 8405 16178 8439
rect 16240 8428 16274 8462
rect 16341 8428 16375 8462
rect 16442 8405 16476 8439
rect 16532 8405 16566 8439
rect 16622 8405 16656 8439
rect 16712 8405 16746 8439
rect 16802 8405 16836 8439
rect 16892 8405 16926 8439
rect 16982 8405 17016 8439
rect 17072 8405 17106 8439
rect 17162 8405 17196 8439
rect 17252 8405 17286 8439
rect 17342 8405 17376 8439
rect 17432 8405 17466 8439
rect 17528 8428 17562 8462
rect 17629 8428 17663 8462
rect 17730 8405 17764 8439
rect 17820 8405 17854 8439
rect 17910 8405 17944 8439
rect 18000 8405 18034 8439
rect 18090 8405 18124 8439
rect 18180 8405 18214 8439
rect 18270 8405 18304 8439
rect 18360 8405 18394 8439
rect 18450 8405 18484 8439
rect 18540 8405 18574 8439
rect 18630 8405 18664 8439
rect 18720 8405 18754 8439
rect 18816 8428 18850 8462
rect 12578 8304 12612 8338
rect 12668 8304 12702 8338
rect 12758 8304 12792 8338
rect 12848 8304 12882 8338
rect 12938 8304 12972 8338
rect 13028 8304 13062 8338
rect 13118 8304 13152 8338
rect 13208 8304 13242 8338
rect 13298 8304 13332 8338
rect 13388 8304 13422 8338
rect 13478 8304 13512 8338
rect 13568 8304 13602 8338
rect 13866 8304 13900 8338
rect 13956 8304 13990 8338
rect 14046 8304 14080 8338
rect 14136 8304 14170 8338
rect 14226 8304 14260 8338
rect 14316 8304 14350 8338
rect 14406 8304 14440 8338
rect 14496 8304 14530 8338
rect 14586 8304 14620 8338
rect 14676 8304 14710 8338
rect 14766 8304 14800 8338
rect 14856 8304 14890 8338
rect 15154 8304 15188 8338
rect 15244 8304 15278 8338
rect 15334 8304 15368 8338
rect 15424 8304 15458 8338
rect 15514 8304 15548 8338
rect 15604 8304 15638 8338
rect 15694 8304 15728 8338
rect 15784 8304 15818 8338
rect 15874 8304 15908 8338
rect 15964 8304 15998 8338
rect 16054 8304 16088 8338
rect 16144 8304 16178 8338
rect 16442 8304 16476 8338
rect 16532 8304 16566 8338
rect 16622 8304 16656 8338
rect 16712 8304 16746 8338
rect 16802 8304 16836 8338
rect 16892 8304 16926 8338
rect 16982 8304 17016 8338
rect 17072 8304 17106 8338
rect 17162 8304 17196 8338
rect 17252 8304 17286 8338
rect 17342 8304 17376 8338
rect 17432 8304 17466 8338
rect 17730 8304 17764 8338
rect 17820 8304 17854 8338
rect 17910 8304 17944 8338
rect 18000 8304 18034 8338
rect 18090 8304 18124 8338
rect 18180 8304 18214 8338
rect 18270 8304 18304 8338
rect 18360 8304 18394 8338
rect 18450 8304 18484 8338
rect 18540 8304 18574 8338
rect 18630 8304 18664 8338
rect 18720 8304 18754 8338
rect 12477 8220 12511 8254
rect 13664 8220 13698 8254
rect 13765 8220 13799 8254
rect 12477 8130 12511 8164
rect 12477 8040 12511 8074
rect 12477 7950 12511 7984
rect 12477 7860 12511 7894
rect 12477 7770 12511 7804
rect 12477 7680 12511 7714
rect 12477 7590 12511 7624
rect 12477 7500 12511 7534
rect 12477 7410 12511 7444
rect 12477 7320 12511 7354
rect 12477 7230 12511 7264
rect 14952 8220 14986 8254
rect 15053 8220 15087 8254
rect 13664 8130 13698 8164
rect 13765 8130 13799 8164
rect 13664 8040 13698 8074
rect 13765 8040 13799 8074
rect 13664 7950 13698 7984
rect 13765 7950 13799 7984
rect 13664 7860 13698 7894
rect 13765 7860 13799 7894
rect 13664 7770 13698 7804
rect 13765 7770 13799 7804
rect 13664 7680 13698 7714
rect 13765 7680 13799 7714
rect 13664 7590 13698 7624
rect 13765 7590 13799 7624
rect 13664 7500 13698 7534
rect 13765 7500 13799 7534
rect 13664 7410 13698 7444
rect 13765 7410 13799 7444
rect 13664 7320 13698 7354
rect 13765 7320 13799 7354
rect 13664 7230 13698 7264
rect 13765 7230 13799 7264
rect 16240 8220 16274 8254
rect 16341 8220 16375 8254
rect 14952 8130 14986 8164
rect 15053 8130 15087 8164
rect 14952 8040 14986 8074
rect 15053 8040 15087 8074
rect 14952 7950 14986 7984
rect 15053 7950 15087 7984
rect 14952 7860 14986 7894
rect 15053 7860 15087 7894
rect 14952 7770 14986 7804
rect 15053 7770 15087 7804
rect 14952 7680 14986 7714
rect 15053 7680 15087 7714
rect 14952 7590 14986 7624
rect 15053 7590 15087 7624
rect 14952 7500 14986 7534
rect 15053 7500 15087 7534
rect 14952 7410 14986 7444
rect 15053 7410 15087 7444
rect 14952 7320 14986 7354
rect 15053 7320 15087 7354
rect 14952 7230 14986 7264
rect 15053 7230 15087 7264
rect 17528 8220 17562 8254
rect 17629 8220 17663 8254
rect 16240 8130 16274 8164
rect 16341 8130 16375 8164
rect 16240 8040 16274 8074
rect 16341 8040 16375 8074
rect 16240 7950 16274 7984
rect 16341 7950 16375 7984
rect 16240 7860 16274 7894
rect 16341 7860 16375 7894
rect 16240 7770 16274 7804
rect 16341 7770 16375 7804
rect 16240 7680 16274 7714
rect 16341 7680 16375 7714
rect 16240 7590 16274 7624
rect 16341 7590 16375 7624
rect 16240 7500 16274 7534
rect 16341 7500 16375 7534
rect 16240 7410 16274 7444
rect 16341 7410 16375 7444
rect 16240 7320 16274 7354
rect 16341 7320 16375 7354
rect 16240 7230 16274 7264
rect 16341 7230 16375 7264
rect 18816 8220 18850 8254
rect 17528 8130 17562 8164
rect 17629 8130 17663 8164
rect 17528 8040 17562 8074
rect 17629 8040 17663 8074
rect 17528 7950 17562 7984
rect 17629 7950 17663 7984
rect 17528 7860 17562 7894
rect 17629 7860 17663 7894
rect 17528 7770 17562 7804
rect 17629 7770 17663 7804
rect 17528 7680 17562 7714
rect 17629 7680 17663 7714
rect 17528 7590 17562 7624
rect 17629 7590 17663 7624
rect 17528 7500 17562 7534
rect 17629 7500 17663 7534
rect 17528 7410 17562 7444
rect 17629 7410 17663 7444
rect 17528 7320 17562 7354
rect 17629 7320 17663 7354
rect 17528 7230 17562 7264
rect 17629 7230 17663 7264
rect 18816 8130 18850 8164
rect 18816 8040 18850 8074
rect 18816 7950 18850 7984
rect 18816 7860 18850 7894
rect 18816 7770 18850 7804
rect 18816 7680 18850 7714
rect 18816 7590 18850 7624
rect 18816 7500 18850 7534
rect 18816 7410 18850 7444
rect 18816 7320 18850 7354
rect 18816 7230 18850 7264
rect 12477 7140 12511 7174
rect 12578 7117 12612 7151
rect 12668 7117 12702 7151
rect 12758 7117 12792 7151
rect 12848 7117 12882 7151
rect 12938 7117 12972 7151
rect 13028 7117 13062 7151
rect 13118 7117 13152 7151
rect 13208 7117 13242 7151
rect 13298 7117 13332 7151
rect 13388 7117 13422 7151
rect 13478 7117 13512 7151
rect 13568 7117 13602 7151
rect 13664 7140 13698 7174
rect 13765 7140 13799 7174
rect 13866 7117 13900 7151
rect 13956 7117 13990 7151
rect 14046 7117 14080 7151
rect 14136 7117 14170 7151
rect 14226 7117 14260 7151
rect 14316 7117 14350 7151
rect 14406 7117 14440 7151
rect 14496 7117 14530 7151
rect 14586 7117 14620 7151
rect 14676 7117 14710 7151
rect 14766 7117 14800 7151
rect 14856 7117 14890 7151
rect 14952 7140 14986 7174
rect 15053 7140 15087 7174
rect 15154 7117 15188 7151
rect 15244 7117 15278 7151
rect 15334 7117 15368 7151
rect 15424 7117 15458 7151
rect 15514 7117 15548 7151
rect 15604 7117 15638 7151
rect 15694 7117 15728 7151
rect 15784 7117 15818 7151
rect 15874 7117 15908 7151
rect 15964 7117 15998 7151
rect 16054 7117 16088 7151
rect 16144 7117 16178 7151
rect 16240 7140 16274 7174
rect 16341 7140 16375 7174
rect 16442 7117 16476 7151
rect 16532 7117 16566 7151
rect 16622 7117 16656 7151
rect 16712 7117 16746 7151
rect 16802 7117 16836 7151
rect 16892 7117 16926 7151
rect 16982 7117 17016 7151
rect 17072 7117 17106 7151
rect 17162 7117 17196 7151
rect 17252 7117 17286 7151
rect 17342 7117 17376 7151
rect 17432 7117 17466 7151
rect 17528 7140 17562 7174
rect 17629 7140 17663 7174
rect 17730 7117 17764 7151
rect 17820 7117 17854 7151
rect 17910 7117 17944 7151
rect 18000 7117 18034 7151
rect 18090 7117 18124 7151
rect 18180 7117 18214 7151
rect 18270 7117 18304 7151
rect 18360 7117 18394 7151
rect 18450 7117 18484 7151
rect 18540 7117 18574 7151
rect 18630 7117 18664 7151
rect 18720 7117 18754 7151
rect 18816 7140 18850 7174
rect 12578 7016 12612 7050
rect 12668 7016 12702 7050
rect 12758 7016 12792 7050
rect 12848 7016 12882 7050
rect 12938 7016 12972 7050
rect 13028 7016 13062 7050
rect 13118 7016 13152 7050
rect 13208 7016 13242 7050
rect 13298 7016 13332 7050
rect 13388 7016 13422 7050
rect 13478 7016 13512 7050
rect 13568 7016 13602 7050
rect 13866 7016 13900 7050
rect 13956 7016 13990 7050
rect 14046 7016 14080 7050
rect 14136 7016 14170 7050
rect 14226 7016 14260 7050
rect 14316 7016 14350 7050
rect 14406 7016 14440 7050
rect 14496 7016 14530 7050
rect 14586 7016 14620 7050
rect 14676 7016 14710 7050
rect 14766 7016 14800 7050
rect 14856 7016 14890 7050
rect 15154 7016 15188 7050
rect 15244 7016 15278 7050
rect 15334 7016 15368 7050
rect 15424 7016 15458 7050
rect 15514 7016 15548 7050
rect 15604 7016 15638 7050
rect 15694 7016 15728 7050
rect 15784 7016 15818 7050
rect 15874 7016 15908 7050
rect 15964 7016 15998 7050
rect 16054 7016 16088 7050
rect 16144 7016 16178 7050
rect 16442 7016 16476 7050
rect 16532 7016 16566 7050
rect 16622 7016 16656 7050
rect 16712 7016 16746 7050
rect 16802 7016 16836 7050
rect 16892 7016 16926 7050
rect 16982 7016 17016 7050
rect 17072 7016 17106 7050
rect 17162 7016 17196 7050
rect 17252 7016 17286 7050
rect 17342 7016 17376 7050
rect 17432 7016 17466 7050
rect 17730 7016 17764 7050
rect 17820 7016 17854 7050
rect 17910 7016 17944 7050
rect 18000 7016 18034 7050
rect 18090 7016 18124 7050
rect 18180 7016 18214 7050
rect 18270 7016 18304 7050
rect 18360 7016 18394 7050
rect 18450 7016 18484 7050
rect 18540 7016 18574 7050
rect 18630 7016 18664 7050
rect 18720 7016 18754 7050
rect 12477 6932 12511 6966
rect 13664 6932 13698 6966
rect 13765 6932 13799 6966
rect 12477 6842 12511 6876
rect 12477 6752 12511 6786
rect 12477 6662 12511 6696
rect 12477 6572 12511 6606
rect 12477 6482 12511 6516
rect 12477 6392 12511 6426
rect 12477 6302 12511 6336
rect 12477 6212 12511 6246
rect 12477 6122 12511 6156
rect 12477 6032 12511 6066
rect 12477 5942 12511 5976
rect 14952 6932 14986 6966
rect 15053 6932 15087 6966
rect 13664 6842 13698 6876
rect 13765 6842 13799 6876
rect 13664 6752 13698 6786
rect 13765 6752 13799 6786
rect 13664 6662 13698 6696
rect 13765 6662 13799 6696
rect 13664 6572 13698 6606
rect 13765 6572 13799 6606
rect 13664 6482 13698 6516
rect 13765 6482 13799 6516
rect 13664 6392 13698 6426
rect 13765 6392 13799 6426
rect 13664 6302 13698 6336
rect 13765 6302 13799 6336
rect 13664 6212 13698 6246
rect 13765 6212 13799 6246
rect 13664 6122 13698 6156
rect 13765 6122 13799 6156
rect 13664 6032 13698 6066
rect 13765 6032 13799 6066
rect 13664 5942 13698 5976
rect 13765 5942 13799 5976
rect 16240 6932 16274 6966
rect 16341 6932 16375 6966
rect 14952 6842 14986 6876
rect 15053 6842 15087 6876
rect 14952 6752 14986 6786
rect 15053 6752 15087 6786
rect 14952 6662 14986 6696
rect 15053 6662 15087 6696
rect 14952 6572 14986 6606
rect 15053 6572 15087 6606
rect 14952 6482 14986 6516
rect 15053 6482 15087 6516
rect 14952 6392 14986 6426
rect 15053 6392 15087 6426
rect 14952 6302 14986 6336
rect 15053 6302 15087 6336
rect 14952 6212 14986 6246
rect 15053 6212 15087 6246
rect 14952 6122 14986 6156
rect 15053 6122 15087 6156
rect 14952 6032 14986 6066
rect 15053 6032 15087 6066
rect 14952 5942 14986 5976
rect 15053 5942 15087 5976
rect 17528 6932 17562 6966
rect 17629 6932 17663 6966
rect 16240 6842 16274 6876
rect 16341 6842 16375 6876
rect 16240 6752 16274 6786
rect 16341 6752 16375 6786
rect 16240 6662 16274 6696
rect 16341 6662 16375 6696
rect 16240 6572 16274 6606
rect 16341 6572 16375 6606
rect 16240 6482 16274 6516
rect 16341 6482 16375 6516
rect 16240 6392 16274 6426
rect 16341 6392 16375 6426
rect 16240 6302 16274 6336
rect 16341 6302 16375 6336
rect 16240 6212 16274 6246
rect 16341 6212 16375 6246
rect 16240 6122 16274 6156
rect 16341 6122 16375 6156
rect 16240 6032 16274 6066
rect 16341 6032 16375 6066
rect 16240 5942 16274 5976
rect 16341 5942 16375 5976
rect 18816 6932 18850 6966
rect 17528 6842 17562 6876
rect 17629 6842 17663 6876
rect 17528 6752 17562 6786
rect 17629 6752 17663 6786
rect 17528 6662 17562 6696
rect 17629 6662 17663 6696
rect 17528 6572 17562 6606
rect 17629 6572 17663 6606
rect 17528 6482 17562 6516
rect 17629 6482 17663 6516
rect 17528 6392 17562 6426
rect 17629 6392 17663 6426
rect 17528 6302 17562 6336
rect 17629 6302 17663 6336
rect 17528 6212 17562 6246
rect 17629 6212 17663 6246
rect 17528 6122 17562 6156
rect 17629 6122 17663 6156
rect 17528 6032 17562 6066
rect 17629 6032 17663 6066
rect 17528 5942 17562 5976
rect 17629 5942 17663 5976
rect 18816 6842 18850 6876
rect 18816 6752 18850 6786
rect 18816 6662 18850 6696
rect 18816 6572 18850 6606
rect 18816 6482 18850 6516
rect 18816 6392 18850 6426
rect 18816 6302 18850 6336
rect 18816 6212 18850 6246
rect 18816 6122 18850 6156
rect 18816 6032 18850 6066
rect 18816 5942 18850 5976
rect 12477 5852 12511 5886
rect 12578 5829 12612 5863
rect 12668 5829 12702 5863
rect 12758 5829 12792 5863
rect 12848 5829 12882 5863
rect 12938 5829 12972 5863
rect 13028 5829 13062 5863
rect 13118 5829 13152 5863
rect 13208 5829 13242 5863
rect 13298 5829 13332 5863
rect 13388 5829 13422 5863
rect 13478 5829 13512 5863
rect 13568 5829 13602 5863
rect 13664 5852 13698 5886
rect 13765 5852 13799 5886
rect 13866 5829 13900 5863
rect 13956 5829 13990 5863
rect 14046 5829 14080 5863
rect 14136 5829 14170 5863
rect 14226 5829 14260 5863
rect 14316 5829 14350 5863
rect 14406 5829 14440 5863
rect 14496 5829 14530 5863
rect 14586 5829 14620 5863
rect 14676 5829 14710 5863
rect 14766 5829 14800 5863
rect 14856 5829 14890 5863
rect 14952 5852 14986 5886
rect 15053 5852 15087 5886
rect 15154 5829 15188 5863
rect 15244 5829 15278 5863
rect 15334 5829 15368 5863
rect 15424 5829 15458 5863
rect 15514 5829 15548 5863
rect 15604 5829 15638 5863
rect 15694 5829 15728 5863
rect 15784 5829 15818 5863
rect 15874 5829 15908 5863
rect 15964 5829 15998 5863
rect 16054 5829 16088 5863
rect 16144 5829 16178 5863
rect 16240 5852 16274 5886
rect 16341 5852 16375 5886
rect 16442 5829 16476 5863
rect 16532 5829 16566 5863
rect 16622 5829 16656 5863
rect 16712 5829 16746 5863
rect 16802 5829 16836 5863
rect 16892 5829 16926 5863
rect 16982 5829 17016 5863
rect 17072 5829 17106 5863
rect 17162 5829 17196 5863
rect 17252 5829 17286 5863
rect 17342 5829 17376 5863
rect 17432 5829 17466 5863
rect 17528 5852 17562 5886
rect 17629 5852 17663 5886
rect 17730 5829 17764 5863
rect 17820 5829 17854 5863
rect 17910 5829 17944 5863
rect 18000 5829 18034 5863
rect 18090 5829 18124 5863
rect 18180 5829 18214 5863
rect 18270 5829 18304 5863
rect 18360 5829 18394 5863
rect 18450 5829 18484 5863
rect 18540 5829 18574 5863
rect 18630 5829 18664 5863
rect 18720 5829 18754 5863
rect 18816 5852 18850 5886
rect 12578 5728 12612 5762
rect 12668 5728 12702 5762
rect 12758 5728 12792 5762
rect 12848 5728 12882 5762
rect 12938 5728 12972 5762
rect 13028 5728 13062 5762
rect 13118 5728 13152 5762
rect 13208 5728 13242 5762
rect 13298 5728 13332 5762
rect 13388 5728 13422 5762
rect 13478 5728 13512 5762
rect 13568 5728 13602 5762
rect 13866 5728 13900 5762
rect 13956 5728 13990 5762
rect 14046 5728 14080 5762
rect 14136 5728 14170 5762
rect 14226 5728 14260 5762
rect 14316 5728 14350 5762
rect 14406 5728 14440 5762
rect 14496 5728 14530 5762
rect 14586 5728 14620 5762
rect 14676 5728 14710 5762
rect 14766 5728 14800 5762
rect 14856 5728 14890 5762
rect 15154 5728 15188 5762
rect 15244 5728 15278 5762
rect 15334 5728 15368 5762
rect 15424 5728 15458 5762
rect 15514 5728 15548 5762
rect 15604 5728 15638 5762
rect 15694 5728 15728 5762
rect 15784 5728 15818 5762
rect 15874 5728 15908 5762
rect 15964 5728 15998 5762
rect 16054 5728 16088 5762
rect 16144 5728 16178 5762
rect 16442 5728 16476 5762
rect 16532 5728 16566 5762
rect 16622 5728 16656 5762
rect 16712 5728 16746 5762
rect 16802 5728 16836 5762
rect 16892 5728 16926 5762
rect 16982 5728 17016 5762
rect 17072 5728 17106 5762
rect 17162 5728 17196 5762
rect 17252 5728 17286 5762
rect 17342 5728 17376 5762
rect 17432 5728 17466 5762
rect 17730 5728 17764 5762
rect 17820 5728 17854 5762
rect 17910 5728 17944 5762
rect 18000 5728 18034 5762
rect 18090 5728 18124 5762
rect 18180 5728 18214 5762
rect 18270 5728 18304 5762
rect 18360 5728 18394 5762
rect 18450 5728 18484 5762
rect 18540 5728 18574 5762
rect 18630 5728 18664 5762
rect 18720 5728 18754 5762
rect 12477 5644 12511 5678
rect 13664 5644 13698 5678
rect 13765 5644 13799 5678
rect 12477 5554 12511 5588
rect 12477 5464 12511 5498
rect 12477 5374 12511 5408
rect 12477 5284 12511 5318
rect 12477 5194 12511 5228
rect 12477 5104 12511 5138
rect 12477 5014 12511 5048
rect 12477 4924 12511 4958
rect 12477 4834 12511 4868
rect 12477 4744 12511 4778
rect 12477 4654 12511 4688
rect 14952 5644 14986 5678
rect 15053 5644 15087 5678
rect 13664 5554 13698 5588
rect 13765 5554 13799 5588
rect 13664 5464 13698 5498
rect 13765 5464 13799 5498
rect 13664 5374 13698 5408
rect 13765 5374 13799 5408
rect 13664 5284 13698 5318
rect 13765 5284 13799 5318
rect 13664 5194 13698 5228
rect 13765 5194 13799 5228
rect 13664 5104 13698 5138
rect 13765 5104 13799 5138
rect 13664 5014 13698 5048
rect 13765 5014 13799 5048
rect 13664 4924 13698 4958
rect 13765 4924 13799 4958
rect 13664 4834 13698 4868
rect 13765 4834 13799 4868
rect 13664 4744 13698 4778
rect 13765 4744 13799 4778
rect 13664 4654 13698 4688
rect 13765 4654 13799 4688
rect 16240 5644 16274 5678
rect 16341 5644 16375 5678
rect 14952 5554 14986 5588
rect 15053 5554 15087 5588
rect 14952 5464 14986 5498
rect 15053 5464 15087 5498
rect 14952 5374 14986 5408
rect 15053 5374 15087 5408
rect 14952 5284 14986 5318
rect 15053 5284 15087 5318
rect 14952 5194 14986 5228
rect 15053 5194 15087 5228
rect 14952 5104 14986 5138
rect 15053 5104 15087 5138
rect 14952 5014 14986 5048
rect 15053 5014 15087 5048
rect 14952 4924 14986 4958
rect 15053 4924 15087 4958
rect 14952 4834 14986 4868
rect 15053 4834 15087 4868
rect 14952 4744 14986 4778
rect 15053 4744 15087 4778
rect 14952 4654 14986 4688
rect 15053 4654 15087 4688
rect 17528 5644 17562 5678
rect 17629 5644 17663 5678
rect 16240 5554 16274 5588
rect 16341 5554 16375 5588
rect 16240 5464 16274 5498
rect 16341 5464 16375 5498
rect 16240 5374 16274 5408
rect 16341 5374 16375 5408
rect 16240 5284 16274 5318
rect 16341 5284 16375 5318
rect 16240 5194 16274 5228
rect 16341 5194 16375 5228
rect 16240 5104 16274 5138
rect 16341 5104 16375 5138
rect 16240 5014 16274 5048
rect 16341 5014 16375 5048
rect 16240 4924 16274 4958
rect 16341 4924 16375 4958
rect 16240 4834 16274 4868
rect 16341 4834 16375 4868
rect 16240 4744 16274 4778
rect 16341 4744 16375 4778
rect 16240 4654 16274 4688
rect 16341 4654 16375 4688
rect 18816 5644 18850 5678
rect 17528 5554 17562 5588
rect 17629 5554 17663 5588
rect 17528 5464 17562 5498
rect 17629 5464 17663 5498
rect 17528 5374 17562 5408
rect 17629 5374 17663 5408
rect 17528 5284 17562 5318
rect 17629 5284 17663 5318
rect 17528 5194 17562 5228
rect 17629 5194 17663 5228
rect 17528 5104 17562 5138
rect 17629 5104 17663 5138
rect 17528 5014 17562 5048
rect 17629 5014 17663 5048
rect 17528 4924 17562 4958
rect 17629 4924 17663 4958
rect 17528 4834 17562 4868
rect 17629 4834 17663 4868
rect 17528 4744 17562 4778
rect 17629 4744 17663 4778
rect 17528 4654 17562 4688
rect 17629 4654 17663 4688
rect 18816 5554 18850 5588
rect 18816 5464 18850 5498
rect 18816 5374 18850 5408
rect 18816 5284 18850 5318
rect 18816 5194 18850 5228
rect 18816 5104 18850 5138
rect 18816 5014 18850 5048
rect 18816 4924 18850 4958
rect 18816 4834 18850 4868
rect 18816 4744 18850 4778
rect 18816 4654 18850 4688
rect 12477 4564 12511 4598
rect 12578 4541 12612 4575
rect 12668 4541 12702 4575
rect 12758 4541 12792 4575
rect 12848 4541 12882 4575
rect 12938 4541 12972 4575
rect 13028 4541 13062 4575
rect 13118 4541 13152 4575
rect 13208 4541 13242 4575
rect 13298 4541 13332 4575
rect 13388 4541 13422 4575
rect 13478 4541 13512 4575
rect 13568 4541 13602 4575
rect 13664 4564 13698 4598
rect 13765 4564 13799 4598
rect 13866 4541 13900 4575
rect 13956 4541 13990 4575
rect 14046 4541 14080 4575
rect 14136 4541 14170 4575
rect 14226 4541 14260 4575
rect 14316 4541 14350 4575
rect 14406 4541 14440 4575
rect 14496 4541 14530 4575
rect 14586 4541 14620 4575
rect 14676 4541 14710 4575
rect 14766 4541 14800 4575
rect 14856 4541 14890 4575
rect 14952 4564 14986 4598
rect 15053 4564 15087 4598
rect 15154 4541 15188 4575
rect 15244 4541 15278 4575
rect 15334 4541 15368 4575
rect 15424 4541 15458 4575
rect 15514 4541 15548 4575
rect 15604 4541 15638 4575
rect 15694 4541 15728 4575
rect 15784 4541 15818 4575
rect 15874 4541 15908 4575
rect 15964 4541 15998 4575
rect 16054 4541 16088 4575
rect 16144 4541 16178 4575
rect 16240 4564 16274 4598
rect 16341 4564 16375 4598
rect 16442 4541 16476 4575
rect 16532 4541 16566 4575
rect 16622 4541 16656 4575
rect 16712 4541 16746 4575
rect 16802 4541 16836 4575
rect 16892 4541 16926 4575
rect 16982 4541 17016 4575
rect 17072 4541 17106 4575
rect 17162 4541 17196 4575
rect 17252 4541 17286 4575
rect 17342 4541 17376 4575
rect 17432 4541 17466 4575
rect 17528 4564 17562 4598
rect 17629 4564 17663 4598
rect 17730 4541 17764 4575
rect 17820 4541 17854 4575
rect 17910 4541 17944 4575
rect 18000 4541 18034 4575
rect 18090 4541 18124 4575
rect 18180 4541 18214 4575
rect 18270 4541 18304 4575
rect 18360 4541 18394 4575
rect 18450 4541 18484 4575
rect 18540 4541 18574 4575
rect 18630 4541 18664 4575
rect 18720 4541 18754 4575
rect 18816 4564 18850 4598
rect 12578 4440 12612 4474
rect 12668 4440 12702 4474
rect 12758 4440 12792 4474
rect 12848 4440 12882 4474
rect 12938 4440 12972 4474
rect 13028 4440 13062 4474
rect 13118 4440 13152 4474
rect 13208 4440 13242 4474
rect 13298 4440 13332 4474
rect 13388 4440 13422 4474
rect 13478 4440 13512 4474
rect 13568 4440 13602 4474
rect 13866 4440 13900 4474
rect 13956 4440 13990 4474
rect 14046 4440 14080 4474
rect 14136 4440 14170 4474
rect 14226 4440 14260 4474
rect 14316 4440 14350 4474
rect 14406 4440 14440 4474
rect 14496 4440 14530 4474
rect 14586 4440 14620 4474
rect 14676 4440 14710 4474
rect 14766 4440 14800 4474
rect 14856 4440 14890 4474
rect 15154 4440 15188 4474
rect 15244 4440 15278 4474
rect 15334 4440 15368 4474
rect 15424 4440 15458 4474
rect 15514 4440 15548 4474
rect 15604 4440 15638 4474
rect 15694 4440 15728 4474
rect 15784 4440 15818 4474
rect 15874 4440 15908 4474
rect 15964 4440 15998 4474
rect 16054 4440 16088 4474
rect 16144 4440 16178 4474
rect 16442 4440 16476 4474
rect 16532 4440 16566 4474
rect 16622 4440 16656 4474
rect 16712 4440 16746 4474
rect 16802 4440 16836 4474
rect 16892 4440 16926 4474
rect 16982 4440 17016 4474
rect 17072 4440 17106 4474
rect 17162 4440 17196 4474
rect 17252 4440 17286 4474
rect 17342 4440 17376 4474
rect 17432 4440 17466 4474
rect 17730 4440 17764 4474
rect 17820 4440 17854 4474
rect 17910 4440 17944 4474
rect 18000 4440 18034 4474
rect 18090 4440 18124 4474
rect 18180 4440 18214 4474
rect 18270 4440 18304 4474
rect 18360 4440 18394 4474
rect 18450 4440 18484 4474
rect 18540 4440 18574 4474
rect 18630 4440 18664 4474
rect 18720 4440 18754 4474
rect 12477 4356 12511 4390
rect 13664 4356 13698 4390
rect 13765 4356 13799 4390
rect 12477 4266 12511 4300
rect 12477 4176 12511 4210
rect 12477 4086 12511 4120
rect 12477 3996 12511 4030
rect 12477 3906 12511 3940
rect 12477 3816 12511 3850
rect 12477 3726 12511 3760
rect 12477 3636 12511 3670
rect 12477 3546 12511 3580
rect 12477 3456 12511 3490
rect 12477 3366 12511 3400
rect 14952 4356 14986 4390
rect 15053 4356 15087 4390
rect 13664 4266 13698 4300
rect 13765 4266 13799 4300
rect 13664 4176 13698 4210
rect 13765 4176 13799 4210
rect 13664 4086 13698 4120
rect 13765 4086 13799 4120
rect 13664 3996 13698 4030
rect 13765 3996 13799 4030
rect 13664 3906 13698 3940
rect 13765 3906 13799 3940
rect 13664 3816 13698 3850
rect 13765 3816 13799 3850
rect 13664 3726 13698 3760
rect 13765 3726 13799 3760
rect 13664 3636 13698 3670
rect 13765 3636 13799 3670
rect 13664 3546 13698 3580
rect 13765 3546 13799 3580
rect 13664 3456 13698 3490
rect 13765 3456 13799 3490
rect 13664 3366 13698 3400
rect 13765 3366 13799 3400
rect 16240 4356 16274 4390
rect 16341 4356 16375 4390
rect 14952 4266 14986 4300
rect 15053 4266 15087 4300
rect 14952 4176 14986 4210
rect 15053 4176 15087 4210
rect 14952 4086 14986 4120
rect 15053 4086 15087 4120
rect 14952 3996 14986 4030
rect 15053 3996 15087 4030
rect 14952 3906 14986 3940
rect 15053 3906 15087 3940
rect 14952 3816 14986 3850
rect 15053 3816 15087 3850
rect 14952 3726 14986 3760
rect 15053 3726 15087 3760
rect 14952 3636 14986 3670
rect 15053 3636 15087 3670
rect 14952 3546 14986 3580
rect 15053 3546 15087 3580
rect 14952 3456 14986 3490
rect 15053 3456 15087 3490
rect 14952 3366 14986 3400
rect 15053 3366 15087 3400
rect 17528 4356 17562 4390
rect 17629 4356 17663 4390
rect 16240 4266 16274 4300
rect 16341 4266 16375 4300
rect 16240 4176 16274 4210
rect 16341 4176 16375 4210
rect 16240 4086 16274 4120
rect 16341 4086 16375 4120
rect 16240 3996 16274 4030
rect 16341 3996 16375 4030
rect 16240 3906 16274 3940
rect 16341 3906 16375 3940
rect 16240 3816 16274 3850
rect 16341 3816 16375 3850
rect 16240 3726 16274 3760
rect 16341 3726 16375 3760
rect 16240 3636 16274 3670
rect 16341 3636 16375 3670
rect 16240 3546 16274 3580
rect 16341 3546 16375 3580
rect 16240 3456 16274 3490
rect 16341 3456 16375 3490
rect 16240 3366 16274 3400
rect 16341 3366 16375 3400
rect 18816 4356 18850 4390
rect 17528 4266 17562 4300
rect 17629 4266 17663 4300
rect 17528 4176 17562 4210
rect 17629 4176 17663 4210
rect 17528 4086 17562 4120
rect 17629 4086 17663 4120
rect 17528 3996 17562 4030
rect 17629 3996 17663 4030
rect 17528 3906 17562 3940
rect 17629 3906 17663 3940
rect 17528 3816 17562 3850
rect 17629 3816 17663 3850
rect 17528 3726 17562 3760
rect 17629 3726 17663 3760
rect 17528 3636 17562 3670
rect 17629 3636 17663 3670
rect 17528 3546 17562 3580
rect 17629 3546 17663 3580
rect 17528 3456 17562 3490
rect 17629 3456 17663 3490
rect 17528 3366 17562 3400
rect 17629 3366 17663 3400
rect 18816 4266 18850 4300
rect 18816 4176 18850 4210
rect 18816 4086 18850 4120
rect 18816 3996 18850 4030
rect 18816 3906 18850 3940
rect 18816 3816 18850 3850
rect 18816 3726 18850 3760
rect 18816 3636 18850 3670
rect 18816 3546 18850 3580
rect 18816 3456 18850 3490
rect 18816 3366 18850 3400
rect 12477 3276 12511 3310
rect 12578 3253 12612 3287
rect 12668 3253 12702 3287
rect 12758 3253 12792 3287
rect 12848 3253 12882 3287
rect 12938 3253 12972 3287
rect 13028 3253 13062 3287
rect 13118 3253 13152 3287
rect 13208 3253 13242 3287
rect 13298 3253 13332 3287
rect 13388 3253 13422 3287
rect 13478 3253 13512 3287
rect 13568 3253 13602 3287
rect 13664 3276 13698 3310
rect 13765 3276 13799 3310
rect 13866 3253 13900 3287
rect 13956 3253 13990 3287
rect 14046 3253 14080 3287
rect 14136 3253 14170 3287
rect 14226 3253 14260 3287
rect 14316 3253 14350 3287
rect 14406 3253 14440 3287
rect 14496 3253 14530 3287
rect 14586 3253 14620 3287
rect 14676 3253 14710 3287
rect 14766 3253 14800 3287
rect 14856 3253 14890 3287
rect 14952 3276 14986 3310
rect 15053 3276 15087 3310
rect 15154 3253 15188 3287
rect 15244 3253 15278 3287
rect 15334 3253 15368 3287
rect 15424 3253 15458 3287
rect 15514 3253 15548 3287
rect 15604 3253 15638 3287
rect 15694 3253 15728 3287
rect 15784 3253 15818 3287
rect 15874 3253 15908 3287
rect 15964 3253 15998 3287
rect 16054 3253 16088 3287
rect 16144 3253 16178 3287
rect 16240 3276 16274 3310
rect 16341 3276 16375 3310
rect 16442 3253 16476 3287
rect 16532 3253 16566 3287
rect 16622 3253 16656 3287
rect 16712 3253 16746 3287
rect 16802 3253 16836 3287
rect 16892 3253 16926 3287
rect 16982 3253 17016 3287
rect 17072 3253 17106 3287
rect 17162 3253 17196 3287
rect 17252 3253 17286 3287
rect 17342 3253 17376 3287
rect 17432 3253 17466 3287
rect 17528 3276 17562 3310
rect 17629 3276 17663 3310
rect 17730 3253 17764 3287
rect 17820 3253 17854 3287
rect 17910 3253 17944 3287
rect 18000 3253 18034 3287
rect 18090 3253 18124 3287
rect 18180 3253 18214 3287
rect 18270 3253 18304 3287
rect 18360 3253 18394 3287
rect 18450 3253 18484 3287
rect 18540 3253 18574 3287
rect 18630 3253 18664 3287
rect 18720 3253 18754 3287
rect 18816 3276 18850 3310
rect 12578 3152 12612 3186
rect 12668 3152 12702 3186
rect 12758 3152 12792 3186
rect 12848 3152 12882 3186
rect 12938 3152 12972 3186
rect 13028 3152 13062 3186
rect 13118 3152 13152 3186
rect 13208 3152 13242 3186
rect 13298 3152 13332 3186
rect 13388 3152 13422 3186
rect 13478 3152 13512 3186
rect 13568 3152 13602 3186
rect 13866 3152 13900 3186
rect 13956 3152 13990 3186
rect 14046 3152 14080 3186
rect 14136 3152 14170 3186
rect 14226 3152 14260 3186
rect 14316 3152 14350 3186
rect 14406 3152 14440 3186
rect 14496 3152 14530 3186
rect 14586 3152 14620 3186
rect 14676 3152 14710 3186
rect 14766 3152 14800 3186
rect 14856 3152 14890 3186
rect 15154 3152 15188 3186
rect 15244 3152 15278 3186
rect 15334 3152 15368 3186
rect 15424 3152 15458 3186
rect 15514 3152 15548 3186
rect 15604 3152 15638 3186
rect 15694 3152 15728 3186
rect 15784 3152 15818 3186
rect 15874 3152 15908 3186
rect 15964 3152 15998 3186
rect 16054 3152 16088 3186
rect 16144 3152 16178 3186
rect 16442 3152 16476 3186
rect 16532 3152 16566 3186
rect 16622 3152 16656 3186
rect 16712 3152 16746 3186
rect 16802 3152 16836 3186
rect 16892 3152 16926 3186
rect 16982 3152 17016 3186
rect 17072 3152 17106 3186
rect 17162 3152 17196 3186
rect 17252 3152 17286 3186
rect 17342 3152 17376 3186
rect 17432 3152 17466 3186
rect 17730 3152 17764 3186
rect 17820 3152 17854 3186
rect 17910 3152 17944 3186
rect 18000 3152 18034 3186
rect 18090 3152 18124 3186
rect 18180 3152 18214 3186
rect 18270 3152 18304 3186
rect 18360 3152 18394 3186
rect 18450 3152 18484 3186
rect 18540 3152 18574 3186
rect 18630 3152 18664 3186
rect 18720 3152 18754 3186
rect 12477 3068 12511 3102
rect 13664 3068 13698 3102
rect 13765 3068 13799 3102
rect 12477 2978 12511 3012
rect 12477 2888 12511 2922
rect 12477 2798 12511 2832
rect 12477 2708 12511 2742
rect 12477 2618 12511 2652
rect 12477 2528 12511 2562
rect 12477 2438 12511 2472
rect 12477 2348 12511 2382
rect 12477 2258 12511 2292
rect 12477 2168 12511 2202
rect 12477 2078 12511 2112
rect 14952 3068 14986 3102
rect 15053 3068 15087 3102
rect 13664 2978 13698 3012
rect 13765 2978 13799 3012
rect 13664 2888 13698 2922
rect 13765 2888 13799 2922
rect 13664 2798 13698 2832
rect 13765 2798 13799 2832
rect 13664 2708 13698 2742
rect 13765 2708 13799 2742
rect 13664 2618 13698 2652
rect 13765 2618 13799 2652
rect 13664 2528 13698 2562
rect 13765 2528 13799 2562
rect 13664 2438 13698 2472
rect 13765 2438 13799 2472
rect 13664 2348 13698 2382
rect 13765 2348 13799 2382
rect 13664 2258 13698 2292
rect 13765 2258 13799 2292
rect 13664 2168 13698 2202
rect 13765 2168 13799 2202
rect 13664 2078 13698 2112
rect 13765 2078 13799 2112
rect 16240 3068 16274 3102
rect 16341 3068 16375 3102
rect 14952 2978 14986 3012
rect 15053 2978 15087 3012
rect 14952 2888 14986 2922
rect 15053 2888 15087 2922
rect 14952 2798 14986 2832
rect 15053 2798 15087 2832
rect 14952 2708 14986 2742
rect 15053 2708 15087 2742
rect 14952 2618 14986 2652
rect 15053 2618 15087 2652
rect 14952 2528 14986 2562
rect 15053 2528 15087 2562
rect 14952 2438 14986 2472
rect 15053 2438 15087 2472
rect 14952 2348 14986 2382
rect 15053 2348 15087 2382
rect 14952 2258 14986 2292
rect 15053 2258 15087 2292
rect 14952 2168 14986 2202
rect 15053 2168 15087 2202
rect 14952 2078 14986 2112
rect 15053 2078 15087 2112
rect 17528 3068 17562 3102
rect 17629 3068 17663 3102
rect 16240 2978 16274 3012
rect 16341 2978 16375 3012
rect 16240 2888 16274 2922
rect 16341 2888 16375 2922
rect 16240 2798 16274 2832
rect 16341 2798 16375 2832
rect 16240 2708 16274 2742
rect 16341 2708 16375 2742
rect 16240 2618 16274 2652
rect 16341 2618 16375 2652
rect 16240 2528 16274 2562
rect 16341 2528 16375 2562
rect 16240 2438 16274 2472
rect 16341 2438 16375 2472
rect 16240 2348 16274 2382
rect 16341 2348 16375 2382
rect 16240 2258 16274 2292
rect 16341 2258 16375 2292
rect 16240 2168 16274 2202
rect 16341 2168 16375 2202
rect 16240 2078 16274 2112
rect 16341 2078 16375 2112
rect 18816 3068 18850 3102
rect 17528 2978 17562 3012
rect 17629 2978 17663 3012
rect 17528 2888 17562 2922
rect 17629 2888 17663 2922
rect 17528 2798 17562 2832
rect 17629 2798 17663 2832
rect 17528 2708 17562 2742
rect 17629 2708 17663 2742
rect 17528 2618 17562 2652
rect 17629 2618 17663 2652
rect 17528 2528 17562 2562
rect 17629 2528 17663 2562
rect 17528 2438 17562 2472
rect 17629 2438 17663 2472
rect 17528 2348 17562 2382
rect 17629 2348 17663 2382
rect 17528 2258 17562 2292
rect 17629 2258 17663 2292
rect 17528 2168 17562 2202
rect 17629 2168 17663 2202
rect 17528 2078 17562 2112
rect 17629 2078 17663 2112
rect 18816 2978 18850 3012
rect 18816 2888 18850 2922
rect 18816 2798 18850 2832
rect 18816 2708 18850 2742
rect 18816 2618 18850 2652
rect 18816 2528 18850 2562
rect 18816 2438 18850 2472
rect 18816 2348 18850 2382
rect 18816 2258 18850 2292
rect 18816 2168 18850 2202
rect 18816 2078 18850 2112
rect 12477 1988 12511 2022
rect 12578 1965 12612 1999
rect 12668 1965 12702 1999
rect 12758 1965 12792 1999
rect 12848 1965 12882 1999
rect 12938 1965 12972 1999
rect 13028 1965 13062 1999
rect 13118 1965 13152 1999
rect 13208 1965 13242 1999
rect 13298 1965 13332 1999
rect 13388 1965 13422 1999
rect 13478 1965 13512 1999
rect 13568 1965 13602 1999
rect 13664 1988 13698 2022
rect 13765 1988 13799 2022
rect 13866 1965 13900 1999
rect 13956 1965 13990 1999
rect 14046 1965 14080 1999
rect 14136 1965 14170 1999
rect 14226 1965 14260 1999
rect 14316 1965 14350 1999
rect 14406 1965 14440 1999
rect 14496 1965 14530 1999
rect 14586 1965 14620 1999
rect 14676 1965 14710 1999
rect 14766 1965 14800 1999
rect 14856 1965 14890 1999
rect 14952 1988 14986 2022
rect 15053 1988 15087 2022
rect 15154 1965 15188 1999
rect 15244 1965 15278 1999
rect 15334 1965 15368 1999
rect 15424 1965 15458 1999
rect 15514 1965 15548 1999
rect 15604 1965 15638 1999
rect 15694 1965 15728 1999
rect 15784 1965 15818 1999
rect 15874 1965 15908 1999
rect 15964 1965 15998 1999
rect 16054 1965 16088 1999
rect 16144 1965 16178 1999
rect 16240 1988 16274 2022
rect 16341 1988 16375 2022
rect 16442 1965 16476 1999
rect 16532 1965 16566 1999
rect 16622 1965 16656 1999
rect 16712 1965 16746 1999
rect 16802 1965 16836 1999
rect 16892 1965 16926 1999
rect 16982 1965 17016 1999
rect 17072 1965 17106 1999
rect 17162 1965 17196 1999
rect 17252 1965 17286 1999
rect 17342 1965 17376 1999
rect 17432 1965 17466 1999
rect 17528 1988 17562 2022
rect 17629 1988 17663 2022
rect 17730 1965 17764 1999
rect 17820 1965 17854 1999
rect 17910 1965 17944 1999
rect 18000 1965 18034 1999
rect 18090 1965 18124 1999
rect 18180 1965 18214 1999
rect 18270 1965 18304 1999
rect 18360 1965 18394 1999
rect 18450 1965 18484 1999
rect 18540 1965 18574 1999
rect 18630 1965 18664 1999
rect 18720 1965 18754 1999
rect 18816 1988 18850 2022
<< nsubdiffcont >>
rect 12718 12018 12752 12052
rect 12808 12018 12842 12052
rect 12898 12018 12932 12052
rect 12988 12018 13022 12052
rect 13078 12018 13112 12052
rect 13168 12018 13202 12052
rect 13258 12018 13292 12052
rect 13348 12018 13382 12052
rect 13438 12018 13472 12052
rect 12626 11924 12660 11958
rect 12626 11834 12660 11868
rect 12626 11744 12660 11778
rect 12626 11654 12660 11688
rect 12626 11564 12660 11598
rect 12626 11474 12660 11508
rect 12626 11384 12660 11418
rect 12626 11294 12660 11328
rect 13516 11905 13550 11939
rect 13516 11815 13550 11849
rect 13516 11725 13550 11759
rect 13516 11635 13550 11669
rect 13516 11545 13550 11579
rect 13516 11455 13550 11489
rect 13516 11365 13550 11399
rect 13516 11275 13550 11309
rect 12626 11204 12660 11238
rect 13516 11185 13550 11219
rect 12684 11128 12718 11162
rect 12774 11128 12808 11162
rect 12864 11128 12898 11162
rect 12954 11128 12988 11162
rect 13044 11128 13078 11162
rect 13134 11128 13168 11162
rect 13224 11128 13258 11162
rect 13314 11128 13348 11162
rect 13404 11128 13438 11162
rect 14006 12018 14040 12052
rect 14096 12018 14130 12052
rect 14186 12018 14220 12052
rect 14276 12018 14310 12052
rect 14366 12018 14400 12052
rect 14456 12018 14490 12052
rect 14546 12018 14580 12052
rect 14636 12018 14670 12052
rect 14726 12018 14760 12052
rect 13914 11924 13948 11958
rect 13914 11834 13948 11868
rect 13914 11744 13948 11778
rect 13914 11654 13948 11688
rect 13914 11564 13948 11598
rect 13914 11474 13948 11508
rect 13914 11384 13948 11418
rect 13914 11294 13948 11328
rect 14804 11905 14838 11939
rect 14804 11815 14838 11849
rect 14804 11725 14838 11759
rect 14804 11635 14838 11669
rect 14804 11545 14838 11579
rect 14804 11455 14838 11489
rect 14804 11365 14838 11399
rect 14804 11275 14838 11309
rect 13914 11204 13948 11238
rect 14804 11185 14838 11219
rect 13972 11128 14006 11162
rect 14062 11128 14096 11162
rect 14152 11128 14186 11162
rect 14242 11128 14276 11162
rect 14332 11128 14366 11162
rect 14422 11128 14456 11162
rect 14512 11128 14546 11162
rect 14602 11128 14636 11162
rect 14692 11128 14726 11162
rect 15294 12018 15328 12052
rect 15384 12018 15418 12052
rect 15474 12018 15508 12052
rect 15564 12018 15598 12052
rect 15654 12018 15688 12052
rect 15744 12018 15778 12052
rect 15834 12018 15868 12052
rect 15924 12018 15958 12052
rect 16014 12018 16048 12052
rect 15202 11924 15236 11958
rect 15202 11834 15236 11868
rect 15202 11744 15236 11778
rect 15202 11654 15236 11688
rect 15202 11564 15236 11598
rect 15202 11474 15236 11508
rect 15202 11384 15236 11418
rect 15202 11294 15236 11328
rect 16092 11905 16126 11939
rect 16092 11815 16126 11849
rect 16092 11725 16126 11759
rect 16092 11635 16126 11669
rect 16092 11545 16126 11579
rect 16092 11455 16126 11489
rect 16092 11365 16126 11399
rect 16092 11275 16126 11309
rect 15202 11204 15236 11238
rect 16092 11185 16126 11219
rect 15260 11128 15294 11162
rect 15350 11128 15384 11162
rect 15440 11128 15474 11162
rect 15530 11128 15564 11162
rect 15620 11128 15654 11162
rect 15710 11128 15744 11162
rect 15800 11128 15834 11162
rect 15890 11128 15924 11162
rect 15980 11128 16014 11162
rect 16582 12018 16616 12052
rect 16672 12018 16706 12052
rect 16762 12018 16796 12052
rect 16852 12018 16886 12052
rect 16942 12018 16976 12052
rect 17032 12018 17066 12052
rect 17122 12018 17156 12052
rect 17212 12018 17246 12052
rect 17302 12018 17336 12052
rect 16490 11924 16524 11958
rect 16490 11834 16524 11868
rect 16490 11744 16524 11778
rect 16490 11654 16524 11688
rect 16490 11564 16524 11598
rect 16490 11474 16524 11508
rect 16490 11384 16524 11418
rect 16490 11294 16524 11328
rect 17380 11905 17414 11939
rect 17380 11815 17414 11849
rect 17380 11725 17414 11759
rect 17380 11635 17414 11669
rect 17380 11545 17414 11579
rect 17380 11455 17414 11489
rect 17380 11365 17414 11399
rect 17380 11275 17414 11309
rect 16490 11204 16524 11238
rect 17380 11185 17414 11219
rect 16548 11128 16582 11162
rect 16638 11128 16672 11162
rect 16728 11128 16762 11162
rect 16818 11128 16852 11162
rect 16908 11128 16942 11162
rect 16998 11128 17032 11162
rect 17088 11128 17122 11162
rect 17178 11128 17212 11162
rect 17268 11128 17302 11162
rect 17870 12018 17904 12052
rect 17960 12018 17994 12052
rect 18050 12018 18084 12052
rect 18140 12018 18174 12052
rect 18230 12018 18264 12052
rect 18320 12018 18354 12052
rect 18410 12018 18444 12052
rect 18500 12018 18534 12052
rect 18590 12018 18624 12052
rect 17778 11924 17812 11958
rect 17778 11834 17812 11868
rect 17778 11744 17812 11778
rect 17778 11654 17812 11688
rect 17778 11564 17812 11598
rect 17778 11474 17812 11508
rect 17778 11384 17812 11418
rect 17778 11294 17812 11328
rect 18668 11905 18702 11939
rect 18668 11815 18702 11849
rect 18668 11725 18702 11759
rect 18668 11635 18702 11669
rect 18668 11545 18702 11579
rect 18668 11455 18702 11489
rect 18668 11365 18702 11399
rect 18668 11275 18702 11309
rect 17778 11204 17812 11238
rect 18668 11185 18702 11219
rect 17836 11128 17870 11162
rect 17926 11128 17960 11162
rect 18016 11128 18050 11162
rect 18106 11128 18140 11162
rect 18196 11128 18230 11162
rect 18286 11128 18320 11162
rect 18376 11128 18410 11162
rect 18466 11128 18500 11162
rect 18556 11128 18590 11162
rect 12718 10730 12752 10764
rect 12808 10730 12842 10764
rect 12898 10730 12932 10764
rect 12988 10730 13022 10764
rect 13078 10730 13112 10764
rect 13168 10730 13202 10764
rect 13258 10730 13292 10764
rect 13348 10730 13382 10764
rect 13438 10730 13472 10764
rect 12626 10636 12660 10670
rect 12626 10546 12660 10580
rect 12626 10456 12660 10490
rect 12626 10366 12660 10400
rect 12626 10276 12660 10310
rect 12626 10186 12660 10220
rect 12626 10096 12660 10130
rect 12626 10006 12660 10040
rect 13516 10617 13550 10651
rect 13516 10527 13550 10561
rect 13516 10437 13550 10471
rect 13516 10347 13550 10381
rect 13516 10257 13550 10291
rect 13516 10167 13550 10201
rect 13516 10077 13550 10111
rect 13516 9987 13550 10021
rect 12626 9916 12660 9950
rect 13516 9897 13550 9931
rect 12684 9840 12718 9874
rect 12774 9840 12808 9874
rect 12864 9840 12898 9874
rect 12954 9840 12988 9874
rect 13044 9840 13078 9874
rect 13134 9840 13168 9874
rect 13224 9840 13258 9874
rect 13314 9840 13348 9874
rect 13404 9840 13438 9874
rect 14006 10730 14040 10764
rect 14096 10730 14130 10764
rect 14186 10730 14220 10764
rect 14276 10730 14310 10764
rect 14366 10730 14400 10764
rect 14456 10730 14490 10764
rect 14546 10730 14580 10764
rect 14636 10730 14670 10764
rect 14726 10730 14760 10764
rect 13914 10636 13948 10670
rect 13914 10546 13948 10580
rect 13914 10456 13948 10490
rect 13914 10366 13948 10400
rect 13914 10276 13948 10310
rect 13914 10186 13948 10220
rect 13914 10096 13948 10130
rect 13914 10006 13948 10040
rect 14804 10617 14838 10651
rect 14804 10527 14838 10561
rect 14804 10437 14838 10471
rect 14804 10347 14838 10381
rect 14804 10257 14838 10291
rect 14804 10167 14838 10201
rect 14804 10077 14838 10111
rect 14804 9987 14838 10021
rect 13914 9916 13948 9950
rect 14804 9897 14838 9931
rect 13972 9840 14006 9874
rect 14062 9840 14096 9874
rect 14152 9840 14186 9874
rect 14242 9840 14276 9874
rect 14332 9840 14366 9874
rect 14422 9840 14456 9874
rect 14512 9840 14546 9874
rect 14602 9840 14636 9874
rect 14692 9840 14726 9874
rect 15294 10730 15328 10764
rect 15384 10730 15418 10764
rect 15474 10730 15508 10764
rect 15564 10730 15598 10764
rect 15654 10730 15688 10764
rect 15744 10730 15778 10764
rect 15834 10730 15868 10764
rect 15924 10730 15958 10764
rect 16014 10730 16048 10764
rect 15202 10636 15236 10670
rect 15202 10546 15236 10580
rect 15202 10456 15236 10490
rect 15202 10366 15236 10400
rect 15202 10276 15236 10310
rect 15202 10186 15236 10220
rect 15202 10096 15236 10130
rect 15202 10006 15236 10040
rect 16092 10617 16126 10651
rect 16092 10527 16126 10561
rect 16092 10437 16126 10471
rect 16092 10347 16126 10381
rect 16092 10257 16126 10291
rect 16092 10167 16126 10201
rect 16092 10077 16126 10111
rect 16092 9987 16126 10021
rect 15202 9916 15236 9950
rect 16092 9897 16126 9931
rect 15260 9840 15294 9874
rect 15350 9840 15384 9874
rect 15440 9840 15474 9874
rect 15530 9840 15564 9874
rect 15620 9840 15654 9874
rect 15710 9840 15744 9874
rect 15800 9840 15834 9874
rect 15890 9840 15924 9874
rect 15980 9840 16014 9874
rect 16582 10730 16616 10764
rect 16672 10730 16706 10764
rect 16762 10730 16796 10764
rect 16852 10730 16886 10764
rect 16942 10730 16976 10764
rect 17032 10730 17066 10764
rect 17122 10730 17156 10764
rect 17212 10730 17246 10764
rect 17302 10730 17336 10764
rect 16490 10636 16524 10670
rect 16490 10546 16524 10580
rect 16490 10456 16524 10490
rect 16490 10366 16524 10400
rect 16490 10276 16524 10310
rect 16490 10186 16524 10220
rect 16490 10096 16524 10130
rect 16490 10006 16524 10040
rect 17380 10617 17414 10651
rect 17380 10527 17414 10561
rect 17380 10437 17414 10471
rect 17380 10347 17414 10381
rect 17380 10257 17414 10291
rect 17380 10167 17414 10201
rect 17380 10077 17414 10111
rect 17380 9987 17414 10021
rect 16490 9916 16524 9950
rect 17380 9897 17414 9931
rect 16548 9840 16582 9874
rect 16638 9840 16672 9874
rect 16728 9840 16762 9874
rect 16818 9840 16852 9874
rect 16908 9840 16942 9874
rect 16998 9840 17032 9874
rect 17088 9840 17122 9874
rect 17178 9840 17212 9874
rect 17268 9840 17302 9874
rect 17870 10730 17904 10764
rect 17960 10730 17994 10764
rect 18050 10730 18084 10764
rect 18140 10730 18174 10764
rect 18230 10730 18264 10764
rect 18320 10730 18354 10764
rect 18410 10730 18444 10764
rect 18500 10730 18534 10764
rect 18590 10730 18624 10764
rect 17778 10636 17812 10670
rect 17778 10546 17812 10580
rect 17778 10456 17812 10490
rect 17778 10366 17812 10400
rect 17778 10276 17812 10310
rect 17778 10186 17812 10220
rect 17778 10096 17812 10130
rect 17778 10006 17812 10040
rect 18668 10617 18702 10651
rect 18668 10527 18702 10561
rect 18668 10437 18702 10471
rect 18668 10347 18702 10381
rect 18668 10257 18702 10291
rect 18668 10167 18702 10201
rect 18668 10077 18702 10111
rect 18668 9987 18702 10021
rect 17778 9916 17812 9950
rect 18668 9897 18702 9931
rect 17836 9840 17870 9874
rect 17926 9840 17960 9874
rect 18016 9840 18050 9874
rect 18106 9840 18140 9874
rect 18196 9840 18230 9874
rect 18286 9840 18320 9874
rect 18376 9840 18410 9874
rect 18466 9840 18500 9874
rect 18556 9840 18590 9874
rect -19250 1800 -19150 4142
rect -10122 1800 -10022 4142
rect -9300 2102 -9100 9102
rect -3390 2102 -3190 9102
rect 2110 2102 2310 9102
rect 8066 2100 8266 9100
rect 12718 9442 12752 9476
rect 12808 9442 12842 9476
rect 12898 9442 12932 9476
rect 12988 9442 13022 9476
rect 13078 9442 13112 9476
rect 13168 9442 13202 9476
rect 13258 9442 13292 9476
rect 13348 9442 13382 9476
rect 13438 9442 13472 9476
rect 12626 9348 12660 9382
rect 12626 9258 12660 9292
rect 12626 9168 12660 9202
rect 12626 9078 12660 9112
rect 12626 8988 12660 9022
rect 12626 8898 12660 8932
rect 12626 8808 12660 8842
rect 12626 8718 12660 8752
rect 13516 9329 13550 9363
rect 13516 9239 13550 9273
rect 13516 9149 13550 9183
rect 13516 9059 13550 9093
rect 13516 8969 13550 9003
rect 13516 8879 13550 8913
rect 13516 8789 13550 8823
rect 13516 8699 13550 8733
rect 12626 8628 12660 8662
rect 13516 8609 13550 8643
rect 12684 8552 12718 8586
rect 12774 8552 12808 8586
rect 12864 8552 12898 8586
rect 12954 8552 12988 8586
rect 13044 8552 13078 8586
rect 13134 8552 13168 8586
rect 13224 8552 13258 8586
rect 13314 8552 13348 8586
rect 13404 8552 13438 8586
rect 14006 9442 14040 9476
rect 14096 9442 14130 9476
rect 14186 9442 14220 9476
rect 14276 9442 14310 9476
rect 14366 9442 14400 9476
rect 14456 9442 14490 9476
rect 14546 9442 14580 9476
rect 14636 9442 14670 9476
rect 14726 9442 14760 9476
rect 13914 9348 13948 9382
rect 13914 9258 13948 9292
rect 13914 9168 13948 9202
rect 13914 9078 13948 9112
rect 13914 8988 13948 9022
rect 13914 8898 13948 8932
rect 13914 8808 13948 8842
rect 13914 8718 13948 8752
rect 14804 9329 14838 9363
rect 14804 9239 14838 9273
rect 14804 9149 14838 9183
rect 14804 9059 14838 9093
rect 14804 8969 14838 9003
rect 14804 8879 14838 8913
rect 14804 8789 14838 8823
rect 14804 8699 14838 8733
rect 13914 8628 13948 8662
rect 14804 8609 14838 8643
rect 13972 8552 14006 8586
rect 14062 8552 14096 8586
rect 14152 8552 14186 8586
rect 14242 8552 14276 8586
rect 14332 8552 14366 8586
rect 14422 8552 14456 8586
rect 14512 8552 14546 8586
rect 14602 8552 14636 8586
rect 14692 8552 14726 8586
rect 15294 9442 15328 9476
rect 15384 9442 15418 9476
rect 15474 9442 15508 9476
rect 15564 9442 15598 9476
rect 15654 9442 15688 9476
rect 15744 9442 15778 9476
rect 15834 9442 15868 9476
rect 15924 9442 15958 9476
rect 16014 9442 16048 9476
rect 15202 9348 15236 9382
rect 15202 9258 15236 9292
rect 15202 9168 15236 9202
rect 15202 9078 15236 9112
rect 15202 8988 15236 9022
rect 15202 8898 15236 8932
rect 15202 8808 15236 8842
rect 15202 8718 15236 8752
rect 16092 9329 16126 9363
rect 16092 9239 16126 9273
rect 16092 9149 16126 9183
rect 16092 9059 16126 9093
rect 16092 8969 16126 9003
rect 16092 8879 16126 8913
rect 16092 8789 16126 8823
rect 16092 8699 16126 8733
rect 15202 8628 15236 8662
rect 16092 8609 16126 8643
rect 15260 8552 15294 8586
rect 15350 8552 15384 8586
rect 15440 8552 15474 8586
rect 15530 8552 15564 8586
rect 15620 8552 15654 8586
rect 15710 8552 15744 8586
rect 15800 8552 15834 8586
rect 15890 8552 15924 8586
rect 15980 8552 16014 8586
rect 16582 9442 16616 9476
rect 16672 9442 16706 9476
rect 16762 9442 16796 9476
rect 16852 9442 16886 9476
rect 16942 9442 16976 9476
rect 17032 9442 17066 9476
rect 17122 9442 17156 9476
rect 17212 9442 17246 9476
rect 17302 9442 17336 9476
rect 16490 9348 16524 9382
rect 16490 9258 16524 9292
rect 16490 9168 16524 9202
rect 16490 9078 16524 9112
rect 16490 8988 16524 9022
rect 16490 8898 16524 8932
rect 16490 8808 16524 8842
rect 16490 8718 16524 8752
rect 17380 9329 17414 9363
rect 17380 9239 17414 9273
rect 17380 9149 17414 9183
rect 17380 9059 17414 9093
rect 17380 8969 17414 9003
rect 17380 8879 17414 8913
rect 17380 8789 17414 8823
rect 17380 8699 17414 8733
rect 16490 8628 16524 8662
rect 17380 8609 17414 8643
rect 16548 8552 16582 8586
rect 16638 8552 16672 8586
rect 16728 8552 16762 8586
rect 16818 8552 16852 8586
rect 16908 8552 16942 8586
rect 16998 8552 17032 8586
rect 17088 8552 17122 8586
rect 17178 8552 17212 8586
rect 17268 8552 17302 8586
rect 17870 9442 17904 9476
rect 17960 9442 17994 9476
rect 18050 9442 18084 9476
rect 18140 9442 18174 9476
rect 18230 9442 18264 9476
rect 18320 9442 18354 9476
rect 18410 9442 18444 9476
rect 18500 9442 18534 9476
rect 18590 9442 18624 9476
rect 17778 9348 17812 9382
rect 17778 9258 17812 9292
rect 17778 9168 17812 9202
rect 17778 9078 17812 9112
rect 17778 8988 17812 9022
rect 17778 8898 17812 8932
rect 17778 8808 17812 8842
rect 17778 8718 17812 8752
rect 18668 9329 18702 9363
rect 18668 9239 18702 9273
rect 18668 9149 18702 9183
rect 18668 9059 18702 9093
rect 18668 8969 18702 9003
rect 18668 8879 18702 8913
rect 18668 8789 18702 8823
rect 18668 8699 18702 8733
rect 17778 8628 17812 8662
rect 18668 8609 18702 8643
rect 17836 8552 17870 8586
rect 17926 8552 17960 8586
rect 18016 8552 18050 8586
rect 18106 8552 18140 8586
rect 18196 8552 18230 8586
rect 18286 8552 18320 8586
rect 18376 8552 18410 8586
rect 18466 8552 18500 8586
rect 18556 8552 18590 8586
rect 12718 8154 12752 8188
rect 12808 8154 12842 8188
rect 12898 8154 12932 8188
rect 12988 8154 13022 8188
rect 13078 8154 13112 8188
rect 13168 8154 13202 8188
rect 13258 8154 13292 8188
rect 13348 8154 13382 8188
rect 13438 8154 13472 8188
rect 12626 8060 12660 8094
rect 12626 7970 12660 8004
rect 12626 7880 12660 7914
rect 12626 7790 12660 7824
rect 12626 7700 12660 7734
rect 12626 7610 12660 7644
rect 12626 7520 12660 7554
rect 12626 7430 12660 7464
rect 13516 8041 13550 8075
rect 13516 7951 13550 7985
rect 13516 7861 13550 7895
rect 13516 7771 13550 7805
rect 13516 7681 13550 7715
rect 13516 7591 13550 7625
rect 13516 7501 13550 7535
rect 13516 7411 13550 7445
rect 12626 7340 12660 7374
rect 13516 7321 13550 7355
rect 12684 7264 12718 7298
rect 12774 7264 12808 7298
rect 12864 7264 12898 7298
rect 12954 7264 12988 7298
rect 13044 7264 13078 7298
rect 13134 7264 13168 7298
rect 13224 7264 13258 7298
rect 13314 7264 13348 7298
rect 13404 7264 13438 7298
rect 14006 8154 14040 8188
rect 14096 8154 14130 8188
rect 14186 8154 14220 8188
rect 14276 8154 14310 8188
rect 14366 8154 14400 8188
rect 14456 8154 14490 8188
rect 14546 8154 14580 8188
rect 14636 8154 14670 8188
rect 14726 8154 14760 8188
rect 13914 8060 13948 8094
rect 13914 7970 13948 8004
rect 13914 7880 13948 7914
rect 13914 7790 13948 7824
rect 13914 7700 13948 7734
rect 13914 7610 13948 7644
rect 13914 7520 13948 7554
rect 13914 7430 13948 7464
rect 14804 8041 14838 8075
rect 14804 7951 14838 7985
rect 14804 7861 14838 7895
rect 14804 7771 14838 7805
rect 14804 7681 14838 7715
rect 14804 7591 14838 7625
rect 14804 7501 14838 7535
rect 14804 7411 14838 7445
rect 13914 7340 13948 7374
rect 14804 7321 14838 7355
rect 13972 7264 14006 7298
rect 14062 7264 14096 7298
rect 14152 7264 14186 7298
rect 14242 7264 14276 7298
rect 14332 7264 14366 7298
rect 14422 7264 14456 7298
rect 14512 7264 14546 7298
rect 14602 7264 14636 7298
rect 14692 7264 14726 7298
rect 15294 8154 15328 8188
rect 15384 8154 15418 8188
rect 15474 8154 15508 8188
rect 15564 8154 15598 8188
rect 15654 8154 15688 8188
rect 15744 8154 15778 8188
rect 15834 8154 15868 8188
rect 15924 8154 15958 8188
rect 16014 8154 16048 8188
rect 15202 8060 15236 8094
rect 15202 7970 15236 8004
rect 15202 7880 15236 7914
rect 15202 7790 15236 7824
rect 15202 7700 15236 7734
rect 15202 7610 15236 7644
rect 15202 7520 15236 7554
rect 15202 7430 15236 7464
rect 16092 8041 16126 8075
rect 16092 7951 16126 7985
rect 16092 7861 16126 7895
rect 16092 7771 16126 7805
rect 16092 7681 16126 7715
rect 16092 7591 16126 7625
rect 16092 7501 16126 7535
rect 16092 7411 16126 7445
rect 15202 7340 15236 7374
rect 16092 7321 16126 7355
rect 15260 7264 15294 7298
rect 15350 7264 15384 7298
rect 15440 7264 15474 7298
rect 15530 7264 15564 7298
rect 15620 7264 15654 7298
rect 15710 7264 15744 7298
rect 15800 7264 15834 7298
rect 15890 7264 15924 7298
rect 15980 7264 16014 7298
rect 16582 8154 16616 8188
rect 16672 8154 16706 8188
rect 16762 8154 16796 8188
rect 16852 8154 16886 8188
rect 16942 8154 16976 8188
rect 17032 8154 17066 8188
rect 17122 8154 17156 8188
rect 17212 8154 17246 8188
rect 17302 8154 17336 8188
rect 16490 8060 16524 8094
rect 16490 7970 16524 8004
rect 16490 7880 16524 7914
rect 16490 7790 16524 7824
rect 16490 7700 16524 7734
rect 16490 7610 16524 7644
rect 16490 7520 16524 7554
rect 16490 7430 16524 7464
rect 17380 8041 17414 8075
rect 17380 7951 17414 7985
rect 17380 7861 17414 7895
rect 17380 7771 17414 7805
rect 17380 7681 17414 7715
rect 17380 7591 17414 7625
rect 17380 7501 17414 7535
rect 17380 7411 17414 7445
rect 16490 7340 16524 7374
rect 17380 7321 17414 7355
rect 16548 7264 16582 7298
rect 16638 7264 16672 7298
rect 16728 7264 16762 7298
rect 16818 7264 16852 7298
rect 16908 7264 16942 7298
rect 16998 7264 17032 7298
rect 17088 7264 17122 7298
rect 17178 7264 17212 7298
rect 17268 7264 17302 7298
rect 17870 8154 17904 8188
rect 17960 8154 17994 8188
rect 18050 8154 18084 8188
rect 18140 8154 18174 8188
rect 18230 8154 18264 8188
rect 18320 8154 18354 8188
rect 18410 8154 18444 8188
rect 18500 8154 18534 8188
rect 18590 8154 18624 8188
rect 17778 8060 17812 8094
rect 17778 7970 17812 8004
rect 17778 7880 17812 7914
rect 17778 7790 17812 7824
rect 17778 7700 17812 7734
rect 17778 7610 17812 7644
rect 17778 7520 17812 7554
rect 17778 7430 17812 7464
rect 18668 8041 18702 8075
rect 18668 7951 18702 7985
rect 18668 7861 18702 7895
rect 18668 7771 18702 7805
rect 18668 7681 18702 7715
rect 18668 7591 18702 7625
rect 18668 7501 18702 7535
rect 18668 7411 18702 7445
rect 17778 7340 17812 7374
rect 18668 7321 18702 7355
rect 17836 7264 17870 7298
rect 17926 7264 17960 7298
rect 18016 7264 18050 7298
rect 18106 7264 18140 7298
rect 18196 7264 18230 7298
rect 18286 7264 18320 7298
rect 18376 7264 18410 7298
rect 18466 7264 18500 7298
rect 18556 7264 18590 7298
rect 12718 6866 12752 6900
rect 12808 6866 12842 6900
rect 12898 6866 12932 6900
rect 12988 6866 13022 6900
rect 13078 6866 13112 6900
rect 13168 6866 13202 6900
rect 13258 6866 13292 6900
rect 13348 6866 13382 6900
rect 13438 6866 13472 6900
rect 12626 6772 12660 6806
rect 12626 6682 12660 6716
rect 12626 6592 12660 6626
rect 12626 6502 12660 6536
rect 12626 6412 12660 6446
rect 12626 6322 12660 6356
rect 12626 6232 12660 6266
rect 12626 6142 12660 6176
rect 13516 6753 13550 6787
rect 13516 6663 13550 6697
rect 13516 6573 13550 6607
rect 13516 6483 13550 6517
rect 13516 6393 13550 6427
rect 13516 6303 13550 6337
rect 13516 6213 13550 6247
rect 13516 6123 13550 6157
rect 12626 6052 12660 6086
rect 13516 6033 13550 6067
rect 12684 5976 12718 6010
rect 12774 5976 12808 6010
rect 12864 5976 12898 6010
rect 12954 5976 12988 6010
rect 13044 5976 13078 6010
rect 13134 5976 13168 6010
rect 13224 5976 13258 6010
rect 13314 5976 13348 6010
rect 13404 5976 13438 6010
rect 14006 6866 14040 6900
rect 14096 6866 14130 6900
rect 14186 6866 14220 6900
rect 14276 6866 14310 6900
rect 14366 6866 14400 6900
rect 14456 6866 14490 6900
rect 14546 6866 14580 6900
rect 14636 6866 14670 6900
rect 14726 6866 14760 6900
rect 13914 6772 13948 6806
rect 13914 6682 13948 6716
rect 13914 6592 13948 6626
rect 13914 6502 13948 6536
rect 13914 6412 13948 6446
rect 13914 6322 13948 6356
rect 13914 6232 13948 6266
rect 13914 6142 13948 6176
rect 14804 6753 14838 6787
rect 14804 6663 14838 6697
rect 14804 6573 14838 6607
rect 14804 6483 14838 6517
rect 14804 6393 14838 6427
rect 14804 6303 14838 6337
rect 14804 6213 14838 6247
rect 14804 6123 14838 6157
rect 13914 6052 13948 6086
rect 14804 6033 14838 6067
rect 13972 5976 14006 6010
rect 14062 5976 14096 6010
rect 14152 5976 14186 6010
rect 14242 5976 14276 6010
rect 14332 5976 14366 6010
rect 14422 5976 14456 6010
rect 14512 5976 14546 6010
rect 14602 5976 14636 6010
rect 14692 5976 14726 6010
rect 15294 6866 15328 6900
rect 15384 6866 15418 6900
rect 15474 6866 15508 6900
rect 15564 6866 15598 6900
rect 15654 6866 15688 6900
rect 15744 6866 15778 6900
rect 15834 6866 15868 6900
rect 15924 6866 15958 6900
rect 16014 6866 16048 6900
rect 15202 6772 15236 6806
rect 15202 6682 15236 6716
rect 15202 6592 15236 6626
rect 15202 6502 15236 6536
rect 15202 6412 15236 6446
rect 15202 6322 15236 6356
rect 15202 6232 15236 6266
rect 15202 6142 15236 6176
rect 16092 6753 16126 6787
rect 16092 6663 16126 6697
rect 16092 6573 16126 6607
rect 16092 6483 16126 6517
rect 16092 6393 16126 6427
rect 16092 6303 16126 6337
rect 16092 6213 16126 6247
rect 16092 6123 16126 6157
rect 15202 6052 15236 6086
rect 16092 6033 16126 6067
rect 15260 5976 15294 6010
rect 15350 5976 15384 6010
rect 15440 5976 15474 6010
rect 15530 5976 15564 6010
rect 15620 5976 15654 6010
rect 15710 5976 15744 6010
rect 15800 5976 15834 6010
rect 15890 5976 15924 6010
rect 15980 5976 16014 6010
rect 16582 6866 16616 6900
rect 16672 6866 16706 6900
rect 16762 6866 16796 6900
rect 16852 6866 16886 6900
rect 16942 6866 16976 6900
rect 17032 6866 17066 6900
rect 17122 6866 17156 6900
rect 17212 6866 17246 6900
rect 17302 6866 17336 6900
rect 16490 6772 16524 6806
rect 16490 6682 16524 6716
rect 16490 6592 16524 6626
rect 16490 6502 16524 6536
rect 16490 6412 16524 6446
rect 16490 6322 16524 6356
rect 16490 6232 16524 6266
rect 16490 6142 16524 6176
rect 17380 6753 17414 6787
rect 17380 6663 17414 6697
rect 17380 6573 17414 6607
rect 17380 6483 17414 6517
rect 17380 6393 17414 6427
rect 17380 6303 17414 6337
rect 17380 6213 17414 6247
rect 17380 6123 17414 6157
rect 16490 6052 16524 6086
rect 17380 6033 17414 6067
rect 16548 5976 16582 6010
rect 16638 5976 16672 6010
rect 16728 5976 16762 6010
rect 16818 5976 16852 6010
rect 16908 5976 16942 6010
rect 16998 5976 17032 6010
rect 17088 5976 17122 6010
rect 17178 5976 17212 6010
rect 17268 5976 17302 6010
rect 17870 6866 17904 6900
rect 17960 6866 17994 6900
rect 18050 6866 18084 6900
rect 18140 6866 18174 6900
rect 18230 6866 18264 6900
rect 18320 6866 18354 6900
rect 18410 6866 18444 6900
rect 18500 6866 18534 6900
rect 18590 6866 18624 6900
rect 17778 6772 17812 6806
rect 17778 6682 17812 6716
rect 17778 6592 17812 6626
rect 17778 6502 17812 6536
rect 17778 6412 17812 6446
rect 17778 6322 17812 6356
rect 17778 6232 17812 6266
rect 17778 6142 17812 6176
rect 18668 6753 18702 6787
rect 18668 6663 18702 6697
rect 18668 6573 18702 6607
rect 18668 6483 18702 6517
rect 18668 6393 18702 6427
rect 18668 6303 18702 6337
rect 18668 6213 18702 6247
rect 18668 6123 18702 6157
rect 17778 6052 17812 6086
rect 18668 6033 18702 6067
rect 17836 5976 17870 6010
rect 17926 5976 17960 6010
rect 18016 5976 18050 6010
rect 18106 5976 18140 6010
rect 18196 5976 18230 6010
rect 18286 5976 18320 6010
rect 18376 5976 18410 6010
rect 18466 5976 18500 6010
rect 18556 5976 18590 6010
rect 12718 5578 12752 5612
rect 12808 5578 12842 5612
rect 12898 5578 12932 5612
rect 12988 5578 13022 5612
rect 13078 5578 13112 5612
rect 13168 5578 13202 5612
rect 13258 5578 13292 5612
rect 13348 5578 13382 5612
rect 13438 5578 13472 5612
rect 12626 5484 12660 5518
rect 12626 5394 12660 5428
rect 12626 5304 12660 5338
rect 12626 5214 12660 5248
rect 12626 5124 12660 5158
rect 12626 5034 12660 5068
rect 12626 4944 12660 4978
rect 12626 4854 12660 4888
rect 13516 5465 13550 5499
rect 13516 5375 13550 5409
rect 13516 5285 13550 5319
rect 13516 5195 13550 5229
rect 13516 5105 13550 5139
rect 13516 5015 13550 5049
rect 13516 4925 13550 4959
rect 13516 4835 13550 4869
rect 12626 4764 12660 4798
rect 13516 4745 13550 4779
rect 12684 4688 12718 4722
rect 12774 4688 12808 4722
rect 12864 4688 12898 4722
rect 12954 4688 12988 4722
rect 13044 4688 13078 4722
rect 13134 4688 13168 4722
rect 13224 4688 13258 4722
rect 13314 4688 13348 4722
rect 13404 4688 13438 4722
rect 14006 5578 14040 5612
rect 14096 5578 14130 5612
rect 14186 5578 14220 5612
rect 14276 5578 14310 5612
rect 14366 5578 14400 5612
rect 14456 5578 14490 5612
rect 14546 5578 14580 5612
rect 14636 5578 14670 5612
rect 14726 5578 14760 5612
rect 13914 5484 13948 5518
rect 13914 5394 13948 5428
rect 13914 5304 13948 5338
rect 13914 5214 13948 5248
rect 13914 5124 13948 5158
rect 13914 5034 13948 5068
rect 13914 4944 13948 4978
rect 13914 4854 13948 4888
rect 14804 5465 14838 5499
rect 14804 5375 14838 5409
rect 14804 5285 14838 5319
rect 14804 5195 14838 5229
rect 14804 5105 14838 5139
rect 14804 5015 14838 5049
rect 14804 4925 14838 4959
rect 14804 4835 14838 4869
rect 13914 4764 13948 4798
rect 14804 4745 14838 4779
rect 13972 4688 14006 4722
rect 14062 4688 14096 4722
rect 14152 4688 14186 4722
rect 14242 4688 14276 4722
rect 14332 4688 14366 4722
rect 14422 4688 14456 4722
rect 14512 4688 14546 4722
rect 14602 4688 14636 4722
rect 14692 4688 14726 4722
rect 15294 5578 15328 5612
rect 15384 5578 15418 5612
rect 15474 5578 15508 5612
rect 15564 5578 15598 5612
rect 15654 5578 15688 5612
rect 15744 5578 15778 5612
rect 15834 5578 15868 5612
rect 15924 5578 15958 5612
rect 16014 5578 16048 5612
rect 15202 5484 15236 5518
rect 15202 5394 15236 5428
rect 15202 5304 15236 5338
rect 15202 5214 15236 5248
rect 15202 5124 15236 5158
rect 15202 5034 15236 5068
rect 15202 4944 15236 4978
rect 15202 4854 15236 4888
rect 16092 5465 16126 5499
rect 16092 5375 16126 5409
rect 16092 5285 16126 5319
rect 16092 5195 16126 5229
rect 16092 5105 16126 5139
rect 16092 5015 16126 5049
rect 16092 4925 16126 4959
rect 16092 4835 16126 4869
rect 15202 4764 15236 4798
rect 16092 4745 16126 4779
rect 15260 4688 15294 4722
rect 15350 4688 15384 4722
rect 15440 4688 15474 4722
rect 15530 4688 15564 4722
rect 15620 4688 15654 4722
rect 15710 4688 15744 4722
rect 15800 4688 15834 4722
rect 15890 4688 15924 4722
rect 15980 4688 16014 4722
rect 16582 5578 16616 5612
rect 16672 5578 16706 5612
rect 16762 5578 16796 5612
rect 16852 5578 16886 5612
rect 16942 5578 16976 5612
rect 17032 5578 17066 5612
rect 17122 5578 17156 5612
rect 17212 5578 17246 5612
rect 17302 5578 17336 5612
rect 16490 5484 16524 5518
rect 16490 5394 16524 5428
rect 16490 5304 16524 5338
rect 16490 5214 16524 5248
rect 16490 5124 16524 5158
rect 16490 5034 16524 5068
rect 16490 4944 16524 4978
rect 16490 4854 16524 4888
rect 17380 5465 17414 5499
rect 17380 5375 17414 5409
rect 17380 5285 17414 5319
rect 17380 5195 17414 5229
rect 17380 5105 17414 5139
rect 17380 5015 17414 5049
rect 17380 4925 17414 4959
rect 17380 4835 17414 4869
rect 16490 4764 16524 4798
rect 17380 4745 17414 4779
rect 16548 4688 16582 4722
rect 16638 4688 16672 4722
rect 16728 4688 16762 4722
rect 16818 4688 16852 4722
rect 16908 4688 16942 4722
rect 16998 4688 17032 4722
rect 17088 4688 17122 4722
rect 17178 4688 17212 4722
rect 17268 4688 17302 4722
rect 17870 5578 17904 5612
rect 17960 5578 17994 5612
rect 18050 5578 18084 5612
rect 18140 5578 18174 5612
rect 18230 5578 18264 5612
rect 18320 5578 18354 5612
rect 18410 5578 18444 5612
rect 18500 5578 18534 5612
rect 18590 5578 18624 5612
rect 17778 5484 17812 5518
rect 17778 5394 17812 5428
rect 17778 5304 17812 5338
rect 17778 5214 17812 5248
rect 17778 5124 17812 5158
rect 17778 5034 17812 5068
rect 17778 4944 17812 4978
rect 17778 4854 17812 4888
rect 18668 5465 18702 5499
rect 18668 5375 18702 5409
rect 18668 5285 18702 5319
rect 18668 5195 18702 5229
rect 18668 5105 18702 5139
rect 18668 5015 18702 5049
rect 18668 4925 18702 4959
rect 18668 4835 18702 4869
rect 17778 4764 17812 4798
rect 18668 4745 18702 4779
rect 17836 4688 17870 4722
rect 17926 4688 17960 4722
rect 18016 4688 18050 4722
rect 18106 4688 18140 4722
rect 18196 4688 18230 4722
rect 18286 4688 18320 4722
rect 18376 4688 18410 4722
rect 18466 4688 18500 4722
rect 18556 4688 18590 4722
rect 12718 4290 12752 4324
rect 12808 4290 12842 4324
rect 12898 4290 12932 4324
rect 12988 4290 13022 4324
rect 13078 4290 13112 4324
rect 13168 4290 13202 4324
rect 13258 4290 13292 4324
rect 13348 4290 13382 4324
rect 13438 4290 13472 4324
rect 12626 4196 12660 4230
rect 12626 4106 12660 4140
rect 12626 4016 12660 4050
rect 12626 3926 12660 3960
rect 12626 3836 12660 3870
rect 12626 3746 12660 3780
rect 12626 3656 12660 3690
rect 12626 3566 12660 3600
rect 13516 4177 13550 4211
rect 13516 4087 13550 4121
rect 13516 3997 13550 4031
rect 13516 3907 13550 3941
rect 13516 3817 13550 3851
rect 13516 3727 13550 3761
rect 13516 3637 13550 3671
rect 13516 3547 13550 3581
rect 12626 3476 12660 3510
rect 13516 3457 13550 3491
rect 12684 3400 12718 3434
rect 12774 3400 12808 3434
rect 12864 3400 12898 3434
rect 12954 3400 12988 3434
rect 13044 3400 13078 3434
rect 13134 3400 13168 3434
rect 13224 3400 13258 3434
rect 13314 3400 13348 3434
rect 13404 3400 13438 3434
rect 14006 4290 14040 4324
rect 14096 4290 14130 4324
rect 14186 4290 14220 4324
rect 14276 4290 14310 4324
rect 14366 4290 14400 4324
rect 14456 4290 14490 4324
rect 14546 4290 14580 4324
rect 14636 4290 14670 4324
rect 14726 4290 14760 4324
rect 13914 4196 13948 4230
rect 13914 4106 13948 4140
rect 13914 4016 13948 4050
rect 13914 3926 13948 3960
rect 13914 3836 13948 3870
rect 13914 3746 13948 3780
rect 13914 3656 13948 3690
rect 13914 3566 13948 3600
rect 14804 4177 14838 4211
rect 14804 4087 14838 4121
rect 14804 3997 14838 4031
rect 14804 3907 14838 3941
rect 14804 3817 14838 3851
rect 14804 3727 14838 3761
rect 14804 3637 14838 3671
rect 14804 3547 14838 3581
rect 13914 3476 13948 3510
rect 14804 3457 14838 3491
rect 13972 3400 14006 3434
rect 14062 3400 14096 3434
rect 14152 3400 14186 3434
rect 14242 3400 14276 3434
rect 14332 3400 14366 3434
rect 14422 3400 14456 3434
rect 14512 3400 14546 3434
rect 14602 3400 14636 3434
rect 14692 3400 14726 3434
rect 15294 4290 15328 4324
rect 15384 4290 15418 4324
rect 15474 4290 15508 4324
rect 15564 4290 15598 4324
rect 15654 4290 15688 4324
rect 15744 4290 15778 4324
rect 15834 4290 15868 4324
rect 15924 4290 15958 4324
rect 16014 4290 16048 4324
rect 15202 4196 15236 4230
rect 15202 4106 15236 4140
rect 15202 4016 15236 4050
rect 15202 3926 15236 3960
rect 15202 3836 15236 3870
rect 15202 3746 15236 3780
rect 15202 3656 15236 3690
rect 15202 3566 15236 3600
rect 16092 4177 16126 4211
rect 16092 4087 16126 4121
rect 16092 3997 16126 4031
rect 16092 3907 16126 3941
rect 16092 3817 16126 3851
rect 16092 3727 16126 3761
rect 16092 3637 16126 3671
rect 16092 3547 16126 3581
rect 15202 3476 15236 3510
rect 16092 3457 16126 3491
rect 15260 3400 15294 3434
rect 15350 3400 15384 3434
rect 15440 3400 15474 3434
rect 15530 3400 15564 3434
rect 15620 3400 15654 3434
rect 15710 3400 15744 3434
rect 15800 3400 15834 3434
rect 15890 3400 15924 3434
rect 15980 3400 16014 3434
rect 16582 4290 16616 4324
rect 16672 4290 16706 4324
rect 16762 4290 16796 4324
rect 16852 4290 16886 4324
rect 16942 4290 16976 4324
rect 17032 4290 17066 4324
rect 17122 4290 17156 4324
rect 17212 4290 17246 4324
rect 17302 4290 17336 4324
rect 16490 4196 16524 4230
rect 16490 4106 16524 4140
rect 16490 4016 16524 4050
rect 16490 3926 16524 3960
rect 16490 3836 16524 3870
rect 16490 3746 16524 3780
rect 16490 3656 16524 3690
rect 16490 3566 16524 3600
rect 17380 4177 17414 4211
rect 17380 4087 17414 4121
rect 17380 3997 17414 4031
rect 17380 3907 17414 3941
rect 17380 3817 17414 3851
rect 17380 3727 17414 3761
rect 17380 3637 17414 3671
rect 17380 3547 17414 3581
rect 16490 3476 16524 3510
rect 17380 3457 17414 3491
rect 16548 3400 16582 3434
rect 16638 3400 16672 3434
rect 16728 3400 16762 3434
rect 16818 3400 16852 3434
rect 16908 3400 16942 3434
rect 16998 3400 17032 3434
rect 17088 3400 17122 3434
rect 17178 3400 17212 3434
rect 17268 3400 17302 3434
rect 17870 4290 17904 4324
rect 17960 4290 17994 4324
rect 18050 4290 18084 4324
rect 18140 4290 18174 4324
rect 18230 4290 18264 4324
rect 18320 4290 18354 4324
rect 18410 4290 18444 4324
rect 18500 4290 18534 4324
rect 18590 4290 18624 4324
rect 17778 4196 17812 4230
rect 17778 4106 17812 4140
rect 17778 4016 17812 4050
rect 17778 3926 17812 3960
rect 17778 3836 17812 3870
rect 17778 3746 17812 3780
rect 17778 3656 17812 3690
rect 17778 3566 17812 3600
rect 18668 4177 18702 4211
rect 18668 4087 18702 4121
rect 18668 3997 18702 4031
rect 18668 3907 18702 3941
rect 18668 3817 18702 3851
rect 18668 3727 18702 3761
rect 18668 3637 18702 3671
rect 18668 3547 18702 3581
rect 17778 3476 17812 3510
rect 18668 3457 18702 3491
rect 17836 3400 17870 3434
rect 17926 3400 17960 3434
rect 18016 3400 18050 3434
rect 18106 3400 18140 3434
rect 18196 3400 18230 3434
rect 18286 3400 18320 3434
rect 18376 3400 18410 3434
rect 18466 3400 18500 3434
rect 18556 3400 18590 3434
rect 12718 3002 12752 3036
rect 12808 3002 12842 3036
rect 12898 3002 12932 3036
rect 12988 3002 13022 3036
rect 13078 3002 13112 3036
rect 13168 3002 13202 3036
rect 13258 3002 13292 3036
rect 13348 3002 13382 3036
rect 13438 3002 13472 3036
rect 12626 2908 12660 2942
rect 12626 2818 12660 2852
rect 12626 2728 12660 2762
rect 12626 2638 12660 2672
rect 12626 2548 12660 2582
rect 12626 2458 12660 2492
rect 12626 2368 12660 2402
rect 12626 2278 12660 2312
rect 13516 2889 13550 2923
rect 13516 2799 13550 2833
rect 13516 2709 13550 2743
rect 13516 2619 13550 2653
rect 13516 2529 13550 2563
rect 13516 2439 13550 2473
rect 13516 2349 13550 2383
rect 13516 2259 13550 2293
rect 12626 2188 12660 2222
rect 13516 2169 13550 2203
rect 12684 2112 12718 2146
rect 12774 2112 12808 2146
rect 12864 2112 12898 2146
rect 12954 2112 12988 2146
rect 13044 2112 13078 2146
rect 13134 2112 13168 2146
rect 13224 2112 13258 2146
rect 13314 2112 13348 2146
rect 13404 2112 13438 2146
rect 14006 3002 14040 3036
rect 14096 3002 14130 3036
rect 14186 3002 14220 3036
rect 14276 3002 14310 3036
rect 14366 3002 14400 3036
rect 14456 3002 14490 3036
rect 14546 3002 14580 3036
rect 14636 3002 14670 3036
rect 14726 3002 14760 3036
rect 13914 2908 13948 2942
rect 13914 2818 13948 2852
rect 13914 2728 13948 2762
rect 13914 2638 13948 2672
rect 13914 2548 13948 2582
rect 13914 2458 13948 2492
rect 13914 2368 13948 2402
rect 13914 2278 13948 2312
rect 14804 2889 14838 2923
rect 14804 2799 14838 2833
rect 14804 2709 14838 2743
rect 14804 2619 14838 2653
rect 14804 2529 14838 2563
rect 14804 2439 14838 2473
rect 14804 2349 14838 2383
rect 14804 2259 14838 2293
rect 13914 2188 13948 2222
rect 14804 2169 14838 2203
rect 13972 2112 14006 2146
rect 14062 2112 14096 2146
rect 14152 2112 14186 2146
rect 14242 2112 14276 2146
rect 14332 2112 14366 2146
rect 14422 2112 14456 2146
rect 14512 2112 14546 2146
rect 14602 2112 14636 2146
rect 14692 2112 14726 2146
rect 15294 3002 15328 3036
rect 15384 3002 15418 3036
rect 15474 3002 15508 3036
rect 15564 3002 15598 3036
rect 15654 3002 15688 3036
rect 15744 3002 15778 3036
rect 15834 3002 15868 3036
rect 15924 3002 15958 3036
rect 16014 3002 16048 3036
rect 15202 2908 15236 2942
rect 15202 2818 15236 2852
rect 15202 2728 15236 2762
rect 15202 2638 15236 2672
rect 15202 2548 15236 2582
rect 15202 2458 15236 2492
rect 15202 2368 15236 2402
rect 15202 2278 15236 2312
rect 16092 2889 16126 2923
rect 16092 2799 16126 2833
rect 16092 2709 16126 2743
rect 16092 2619 16126 2653
rect 16092 2529 16126 2563
rect 16092 2439 16126 2473
rect 16092 2349 16126 2383
rect 16092 2259 16126 2293
rect 15202 2188 15236 2222
rect 16092 2169 16126 2203
rect 15260 2112 15294 2146
rect 15350 2112 15384 2146
rect 15440 2112 15474 2146
rect 15530 2112 15564 2146
rect 15620 2112 15654 2146
rect 15710 2112 15744 2146
rect 15800 2112 15834 2146
rect 15890 2112 15924 2146
rect 15980 2112 16014 2146
rect 16582 3002 16616 3036
rect 16672 3002 16706 3036
rect 16762 3002 16796 3036
rect 16852 3002 16886 3036
rect 16942 3002 16976 3036
rect 17032 3002 17066 3036
rect 17122 3002 17156 3036
rect 17212 3002 17246 3036
rect 17302 3002 17336 3036
rect 16490 2908 16524 2942
rect 16490 2818 16524 2852
rect 16490 2728 16524 2762
rect 16490 2638 16524 2672
rect 16490 2548 16524 2582
rect 16490 2458 16524 2492
rect 16490 2368 16524 2402
rect 16490 2278 16524 2312
rect 17380 2889 17414 2923
rect 17380 2799 17414 2833
rect 17380 2709 17414 2743
rect 17380 2619 17414 2653
rect 17380 2529 17414 2563
rect 17380 2439 17414 2473
rect 17380 2349 17414 2383
rect 17380 2259 17414 2293
rect 16490 2188 16524 2222
rect 17380 2169 17414 2203
rect 16548 2112 16582 2146
rect 16638 2112 16672 2146
rect 16728 2112 16762 2146
rect 16818 2112 16852 2146
rect 16908 2112 16942 2146
rect 16998 2112 17032 2146
rect 17088 2112 17122 2146
rect 17178 2112 17212 2146
rect 17268 2112 17302 2146
rect 17870 3002 17904 3036
rect 17960 3002 17994 3036
rect 18050 3002 18084 3036
rect 18140 3002 18174 3036
rect 18230 3002 18264 3036
rect 18320 3002 18354 3036
rect 18410 3002 18444 3036
rect 18500 3002 18534 3036
rect 18590 3002 18624 3036
rect 17778 2908 17812 2942
rect 17778 2818 17812 2852
rect 17778 2728 17812 2762
rect 17778 2638 17812 2672
rect 17778 2548 17812 2582
rect 17778 2458 17812 2492
rect 17778 2368 17812 2402
rect 17778 2278 17812 2312
rect 18668 2889 18702 2923
rect 18668 2799 18702 2833
rect 18668 2709 18702 2743
rect 18668 2619 18702 2653
rect 18668 2529 18702 2563
rect 18668 2439 18702 2473
rect 18668 2349 18702 2383
rect 18668 2259 18702 2293
rect 17778 2188 17812 2222
rect 18668 2169 18702 2203
rect 17836 2112 17870 2146
rect 17926 2112 17960 2146
rect 18016 2112 18050 2146
rect 18106 2112 18140 2146
rect 18196 2112 18230 2146
rect 18286 2112 18320 2146
rect 18376 2112 18410 2146
rect 18466 2112 18500 2146
rect 18556 2112 18590 2146
rect -15668 1196 -13326 1296
<< poly >>
rect -8754 9440 -8354 9466
rect -8296 9440 -7896 9466
rect -7838 9440 -7438 9466
rect -7380 9440 -6980 9466
rect -6922 9440 -6522 9466
rect -6464 9440 -6064 9466
rect -6006 9440 -5606 9466
rect -5548 9440 -5148 9466
rect -5090 9440 -4690 9466
rect -4632 9440 -4232 9466
rect -4174 9440 -3774 9466
rect -2796 9440 -2396 9466
rect -2338 9440 -1938 9466
rect -1880 9440 -1480 9466
rect -1422 9440 -1022 9466
rect -964 9440 -564 9466
rect -506 9440 -106 9466
rect -48 9440 352 9466
rect 410 9440 810 9466
rect 868 9440 1268 9466
rect 1326 9440 1726 9466
rect 2704 9440 3104 9466
rect 3162 9440 3562 9466
rect 3620 9440 4020 9466
rect 4078 9440 4478 9466
rect 4536 9440 4936 9466
rect 4994 9440 5394 9466
rect 5452 9440 5852 9466
rect 5910 9440 6310 9466
rect 6368 9440 6768 9466
rect 6826 9440 7226 9466
rect 7284 9440 7684 9466
rect -17264 8790 -17176 8806
rect -17264 8422 -17248 8790
rect -17214 8422 -17176 8790
rect -17264 8406 -17176 8422
rect -11776 8406 -11750 8806
rect -16836 6726 -16436 6742
rect -16836 6692 -16820 6726
rect -16452 6692 -16436 6726
rect -16836 6654 -16436 6692
rect -16264 6726 -15864 6742
rect -16264 6692 -16248 6726
rect -15880 6692 -15864 6726
rect -16264 6654 -15864 6692
rect -15692 6726 -15292 6742
rect -15692 6692 -15676 6726
rect -15308 6692 -15292 6726
rect -15692 6654 -15292 6692
rect -15120 6726 -14720 6742
rect -15120 6692 -15104 6726
rect -14736 6692 -14720 6726
rect -15120 6654 -14720 6692
rect -14548 6726 -14148 6742
rect -14548 6692 -14532 6726
rect -14164 6692 -14148 6726
rect -14548 6654 -14148 6692
rect -13976 6726 -13576 6742
rect -13976 6692 -13960 6726
rect -13592 6692 -13576 6726
rect -13976 6654 -13576 6692
rect -13404 6726 -13004 6742
rect -13404 6692 -13388 6726
rect -13020 6692 -13004 6726
rect -13404 6654 -13004 6692
rect -12832 6726 -12432 6742
rect -12832 6692 -12816 6726
rect -12448 6692 -12432 6726
rect -12832 6654 -12432 6692
rect -21766 5604 -21366 5620
rect -21766 5570 -21750 5604
rect -21382 5570 -21366 5604
rect -21766 5532 -21366 5570
rect -21308 5604 -20908 5620
rect -21308 5570 -21292 5604
rect -20924 5570 -20908 5604
rect -21308 5532 -20908 5570
rect -20850 5604 -20450 5620
rect -20850 5570 -20834 5604
rect -20466 5570 -20450 5604
rect -20850 5532 -20450 5570
rect -20392 5604 -19992 5620
rect -20392 5570 -20376 5604
rect -20008 5570 -19992 5604
rect -20392 5532 -19992 5570
rect -19934 5604 -19534 5620
rect -19934 5570 -19918 5604
rect -19550 5570 -19534 5604
rect -19934 5532 -19534 5570
rect -19476 5604 -19076 5620
rect -19476 5570 -19460 5604
rect -19092 5570 -19076 5604
rect -19476 5532 -19076 5570
rect -21766 5106 -21366 5132
rect -21308 5106 -20908 5132
rect -20850 5106 -20450 5132
rect -20392 5106 -19992 5132
rect -19934 5106 -19534 5132
rect -19476 5106 -19076 5132
rect -16836 4828 -16436 4854
rect -16264 4828 -15864 4854
rect -15692 4828 -15292 4854
rect -15120 4828 -14720 4854
rect -14548 4828 -14148 4854
rect -13976 4828 -13576 4854
rect -13404 4828 -13004 4854
rect -12832 4828 -12432 4854
rect -18562 4323 -18162 4339
rect -18562 4289 -18546 4323
rect -18178 4289 -18162 4323
rect -18562 4242 -18162 4289
rect -17990 4323 -17590 4339
rect -17990 4289 -17974 4323
rect -17606 4289 -17590 4323
rect -17990 4242 -17590 4289
rect -17418 4323 -17018 4339
rect -17418 4289 -17402 4323
rect -17034 4289 -17018 4323
rect -17418 4242 -17018 4289
rect -16846 4323 -16446 4339
rect -16846 4289 -16830 4323
rect -16462 4289 -16446 4323
rect -16846 4242 -16446 4289
rect -16274 4323 -15874 4339
rect -16274 4289 -16258 4323
rect -15890 4289 -15874 4323
rect -16274 4242 -15874 4289
rect -15702 4323 -15302 4339
rect -15702 4289 -15686 4323
rect -15318 4289 -15302 4323
rect -15702 4242 -15302 4289
rect -15130 4323 -14730 4339
rect -15130 4289 -15114 4323
rect -14746 4289 -14730 4323
rect -15130 4242 -14730 4289
rect -14558 4323 -14158 4339
rect -14558 4289 -14542 4323
rect -14174 4289 -14158 4323
rect -14558 4242 -14158 4289
rect -13986 4323 -13586 4339
rect -13986 4289 -13970 4323
rect -13602 4289 -13586 4323
rect -13986 4242 -13586 4289
rect -13414 4323 -13014 4339
rect -13414 4289 -13398 4323
rect -13030 4289 -13014 4323
rect -13414 4242 -13014 4289
rect -12842 4323 -12442 4339
rect -12842 4289 -12826 4323
rect -12458 4289 -12442 4323
rect -12842 4242 -12442 4289
rect -12270 4323 -11870 4339
rect -12270 4289 -12254 4323
rect -11886 4289 -11870 4323
rect -12270 4242 -11870 4289
rect -11698 4323 -11298 4339
rect -11698 4289 -11682 4323
rect -11314 4289 -11298 4323
rect -11698 4242 -11298 4289
rect -11126 4323 -10726 4339
rect -11126 4289 -11110 4323
rect -10742 4289 -10726 4323
rect -11126 4242 -10726 4289
rect -18562 1636 -18162 1662
rect -17990 1636 -17590 1662
rect -17418 1636 -17018 1662
rect -16846 1636 -16446 1662
rect -16274 1636 -15874 1662
rect -15702 1636 -15302 1662
rect -15130 1636 -14730 1662
rect -14558 1636 -14158 1662
rect -13986 1636 -13586 1662
rect -13414 1636 -13014 1662
rect -12842 1636 -12442 1662
rect -12270 1636 -11870 1662
rect -11698 1636 -11298 1662
rect -11126 1636 -10726 1662
rect -8754 1653 -8354 1700
rect -8754 1619 -8738 1653
rect -8370 1619 -8354 1653
rect -8754 1603 -8354 1619
rect -8296 1653 -7896 1700
rect -8296 1619 -8280 1653
rect -7912 1619 -7896 1653
rect -8296 1603 -7896 1619
rect -7838 1653 -7438 1700
rect -7838 1619 -7822 1653
rect -7454 1619 -7438 1653
rect -7838 1603 -7438 1619
rect -7380 1653 -6980 1700
rect -7380 1619 -7364 1653
rect -6996 1619 -6980 1653
rect -7380 1603 -6980 1619
rect -6922 1653 -6522 1700
rect -6922 1619 -6906 1653
rect -6538 1619 -6522 1653
rect -6922 1603 -6522 1619
rect -6464 1653 -6064 1700
rect -6464 1619 -6448 1653
rect -6080 1619 -6064 1653
rect -6464 1603 -6064 1619
rect -6006 1653 -5606 1700
rect -6006 1619 -5990 1653
rect -5622 1619 -5606 1653
rect -6006 1603 -5606 1619
rect -5548 1653 -5148 1700
rect -5548 1619 -5532 1653
rect -5164 1619 -5148 1653
rect -5548 1603 -5148 1619
rect -5090 1653 -4690 1700
rect -5090 1619 -5074 1653
rect -4706 1619 -4690 1653
rect -5090 1603 -4690 1619
rect -4632 1653 -4232 1700
rect -4632 1619 -4616 1653
rect -4248 1619 -4232 1653
rect -4632 1603 -4232 1619
rect -4174 1653 -3774 1700
rect -4174 1619 -4158 1653
rect -3790 1619 -3774 1653
rect -4174 1603 -3774 1619
rect -2796 1653 -2396 1700
rect -2796 1619 -2780 1653
rect -2412 1619 -2396 1653
rect -2796 1603 -2396 1619
rect -2338 1653 -1938 1700
rect -2338 1619 -2322 1653
rect -1954 1619 -1938 1653
rect -2338 1603 -1938 1619
rect -1880 1653 -1480 1700
rect -1880 1619 -1864 1653
rect -1496 1619 -1480 1653
rect -1880 1603 -1480 1619
rect -1422 1653 -1022 1700
rect -1422 1619 -1406 1653
rect -1038 1619 -1022 1653
rect -1422 1603 -1022 1619
rect -964 1653 -564 1700
rect -964 1619 -948 1653
rect -580 1619 -564 1653
rect -964 1603 -564 1619
rect -506 1653 -106 1700
rect -506 1619 -490 1653
rect -122 1619 -106 1653
rect -506 1603 -106 1619
rect -48 1653 352 1700
rect -48 1619 -32 1653
rect 336 1619 352 1653
rect -48 1603 352 1619
rect 410 1653 810 1700
rect 410 1619 426 1653
rect 794 1619 810 1653
rect 410 1603 810 1619
rect 868 1653 1268 1700
rect 868 1619 884 1653
rect 1252 1619 1268 1653
rect 868 1603 1268 1619
rect 1326 1653 1726 1700
rect 1326 1619 1342 1653
rect 1710 1619 1726 1653
rect 1326 1603 1726 1619
rect 2704 1653 3104 1700
rect 2704 1619 2720 1653
rect 3088 1619 3104 1653
rect 2704 1603 3104 1619
rect 3162 1653 3562 1700
rect 3162 1619 3178 1653
rect 3546 1619 3562 1653
rect 3162 1603 3562 1619
rect 3620 1653 4020 1700
rect 3620 1619 3636 1653
rect 4004 1619 4020 1653
rect 3620 1603 4020 1619
rect 4078 1653 4478 1700
rect 4078 1619 4094 1653
rect 4462 1619 4478 1653
rect 4078 1603 4478 1619
rect 4536 1653 4936 1700
rect 4536 1619 4552 1653
rect 4920 1619 4936 1653
rect 4536 1603 4936 1619
rect 4994 1653 5394 1700
rect 4994 1619 5010 1653
rect 5378 1619 5394 1653
rect 4994 1603 5394 1619
rect 5452 1653 5852 1700
rect 5452 1619 5468 1653
rect 5836 1619 5852 1653
rect 5452 1603 5852 1619
rect 5910 1653 6310 1700
rect 5910 1619 5926 1653
rect 6294 1619 6310 1653
rect 5910 1603 6310 1619
rect 6368 1653 6768 1700
rect 6368 1619 6384 1653
rect 6752 1619 6768 1653
rect 6368 1603 6768 1619
rect 6826 1653 7226 1700
rect 6826 1619 6842 1653
rect 7210 1619 7226 1653
rect 6826 1603 7226 1619
rect 7284 1653 7684 1700
rect 7284 1619 7300 1653
rect 7668 1619 7684 1653
rect 7284 1603 7684 1619
<< polycont >>
rect -17248 8422 -17214 8790
rect -16820 6692 -16452 6726
rect -16248 6692 -15880 6726
rect -15676 6692 -15308 6726
rect -15104 6692 -14736 6726
rect -14532 6692 -14164 6726
rect -13960 6692 -13592 6726
rect -13388 6692 -13020 6726
rect -12816 6692 -12448 6726
rect -21750 5570 -21382 5604
rect -21292 5570 -20924 5604
rect -20834 5570 -20466 5604
rect -20376 5570 -20008 5604
rect -19918 5570 -19550 5604
rect -19460 5570 -19092 5604
rect -18546 4289 -18178 4323
rect -17974 4289 -17606 4323
rect -17402 4289 -17034 4323
rect -16830 4289 -16462 4323
rect -16258 4289 -15890 4323
rect -15686 4289 -15318 4323
rect -15114 4289 -14746 4323
rect -14542 4289 -14174 4323
rect -13970 4289 -13602 4323
rect -13398 4289 -13030 4323
rect -12826 4289 -12458 4323
rect -12254 4289 -11886 4323
rect -11682 4289 -11314 4323
rect -11110 4289 -10742 4323
rect -8738 1619 -8370 1653
rect -8280 1619 -7912 1653
rect -7822 1619 -7454 1653
rect -7364 1619 -6996 1653
rect -6906 1619 -6538 1653
rect -6448 1619 -6080 1653
rect -5990 1619 -5622 1653
rect -5532 1619 -5164 1653
rect -5074 1619 -4706 1653
rect -4616 1619 -4248 1653
rect -4158 1619 -3790 1653
rect -2780 1619 -2412 1653
rect -2322 1619 -1954 1653
rect -1864 1619 -1496 1653
rect -1406 1619 -1038 1653
rect -948 1619 -580 1653
rect -490 1619 -122 1653
rect -32 1619 336 1653
rect 426 1619 794 1653
rect 884 1619 1252 1653
rect 1342 1619 1710 1653
rect 2720 1619 3088 1653
rect 3178 1619 3546 1653
rect 3636 1619 4004 1653
rect 4094 1619 4462 1653
rect 4552 1619 4920 1653
rect 5010 1619 5378 1653
rect 5468 1619 5836 1653
rect 5926 1619 6294 1653
rect 6384 1619 6752 1653
rect 6842 1619 7210 1653
rect 7300 1619 7668 1653
<< xpolycontact >>
rect -5660 21562 -5090 21994
rect -8932 20176 -8362 20608
rect -8932 16420 -8362 16852
rect -8114 20176 -7544 20608
rect -8114 16420 -7544 16852
rect -7296 20176 -6726 20608
rect -7296 16420 -6726 16852
rect -5660 16830 -5090 17262
rect -4842 21562 -4272 21994
rect -4842 16830 -4272 17262
rect -4024 21562 -3454 21994
rect -4024 16830 -3454 17262
rect -3206 21562 -2636 21994
rect -3206 16830 -2636 17262
rect -752 21500 -182 21932
rect -752 14764 -182 15196
rect 66 21500 636 21932
rect 66 14764 636 15196
rect 884 21500 1454 21932
rect 884 14764 1454 15196
rect 1702 21500 2272 21932
rect 1702 14764 2272 15196
rect 2520 21500 3090 21932
rect 2520 14764 3090 15196
rect 3338 21500 3908 21932
rect 3338 14764 3908 15196
rect 4156 21500 4726 21932
rect 4156 14764 4726 15196
rect 4974 21500 5544 21932
rect 4974 14764 5544 15196
rect 5792 21500 6362 21932
rect 5792 14764 6362 15196
rect 6610 21500 7180 21932
rect 6610 14764 7180 15196
rect 7428 21500 7998 21932
rect 7428 14764 7998 15196
rect 8246 21500 8816 21932
rect 8246 14764 8816 15196
rect 9064 21500 9634 21932
rect 9064 14764 9634 15196
rect 9882 21500 10452 21932
rect 9882 14764 10452 15196
rect 10700 21500 11270 21932
rect 10700 14764 11270 15196
rect 11518 21500 12088 21932
rect 11518 14764 12088 15196
rect 12336 21500 12906 21932
rect 12336 14764 12906 15196
<< xpolyres >>
rect -8932 16852 -8362 20176
rect -8114 16852 -7544 20176
rect -7296 16852 -6726 20176
rect -5660 17262 -5090 21562
rect -4842 17262 -4272 21562
rect -4024 17262 -3454 21562
rect -3206 17262 -2636 21562
rect -752 15196 -182 21500
rect 66 15196 636 21500
rect 884 15196 1454 21500
rect 1702 15196 2272 21500
rect 2520 15196 3090 21500
rect 3338 15196 3908 21500
rect 4156 15196 4726 21500
rect 4974 15196 5544 21500
rect 5792 15196 6362 21500
rect 6610 15196 7180 21500
rect 7428 15196 7998 21500
rect 8246 15196 8816 21500
rect 9064 15196 9634 21500
rect 9882 15196 10452 21500
rect 10700 15196 11270 21500
rect 11518 15196 12088 21500
rect 12336 15196 12906 21500
<< locali >>
rect -6534 21562 -5660 21994
rect -2636 21932 -1236 21994
rect -2636 21562 -752 21932
rect -6534 21516 -5930 21562
rect -3206 21558 -752 21562
rect -9772 21500 -9170 21516
rect -9772 20608 -9756 21500
rect -9782 20166 -9756 20608
rect -9772 16106 -9756 20166
rect -9776 15602 -9756 16106
rect -9772 15196 -9756 15602
rect -9186 20608 -9170 21500
rect -6534 21500 -5926 21516
rect -1576 21500 -752 21558
rect 12906 21500 13730 21932
rect -6534 21004 -6512 21500
rect -6528 20608 -6512 21004
rect -9186 20176 -8932 20608
rect -8362 20176 -8114 20608
rect -7544 20176 -7296 20608
rect -6726 20176 -6512 20608
rect -9186 20166 -6512 20176
rect -9186 16106 -9170 20166
rect -6528 16852 -6512 20166
rect -6726 16420 -6512 16852
rect -8932 16110 -8362 16420
rect -6528 16110 -6512 16420
rect -8932 16106 -8104 16110
rect -9186 15602 -8104 16106
rect -7556 15602 -6512 16110
rect -9186 15196 -9170 15602
rect -9772 15180 -9170 15196
rect -6528 15196 -6512 15602
rect -5942 17258 -5926 21500
rect -1568 17262 -1552 21500
rect -5942 16830 -5660 17258
rect -5090 16830 -4842 17262
rect -4272 16830 -4024 17262
rect -3454 16830 -3206 17262
rect -2636 16830 -1552 17262
rect -5942 16732 -1552 16830
rect -5942 16110 -5926 16732
rect -5942 15602 -5916 16110
rect -5942 15196 -5926 15602
rect -1568 15196 -1552 16732
rect -982 15196 -966 21500
rect 13120 15196 13136 21500
rect 13706 15196 13722 21500
rect -6528 15180 -5926 15196
rect -1576 14764 -752 15196
rect 12906 14764 13730 15196
rect 12444 12202 18884 12234
rect 12444 12168 12578 12202
rect 12612 12168 12668 12202
rect 12702 12168 12758 12202
rect 12792 12168 12848 12202
rect 12882 12168 12938 12202
rect 12972 12168 13028 12202
rect 13062 12168 13118 12202
rect 13152 12168 13208 12202
rect 13242 12168 13298 12202
rect 13332 12168 13388 12202
rect 13422 12168 13478 12202
rect 13512 12168 13568 12202
rect 13602 12168 13866 12202
rect 13900 12168 13956 12202
rect 13990 12168 14046 12202
rect 14080 12168 14136 12202
rect 14170 12168 14226 12202
rect 14260 12168 14316 12202
rect 14350 12168 14406 12202
rect 14440 12168 14496 12202
rect 14530 12168 14586 12202
rect 14620 12168 14676 12202
rect 14710 12168 14766 12202
rect 14800 12168 14856 12202
rect 14890 12168 15154 12202
rect 15188 12168 15244 12202
rect 15278 12168 15334 12202
rect 15368 12168 15424 12202
rect 15458 12168 15514 12202
rect 15548 12168 15604 12202
rect 15638 12168 15694 12202
rect 15728 12168 15784 12202
rect 15818 12168 15874 12202
rect 15908 12168 15964 12202
rect 15998 12168 16054 12202
rect 16088 12168 16144 12202
rect 16178 12168 16442 12202
rect 16476 12168 16532 12202
rect 16566 12168 16622 12202
rect 16656 12168 16712 12202
rect 16746 12168 16802 12202
rect 16836 12168 16892 12202
rect 16926 12168 16982 12202
rect 17016 12168 17072 12202
rect 17106 12168 17162 12202
rect 17196 12168 17252 12202
rect 17286 12168 17342 12202
rect 17376 12168 17432 12202
rect 17466 12168 17730 12202
rect 17764 12168 17820 12202
rect 17854 12168 17910 12202
rect 17944 12168 18000 12202
rect 18034 12168 18090 12202
rect 18124 12168 18180 12202
rect 18214 12168 18270 12202
rect 18304 12168 18360 12202
rect 18394 12168 18450 12202
rect 18484 12168 18540 12202
rect 18574 12168 18630 12202
rect 18664 12168 18720 12202
rect 18754 12168 18884 12202
rect 12444 12135 18884 12168
rect 12444 12118 12684 12135
rect 12444 12084 12477 12118
rect 12511 12084 12684 12118
rect 12444 12071 12684 12084
rect 13484 12118 13984 12135
rect 13484 12084 13664 12118
rect 13698 12084 13765 12118
rect 13799 12084 13984 12118
rect 13484 12071 13984 12084
rect 14784 12118 15184 12135
rect 14784 12084 14952 12118
rect 14986 12084 15053 12118
rect 15087 12084 15184 12118
rect 14784 12071 15184 12084
rect 16084 12118 16484 12135
rect 16084 12084 16240 12118
rect 16274 12084 16341 12118
rect 16375 12084 16484 12118
rect 16084 12071 16484 12084
rect 17384 12118 17784 12135
rect 17384 12084 17528 12118
rect 17562 12084 17629 12118
rect 17663 12084 17784 12118
rect 17384 12071 17784 12084
rect 18684 12118 18884 12135
rect 18684 12084 18816 12118
rect 18850 12084 18884 12118
rect 18684 12071 18884 12084
rect 12444 12052 18884 12071
rect 12444 12028 12718 12052
rect 12444 11994 12477 12028
rect 12511 12018 12718 12028
rect 12752 12018 12808 12052
rect 12842 12018 12898 12052
rect 12932 12018 12988 12052
rect 13022 12018 13078 12052
rect 13112 12018 13168 12052
rect 13202 12018 13258 12052
rect 13292 12018 13348 12052
rect 13382 12018 13438 12052
rect 13472 12028 14006 12052
rect 13472 12018 13664 12028
rect 12511 11999 13664 12018
rect 12511 11994 12684 11999
rect 12444 11958 12684 11994
rect 12444 11938 12626 11958
rect 12444 11904 12477 11938
rect 12511 11924 12626 11938
rect 12660 11924 12684 11958
rect 13484 11994 13664 11999
rect 13698 11994 13765 12028
rect 13799 12018 14006 12028
rect 14040 12018 14096 12052
rect 14130 12018 14186 12052
rect 14220 12018 14276 12052
rect 14310 12018 14366 12052
rect 14400 12018 14456 12052
rect 14490 12018 14546 12052
rect 14580 12018 14636 12052
rect 14670 12018 14726 12052
rect 14760 12028 15294 12052
rect 14760 12018 14952 12028
rect 13799 11999 14952 12018
rect 13799 11994 13984 11999
rect 13484 11958 13984 11994
rect 13484 11939 13914 11958
rect 12511 11904 12684 11924
rect 12444 11868 12684 11904
rect 12444 11848 12626 11868
rect 12444 11814 12477 11848
rect 12511 11834 12626 11848
rect 12660 11834 12684 11868
rect 12511 11814 12684 11834
rect 12444 11778 12684 11814
rect 12444 11758 12626 11778
rect 12444 11724 12477 11758
rect 12511 11744 12626 11758
rect 12660 11744 12684 11778
rect 12511 11724 12684 11744
rect 12444 11688 12684 11724
rect 12444 11668 12626 11688
rect 12444 11634 12477 11668
rect 12511 11654 12626 11668
rect 12660 11654 12684 11688
rect 12511 11634 12684 11654
rect 12444 11598 12684 11634
rect 12444 11578 12626 11598
rect 12444 11544 12477 11578
rect 12511 11564 12626 11578
rect 12660 11564 12684 11598
rect 12511 11544 12684 11564
rect 12444 11508 12684 11544
rect 12444 11488 12626 11508
rect 12444 11454 12477 11488
rect 12511 11474 12626 11488
rect 12660 11474 12684 11508
rect 12511 11454 12684 11474
rect 12444 11418 12684 11454
rect 12444 11398 12626 11418
rect 12444 11364 12477 11398
rect 12511 11384 12626 11398
rect 12660 11384 12684 11418
rect 12511 11364 12684 11384
rect 12444 11328 12684 11364
rect 12444 11308 12626 11328
rect 12444 11274 12477 11308
rect 12511 11294 12626 11308
rect 12660 11294 12684 11328
rect 12511 11274 12684 11294
rect 12444 11238 12684 11274
rect 12741 11876 13435 11937
rect 12741 11842 12800 11876
rect 12834 11864 12890 11876
rect 12862 11842 12890 11864
rect 12924 11864 12980 11876
rect 12924 11842 12928 11864
rect 12741 11830 12828 11842
rect 12862 11830 12928 11842
rect 12962 11842 12980 11864
rect 13014 11864 13070 11876
rect 13014 11842 13028 11864
rect 12962 11830 13028 11842
rect 13062 11842 13070 11864
rect 13104 11864 13160 11876
rect 13194 11864 13250 11876
rect 13284 11864 13340 11876
rect 13104 11842 13128 11864
rect 13194 11842 13228 11864
rect 13284 11842 13328 11864
rect 13374 11842 13435 11876
rect 13062 11830 13128 11842
rect 13162 11830 13228 11842
rect 13262 11830 13328 11842
rect 13362 11830 13435 11842
rect 12741 11786 13435 11830
rect 12741 11752 12800 11786
rect 12834 11764 12890 11786
rect 12862 11752 12890 11764
rect 12924 11764 12980 11786
rect 12924 11752 12928 11764
rect 12741 11730 12828 11752
rect 12862 11730 12928 11752
rect 12962 11752 12980 11764
rect 13014 11764 13070 11786
rect 13014 11752 13028 11764
rect 12962 11730 13028 11752
rect 13062 11752 13070 11764
rect 13104 11764 13160 11786
rect 13194 11764 13250 11786
rect 13284 11764 13340 11786
rect 13104 11752 13128 11764
rect 13194 11752 13228 11764
rect 13284 11752 13328 11764
rect 13374 11752 13435 11786
rect 13062 11730 13128 11752
rect 13162 11730 13228 11752
rect 13262 11730 13328 11752
rect 13362 11730 13435 11752
rect 12741 11696 13435 11730
rect 12741 11662 12800 11696
rect 12834 11664 12890 11696
rect 12862 11662 12890 11664
rect 12924 11664 12980 11696
rect 12924 11662 12928 11664
rect 12741 11630 12828 11662
rect 12862 11630 12928 11662
rect 12962 11662 12980 11664
rect 13014 11664 13070 11696
rect 13014 11662 13028 11664
rect 12962 11630 13028 11662
rect 13062 11662 13070 11664
rect 13104 11664 13160 11696
rect 13194 11664 13250 11696
rect 13284 11664 13340 11696
rect 13104 11662 13128 11664
rect 13194 11662 13228 11664
rect 13284 11662 13328 11664
rect 13374 11662 13435 11696
rect 13062 11630 13128 11662
rect 13162 11630 13228 11662
rect 13262 11630 13328 11662
rect 13362 11630 13435 11662
rect 12741 11606 13435 11630
rect 12741 11572 12800 11606
rect 12834 11572 12890 11606
rect 12924 11572 12980 11606
rect 13014 11572 13070 11606
rect 13104 11572 13160 11606
rect 13194 11572 13250 11606
rect 13284 11572 13340 11606
rect 13374 11572 13435 11606
rect 12741 11564 13435 11572
rect 12741 11530 12828 11564
rect 12862 11530 12928 11564
rect 12962 11530 13028 11564
rect 13062 11530 13128 11564
rect 13162 11530 13228 11564
rect 13262 11530 13328 11564
rect 13362 11530 13435 11564
rect 12741 11516 13435 11530
rect 12741 11482 12800 11516
rect 12834 11482 12890 11516
rect 12924 11482 12980 11516
rect 13014 11482 13070 11516
rect 13104 11482 13160 11516
rect 13194 11482 13250 11516
rect 13284 11482 13340 11516
rect 13374 11482 13435 11516
rect 12741 11464 13435 11482
rect 12741 11430 12828 11464
rect 12862 11430 12928 11464
rect 12962 11430 13028 11464
rect 13062 11430 13128 11464
rect 13162 11430 13228 11464
rect 13262 11430 13328 11464
rect 13362 11430 13435 11464
rect 12741 11426 13435 11430
rect 12741 11392 12800 11426
rect 12834 11392 12890 11426
rect 12924 11392 12980 11426
rect 13014 11392 13070 11426
rect 13104 11392 13160 11426
rect 13194 11392 13250 11426
rect 13284 11392 13340 11426
rect 13374 11392 13435 11426
rect 12741 11364 13435 11392
rect 12741 11336 12828 11364
rect 12862 11336 12928 11364
rect 12741 11302 12800 11336
rect 12862 11330 12890 11336
rect 12834 11302 12890 11330
rect 12924 11330 12928 11336
rect 12962 11336 13028 11364
rect 12962 11330 12980 11336
rect 12924 11302 12980 11330
rect 13014 11330 13028 11336
rect 13062 11336 13128 11364
rect 13162 11336 13228 11364
rect 13262 11336 13328 11364
rect 13362 11336 13435 11364
rect 13062 11330 13070 11336
rect 13014 11302 13070 11330
rect 13104 11330 13128 11336
rect 13194 11330 13228 11336
rect 13284 11330 13328 11336
rect 13104 11302 13160 11330
rect 13194 11302 13250 11330
rect 13284 11302 13340 11330
rect 13374 11302 13435 11336
rect 12741 11243 13435 11302
rect 13484 11905 13516 11939
rect 13550 11938 13914 11939
rect 13550 11905 13664 11938
rect 13484 11904 13664 11905
rect 13698 11904 13765 11938
rect 13799 11924 13914 11938
rect 13948 11924 13984 11958
rect 14784 11994 14952 11999
rect 14986 11994 15053 12028
rect 15087 12018 15294 12028
rect 15328 12018 15384 12052
rect 15418 12018 15474 12052
rect 15508 12018 15564 12052
rect 15598 12018 15654 12052
rect 15688 12018 15744 12052
rect 15778 12018 15834 12052
rect 15868 12018 15924 12052
rect 15958 12018 16014 12052
rect 16048 12028 16582 12052
rect 16048 12018 16240 12028
rect 15087 11999 16240 12018
rect 15087 11994 15255 11999
rect 14784 11958 15255 11994
rect 14784 11939 15202 11958
rect 13799 11904 13984 11924
rect 13484 11868 13984 11904
rect 13484 11849 13914 11868
rect 13484 11815 13516 11849
rect 13550 11848 13914 11849
rect 13550 11815 13664 11848
rect 13484 11814 13664 11815
rect 13698 11814 13765 11848
rect 13799 11834 13914 11848
rect 13948 11834 13984 11868
rect 13799 11814 13984 11834
rect 13484 11778 13984 11814
rect 13484 11759 13914 11778
rect 13484 11725 13516 11759
rect 13550 11758 13914 11759
rect 13550 11725 13664 11758
rect 13484 11724 13664 11725
rect 13698 11724 13765 11758
rect 13799 11744 13914 11758
rect 13948 11744 13984 11778
rect 13799 11724 13984 11744
rect 13484 11688 13984 11724
rect 13484 11669 13914 11688
rect 13484 11635 13516 11669
rect 13550 11668 13914 11669
rect 13550 11635 13664 11668
rect 13484 11634 13664 11635
rect 13698 11634 13765 11668
rect 13799 11654 13914 11668
rect 13948 11654 13984 11688
rect 13799 11634 13984 11654
rect 13484 11598 13984 11634
rect 13484 11579 13914 11598
rect 13484 11545 13516 11579
rect 13550 11578 13914 11579
rect 13550 11545 13664 11578
rect 13484 11544 13664 11545
rect 13698 11544 13765 11578
rect 13799 11564 13914 11578
rect 13948 11564 13984 11598
rect 13799 11544 13984 11564
rect 13484 11508 13984 11544
rect 13484 11489 13914 11508
rect 13484 11455 13516 11489
rect 13550 11488 13914 11489
rect 13550 11455 13664 11488
rect 13484 11454 13664 11455
rect 13698 11454 13765 11488
rect 13799 11474 13914 11488
rect 13948 11474 13984 11508
rect 13799 11454 13984 11474
rect 13484 11418 13984 11454
rect 13484 11399 13914 11418
rect 13484 11365 13516 11399
rect 13550 11398 13914 11399
rect 13550 11365 13664 11398
rect 13484 11364 13664 11365
rect 13698 11364 13765 11398
rect 13799 11384 13914 11398
rect 13948 11384 13984 11418
rect 13799 11364 13984 11384
rect 13484 11328 13984 11364
rect 13484 11309 13914 11328
rect 13484 11275 13516 11309
rect 13550 11308 13914 11309
rect 13550 11275 13664 11308
rect 13484 11274 13664 11275
rect 13698 11274 13765 11308
rect 13799 11294 13914 11308
rect 13948 11294 13984 11328
rect 13799 11274 13984 11294
rect 12444 11218 12626 11238
rect 12444 11184 12477 11218
rect 12511 11204 12626 11218
rect 12660 11204 12684 11238
rect 12511 11184 12684 11204
rect 12444 11181 12684 11184
rect 13484 11238 13984 11274
rect 14029 11876 14723 11937
rect 14029 11842 14088 11876
rect 14122 11864 14178 11876
rect 14150 11842 14178 11864
rect 14212 11864 14268 11876
rect 14212 11842 14216 11864
rect 14029 11830 14116 11842
rect 14150 11830 14216 11842
rect 14250 11842 14268 11864
rect 14302 11864 14358 11876
rect 14302 11842 14316 11864
rect 14250 11830 14316 11842
rect 14350 11842 14358 11864
rect 14392 11864 14448 11876
rect 14482 11864 14538 11876
rect 14572 11864 14628 11876
rect 14392 11842 14416 11864
rect 14482 11842 14516 11864
rect 14572 11842 14616 11864
rect 14662 11842 14723 11876
rect 14350 11830 14416 11842
rect 14450 11830 14516 11842
rect 14550 11830 14616 11842
rect 14650 11830 14723 11842
rect 14029 11786 14723 11830
rect 14029 11752 14088 11786
rect 14122 11764 14178 11786
rect 14150 11752 14178 11764
rect 14212 11764 14268 11786
rect 14212 11752 14216 11764
rect 14029 11730 14116 11752
rect 14150 11730 14216 11752
rect 14250 11752 14268 11764
rect 14302 11764 14358 11786
rect 14302 11752 14316 11764
rect 14250 11730 14316 11752
rect 14350 11752 14358 11764
rect 14392 11764 14448 11786
rect 14482 11764 14538 11786
rect 14572 11764 14628 11786
rect 14392 11752 14416 11764
rect 14482 11752 14516 11764
rect 14572 11752 14616 11764
rect 14662 11752 14723 11786
rect 14350 11730 14416 11752
rect 14450 11730 14516 11752
rect 14550 11730 14616 11752
rect 14650 11730 14723 11752
rect 14029 11696 14723 11730
rect 14029 11662 14088 11696
rect 14122 11664 14178 11696
rect 14150 11662 14178 11664
rect 14212 11664 14268 11696
rect 14212 11662 14216 11664
rect 14029 11630 14116 11662
rect 14150 11630 14216 11662
rect 14250 11662 14268 11664
rect 14302 11664 14358 11696
rect 14302 11662 14316 11664
rect 14250 11630 14316 11662
rect 14350 11662 14358 11664
rect 14392 11664 14448 11696
rect 14482 11664 14538 11696
rect 14572 11664 14628 11696
rect 14392 11662 14416 11664
rect 14482 11662 14516 11664
rect 14572 11662 14616 11664
rect 14662 11662 14723 11696
rect 14350 11630 14416 11662
rect 14450 11630 14516 11662
rect 14550 11630 14616 11662
rect 14650 11630 14723 11662
rect 14029 11606 14723 11630
rect 14029 11572 14088 11606
rect 14122 11572 14178 11606
rect 14212 11572 14268 11606
rect 14302 11572 14358 11606
rect 14392 11572 14448 11606
rect 14482 11572 14538 11606
rect 14572 11572 14628 11606
rect 14662 11572 14723 11606
rect 14029 11564 14723 11572
rect 14029 11530 14116 11564
rect 14150 11530 14216 11564
rect 14250 11530 14316 11564
rect 14350 11530 14416 11564
rect 14450 11530 14516 11564
rect 14550 11530 14616 11564
rect 14650 11530 14723 11564
rect 14029 11516 14723 11530
rect 14029 11482 14088 11516
rect 14122 11482 14178 11516
rect 14212 11482 14268 11516
rect 14302 11482 14358 11516
rect 14392 11482 14448 11516
rect 14482 11482 14538 11516
rect 14572 11482 14628 11516
rect 14662 11482 14723 11516
rect 14029 11464 14723 11482
rect 14029 11430 14116 11464
rect 14150 11430 14216 11464
rect 14250 11430 14316 11464
rect 14350 11430 14416 11464
rect 14450 11430 14516 11464
rect 14550 11430 14616 11464
rect 14650 11430 14723 11464
rect 14029 11426 14723 11430
rect 14029 11392 14088 11426
rect 14122 11392 14178 11426
rect 14212 11392 14268 11426
rect 14302 11392 14358 11426
rect 14392 11392 14448 11426
rect 14482 11392 14538 11426
rect 14572 11392 14628 11426
rect 14662 11392 14723 11426
rect 14029 11364 14723 11392
rect 14029 11336 14116 11364
rect 14150 11336 14216 11364
rect 14029 11302 14088 11336
rect 14150 11330 14178 11336
rect 14122 11302 14178 11330
rect 14212 11330 14216 11336
rect 14250 11336 14316 11364
rect 14250 11330 14268 11336
rect 14212 11302 14268 11330
rect 14302 11330 14316 11336
rect 14350 11336 14416 11364
rect 14450 11336 14516 11364
rect 14550 11336 14616 11364
rect 14650 11336 14723 11364
rect 14350 11330 14358 11336
rect 14302 11302 14358 11330
rect 14392 11330 14416 11336
rect 14482 11330 14516 11336
rect 14572 11330 14616 11336
rect 14392 11302 14448 11330
rect 14482 11302 14538 11330
rect 14572 11302 14628 11330
rect 14662 11302 14723 11336
rect 14029 11243 14723 11302
rect 14784 11905 14804 11939
rect 14838 11938 15202 11939
rect 14838 11905 14952 11938
rect 14784 11904 14952 11905
rect 14986 11904 15053 11938
rect 15087 11924 15202 11938
rect 15236 11924 15255 11958
rect 16073 11994 16240 11999
rect 16274 11994 16341 12028
rect 16375 12018 16582 12028
rect 16616 12018 16672 12052
rect 16706 12018 16762 12052
rect 16796 12018 16852 12052
rect 16886 12018 16942 12052
rect 16976 12018 17032 12052
rect 17066 12018 17122 12052
rect 17156 12018 17212 12052
rect 17246 12018 17302 12052
rect 17336 12028 17870 12052
rect 17336 12018 17528 12028
rect 16375 11999 17528 12018
rect 16375 11994 16543 11999
rect 16073 11958 16543 11994
rect 16073 11939 16490 11958
rect 15087 11904 15255 11924
rect 14784 11868 15255 11904
rect 14784 11849 15202 11868
rect 14784 11815 14804 11849
rect 14838 11848 15202 11849
rect 14838 11815 14952 11848
rect 14784 11814 14952 11815
rect 14986 11814 15053 11848
rect 15087 11834 15202 11848
rect 15236 11834 15255 11868
rect 15087 11814 15255 11834
rect 14784 11778 15255 11814
rect 14784 11759 15202 11778
rect 14784 11725 14804 11759
rect 14838 11758 15202 11759
rect 14838 11725 14952 11758
rect 14784 11724 14952 11725
rect 14986 11724 15053 11758
rect 15087 11744 15202 11758
rect 15236 11744 15255 11778
rect 15087 11724 15255 11744
rect 14784 11688 15255 11724
rect 14784 11669 15202 11688
rect 14784 11635 14804 11669
rect 14838 11668 15202 11669
rect 14838 11635 14952 11668
rect 14784 11634 14952 11635
rect 14986 11634 15053 11668
rect 15087 11654 15202 11668
rect 15236 11654 15255 11688
rect 15087 11634 15255 11654
rect 14784 11598 15255 11634
rect 14784 11579 15202 11598
rect 14784 11545 14804 11579
rect 14838 11578 15202 11579
rect 14838 11545 14952 11578
rect 14784 11544 14952 11545
rect 14986 11544 15053 11578
rect 15087 11564 15202 11578
rect 15236 11564 15255 11598
rect 15087 11544 15255 11564
rect 14784 11508 15255 11544
rect 14784 11489 15202 11508
rect 14784 11455 14804 11489
rect 14838 11488 15202 11489
rect 14838 11455 14952 11488
rect 14784 11454 14952 11455
rect 14986 11454 15053 11488
rect 15087 11474 15202 11488
rect 15236 11474 15255 11508
rect 15087 11454 15255 11474
rect 14784 11418 15255 11454
rect 14784 11399 15202 11418
rect 14784 11365 14804 11399
rect 14838 11398 15202 11399
rect 14838 11365 14952 11398
rect 14784 11364 14952 11365
rect 14986 11364 15053 11398
rect 15087 11384 15202 11398
rect 15236 11384 15255 11418
rect 15087 11364 15255 11384
rect 14784 11328 15255 11364
rect 14784 11309 15202 11328
rect 14784 11275 14804 11309
rect 14838 11308 15202 11309
rect 14838 11275 14952 11308
rect 14784 11274 14952 11275
rect 14986 11274 15053 11308
rect 15087 11294 15202 11308
rect 15236 11294 15255 11328
rect 15087 11274 15255 11294
rect 13484 11219 13914 11238
rect 13484 11185 13516 11219
rect 13550 11218 13914 11219
rect 13550 11185 13664 11218
rect 13484 11184 13664 11185
rect 13698 11184 13765 11218
rect 13799 11204 13914 11218
rect 13948 11204 13984 11238
rect 13799 11184 13984 11204
rect 13484 11181 13984 11184
rect 14784 11238 15255 11274
rect 15317 11876 16011 11937
rect 15317 11842 15376 11876
rect 15410 11864 15466 11876
rect 15438 11842 15466 11864
rect 15500 11864 15556 11876
rect 15500 11842 15504 11864
rect 15317 11830 15404 11842
rect 15438 11830 15504 11842
rect 15538 11842 15556 11864
rect 15590 11864 15646 11876
rect 15590 11842 15604 11864
rect 15538 11830 15604 11842
rect 15638 11842 15646 11864
rect 15680 11864 15736 11876
rect 15770 11864 15826 11876
rect 15860 11864 15916 11876
rect 15680 11842 15704 11864
rect 15770 11842 15804 11864
rect 15860 11842 15904 11864
rect 15950 11842 16011 11876
rect 15638 11830 15704 11842
rect 15738 11830 15804 11842
rect 15838 11830 15904 11842
rect 15938 11830 16011 11842
rect 15317 11786 16011 11830
rect 15317 11752 15376 11786
rect 15410 11764 15466 11786
rect 15438 11752 15466 11764
rect 15500 11764 15556 11786
rect 15500 11752 15504 11764
rect 15317 11730 15404 11752
rect 15438 11730 15504 11752
rect 15538 11752 15556 11764
rect 15590 11764 15646 11786
rect 15590 11752 15604 11764
rect 15538 11730 15604 11752
rect 15638 11752 15646 11764
rect 15680 11764 15736 11786
rect 15770 11764 15826 11786
rect 15860 11764 15916 11786
rect 15680 11752 15704 11764
rect 15770 11752 15804 11764
rect 15860 11752 15904 11764
rect 15950 11752 16011 11786
rect 15638 11730 15704 11752
rect 15738 11730 15804 11752
rect 15838 11730 15904 11752
rect 15938 11730 16011 11752
rect 15317 11696 16011 11730
rect 15317 11662 15376 11696
rect 15410 11664 15466 11696
rect 15438 11662 15466 11664
rect 15500 11664 15556 11696
rect 15500 11662 15504 11664
rect 15317 11630 15404 11662
rect 15438 11630 15504 11662
rect 15538 11662 15556 11664
rect 15590 11664 15646 11696
rect 15590 11662 15604 11664
rect 15538 11630 15604 11662
rect 15638 11662 15646 11664
rect 15680 11664 15736 11696
rect 15770 11664 15826 11696
rect 15860 11664 15916 11696
rect 15680 11662 15704 11664
rect 15770 11662 15804 11664
rect 15860 11662 15904 11664
rect 15950 11662 16011 11696
rect 15638 11630 15704 11662
rect 15738 11630 15804 11662
rect 15838 11630 15904 11662
rect 15938 11630 16011 11662
rect 15317 11606 16011 11630
rect 15317 11572 15376 11606
rect 15410 11572 15466 11606
rect 15500 11572 15556 11606
rect 15590 11572 15646 11606
rect 15680 11572 15736 11606
rect 15770 11572 15826 11606
rect 15860 11572 15916 11606
rect 15950 11572 16011 11606
rect 15317 11564 16011 11572
rect 15317 11530 15404 11564
rect 15438 11530 15504 11564
rect 15538 11530 15604 11564
rect 15638 11530 15704 11564
rect 15738 11530 15804 11564
rect 15838 11530 15904 11564
rect 15938 11530 16011 11564
rect 15317 11516 16011 11530
rect 15317 11482 15376 11516
rect 15410 11482 15466 11516
rect 15500 11482 15556 11516
rect 15590 11482 15646 11516
rect 15680 11482 15736 11516
rect 15770 11482 15826 11516
rect 15860 11482 15916 11516
rect 15950 11482 16011 11516
rect 15317 11464 16011 11482
rect 15317 11430 15404 11464
rect 15438 11430 15504 11464
rect 15538 11430 15604 11464
rect 15638 11430 15704 11464
rect 15738 11430 15804 11464
rect 15838 11430 15904 11464
rect 15938 11430 16011 11464
rect 15317 11426 16011 11430
rect 15317 11392 15376 11426
rect 15410 11392 15466 11426
rect 15500 11392 15556 11426
rect 15590 11392 15646 11426
rect 15680 11392 15736 11426
rect 15770 11392 15826 11426
rect 15860 11392 15916 11426
rect 15950 11392 16011 11426
rect 15317 11364 16011 11392
rect 15317 11336 15404 11364
rect 15438 11336 15504 11364
rect 15317 11302 15376 11336
rect 15438 11330 15466 11336
rect 15410 11302 15466 11330
rect 15500 11330 15504 11336
rect 15538 11336 15604 11364
rect 15538 11330 15556 11336
rect 15500 11302 15556 11330
rect 15590 11330 15604 11336
rect 15638 11336 15704 11364
rect 15738 11336 15804 11364
rect 15838 11336 15904 11364
rect 15938 11336 16011 11364
rect 15638 11330 15646 11336
rect 15590 11302 15646 11330
rect 15680 11330 15704 11336
rect 15770 11330 15804 11336
rect 15860 11330 15904 11336
rect 15680 11302 15736 11330
rect 15770 11302 15826 11330
rect 15860 11302 15916 11330
rect 15950 11302 16011 11336
rect 15317 11243 16011 11302
rect 16073 11905 16092 11939
rect 16126 11938 16490 11939
rect 16126 11905 16240 11938
rect 16073 11904 16240 11905
rect 16274 11904 16341 11938
rect 16375 11924 16490 11938
rect 16524 11924 16543 11958
rect 17361 11994 17528 11999
rect 17562 11994 17629 12028
rect 17663 12018 17870 12028
rect 17904 12018 17960 12052
rect 17994 12018 18050 12052
rect 18084 12018 18140 12052
rect 18174 12018 18230 12052
rect 18264 12018 18320 12052
rect 18354 12018 18410 12052
rect 18444 12018 18500 12052
rect 18534 12018 18590 12052
rect 18624 12028 18884 12052
rect 18624 12018 18816 12028
rect 17663 11999 18816 12018
rect 17663 11994 17831 11999
rect 17361 11958 17831 11994
rect 17361 11939 17778 11958
rect 16375 11904 16543 11924
rect 16073 11868 16543 11904
rect 16073 11849 16490 11868
rect 16073 11815 16092 11849
rect 16126 11848 16490 11849
rect 16126 11815 16240 11848
rect 16073 11814 16240 11815
rect 16274 11814 16341 11848
rect 16375 11834 16490 11848
rect 16524 11834 16543 11868
rect 16375 11814 16543 11834
rect 16073 11778 16543 11814
rect 16073 11759 16490 11778
rect 16073 11725 16092 11759
rect 16126 11758 16490 11759
rect 16126 11725 16240 11758
rect 16073 11724 16240 11725
rect 16274 11724 16341 11758
rect 16375 11744 16490 11758
rect 16524 11744 16543 11778
rect 16375 11724 16543 11744
rect 16073 11688 16543 11724
rect 16073 11669 16490 11688
rect 16073 11635 16092 11669
rect 16126 11668 16490 11669
rect 16126 11635 16240 11668
rect 16073 11634 16240 11635
rect 16274 11634 16341 11668
rect 16375 11654 16490 11668
rect 16524 11654 16543 11688
rect 16375 11634 16543 11654
rect 16073 11598 16543 11634
rect 16073 11579 16490 11598
rect 16073 11545 16092 11579
rect 16126 11578 16490 11579
rect 16126 11545 16240 11578
rect 16073 11544 16240 11545
rect 16274 11544 16341 11578
rect 16375 11564 16490 11578
rect 16524 11564 16543 11598
rect 16375 11544 16543 11564
rect 16073 11508 16543 11544
rect 16073 11489 16490 11508
rect 16073 11455 16092 11489
rect 16126 11488 16490 11489
rect 16126 11455 16240 11488
rect 16073 11454 16240 11455
rect 16274 11454 16341 11488
rect 16375 11474 16490 11488
rect 16524 11474 16543 11508
rect 16375 11454 16543 11474
rect 16073 11418 16543 11454
rect 16073 11399 16490 11418
rect 16073 11365 16092 11399
rect 16126 11398 16490 11399
rect 16126 11365 16240 11398
rect 16073 11364 16240 11365
rect 16274 11364 16341 11398
rect 16375 11384 16490 11398
rect 16524 11384 16543 11418
rect 16375 11364 16543 11384
rect 16073 11328 16543 11364
rect 16073 11309 16490 11328
rect 16073 11275 16092 11309
rect 16126 11308 16490 11309
rect 16126 11275 16240 11308
rect 16073 11274 16240 11275
rect 16274 11274 16341 11308
rect 16375 11294 16490 11308
rect 16524 11294 16543 11328
rect 16375 11274 16543 11294
rect 14784 11219 15202 11238
rect 14784 11185 14804 11219
rect 14838 11218 15202 11219
rect 14838 11185 14952 11218
rect 14784 11184 14952 11185
rect 14986 11184 15053 11218
rect 15087 11204 15202 11218
rect 15236 11204 15255 11238
rect 15087 11184 15255 11204
rect 14784 11181 15255 11184
rect 16073 11238 16543 11274
rect 16605 11876 17299 11937
rect 16605 11842 16664 11876
rect 16698 11864 16754 11876
rect 16726 11842 16754 11864
rect 16788 11864 16844 11876
rect 16788 11842 16792 11864
rect 16605 11830 16692 11842
rect 16726 11830 16792 11842
rect 16826 11842 16844 11864
rect 16878 11864 16934 11876
rect 16878 11842 16892 11864
rect 16826 11830 16892 11842
rect 16926 11842 16934 11864
rect 16968 11864 17024 11876
rect 17058 11864 17114 11876
rect 17148 11864 17204 11876
rect 16968 11842 16992 11864
rect 17058 11842 17092 11864
rect 17148 11842 17192 11864
rect 17238 11842 17299 11876
rect 16926 11830 16992 11842
rect 17026 11830 17092 11842
rect 17126 11830 17192 11842
rect 17226 11830 17299 11842
rect 16605 11786 17299 11830
rect 16605 11752 16664 11786
rect 16698 11764 16754 11786
rect 16726 11752 16754 11764
rect 16788 11764 16844 11786
rect 16788 11752 16792 11764
rect 16605 11730 16692 11752
rect 16726 11730 16792 11752
rect 16826 11752 16844 11764
rect 16878 11764 16934 11786
rect 16878 11752 16892 11764
rect 16826 11730 16892 11752
rect 16926 11752 16934 11764
rect 16968 11764 17024 11786
rect 17058 11764 17114 11786
rect 17148 11764 17204 11786
rect 16968 11752 16992 11764
rect 17058 11752 17092 11764
rect 17148 11752 17192 11764
rect 17238 11752 17299 11786
rect 16926 11730 16992 11752
rect 17026 11730 17092 11752
rect 17126 11730 17192 11752
rect 17226 11730 17299 11752
rect 16605 11696 17299 11730
rect 16605 11662 16664 11696
rect 16698 11664 16754 11696
rect 16726 11662 16754 11664
rect 16788 11664 16844 11696
rect 16788 11662 16792 11664
rect 16605 11630 16692 11662
rect 16726 11630 16792 11662
rect 16826 11662 16844 11664
rect 16878 11664 16934 11696
rect 16878 11662 16892 11664
rect 16826 11630 16892 11662
rect 16926 11662 16934 11664
rect 16968 11664 17024 11696
rect 17058 11664 17114 11696
rect 17148 11664 17204 11696
rect 16968 11662 16992 11664
rect 17058 11662 17092 11664
rect 17148 11662 17192 11664
rect 17238 11662 17299 11696
rect 16926 11630 16992 11662
rect 17026 11630 17092 11662
rect 17126 11630 17192 11662
rect 17226 11630 17299 11662
rect 16605 11606 17299 11630
rect 16605 11572 16664 11606
rect 16698 11572 16754 11606
rect 16788 11572 16844 11606
rect 16878 11572 16934 11606
rect 16968 11572 17024 11606
rect 17058 11572 17114 11606
rect 17148 11572 17204 11606
rect 17238 11572 17299 11606
rect 16605 11564 17299 11572
rect 16605 11530 16692 11564
rect 16726 11530 16792 11564
rect 16826 11530 16892 11564
rect 16926 11530 16992 11564
rect 17026 11530 17092 11564
rect 17126 11530 17192 11564
rect 17226 11530 17299 11564
rect 16605 11516 17299 11530
rect 16605 11482 16664 11516
rect 16698 11482 16754 11516
rect 16788 11482 16844 11516
rect 16878 11482 16934 11516
rect 16968 11482 17024 11516
rect 17058 11482 17114 11516
rect 17148 11482 17204 11516
rect 17238 11482 17299 11516
rect 16605 11464 17299 11482
rect 16605 11430 16692 11464
rect 16726 11430 16792 11464
rect 16826 11430 16892 11464
rect 16926 11430 16992 11464
rect 17026 11430 17092 11464
rect 17126 11430 17192 11464
rect 17226 11430 17299 11464
rect 16605 11426 17299 11430
rect 16605 11392 16664 11426
rect 16698 11392 16754 11426
rect 16788 11392 16844 11426
rect 16878 11392 16934 11426
rect 16968 11392 17024 11426
rect 17058 11392 17114 11426
rect 17148 11392 17204 11426
rect 17238 11392 17299 11426
rect 16605 11364 17299 11392
rect 16605 11336 16692 11364
rect 16726 11336 16792 11364
rect 16605 11302 16664 11336
rect 16726 11330 16754 11336
rect 16698 11302 16754 11330
rect 16788 11330 16792 11336
rect 16826 11336 16892 11364
rect 16826 11330 16844 11336
rect 16788 11302 16844 11330
rect 16878 11330 16892 11336
rect 16926 11336 16992 11364
rect 17026 11336 17092 11364
rect 17126 11336 17192 11364
rect 17226 11336 17299 11364
rect 16926 11330 16934 11336
rect 16878 11302 16934 11330
rect 16968 11330 16992 11336
rect 17058 11330 17092 11336
rect 17148 11330 17192 11336
rect 16968 11302 17024 11330
rect 17058 11302 17114 11330
rect 17148 11302 17204 11330
rect 17238 11302 17299 11336
rect 16605 11243 17299 11302
rect 17361 11905 17380 11939
rect 17414 11938 17778 11939
rect 17414 11905 17528 11938
rect 17361 11904 17528 11905
rect 17562 11904 17629 11938
rect 17663 11924 17778 11938
rect 17812 11924 17831 11958
rect 18649 11994 18816 11999
rect 18850 11994 18884 12028
rect 18649 11939 18884 11994
rect 17663 11904 17831 11924
rect 17361 11868 17831 11904
rect 17361 11849 17778 11868
rect 17361 11815 17380 11849
rect 17414 11848 17778 11849
rect 17414 11815 17528 11848
rect 17361 11814 17528 11815
rect 17562 11814 17629 11848
rect 17663 11834 17778 11848
rect 17812 11834 17831 11868
rect 17663 11814 17831 11834
rect 17361 11778 17831 11814
rect 17361 11759 17778 11778
rect 17361 11725 17380 11759
rect 17414 11758 17778 11759
rect 17414 11725 17528 11758
rect 17361 11724 17528 11725
rect 17562 11724 17629 11758
rect 17663 11744 17778 11758
rect 17812 11744 17831 11778
rect 17663 11724 17831 11744
rect 17361 11688 17831 11724
rect 17361 11669 17778 11688
rect 17361 11635 17380 11669
rect 17414 11668 17778 11669
rect 17414 11635 17528 11668
rect 17361 11634 17528 11635
rect 17562 11634 17629 11668
rect 17663 11654 17778 11668
rect 17812 11654 17831 11688
rect 17663 11634 17831 11654
rect 17361 11598 17831 11634
rect 17361 11579 17778 11598
rect 17361 11545 17380 11579
rect 17414 11578 17778 11579
rect 17414 11545 17528 11578
rect 17361 11544 17528 11545
rect 17562 11544 17629 11578
rect 17663 11564 17778 11578
rect 17812 11564 17831 11598
rect 17663 11544 17831 11564
rect 17361 11508 17831 11544
rect 17361 11489 17778 11508
rect 17361 11455 17380 11489
rect 17414 11488 17778 11489
rect 17414 11455 17528 11488
rect 17361 11454 17528 11455
rect 17562 11454 17629 11488
rect 17663 11474 17778 11488
rect 17812 11474 17831 11508
rect 17663 11454 17831 11474
rect 17361 11418 17831 11454
rect 17361 11399 17778 11418
rect 17361 11365 17380 11399
rect 17414 11398 17778 11399
rect 17414 11365 17528 11398
rect 17361 11364 17528 11365
rect 17562 11364 17629 11398
rect 17663 11384 17778 11398
rect 17812 11384 17831 11418
rect 17663 11364 17831 11384
rect 17361 11328 17831 11364
rect 17361 11309 17778 11328
rect 17361 11275 17380 11309
rect 17414 11308 17778 11309
rect 17414 11275 17528 11308
rect 17361 11274 17528 11275
rect 17562 11274 17629 11308
rect 17663 11294 17778 11308
rect 17812 11294 17831 11328
rect 17663 11274 17831 11294
rect 16073 11219 16490 11238
rect 16073 11185 16092 11219
rect 16126 11218 16490 11219
rect 16126 11185 16240 11218
rect 16073 11184 16240 11185
rect 16274 11184 16341 11218
rect 16375 11204 16490 11218
rect 16524 11204 16543 11238
rect 16375 11184 16543 11204
rect 16073 11181 16543 11184
rect 17361 11238 17831 11274
rect 17893 11876 18587 11937
rect 17893 11842 17952 11876
rect 17986 11864 18042 11876
rect 18014 11842 18042 11864
rect 18076 11864 18132 11876
rect 18076 11842 18080 11864
rect 17893 11830 17980 11842
rect 18014 11830 18080 11842
rect 18114 11842 18132 11864
rect 18166 11864 18222 11876
rect 18166 11842 18180 11864
rect 18114 11830 18180 11842
rect 18214 11842 18222 11864
rect 18256 11864 18312 11876
rect 18346 11864 18402 11876
rect 18436 11864 18492 11876
rect 18256 11842 18280 11864
rect 18346 11842 18380 11864
rect 18436 11842 18480 11864
rect 18526 11842 18587 11876
rect 18214 11830 18280 11842
rect 18314 11830 18380 11842
rect 18414 11830 18480 11842
rect 18514 11830 18587 11842
rect 17893 11786 18587 11830
rect 17893 11752 17952 11786
rect 17986 11764 18042 11786
rect 18014 11752 18042 11764
rect 18076 11764 18132 11786
rect 18076 11752 18080 11764
rect 17893 11730 17980 11752
rect 18014 11730 18080 11752
rect 18114 11752 18132 11764
rect 18166 11764 18222 11786
rect 18166 11752 18180 11764
rect 18114 11730 18180 11752
rect 18214 11752 18222 11764
rect 18256 11764 18312 11786
rect 18346 11764 18402 11786
rect 18436 11764 18492 11786
rect 18256 11752 18280 11764
rect 18346 11752 18380 11764
rect 18436 11752 18480 11764
rect 18526 11752 18587 11786
rect 18214 11730 18280 11752
rect 18314 11730 18380 11752
rect 18414 11730 18480 11752
rect 18514 11730 18587 11752
rect 17893 11696 18587 11730
rect 17893 11662 17952 11696
rect 17986 11664 18042 11696
rect 18014 11662 18042 11664
rect 18076 11664 18132 11696
rect 18076 11662 18080 11664
rect 17893 11630 17980 11662
rect 18014 11630 18080 11662
rect 18114 11662 18132 11664
rect 18166 11664 18222 11696
rect 18166 11662 18180 11664
rect 18114 11630 18180 11662
rect 18214 11662 18222 11664
rect 18256 11664 18312 11696
rect 18346 11664 18402 11696
rect 18436 11664 18492 11696
rect 18256 11662 18280 11664
rect 18346 11662 18380 11664
rect 18436 11662 18480 11664
rect 18526 11662 18587 11696
rect 18214 11630 18280 11662
rect 18314 11630 18380 11662
rect 18414 11630 18480 11662
rect 18514 11630 18587 11662
rect 17893 11606 18587 11630
rect 17893 11572 17952 11606
rect 17986 11572 18042 11606
rect 18076 11572 18132 11606
rect 18166 11572 18222 11606
rect 18256 11572 18312 11606
rect 18346 11572 18402 11606
rect 18436 11572 18492 11606
rect 18526 11572 18587 11606
rect 17893 11564 18587 11572
rect 17893 11530 17980 11564
rect 18014 11530 18080 11564
rect 18114 11530 18180 11564
rect 18214 11530 18280 11564
rect 18314 11530 18380 11564
rect 18414 11530 18480 11564
rect 18514 11530 18587 11564
rect 17893 11516 18587 11530
rect 17893 11482 17952 11516
rect 17986 11482 18042 11516
rect 18076 11482 18132 11516
rect 18166 11482 18222 11516
rect 18256 11482 18312 11516
rect 18346 11482 18402 11516
rect 18436 11482 18492 11516
rect 18526 11482 18587 11516
rect 17893 11464 18587 11482
rect 17893 11430 17980 11464
rect 18014 11430 18080 11464
rect 18114 11430 18180 11464
rect 18214 11430 18280 11464
rect 18314 11430 18380 11464
rect 18414 11430 18480 11464
rect 18514 11430 18587 11464
rect 17893 11426 18587 11430
rect 17893 11392 17952 11426
rect 17986 11392 18042 11426
rect 18076 11392 18132 11426
rect 18166 11392 18222 11426
rect 18256 11392 18312 11426
rect 18346 11392 18402 11426
rect 18436 11392 18492 11426
rect 18526 11392 18587 11426
rect 17893 11364 18587 11392
rect 17893 11336 17980 11364
rect 18014 11336 18080 11364
rect 17893 11302 17952 11336
rect 18014 11330 18042 11336
rect 17986 11302 18042 11330
rect 18076 11330 18080 11336
rect 18114 11336 18180 11364
rect 18114 11330 18132 11336
rect 18076 11302 18132 11330
rect 18166 11330 18180 11336
rect 18214 11336 18280 11364
rect 18314 11336 18380 11364
rect 18414 11336 18480 11364
rect 18514 11336 18587 11364
rect 18214 11330 18222 11336
rect 18166 11302 18222 11330
rect 18256 11330 18280 11336
rect 18346 11330 18380 11336
rect 18436 11330 18480 11336
rect 18256 11302 18312 11330
rect 18346 11302 18402 11330
rect 18436 11302 18492 11330
rect 18526 11302 18587 11336
rect 17893 11243 18587 11302
rect 18649 11905 18668 11939
rect 18702 11938 18884 11939
rect 18702 11905 18816 11938
rect 18649 11904 18816 11905
rect 18850 11904 18884 11938
rect 18649 11849 18884 11904
rect 18649 11815 18668 11849
rect 18702 11848 18884 11849
rect 18702 11815 18816 11848
rect 18649 11814 18816 11815
rect 18850 11814 18884 11848
rect 18649 11759 18884 11814
rect 18649 11725 18668 11759
rect 18702 11758 18884 11759
rect 18702 11725 18816 11758
rect 18649 11724 18816 11725
rect 18850 11724 18884 11758
rect 18649 11669 18884 11724
rect 18649 11635 18668 11669
rect 18702 11668 18884 11669
rect 18702 11635 18816 11668
rect 18649 11634 18816 11635
rect 18850 11634 18884 11668
rect 18649 11579 18884 11634
rect 18649 11545 18668 11579
rect 18702 11578 18884 11579
rect 18702 11545 18816 11578
rect 18649 11544 18816 11545
rect 18850 11544 18884 11578
rect 18649 11489 18884 11544
rect 18649 11455 18668 11489
rect 18702 11488 18884 11489
rect 18702 11455 18816 11488
rect 18649 11454 18816 11455
rect 18850 11454 18884 11488
rect 18649 11399 18884 11454
rect 18649 11365 18668 11399
rect 18702 11398 18884 11399
rect 18702 11365 18816 11398
rect 18649 11364 18816 11365
rect 18850 11364 18884 11398
rect 18649 11309 18884 11364
rect 18649 11275 18668 11309
rect 18702 11308 18884 11309
rect 18702 11275 18816 11308
rect 18649 11274 18816 11275
rect 18850 11274 18884 11308
rect 17361 11219 17778 11238
rect 17361 11185 17380 11219
rect 17414 11218 17778 11219
rect 17414 11185 17528 11218
rect 17361 11184 17528 11185
rect 17562 11184 17629 11218
rect 17663 11204 17778 11218
rect 17812 11204 17831 11238
rect 17663 11184 17831 11204
rect 17361 11181 17831 11184
rect 18649 11219 18884 11274
rect 18649 11185 18668 11219
rect 18702 11218 18884 11219
rect 18702 11185 18816 11218
rect 18649 11184 18816 11185
rect 18850 11184 18884 11218
rect 18649 11181 18884 11184
rect 12444 11162 18884 11181
rect 12444 11128 12684 11162
rect 12718 11128 12774 11162
rect 12808 11128 12864 11162
rect 12898 11128 12954 11162
rect 12988 11128 13044 11162
rect 13078 11128 13134 11162
rect 13168 11128 13224 11162
rect 13258 11128 13314 11162
rect 13348 11128 13404 11162
rect 13438 11128 13972 11162
rect 14006 11128 14062 11162
rect 14096 11128 14152 11162
rect 14186 11128 14242 11162
rect 14276 11128 14332 11162
rect 14366 11128 14422 11162
rect 14456 11128 14512 11162
rect 14546 11128 14602 11162
rect 14636 11128 14692 11162
rect 14726 11128 15260 11162
rect 15294 11128 15350 11162
rect 15384 11128 15440 11162
rect 15474 11128 15530 11162
rect 15564 11128 15620 11162
rect 15654 11128 15710 11162
rect 15744 11128 15800 11162
rect 15834 11128 15890 11162
rect 15924 11128 15980 11162
rect 16014 11128 16548 11162
rect 16582 11128 16638 11162
rect 16672 11128 16728 11162
rect 16762 11128 16818 11162
rect 16852 11128 16908 11162
rect 16942 11128 16998 11162
rect 17032 11128 17088 11162
rect 17122 11128 17178 11162
rect 17212 11128 17268 11162
rect 17302 11128 17836 11162
rect 17870 11128 17926 11162
rect 17960 11128 18016 11162
rect 18050 11128 18106 11162
rect 18140 11128 18196 11162
rect 18230 11128 18286 11162
rect 18320 11128 18376 11162
rect 18410 11128 18466 11162
rect 18500 11128 18556 11162
rect 18590 11128 18884 11162
rect 12444 11094 12477 11128
rect 12511 11109 13664 11128
rect 12511 11094 12684 11109
rect 12444 11045 12684 11094
rect 13484 11094 13664 11109
rect 13698 11094 13765 11128
rect 13799 11109 14952 11128
rect 13799 11094 13984 11109
rect 13484 11045 13984 11094
rect 14784 11094 14952 11109
rect 14986 11094 15053 11128
rect 15087 11109 16240 11128
rect 15087 11094 15184 11109
rect 14784 11045 15184 11094
rect 16084 11094 16240 11109
rect 16274 11094 16341 11128
rect 16375 11109 17528 11128
rect 16375 11094 16484 11109
rect 16084 11045 16484 11094
rect 17384 11094 17528 11109
rect 17562 11094 17629 11128
rect 17663 11109 18816 11128
rect 17663 11094 17784 11109
rect 17384 11045 17784 11094
rect 18684 11094 18816 11109
rect 18850 11094 18884 11128
rect 18684 11045 18884 11094
rect 12444 11038 18884 11045
rect 12444 11004 12477 11038
rect 12511 11015 13664 11038
rect 12511 11004 12578 11015
rect 12444 10981 12578 11004
rect 12612 10981 12668 11015
rect 12702 10981 12758 11015
rect 12792 10981 12848 11015
rect 12882 10981 12938 11015
rect 12972 10981 13028 11015
rect 13062 10981 13118 11015
rect 13152 10981 13208 11015
rect 13242 10981 13298 11015
rect 13332 10981 13388 11015
rect 13422 10981 13478 11015
rect 13512 10981 13568 11015
rect 13602 11004 13664 11015
rect 13698 11004 13765 11038
rect 13799 11015 14952 11038
rect 13799 11004 13866 11015
rect 13602 10981 13866 11004
rect 13900 10981 13956 11015
rect 13990 10981 14046 11015
rect 14080 10981 14136 11015
rect 14170 10981 14226 11015
rect 14260 10981 14316 11015
rect 14350 10981 14406 11015
rect 14440 10981 14496 11015
rect 14530 10981 14586 11015
rect 14620 10981 14676 11015
rect 14710 10981 14766 11015
rect 14800 10981 14856 11015
rect 14890 11004 14952 11015
rect 14986 11004 15053 11038
rect 15087 11015 16240 11038
rect 15087 11004 15154 11015
rect 14890 10981 15154 11004
rect 15188 10981 15244 11015
rect 15278 10981 15334 11015
rect 15368 10981 15424 11015
rect 15458 10981 15514 11015
rect 15548 10981 15604 11015
rect 15638 10981 15694 11015
rect 15728 10981 15784 11015
rect 15818 10981 15874 11015
rect 15908 10981 15964 11015
rect 15998 10981 16054 11015
rect 16088 10981 16144 11015
rect 16178 11004 16240 11015
rect 16274 11004 16341 11038
rect 16375 11015 17528 11038
rect 16375 11004 16442 11015
rect 16178 10981 16442 11004
rect 16476 10981 16532 11015
rect 16566 10981 16622 11015
rect 16656 10981 16712 11015
rect 16746 10981 16802 11015
rect 16836 10981 16892 11015
rect 16926 10981 16982 11015
rect 17016 10981 17072 11015
rect 17106 10981 17162 11015
rect 17196 10981 17252 11015
rect 17286 10981 17342 11015
rect 17376 10981 17432 11015
rect 17466 11004 17528 11015
rect 17562 11004 17629 11038
rect 17663 11015 18816 11038
rect 17663 11004 17730 11015
rect 17466 10981 17730 11004
rect 17764 10981 17820 11015
rect 17854 10981 17910 11015
rect 17944 10981 18000 11015
rect 18034 10981 18090 11015
rect 18124 10981 18180 11015
rect 18214 10981 18270 11015
rect 18304 10981 18360 11015
rect 18394 10981 18450 11015
rect 18484 10981 18540 11015
rect 18574 10981 18630 11015
rect 18664 10981 18720 11015
rect 18754 11004 18816 11015
rect 18850 11004 18884 11038
rect 18754 10981 18884 11004
rect 12444 10914 18884 10981
rect 12444 10880 12578 10914
rect 12612 10880 12668 10914
rect 12702 10880 12758 10914
rect 12792 10880 12848 10914
rect 12882 10880 12938 10914
rect 12972 10880 13028 10914
rect 13062 10880 13118 10914
rect 13152 10880 13208 10914
rect 13242 10880 13298 10914
rect 13332 10880 13388 10914
rect 13422 10880 13478 10914
rect 13512 10880 13568 10914
rect 13602 10880 13866 10914
rect 13900 10880 13956 10914
rect 13990 10880 14046 10914
rect 14080 10880 14136 10914
rect 14170 10880 14226 10914
rect 14260 10880 14316 10914
rect 14350 10880 14406 10914
rect 14440 10880 14496 10914
rect 14530 10880 14586 10914
rect 14620 10880 14676 10914
rect 14710 10880 14766 10914
rect 14800 10880 14856 10914
rect 14890 10880 15154 10914
rect 15188 10880 15244 10914
rect 15278 10880 15334 10914
rect 15368 10880 15424 10914
rect 15458 10880 15514 10914
rect 15548 10880 15604 10914
rect 15638 10880 15694 10914
rect 15728 10880 15784 10914
rect 15818 10880 15874 10914
rect 15908 10880 15964 10914
rect 15998 10880 16054 10914
rect 16088 10880 16144 10914
rect 16178 10880 16442 10914
rect 16476 10880 16532 10914
rect 16566 10880 16622 10914
rect 16656 10880 16712 10914
rect 16746 10880 16802 10914
rect 16836 10880 16892 10914
rect 16926 10880 16982 10914
rect 17016 10880 17072 10914
rect 17106 10880 17162 10914
rect 17196 10880 17252 10914
rect 17286 10880 17342 10914
rect 17376 10880 17432 10914
rect 17466 10880 17730 10914
rect 17764 10880 17820 10914
rect 17854 10880 17910 10914
rect 17944 10880 18000 10914
rect 18034 10880 18090 10914
rect 18124 10880 18180 10914
rect 18214 10880 18270 10914
rect 18304 10880 18360 10914
rect 18394 10880 18450 10914
rect 18484 10880 18540 10914
rect 18574 10880 18630 10914
rect 18664 10880 18720 10914
rect 18754 10880 18884 10914
rect 12444 10847 18884 10880
rect 12444 10830 12684 10847
rect 12444 10796 12477 10830
rect 12511 10796 12684 10830
rect 12444 10783 12684 10796
rect 13484 10830 13984 10847
rect 13484 10796 13664 10830
rect 13698 10796 13765 10830
rect 13799 10796 13984 10830
rect 13484 10783 13984 10796
rect 14784 10830 15184 10847
rect 14784 10796 14952 10830
rect 14986 10796 15053 10830
rect 15087 10796 15184 10830
rect 14784 10783 15184 10796
rect 16084 10830 16484 10847
rect 16084 10796 16240 10830
rect 16274 10796 16341 10830
rect 16375 10796 16484 10830
rect 16084 10783 16484 10796
rect 17384 10830 17784 10847
rect 17384 10796 17528 10830
rect 17562 10796 17629 10830
rect 17663 10796 17784 10830
rect 17384 10783 17784 10796
rect 18684 10830 18884 10847
rect 18684 10796 18816 10830
rect 18850 10796 18884 10830
rect 18684 10783 18884 10796
rect 12444 10764 18884 10783
rect 12444 10740 12718 10764
rect 12444 10706 12477 10740
rect 12511 10730 12718 10740
rect 12752 10730 12808 10764
rect 12842 10730 12898 10764
rect 12932 10730 12988 10764
rect 13022 10730 13078 10764
rect 13112 10730 13168 10764
rect 13202 10730 13258 10764
rect 13292 10730 13348 10764
rect 13382 10730 13438 10764
rect 13472 10740 14006 10764
rect 13472 10730 13664 10740
rect 12511 10711 13664 10730
rect 12511 10706 12684 10711
rect 12444 10670 12684 10706
rect 12444 10650 12626 10670
rect 12444 10616 12477 10650
rect 12511 10636 12626 10650
rect 12660 10636 12684 10670
rect 13484 10706 13664 10711
rect 13698 10706 13765 10740
rect 13799 10730 14006 10740
rect 14040 10730 14096 10764
rect 14130 10730 14186 10764
rect 14220 10730 14276 10764
rect 14310 10730 14366 10764
rect 14400 10730 14456 10764
rect 14490 10730 14546 10764
rect 14580 10730 14636 10764
rect 14670 10730 14726 10764
rect 14760 10740 15294 10764
rect 14760 10730 14952 10740
rect 13799 10711 14952 10730
rect 13799 10706 13984 10711
rect 13484 10670 13984 10706
rect 13484 10651 13914 10670
rect 12511 10616 12684 10636
rect 12444 10580 12684 10616
rect 12444 10560 12626 10580
rect 12444 10526 12477 10560
rect 12511 10546 12626 10560
rect 12660 10546 12684 10580
rect 12511 10526 12684 10546
rect 12444 10490 12684 10526
rect 12444 10470 12626 10490
rect 12444 10436 12477 10470
rect 12511 10456 12626 10470
rect 12660 10456 12684 10490
rect 12511 10436 12684 10456
rect 12444 10400 12684 10436
rect 12444 10380 12626 10400
rect 12444 10346 12477 10380
rect 12511 10366 12626 10380
rect 12660 10366 12684 10400
rect 12511 10346 12684 10366
rect 12444 10310 12684 10346
rect 12444 10290 12626 10310
rect 12444 10256 12477 10290
rect 12511 10276 12626 10290
rect 12660 10276 12684 10310
rect 12511 10256 12684 10276
rect 12444 10220 12684 10256
rect 12444 10200 12626 10220
rect 12444 10166 12477 10200
rect 12511 10186 12626 10200
rect 12660 10186 12684 10220
rect 12511 10166 12684 10186
rect 12444 10130 12684 10166
rect 12444 10110 12626 10130
rect 12444 10076 12477 10110
rect 12511 10096 12626 10110
rect 12660 10096 12684 10130
rect 12511 10076 12684 10096
rect 12444 10040 12684 10076
rect 12444 10020 12626 10040
rect 12444 9986 12477 10020
rect 12511 10006 12626 10020
rect 12660 10006 12684 10040
rect 12511 9986 12684 10006
rect 12444 9950 12684 9986
rect 12741 10588 13435 10649
rect 12741 10554 12800 10588
rect 12834 10576 12890 10588
rect 12862 10554 12890 10576
rect 12924 10576 12980 10588
rect 12924 10554 12928 10576
rect 12741 10542 12828 10554
rect 12862 10542 12928 10554
rect 12962 10554 12980 10576
rect 13014 10576 13070 10588
rect 13014 10554 13028 10576
rect 12962 10542 13028 10554
rect 13062 10554 13070 10576
rect 13104 10576 13160 10588
rect 13194 10576 13250 10588
rect 13284 10576 13340 10588
rect 13104 10554 13128 10576
rect 13194 10554 13228 10576
rect 13284 10554 13328 10576
rect 13374 10554 13435 10588
rect 13062 10542 13128 10554
rect 13162 10542 13228 10554
rect 13262 10542 13328 10554
rect 13362 10542 13435 10554
rect 12741 10498 13435 10542
rect 12741 10464 12800 10498
rect 12834 10476 12890 10498
rect 12862 10464 12890 10476
rect 12924 10476 12980 10498
rect 12924 10464 12928 10476
rect 12741 10442 12828 10464
rect 12862 10442 12928 10464
rect 12962 10464 12980 10476
rect 13014 10476 13070 10498
rect 13014 10464 13028 10476
rect 12962 10442 13028 10464
rect 13062 10464 13070 10476
rect 13104 10476 13160 10498
rect 13194 10476 13250 10498
rect 13284 10476 13340 10498
rect 13104 10464 13128 10476
rect 13194 10464 13228 10476
rect 13284 10464 13328 10476
rect 13374 10464 13435 10498
rect 13062 10442 13128 10464
rect 13162 10442 13228 10464
rect 13262 10442 13328 10464
rect 13362 10442 13435 10464
rect 12741 10408 13435 10442
rect 12741 10374 12800 10408
rect 12834 10376 12890 10408
rect 12862 10374 12890 10376
rect 12924 10376 12980 10408
rect 12924 10374 12928 10376
rect 12741 10342 12828 10374
rect 12862 10342 12928 10374
rect 12962 10374 12980 10376
rect 13014 10376 13070 10408
rect 13014 10374 13028 10376
rect 12962 10342 13028 10374
rect 13062 10374 13070 10376
rect 13104 10376 13160 10408
rect 13194 10376 13250 10408
rect 13284 10376 13340 10408
rect 13104 10374 13128 10376
rect 13194 10374 13228 10376
rect 13284 10374 13328 10376
rect 13374 10374 13435 10408
rect 13062 10342 13128 10374
rect 13162 10342 13228 10374
rect 13262 10342 13328 10374
rect 13362 10342 13435 10374
rect 12741 10318 13435 10342
rect 12741 10284 12800 10318
rect 12834 10284 12890 10318
rect 12924 10284 12980 10318
rect 13014 10284 13070 10318
rect 13104 10284 13160 10318
rect 13194 10284 13250 10318
rect 13284 10284 13340 10318
rect 13374 10284 13435 10318
rect 12741 10276 13435 10284
rect 12741 10242 12828 10276
rect 12862 10242 12928 10276
rect 12962 10242 13028 10276
rect 13062 10242 13128 10276
rect 13162 10242 13228 10276
rect 13262 10242 13328 10276
rect 13362 10242 13435 10276
rect 12741 10228 13435 10242
rect 12741 10194 12800 10228
rect 12834 10194 12890 10228
rect 12924 10194 12980 10228
rect 13014 10194 13070 10228
rect 13104 10194 13160 10228
rect 13194 10194 13250 10228
rect 13284 10194 13340 10228
rect 13374 10194 13435 10228
rect 12741 10176 13435 10194
rect 12741 10142 12828 10176
rect 12862 10142 12928 10176
rect 12962 10142 13028 10176
rect 13062 10142 13128 10176
rect 13162 10142 13228 10176
rect 13262 10142 13328 10176
rect 13362 10142 13435 10176
rect 12741 10138 13435 10142
rect 12741 10104 12800 10138
rect 12834 10104 12890 10138
rect 12924 10104 12980 10138
rect 13014 10104 13070 10138
rect 13104 10104 13160 10138
rect 13194 10104 13250 10138
rect 13284 10104 13340 10138
rect 13374 10104 13435 10138
rect 12741 10076 13435 10104
rect 12741 10048 12828 10076
rect 12862 10048 12928 10076
rect 12741 10014 12800 10048
rect 12862 10042 12890 10048
rect 12834 10014 12890 10042
rect 12924 10042 12928 10048
rect 12962 10048 13028 10076
rect 12962 10042 12980 10048
rect 12924 10014 12980 10042
rect 13014 10042 13028 10048
rect 13062 10048 13128 10076
rect 13162 10048 13228 10076
rect 13262 10048 13328 10076
rect 13362 10048 13435 10076
rect 13062 10042 13070 10048
rect 13014 10014 13070 10042
rect 13104 10042 13128 10048
rect 13194 10042 13228 10048
rect 13284 10042 13328 10048
rect 13104 10014 13160 10042
rect 13194 10014 13250 10042
rect 13284 10014 13340 10042
rect 13374 10014 13435 10048
rect 12741 9955 13435 10014
rect 13484 10617 13516 10651
rect 13550 10650 13914 10651
rect 13550 10617 13664 10650
rect 13484 10616 13664 10617
rect 13698 10616 13765 10650
rect 13799 10636 13914 10650
rect 13948 10636 13984 10670
rect 14784 10706 14952 10711
rect 14986 10706 15053 10740
rect 15087 10730 15294 10740
rect 15328 10730 15384 10764
rect 15418 10730 15474 10764
rect 15508 10730 15564 10764
rect 15598 10730 15654 10764
rect 15688 10730 15744 10764
rect 15778 10730 15834 10764
rect 15868 10730 15924 10764
rect 15958 10730 16014 10764
rect 16048 10740 16582 10764
rect 16048 10730 16240 10740
rect 15087 10711 16240 10730
rect 15087 10706 15255 10711
rect 14784 10670 15255 10706
rect 14784 10651 15202 10670
rect 13799 10616 13984 10636
rect 13484 10580 13984 10616
rect 13484 10561 13914 10580
rect 13484 10527 13516 10561
rect 13550 10560 13914 10561
rect 13550 10527 13664 10560
rect 13484 10526 13664 10527
rect 13698 10526 13765 10560
rect 13799 10546 13914 10560
rect 13948 10546 13984 10580
rect 13799 10526 13984 10546
rect 13484 10490 13984 10526
rect 13484 10471 13914 10490
rect 13484 10437 13516 10471
rect 13550 10470 13914 10471
rect 13550 10437 13664 10470
rect 13484 10436 13664 10437
rect 13698 10436 13765 10470
rect 13799 10456 13914 10470
rect 13948 10456 13984 10490
rect 13799 10436 13984 10456
rect 13484 10400 13984 10436
rect 13484 10381 13914 10400
rect 13484 10347 13516 10381
rect 13550 10380 13914 10381
rect 13550 10347 13664 10380
rect 13484 10346 13664 10347
rect 13698 10346 13765 10380
rect 13799 10366 13914 10380
rect 13948 10366 13984 10400
rect 13799 10346 13984 10366
rect 13484 10310 13984 10346
rect 13484 10291 13914 10310
rect 13484 10257 13516 10291
rect 13550 10290 13914 10291
rect 13550 10257 13664 10290
rect 13484 10256 13664 10257
rect 13698 10256 13765 10290
rect 13799 10276 13914 10290
rect 13948 10276 13984 10310
rect 13799 10256 13984 10276
rect 13484 10220 13984 10256
rect 13484 10201 13914 10220
rect 13484 10167 13516 10201
rect 13550 10200 13914 10201
rect 13550 10167 13664 10200
rect 13484 10166 13664 10167
rect 13698 10166 13765 10200
rect 13799 10186 13914 10200
rect 13948 10186 13984 10220
rect 13799 10166 13984 10186
rect 13484 10130 13984 10166
rect 13484 10111 13914 10130
rect 13484 10077 13516 10111
rect 13550 10110 13914 10111
rect 13550 10077 13664 10110
rect 13484 10076 13664 10077
rect 13698 10076 13765 10110
rect 13799 10096 13914 10110
rect 13948 10096 13984 10130
rect 13799 10076 13984 10096
rect 13484 10040 13984 10076
rect 13484 10021 13914 10040
rect 13484 9987 13516 10021
rect 13550 10020 13914 10021
rect 13550 9987 13664 10020
rect 13484 9986 13664 9987
rect 13698 9986 13765 10020
rect 13799 10006 13914 10020
rect 13948 10006 13984 10040
rect 13799 9986 13984 10006
rect 12444 9930 12626 9950
rect 12444 9896 12477 9930
rect 12511 9916 12626 9930
rect 12660 9916 12684 9950
rect 12511 9896 12684 9916
rect 12444 9893 12684 9896
rect 13484 9950 13984 9986
rect 14029 10588 14723 10649
rect 14029 10554 14088 10588
rect 14122 10576 14178 10588
rect 14150 10554 14178 10576
rect 14212 10576 14268 10588
rect 14212 10554 14216 10576
rect 14029 10542 14116 10554
rect 14150 10542 14216 10554
rect 14250 10554 14268 10576
rect 14302 10576 14358 10588
rect 14302 10554 14316 10576
rect 14250 10542 14316 10554
rect 14350 10554 14358 10576
rect 14392 10576 14448 10588
rect 14482 10576 14538 10588
rect 14572 10576 14628 10588
rect 14392 10554 14416 10576
rect 14482 10554 14516 10576
rect 14572 10554 14616 10576
rect 14662 10554 14723 10588
rect 14350 10542 14416 10554
rect 14450 10542 14516 10554
rect 14550 10542 14616 10554
rect 14650 10542 14723 10554
rect 14029 10498 14723 10542
rect 14029 10464 14088 10498
rect 14122 10476 14178 10498
rect 14150 10464 14178 10476
rect 14212 10476 14268 10498
rect 14212 10464 14216 10476
rect 14029 10442 14116 10464
rect 14150 10442 14216 10464
rect 14250 10464 14268 10476
rect 14302 10476 14358 10498
rect 14302 10464 14316 10476
rect 14250 10442 14316 10464
rect 14350 10464 14358 10476
rect 14392 10476 14448 10498
rect 14482 10476 14538 10498
rect 14572 10476 14628 10498
rect 14392 10464 14416 10476
rect 14482 10464 14516 10476
rect 14572 10464 14616 10476
rect 14662 10464 14723 10498
rect 14350 10442 14416 10464
rect 14450 10442 14516 10464
rect 14550 10442 14616 10464
rect 14650 10442 14723 10464
rect 14029 10408 14723 10442
rect 14029 10374 14088 10408
rect 14122 10376 14178 10408
rect 14150 10374 14178 10376
rect 14212 10376 14268 10408
rect 14212 10374 14216 10376
rect 14029 10342 14116 10374
rect 14150 10342 14216 10374
rect 14250 10374 14268 10376
rect 14302 10376 14358 10408
rect 14302 10374 14316 10376
rect 14250 10342 14316 10374
rect 14350 10374 14358 10376
rect 14392 10376 14448 10408
rect 14482 10376 14538 10408
rect 14572 10376 14628 10408
rect 14392 10374 14416 10376
rect 14482 10374 14516 10376
rect 14572 10374 14616 10376
rect 14662 10374 14723 10408
rect 14350 10342 14416 10374
rect 14450 10342 14516 10374
rect 14550 10342 14616 10374
rect 14650 10342 14723 10374
rect 14029 10318 14723 10342
rect 14029 10284 14088 10318
rect 14122 10284 14178 10318
rect 14212 10284 14268 10318
rect 14302 10284 14358 10318
rect 14392 10284 14448 10318
rect 14482 10284 14538 10318
rect 14572 10284 14628 10318
rect 14662 10284 14723 10318
rect 14029 10276 14723 10284
rect 14029 10242 14116 10276
rect 14150 10242 14216 10276
rect 14250 10242 14316 10276
rect 14350 10242 14416 10276
rect 14450 10242 14516 10276
rect 14550 10242 14616 10276
rect 14650 10242 14723 10276
rect 14029 10228 14723 10242
rect 14029 10194 14088 10228
rect 14122 10194 14178 10228
rect 14212 10194 14268 10228
rect 14302 10194 14358 10228
rect 14392 10194 14448 10228
rect 14482 10194 14538 10228
rect 14572 10194 14628 10228
rect 14662 10194 14723 10228
rect 14029 10176 14723 10194
rect 14029 10142 14116 10176
rect 14150 10142 14216 10176
rect 14250 10142 14316 10176
rect 14350 10142 14416 10176
rect 14450 10142 14516 10176
rect 14550 10142 14616 10176
rect 14650 10142 14723 10176
rect 14029 10138 14723 10142
rect 14029 10104 14088 10138
rect 14122 10104 14178 10138
rect 14212 10104 14268 10138
rect 14302 10104 14358 10138
rect 14392 10104 14448 10138
rect 14482 10104 14538 10138
rect 14572 10104 14628 10138
rect 14662 10104 14723 10138
rect 14029 10076 14723 10104
rect 14029 10048 14116 10076
rect 14150 10048 14216 10076
rect 14029 10014 14088 10048
rect 14150 10042 14178 10048
rect 14122 10014 14178 10042
rect 14212 10042 14216 10048
rect 14250 10048 14316 10076
rect 14250 10042 14268 10048
rect 14212 10014 14268 10042
rect 14302 10042 14316 10048
rect 14350 10048 14416 10076
rect 14450 10048 14516 10076
rect 14550 10048 14616 10076
rect 14650 10048 14723 10076
rect 14350 10042 14358 10048
rect 14302 10014 14358 10042
rect 14392 10042 14416 10048
rect 14482 10042 14516 10048
rect 14572 10042 14616 10048
rect 14392 10014 14448 10042
rect 14482 10014 14538 10042
rect 14572 10014 14628 10042
rect 14662 10014 14723 10048
rect 14029 9955 14723 10014
rect 14784 10617 14804 10651
rect 14838 10650 15202 10651
rect 14838 10617 14952 10650
rect 14784 10616 14952 10617
rect 14986 10616 15053 10650
rect 15087 10636 15202 10650
rect 15236 10636 15255 10670
rect 16073 10706 16240 10711
rect 16274 10706 16341 10740
rect 16375 10730 16582 10740
rect 16616 10730 16672 10764
rect 16706 10730 16762 10764
rect 16796 10730 16852 10764
rect 16886 10730 16942 10764
rect 16976 10730 17032 10764
rect 17066 10730 17122 10764
rect 17156 10730 17212 10764
rect 17246 10730 17302 10764
rect 17336 10740 17870 10764
rect 17336 10730 17528 10740
rect 16375 10711 17528 10730
rect 16375 10706 16543 10711
rect 16073 10670 16543 10706
rect 16073 10651 16490 10670
rect 15087 10616 15255 10636
rect 14784 10580 15255 10616
rect 14784 10561 15202 10580
rect 14784 10527 14804 10561
rect 14838 10560 15202 10561
rect 14838 10527 14952 10560
rect 14784 10526 14952 10527
rect 14986 10526 15053 10560
rect 15087 10546 15202 10560
rect 15236 10546 15255 10580
rect 15087 10526 15255 10546
rect 14784 10490 15255 10526
rect 14784 10471 15202 10490
rect 14784 10437 14804 10471
rect 14838 10470 15202 10471
rect 14838 10437 14952 10470
rect 14784 10436 14952 10437
rect 14986 10436 15053 10470
rect 15087 10456 15202 10470
rect 15236 10456 15255 10490
rect 15087 10436 15255 10456
rect 14784 10400 15255 10436
rect 14784 10381 15202 10400
rect 14784 10347 14804 10381
rect 14838 10380 15202 10381
rect 14838 10347 14952 10380
rect 14784 10346 14952 10347
rect 14986 10346 15053 10380
rect 15087 10366 15202 10380
rect 15236 10366 15255 10400
rect 15087 10346 15255 10366
rect 14784 10310 15255 10346
rect 14784 10291 15202 10310
rect 14784 10257 14804 10291
rect 14838 10290 15202 10291
rect 14838 10257 14952 10290
rect 14784 10256 14952 10257
rect 14986 10256 15053 10290
rect 15087 10276 15202 10290
rect 15236 10276 15255 10310
rect 15087 10256 15255 10276
rect 14784 10220 15255 10256
rect 14784 10201 15202 10220
rect 14784 10167 14804 10201
rect 14838 10200 15202 10201
rect 14838 10167 14952 10200
rect 14784 10166 14952 10167
rect 14986 10166 15053 10200
rect 15087 10186 15202 10200
rect 15236 10186 15255 10220
rect 15087 10166 15255 10186
rect 14784 10130 15255 10166
rect 14784 10111 15202 10130
rect 14784 10077 14804 10111
rect 14838 10110 15202 10111
rect 14838 10077 14952 10110
rect 14784 10076 14952 10077
rect 14986 10076 15053 10110
rect 15087 10096 15202 10110
rect 15236 10096 15255 10130
rect 15087 10076 15255 10096
rect 14784 10040 15255 10076
rect 14784 10021 15202 10040
rect 14784 9987 14804 10021
rect 14838 10020 15202 10021
rect 14838 9987 14952 10020
rect 14784 9986 14952 9987
rect 14986 9986 15053 10020
rect 15087 10006 15202 10020
rect 15236 10006 15255 10040
rect 15087 9986 15255 10006
rect 13484 9931 13914 9950
rect 13484 9897 13516 9931
rect 13550 9930 13914 9931
rect 13550 9897 13664 9930
rect 13484 9896 13664 9897
rect 13698 9896 13765 9930
rect 13799 9916 13914 9930
rect 13948 9916 13984 9950
rect 13799 9896 13984 9916
rect 13484 9893 13984 9896
rect 14784 9950 15255 9986
rect 15317 10588 16011 10649
rect 15317 10554 15376 10588
rect 15410 10576 15466 10588
rect 15438 10554 15466 10576
rect 15500 10576 15556 10588
rect 15500 10554 15504 10576
rect 15317 10542 15404 10554
rect 15438 10542 15504 10554
rect 15538 10554 15556 10576
rect 15590 10576 15646 10588
rect 15590 10554 15604 10576
rect 15538 10542 15604 10554
rect 15638 10554 15646 10576
rect 15680 10576 15736 10588
rect 15770 10576 15826 10588
rect 15860 10576 15916 10588
rect 15680 10554 15704 10576
rect 15770 10554 15804 10576
rect 15860 10554 15904 10576
rect 15950 10554 16011 10588
rect 15638 10542 15704 10554
rect 15738 10542 15804 10554
rect 15838 10542 15904 10554
rect 15938 10542 16011 10554
rect 15317 10498 16011 10542
rect 15317 10464 15376 10498
rect 15410 10476 15466 10498
rect 15438 10464 15466 10476
rect 15500 10476 15556 10498
rect 15500 10464 15504 10476
rect 15317 10442 15404 10464
rect 15438 10442 15504 10464
rect 15538 10464 15556 10476
rect 15590 10476 15646 10498
rect 15590 10464 15604 10476
rect 15538 10442 15604 10464
rect 15638 10464 15646 10476
rect 15680 10476 15736 10498
rect 15770 10476 15826 10498
rect 15860 10476 15916 10498
rect 15680 10464 15704 10476
rect 15770 10464 15804 10476
rect 15860 10464 15904 10476
rect 15950 10464 16011 10498
rect 15638 10442 15704 10464
rect 15738 10442 15804 10464
rect 15838 10442 15904 10464
rect 15938 10442 16011 10464
rect 15317 10408 16011 10442
rect 15317 10374 15376 10408
rect 15410 10376 15466 10408
rect 15438 10374 15466 10376
rect 15500 10376 15556 10408
rect 15500 10374 15504 10376
rect 15317 10342 15404 10374
rect 15438 10342 15504 10374
rect 15538 10374 15556 10376
rect 15590 10376 15646 10408
rect 15590 10374 15604 10376
rect 15538 10342 15604 10374
rect 15638 10374 15646 10376
rect 15680 10376 15736 10408
rect 15770 10376 15826 10408
rect 15860 10376 15916 10408
rect 15680 10374 15704 10376
rect 15770 10374 15804 10376
rect 15860 10374 15904 10376
rect 15950 10374 16011 10408
rect 15638 10342 15704 10374
rect 15738 10342 15804 10374
rect 15838 10342 15904 10374
rect 15938 10342 16011 10374
rect 15317 10318 16011 10342
rect 15317 10284 15376 10318
rect 15410 10284 15466 10318
rect 15500 10284 15556 10318
rect 15590 10284 15646 10318
rect 15680 10284 15736 10318
rect 15770 10284 15826 10318
rect 15860 10284 15916 10318
rect 15950 10284 16011 10318
rect 15317 10276 16011 10284
rect 15317 10242 15404 10276
rect 15438 10242 15504 10276
rect 15538 10242 15604 10276
rect 15638 10242 15704 10276
rect 15738 10242 15804 10276
rect 15838 10242 15904 10276
rect 15938 10242 16011 10276
rect 15317 10228 16011 10242
rect 15317 10194 15376 10228
rect 15410 10194 15466 10228
rect 15500 10194 15556 10228
rect 15590 10194 15646 10228
rect 15680 10194 15736 10228
rect 15770 10194 15826 10228
rect 15860 10194 15916 10228
rect 15950 10194 16011 10228
rect 15317 10176 16011 10194
rect 15317 10142 15404 10176
rect 15438 10142 15504 10176
rect 15538 10142 15604 10176
rect 15638 10142 15704 10176
rect 15738 10142 15804 10176
rect 15838 10142 15904 10176
rect 15938 10142 16011 10176
rect 15317 10138 16011 10142
rect 15317 10104 15376 10138
rect 15410 10104 15466 10138
rect 15500 10104 15556 10138
rect 15590 10104 15646 10138
rect 15680 10104 15736 10138
rect 15770 10104 15826 10138
rect 15860 10104 15916 10138
rect 15950 10104 16011 10138
rect 15317 10076 16011 10104
rect 15317 10048 15404 10076
rect 15438 10048 15504 10076
rect 15317 10014 15376 10048
rect 15438 10042 15466 10048
rect 15410 10014 15466 10042
rect 15500 10042 15504 10048
rect 15538 10048 15604 10076
rect 15538 10042 15556 10048
rect 15500 10014 15556 10042
rect 15590 10042 15604 10048
rect 15638 10048 15704 10076
rect 15738 10048 15804 10076
rect 15838 10048 15904 10076
rect 15938 10048 16011 10076
rect 15638 10042 15646 10048
rect 15590 10014 15646 10042
rect 15680 10042 15704 10048
rect 15770 10042 15804 10048
rect 15860 10042 15904 10048
rect 15680 10014 15736 10042
rect 15770 10014 15826 10042
rect 15860 10014 15916 10042
rect 15950 10014 16011 10048
rect 15317 9955 16011 10014
rect 16073 10617 16092 10651
rect 16126 10650 16490 10651
rect 16126 10617 16240 10650
rect 16073 10616 16240 10617
rect 16274 10616 16341 10650
rect 16375 10636 16490 10650
rect 16524 10636 16543 10670
rect 17361 10706 17528 10711
rect 17562 10706 17629 10740
rect 17663 10730 17870 10740
rect 17904 10730 17960 10764
rect 17994 10730 18050 10764
rect 18084 10730 18140 10764
rect 18174 10730 18230 10764
rect 18264 10730 18320 10764
rect 18354 10730 18410 10764
rect 18444 10730 18500 10764
rect 18534 10730 18590 10764
rect 18624 10740 18884 10764
rect 18624 10730 18816 10740
rect 17663 10711 18816 10730
rect 17663 10706 17831 10711
rect 17361 10670 17831 10706
rect 17361 10651 17778 10670
rect 16375 10616 16543 10636
rect 16073 10580 16543 10616
rect 16073 10561 16490 10580
rect 16073 10527 16092 10561
rect 16126 10560 16490 10561
rect 16126 10527 16240 10560
rect 16073 10526 16240 10527
rect 16274 10526 16341 10560
rect 16375 10546 16490 10560
rect 16524 10546 16543 10580
rect 16375 10526 16543 10546
rect 16073 10490 16543 10526
rect 16073 10471 16490 10490
rect 16073 10437 16092 10471
rect 16126 10470 16490 10471
rect 16126 10437 16240 10470
rect 16073 10436 16240 10437
rect 16274 10436 16341 10470
rect 16375 10456 16490 10470
rect 16524 10456 16543 10490
rect 16375 10436 16543 10456
rect 16073 10400 16543 10436
rect 16073 10381 16490 10400
rect 16073 10347 16092 10381
rect 16126 10380 16490 10381
rect 16126 10347 16240 10380
rect 16073 10346 16240 10347
rect 16274 10346 16341 10380
rect 16375 10366 16490 10380
rect 16524 10366 16543 10400
rect 16375 10346 16543 10366
rect 16073 10310 16543 10346
rect 16073 10291 16490 10310
rect 16073 10257 16092 10291
rect 16126 10290 16490 10291
rect 16126 10257 16240 10290
rect 16073 10256 16240 10257
rect 16274 10256 16341 10290
rect 16375 10276 16490 10290
rect 16524 10276 16543 10310
rect 16375 10256 16543 10276
rect 16073 10220 16543 10256
rect 16073 10201 16490 10220
rect 16073 10167 16092 10201
rect 16126 10200 16490 10201
rect 16126 10167 16240 10200
rect 16073 10166 16240 10167
rect 16274 10166 16341 10200
rect 16375 10186 16490 10200
rect 16524 10186 16543 10220
rect 16375 10166 16543 10186
rect 16073 10130 16543 10166
rect 16073 10111 16490 10130
rect 16073 10077 16092 10111
rect 16126 10110 16490 10111
rect 16126 10077 16240 10110
rect 16073 10076 16240 10077
rect 16274 10076 16341 10110
rect 16375 10096 16490 10110
rect 16524 10096 16543 10130
rect 16375 10076 16543 10096
rect 16073 10040 16543 10076
rect 16073 10021 16490 10040
rect 16073 9987 16092 10021
rect 16126 10020 16490 10021
rect 16126 9987 16240 10020
rect 16073 9986 16240 9987
rect 16274 9986 16341 10020
rect 16375 10006 16490 10020
rect 16524 10006 16543 10040
rect 16375 9986 16543 10006
rect 14784 9931 15202 9950
rect 14784 9897 14804 9931
rect 14838 9930 15202 9931
rect 14838 9897 14952 9930
rect 14784 9896 14952 9897
rect 14986 9896 15053 9930
rect 15087 9916 15202 9930
rect 15236 9916 15255 9950
rect 15087 9896 15255 9916
rect 14784 9893 15255 9896
rect 16073 9950 16543 9986
rect 16605 10588 17299 10649
rect 16605 10554 16664 10588
rect 16698 10576 16754 10588
rect 16726 10554 16754 10576
rect 16788 10576 16844 10588
rect 16788 10554 16792 10576
rect 16605 10542 16692 10554
rect 16726 10542 16792 10554
rect 16826 10554 16844 10576
rect 16878 10576 16934 10588
rect 16878 10554 16892 10576
rect 16826 10542 16892 10554
rect 16926 10554 16934 10576
rect 16968 10576 17024 10588
rect 17058 10576 17114 10588
rect 17148 10576 17204 10588
rect 16968 10554 16992 10576
rect 17058 10554 17092 10576
rect 17148 10554 17192 10576
rect 17238 10554 17299 10588
rect 16926 10542 16992 10554
rect 17026 10542 17092 10554
rect 17126 10542 17192 10554
rect 17226 10542 17299 10554
rect 16605 10498 17299 10542
rect 16605 10464 16664 10498
rect 16698 10476 16754 10498
rect 16726 10464 16754 10476
rect 16788 10476 16844 10498
rect 16788 10464 16792 10476
rect 16605 10442 16692 10464
rect 16726 10442 16792 10464
rect 16826 10464 16844 10476
rect 16878 10476 16934 10498
rect 16878 10464 16892 10476
rect 16826 10442 16892 10464
rect 16926 10464 16934 10476
rect 16968 10476 17024 10498
rect 17058 10476 17114 10498
rect 17148 10476 17204 10498
rect 16968 10464 16992 10476
rect 17058 10464 17092 10476
rect 17148 10464 17192 10476
rect 17238 10464 17299 10498
rect 16926 10442 16992 10464
rect 17026 10442 17092 10464
rect 17126 10442 17192 10464
rect 17226 10442 17299 10464
rect 16605 10408 17299 10442
rect 16605 10374 16664 10408
rect 16698 10376 16754 10408
rect 16726 10374 16754 10376
rect 16788 10376 16844 10408
rect 16788 10374 16792 10376
rect 16605 10342 16692 10374
rect 16726 10342 16792 10374
rect 16826 10374 16844 10376
rect 16878 10376 16934 10408
rect 16878 10374 16892 10376
rect 16826 10342 16892 10374
rect 16926 10374 16934 10376
rect 16968 10376 17024 10408
rect 17058 10376 17114 10408
rect 17148 10376 17204 10408
rect 16968 10374 16992 10376
rect 17058 10374 17092 10376
rect 17148 10374 17192 10376
rect 17238 10374 17299 10408
rect 16926 10342 16992 10374
rect 17026 10342 17092 10374
rect 17126 10342 17192 10374
rect 17226 10342 17299 10374
rect 16605 10318 17299 10342
rect 16605 10284 16664 10318
rect 16698 10284 16754 10318
rect 16788 10284 16844 10318
rect 16878 10284 16934 10318
rect 16968 10284 17024 10318
rect 17058 10284 17114 10318
rect 17148 10284 17204 10318
rect 17238 10284 17299 10318
rect 16605 10276 17299 10284
rect 16605 10242 16692 10276
rect 16726 10242 16792 10276
rect 16826 10242 16892 10276
rect 16926 10242 16992 10276
rect 17026 10242 17092 10276
rect 17126 10242 17192 10276
rect 17226 10242 17299 10276
rect 16605 10228 17299 10242
rect 16605 10194 16664 10228
rect 16698 10194 16754 10228
rect 16788 10194 16844 10228
rect 16878 10194 16934 10228
rect 16968 10194 17024 10228
rect 17058 10194 17114 10228
rect 17148 10194 17204 10228
rect 17238 10194 17299 10228
rect 16605 10176 17299 10194
rect 16605 10142 16692 10176
rect 16726 10142 16792 10176
rect 16826 10142 16892 10176
rect 16926 10142 16992 10176
rect 17026 10142 17092 10176
rect 17126 10142 17192 10176
rect 17226 10142 17299 10176
rect 16605 10138 17299 10142
rect 16605 10104 16664 10138
rect 16698 10104 16754 10138
rect 16788 10104 16844 10138
rect 16878 10104 16934 10138
rect 16968 10104 17024 10138
rect 17058 10104 17114 10138
rect 17148 10104 17204 10138
rect 17238 10104 17299 10138
rect 16605 10076 17299 10104
rect 16605 10048 16692 10076
rect 16726 10048 16792 10076
rect 16605 10014 16664 10048
rect 16726 10042 16754 10048
rect 16698 10014 16754 10042
rect 16788 10042 16792 10048
rect 16826 10048 16892 10076
rect 16826 10042 16844 10048
rect 16788 10014 16844 10042
rect 16878 10042 16892 10048
rect 16926 10048 16992 10076
rect 17026 10048 17092 10076
rect 17126 10048 17192 10076
rect 17226 10048 17299 10076
rect 16926 10042 16934 10048
rect 16878 10014 16934 10042
rect 16968 10042 16992 10048
rect 17058 10042 17092 10048
rect 17148 10042 17192 10048
rect 16968 10014 17024 10042
rect 17058 10014 17114 10042
rect 17148 10014 17204 10042
rect 17238 10014 17299 10048
rect 16605 9955 17299 10014
rect 17361 10617 17380 10651
rect 17414 10650 17778 10651
rect 17414 10617 17528 10650
rect 17361 10616 17528 10617
rect 17562 10616 17629 10650
rect 17663 10636 17778 10650
rect 17812 10636 17831 10670
rect 18649 10706 18816 10711
rect 18850 10706 18884 10740
rect 18649 10651 18884 10706
rect 17663 10616 17831 10636
rect 17361 10580 17831 10616
rect 17361 10561 17778 10580
rect 17361 10527 17380 10561
rect 17414 10560 17778 10561
rect 17414 10527 17528 10560
rect 17361 10526 17528 10527
rect 17562 10526 17629 10560
rect 17663 10546 17778 10560
rect 17812 10546 17831 10580
rect 17663 10526 17831 10546
rect 17361 10490 17831 10526
rect 17361 10471 17778 10490
rect 17361 10437 17380 10471
rect 17414 10470 17778 10471
rect 17414 10437 17528 10470
rect 17361 10436 17528 10437
rect 17562 10436 17629 10470
rect 17663 10456 17778 10470
rect 17812 10456 17831 10490
rect 17663 10436 17831 10456
rect 17361 10400 17831 10436
rect 17361 10381 17778 10400
rect 17361 10347 17380 10381
rect 17414 10380 17778 10381
rect 17414 10347 17528 10380
rect 17361 10346 17528 10347
rect 17562 10346 17629 10380
rect 17663 10366 17778 10380
rect 17812 10366 17831 10400
rect 17663 10346 17831 10366
rect 17361 10310 17831 10346
rect 17361 10291 17778 10310
rect 17361 10257 17380 10291
rect 17414 10290 17778 10291
rect 17414 10257 17528 10290
rect 17361 10256 17528 10257
rect 17562 10256 17629 10290
rect 17663 10276 17778 10290
rect 17812 10276 17831 10310
rect 17663 10256 17831 10276
rect 17361 10220 17831 10256
rect 17361 10201 17778 10220
rect 17361 10167 17380 10201
rect 17414 10200 17778 10201
rect 17414 10167 17528 10200
rect 17361 10166 17528 10167
rect 17562 10166 17629 10200
rect 17663 10186 17778 10200
rect 17812 10186 17831 10220
rect 17663 10166 17831 10186
rect 17361 10130 17831 10166
rect 17361 10111 17778 10130
rect 17361 10077 17380 10111
rect 17414 10110 17778 10111
rect 17414 10077 17528 10110
rect 17361 10076 17528 10077
rect 17562 10076 17629 10110
rect 17663 10096 17778 10110
rect 17812 10096 17831 10130
rect 17663 10076 17831 10096
rect 17361 10040 17831 10076
rect 17361 10021 17778 10040
rect 17361 9987 17380 10021
rect 17414 10020 17778 10021
rect 17414 9987 17528 10020
rect 17361 9986 17528 9987
rect 17562 9986 17629 10020
rect 17663 10006 17778 10020
rect 17812 10006 17831 10040
rect 17663 9986 17831 10006
rect 16073 9931 16490 9950
rect 16073 9897 16092 9931
rect 16126 9930 16490 9931
rect 16126 9897 16240 9930
rect 16073 9896 16240 9897
rect 16274 9896 16341 9930
rect 16375 9916 16490 9930
rect 16524 9916 16543 9950
rect 16375 9896 16543 9916
rect 16073 9893 16543 9896
rect 17361 9950 17831 9986
rect 17893 10588 18587 10649
rect 17893 10554 17952 10588
rect 17986 10576 18042 10588
rect 18014 10554 18042 10576
rect 18076 10576 18132 10588
rect 18076 10554 18080 10576
rect 17893 10542 17980 10554
rect 18014 10542 18080 10554
rect 18114 10554 18132 10576
rect 18166 10576 18222 10588
rect 18166 10554 18180 10576
rect 18114 10542 18180 10554
rect 18214 10554 18222 10576
rect 18256 10576 18312 10588
rect 18346 10576 18402 10588
rect 18436 10576 18492 10588
rect 18256 10554 18280 10576
rect 18346 10554 18380 10576
rect 18436 10554 18480 10576
rect 18526 10554 18587 10588
rect 18214 10542 18280 10554
rect 18314 10542 18380 10554
rect 18414 10542 18480 10554
rect 18514 10542 18587 10554
rect 17893 10498 18587 10542
rect 17893 10464 17952 10498
rect 17986 10476 18042 10498
rect 18014 10464 18042 10476
rect 18076 10476 18132 10498
rect 18076 10464 18080 10476
rect 17893 10442 17980 10464
rect 18014 10442 18080 10464
rect 18114 10464 18132 10476
rect 18166 10476 18222 10498
rect 18166 10464 18180 10476
rect 18114 10442 18180 10464
rect 18214 10464 18222 10476
rect 18256 10476 18312 10498
rect 18346 10476 18402 10498
rect 18436 10476 18492 10498
rect 18256 10464 18280 10476
rect 18346 10464 18380 10476
rect 18436 10464 18480 10476
rect 18526 10464 18587 10498
rect 18214 10442 18280 10464
rect 18314 10442 18380 10464
rect 18414 10442 18480 10464
rect 18514 10442 18587 10464
rect 17893 10408 18587 10442
rect 17893 10374 17952 10408
rect 17986 10376 18042 10408
rect 18014 10374 18042 10376
rect 18076 10376 18132 10408
rect 18076 10374 18080 10376
rect 17893 10342 17980 10374
rect 18014 10342 18080 10374
rect 18114 10374 18132 10376
rect 18166 10376 18222 10408
rect 18166 10374 18180 10376
rect 18114 10342 18180 10374
rect 18214 10374 18222 10376
rect 18256 10376 18312 10408
rect 18346 10376 18402 10408
rect 18436 10376 18492 10408
rect 18256 10374 18280 10376
rect 18346 10374 18380 10376
rect 18436 10374 18480 10376
rect 18526 10374 18587 10408
rect 18214 10342 18280 10374
rect 18314 10342 18380 10374
rect 18414 10342 18480 10374
rect 18514 10342 18587 10374
rect 17893 10318 18587 10342
rect 17893 10284 17952 10318
rect 17986 10284 18042 10318
rect 18076 10284 18132 10318
rect 18166 10284 18222 10318
rect 18256 10284 18312 10318
rect 18346 10284 18402 10318
rect 18436 10284 18492 10318
rect 18526 10284 18587 10318
rect 17893 10276 18587 10284
rect 17893 10242 17980 10276
rect 18014 10242 18080 10276
rect 18114 10242 18180 10276
rect 18214 10242 18280 10276
rect 18314 10242 18380 10276
rect 18414 10242 18480 10276
rect 18514 10242 18587 10276
rect 17893 10228 18587 10242
rect 17893 10194 17952 10228
rect 17986 10194 18042 10228
rect 18076 10194 18132 10228
rect 18166 10194 18222 10228
rect 18256 10194 18312 10228
rect 18346 10194 18402 10228
rect 18436 10194 18492 10228
rect 18526 10194 18587 10228
rect 17893 10176 18587 10194
rect 17893 10142 17980 10176
rect 18014 10142 18080 10176
rect 18114 10142 18180 10176
rect 18214 10142 18280 10176
rect 18314 10142 18380 10176
rect 18414 10142 18480 10176
rect 18514 10142 18587 10176
rect 17893 10138 18587 10142
rect 17893 10104 17952 10138
rect 17986 10104 18042 10138
rect 18076 10104 18132 10138
rect 18166 10104 18222 10138
rect 18256 10104 18312 10138
rect 18346 10104 18402 10138
rect 18436 10104 18492 10138
rect 18526 10104 18587 10138
rect 17893 10076 18587 10104
rect 17893 10048 17980 10076
rect 18014 10048 18080 10076
rect 17893 10014 17952 10048
rect 18014 10042 18042 10048
rect 17986 10014 18042 10042
rect 18076 10042 18080 10048
rect 18114 10048 18180 10076
rect 18114 10042 18132 10048
rect 18076 10014 18132 10042
rect 18166 10042 18180 10048
rect 18214 10048 18280 10076
rect 18314 10048 18380 10076
rect 18414 10048 18480 10076
rect 18514 10048 18587 10076
rect 18214 10042 18222 10048
rect 18166 10014 18222 10042
rect 18256 10042 18280 10048
rect 18346 10042 18380 10048
rect 18436 10042 18480 10048
rect 18256 10014 18312 10042
rect 18346 10014 18402 10042
rect 18436 10014 18492 10042
rect 18526 10014 18587 10048
rect 17893 9955 18587 10014
rect 18649 10617 18668 10651
rect 18702 10650 18884 10651
rect 18702 10617 18816 10650
rect 18649 10616 18816 10617
rect 18850 10616 18884 10650
rect 18649 10561 18884 10616
rect 18649 10527 18668 10561
rect 18702 10560 18884 10561
rect 18702 10527 18816 10560
rect 18649 10526 18816 10527
rect 18850 10526 18884 10560
rect 18649 10471 18884 10526
rect 18649 10437 18668 10471
rect 18702 10470 18884 10471
rect 18702 10437 18816 10470
rect 18649 10436 18816 10437
rect 18850 10436 18884 10470
rect 18649 10381 18884 10436
rect 18649 10347 18668 10381
rect 18702 10380 18884 10381
rect 18702 10347 18816 10380
rect 18649 10346 18816 10347
rect 18850 10346 18884 10380
rect 18649 10291 18884 10346
rect 18649 10257 18668 10291
rect 18702 10290 18884 10291
rect 18702 10257 18816 10290
rect 18649 10256 18816 10257
rect 18850 10256 18884 10290
rect 18649 10201 18884 10256
rect 18649 10167 18668 10201
rect 18702 10200 18884 10201
rect 18702 10167 18816 10200
rect 18649 10166 18816 10167
rect 18850 10166 18884 10200
rect 18649 10111 18884 10166
rect 18649 10077 18668 10111
rect 18702 10110 18884 10111
rect 18702 10077 18816 10110
rect 18649 10076 18816 10077
rect 18850 10076 18884 10110
rect 18649 10021 18884 10076
rect 18649 9987 18668 10021
rect 18702 10020 18884 10021
rect 18702 9987 18816 10020
rect 18649 9986 18816 9987
rect 18850 9986 18884 10020
rect 17361 9931 17778 9950
rect 17361 9897 17380 9931
rect 17414 9930 17778 9931
rect 17414 9897 17528 9930
rect 17361 9896 17528 9897
rect 17562 9896 17629 9930
rect 17663 9916 17778 9930
rect 17812 9916 17831 9950
rect 17663 9896 17831 9916
rect 17361 9893 17831 9896
rect 18649 9931 18884 9986
rect 18649 9897 18668 9931
rect 18702 9930 18884 9931
rect 18702 9897 18816 9930
rect 18649 9896 18816 9897
rect 18850 9896 18884 9930
rect 18649 9893 18884 9896
rect 12444 9874 18884 9893
rect 12444 9840 12684 9874
rect 12718 9840 12774 9874
rect 12808 9840 12864 9874
rect 12898 9840 12954 9874
rect 12988 9840 13044 9874
rect 13078 9840 13134 9874
rect 13168 9840 13224 9874
rect 13258 9840 13314 9874
rect 13348 9840 13404 9874
rect 13438 9840 13972 9874
rect 14006 9840 14062 9874
rect 14096 9840 14152 9874
rect 14186 9840 14242 9874
rect 14276 9840 14332 9874
rect 14366 9840 14422 9874
rect 14456 9840 14512 9874
rect 14546 9840 14602 9874
rect 14636 9840 14692 9874
rect 14726 9840 15260 9874
rect 15294 9840 15350 9874
rect 15384 9840 15440 9874
rect 15474 9840 15530 9874
rect 15564 9840 15620 9874
rect 15654 9840 15710 9874
rect 15744 9840 15800 9874
rect 15834 9840 15890 9874
rect 15924 9840 15980 9874
rect 16014 9840 16548 9874
rect 16582 9840 16638 9874
rect 16672 9840 16728 9874
rect 16762 9840 16818 9874
rect 16852 9840 16908 9874
rect 16942 9840 16998 9874
rect 17032 9840 17088 9874
rect 17122 9840 17178 9874
rect 17212 9840 17268 9874
rect 17302 9840 17836 9874
rect 17870 9840 17926 9874
rect 17960 9840 18016 9874
rect 18050 9840 18106 9874
rect 18140 9840 18196 9874
rect 18230 9840 18286 9874
rect 18320 9840 18376 9874
rect 18410 9840 18466 9874
rect 18500 9840 18556 9874
rect 18590 9840 18884 9874
rect 12444 9806 12477 9840
rect 12511 9821 13664 9840
rect 12511 9806 12684 9821
rect 12444 9757 12684 9806
rect 13484 9806 13664 9821
rect 13698 9806 13765 9840
rect 13799 9821 14952 9840
rect 13799 9806 13984 9821
rect 13484 9757 13984 9806
rect 14784 9806 14952 9821
rect 14986 9806 15053 9840
rect 15087 9821 16240 9840
rect 15087 9806 15184 9821
rect 14784 9757 15184 9806
rect 16084 9806 16240 9821
rect 16274 9806 16341 9840
rect 16375 9821 17528 9840
rect 16375 9806 16484 9821
rect 16084 9757 16484 9806
rect 17384 9806 17528 9821
rect 17562 9806 17629 9840
rect 17663 9821 18816 9840
rect 17663 9806 17784 9821
rect 17384 9757 17784 9806
rect 18684 9806 18816 9821
rect 18850 9806 18884 9840
rect 18684 9757 18884 9806
rect 12444 9750 18884 9757
rect 12444 9716 12477 9750
rect 12511 9727 13664 9750
rect 12511 9716 12578 9727
rect 12444 9693 12578 9716
rect 12612 9693 12668 9727
rect 12702 9693 12758 9727
rect 12792 9693 12848 9727
rect 12882 9693 12938 9727
rect 12972 9693 13028 9727
rect 13062 9693 13118 9727
rect 13152 9693 13208 9727
rect 13242 9693 13298 9727
rect 13332 9693 13388 9727
rect 13422 9693 13478 9727
rect 13512 9693 13568 9727
rect 13602 9716 13664 9727
rect 13698 9716 13765 9750
rect 13799 9727 14952 9750
rect 13799 9716 13866 9727
rect 13602 9693 13866 9716
rect 13900 9693 13956 9727
rect 13990 9693 14046 9727
rect 14080 9693 14136 9727
rect 14170 9693 14226 9727
rect 14260 9693 14316 9727
rect 14350 9693 14406 9727
rect 14440 9693 14496 9727
rect 14530 9693 14586 9727
rect 14620 9693 14676 9727
rect 14710 9693 14766 9727
rect 14800 9693 14856 9727
rect 14890 9716 14952 9727
rect 14986 9716 15053 9750
rect 15087 9727 16240 9750
rect 15087 9716 15154 9727
rect 14890 9693 15154 9716
rect 15188 9693 15244 9727
rect 15278 9693 15334 9727
rect 15368 9693 15424 9727
rect 15458 9693 15514 9727
rect 15548 9693 15604 9727
rect 15638 9693 15694 9727
rect 15728 9693 15784 9727
rect 15818 9693 15874 9727
rect 15908 9693 15964 9727
rect 15998 9693 16054 9727
rect 16088 9693 16144 9727
rect 16178 9716 16240 9727
rect 16274 9716 16341 9750
rect 16375 9727 17528 9750
rect 16375 9716 16442 9727
rect 16178 9693 16442 9716
rect 16476 9693 16532 9727
rect 16566 9693 16622 9727
rect 16656 9693 16712 9727
rect 16746 9693 16802 9727
rect 16836 9693 16892 9727
rect 16926 9693 16982 9727
rect 17016 9693 17072 9727
rect 17106 9693 17162 9727
rect 17196 9693 17252 9727
rect 17286 9693 17342 9727
rect 17376 9693 17432 9727
rect 17466 9716 17528 9727
rect 17562 9716 17629 9750
rect 17663 9727 18816 9750
rect 17663 9716 17730 9727
rect 17466 9693 17730 9716
rect 17764 9693 17820 9727
rect 17854 9693 17910 9727
rect 17944 9693 18000 9727
rect 18034 9693 18090 9727
rect 18124 9693 18180 9727
rect 18214 9693 18270 9727
rect 18304 9693 18360 9727
rect 18394 9693 18450 9727
rect 18484 9693 18540 9727
rect 18574 9693 18630 9727
rect 18664 9693 18720 9727
rect 18754 9716 18816 9727
rect 18850 9716 18884 9750
rect 18754 9693 18884 9716
rect 12444 9626 18884 9693
rect 12444 9592 12578 9626
rect 12612 9592 12668 9626
rect 12702 9592 12758 9626
rect 12792 9592 12848 9626
rect 12882 9592 12938 9626
rect 12972 9592 13028 9626
rect 13062 9592 13118 9626
rect 13152 9592 13208 9626
rect 13242 9592 13298 9626
rect 13332 9592 13388 9626
rect 13422 9592 13478 9626
rect 13512 9592 13568 9626
rect 13602 9592 13866 9626
rect 13900 9592 13956 9626
rect 13990 9592 14046 9626
rect 14080 9592 14136 9626
rect 14170 9592 14226 9626
rect 14260 9592 14316 9626
rect 14350 9592 14406 9626
rect 14440 9592 14496 9626
rect 14530 9592 14586 9626
rect 14620 9592 14676 9626
rect 14710 9592 14766 9626
rect 14800 9592 14856 9626
rect 14890 9592 15154 9626
rect 15188 9592 15244 9626
rect 15278 9592 15334 9626
rect 15368 9592 15424 9626
rect 15458 9592 15514 9626
rect 15548 9592 15604 9626
rect 15638 9592 15694 9626
rect 15728 9592 15784 9626
rect 15818 9592 15874 9626
rect 15908 9592 15964 9626
rect 15998 9592 16054 9626
rect 16088 9592 16144 9626
rect 16178 9592 16442 9626
rect 16476 9592 16532 9626
rect 16566 9592 16622 9626
rect 16656 9592 16712 9626
rect 16746 9592 16802 9626
rect 16836 9592 16892 9626
rect 16926 9592 16982 9626
rect 17016 9592 17072 9626
rect 17106 9592 17162 9626
rect 17196 9592 17252 9626
rect 17286 9592 17342 9626
rect 17376 9592 17432 9626
rect 17466 9592 17730 9626
rect 17764 9592 17820 9626
rect 17854 9592 17910 9626
rect 17944 9592 18000 9626
rect 18034 9592 18090 9626
rect 18124 9592 18180 9626
rect 18214 9592 18270 9626
rect 18304 9592 18360 9626
rect 18394 9592 18450 9626
rect 18484 9592 18540 9626
rect 18574 9592 18630 9626
rect 18664 9592 18720 9626
rect 18754 9592 18884 9626
rect 12444 9559 18884 9592
rect 12444 9542 12684 9559
rect 12444 9508 12477 9542
rect 12511 9508 12684 9542
rect 12444 9495 12684 9508
rect 13484 9542 13984 9559
rect 13484 9508 13664 9542
rect 13698 9508 13765 9542
rect 13799 9508 13984 9542
rect 13484 9495 13984 9508
rect 14784 9542 15184 9559
rect 14784 9508 14952 9542
rect 14986 9508 15053 9542
rect 15087 9508 15184 9542
rect 14784 9495 15184 9508
rect 16084 9542 16484 9559
rect 16084 9508 16240 9542
rect 16274 9508 16341 9542
rect 16375 9508 16484 9542
rect 16084 9495 16484 9508
rect 17384 9542 17784 9559
rect 17384 9508 17528 9542
rect 17562 9508 17629 9542
rect 17663 9508 17784 9542
rect 17384 9495 17784 9508
rect 18684 9542 18884 9559
rect 18684 9508 18816 9542
rect 18850 9508 18884 9542
rect 18684 9495 18884 9508
rect 12444 9476 18884 9495
rect 12444 9452 12718 9476
rect -8800 9428 -8766 9444
rect -17898 9388 -11414 9398
rect -17898 9044 -17888 9388
rect -11424 9044 -11414 9388
rect -17898 9034 -11414 9044
rect -9500 9102 -8900 9302
rect -17180 8818 -17164 8852
rect -11788 8818 -11772 8852
rect -17248 8790 -17214 8806
rect -17248 8406 -17214 8422
rect -17180 8360 -17164 8394
rect -11788 8360 -11772 8394
rect -16836 6692 -16820 6726
rect -16452 6692 -16436 6726
rect -16264 6692 -16248 6726
rect -15880 6692 -15864 6726
rect -15692 6692 -15676 6726
rect -15308 6692 -15292 6726
rect -15120 6692 -15104 6726
rect -14736 6692 -14720 6726
rect -14548 6692 -14532 6726
rect -14164 6692 -14148 6726
rect -13976 6692 -13960 6726
rect -13592 6692 -13576 6726
rect -13404 6692 -13388 6726
rect -13020 6692 -13004 6726
rect -12832 6692 -12816 6726
rect -12448 6692 -12432 6726
rect -17450 6642 -17318 6658
rect -20934 5836 -19910 5852
rect -20934 5760 -20918 5836
rect -19926 5760 -19910 5836
rect -20934 5720 -19910 5760
rect -22320 5682 -21888 5698
rect -22320 5106 -22304 5682
rect -21904 5604 -21888 5682
rect -20934 5668 -20906 5720
rect -20854 5668 -19990 5720
rect -19938 5668 -19910 5720
rect -20934 5656 -19910 5668
rect -18954 5682 -18522 5698
rect -18954 5604 -18938 5682
rect -21904 5570 -21750 5604
rect -21382 5570 -21366 5604
rect -21308 5570 -21292 5604
rect -20924 5570 -20834 5604
rect -20466 5570 -20376 5604
rect -20008 5570 -19918 5604
rect -19550 5570 -19534 5604
rect -19476 5570 -19460 5604
rect -19092 5570 -18938 5604
rect -21904 5520 -21778 5570
rect -21904 5144 -21812 5520
rect -21904 5128 -21778 5144
rect -21354 5520 -21320 5536
rect -21354 5128 -21320 5144
rect -20896 5520 -20862 5536
rect -20896 5128 -20862 5144
rect -20438 5520 -20404 5536
rect -20438 5128 -20404 5144
rect -19980 5520 -19946 5536
rect -19980 5128 -19946 5144
rect -19522 5520 -19488 5536
rect -19522 5128 -19488 5144
rect -19064 5520 -18938 5570
rect -19030 5144 -18938 5520
rect -19064 5128 -18938 5144
rect -21904 5106 -21888 5128
rect -22320 5090 -21888 5106
rect -18954 5106 -18938 5128
rect -18538 5106 -18522 5682
rect -18954 5090 -18522 5106
rect -17450 5042 -17434 6642
rect -17334 5042 -17318 6642
rect -17450 5026 -17318 5042
rect -16882 6642 -16848 6658
rect -16882 4850 -16848 4866
rect -16424 6642 -16390 6658
rect -16424 4850 -16390 4866
rect -16310 6642 -16276 6658
rect -16310 4850 -16276 4866
rect -15852 6642 -15818 6658
rect -15852 4850 -15818 4866
rect -15738 6642 -15704 6658
rect -15738 4850 -15704 4866
rect -15280 6642 -15246 6658
rect -15280 4850 -15246 4866
rect -15166 6642 -15132 6658
rect -15166 4850 -15132 4866
rect -14708 6642 -14674 6658
rect -14708 4850 -14674 4866
rect -14594 6642 -14560 6658
rect -14594 4850 -14560 4866
rect -14136 6642 -14102 6658
rect -14136 4850 -14102 4866
rect -14022 6642 -13988 6658
rect -14022 4850 -13988 4866
rect -13564 6642 -13530 6658
rect -13564 4850 -13530 4866
rect -13450 6642 -13416 6658
rect -13450 4850 -13416 4866
rect -12992 6642 -12958 6658
rect -12992 4850 -12958 4866
rect -12878 6642 -12844 6658
rect -12878 4850 -12844 4866
rect -12420 6642 -12386 6658
rect -11950 6642 -11818 6658
rect -11950 5042 -11934 6642
rect -11834 5042 -11818 6642
rect -11950 5026 -11818 5042
rect -12420 4850 -12386 4866
rect -18562 4289 -18546 4323
rect -18178 4289 -18162 4323
rect -17990 4289 -17974 4323
rect -17606 4289 -17590 4323
rect -17418 4289 -17402 4323
rect -17034 4289 -17018 4323
rect -16846 4289 -16830 4323
rect -16462 4289 -16446 4323
rect -16274 4289 -16258 4323
rect -15890 4289 -15874 4323
rect -15702 4289 -15686 4323
rect -15318 4289 -15302 4323
rect -15130 4289 -15114 4323
rect -14746 4289 -14730 4323
rect -14558 4289 -14542 4323
rect -14174 4289 -14158 4323
rect -13986 4289 -13970 4323
rect -13602 4289 -13586 4323
rect -13414 4289 -13398 4323
rect -13030 4289 -13014 4323
rect -12842 4289 -12826 4323
rect -12458 4289 -12442 4323
rect -12270 4289 -12254 4323
rect -11886 4289 -11870 4323
rect -11698 4289 -11682 4323
rect -11314 4289 -11298 4323
rect -11126 4289 -11110 4323
rect -10742 4289 -10726 4323
rect -18608 4230 -18574 4246
rect -19266 4142 -19134 4154
rect -19266 1800 -19250 4142
rect -19150 1800 -19134 4142
rect -19266 1784 -19134 1800
rect -18608 1658 -18574 1674
rect -18150 4230 -18116 4246
rect -18150 1658 -18116 1674
rect -18036 4230 -18002 4246
rect -18036 1658 -18002 1674
rect -17578 4230 -17544 4246
rect -17578 1658 -17544 1674
rect -17464 4230 -17430 4246
rect -17464 1658 -17430 1674
rect -17006 4230 -16972 4246
rect -17006 1658 -16972 1674
rect -16892 4230 -16858 4246
rect -16892 1658 -16858 1674
rect -16434 4230 -16400 4246
rect -16434 1658 -16400 1674
rect -16320 4230 -16286 4246
rect -16320 1658 -16286 1674
rect -15862 4230 -15828 4246
rect -15862 1658 -15828 1674
rect -15748 4230 -15714 4246
rect -15748 1658 -15714 1674
rect -15290 4230 -15256 4246
rect -15290 1658 -15256 1674
rect -15176 4230 -15142 4246
rect -15176 1658 -15142 1674
rect -14718 4230 -14684 4246
rect -14718 1658 -14684 1674
rect -14604 4230 -14570 4246
rect -14604 1658 -14570 1674
rect -14146 4230 -14112 4246
rect -14146 1658 -14112 1674
rect -14032 4230 -13998 4246
rect -14032 1658 -13998 1674
rect -13574 4230 -13540 4246
rect -13574 1658 -13540 1674
rect -13460 4230 -13426 4246
rect -13460 1658 -13426 1674
rect -13002 4230 -12968 4246
rect -13002 1658 -12968 1674
rect -12888 4230 -12854 4246
rect -12888 1658 -12854 1674
rect -12430 4230 -12396 4246
rect -12430 1658 -12396 1674
rect -12316 4230 -12282 4246
rect -12316 1658 -12282 1674
rect -11858 4230 -11824 4246
rect -11858 1658 -11824 1674
rect -11744 4230 -11710 4246
rect -11744 1658 -11710 1674
rect -11286 4230 -11252 4246
rect -11286 1658 -11252 1674
rect -11172 4230 -11138 4246
rect -11172 1658 -11138 1674
rect -10714 4230 -10680 4246
rect -10138 4142 -10006 4154
rect -10138 1800 -10122 4142
rect -10022 1800 -10006 4142
rect -10138 1784 -10006 1800
rect -9500 2102 -9300 9102
rect -9100 2102 -8900 9102
rect -10714 1658 -10680 1674
rect -15680 1296 -13310 1312
rect -15680 1196 -15668 1296
rect -13326 1196 -13310 1296
rect -15680 1180 -13310 1196
rect -9500 1202 -8900 2102
rect -8800 1696 -8766 1712
rect -8342 9428 -8308 9444
rect -8342 1696 -8308 1712
rect -7884 9428 -7850 9444
rect -7884 1696 -7850 1712
rect -7426 9428 -7392 9444
rect -7426 1696 -7392 1712
rect -6968 9428 -6934 9444
rect -6968 1696 -6934 1712
rect -6510 9428 -6476 9444
rect -6510 1696 -6476 1712
rect -6052 9428 -6018 9444
rect -6052 1696 -6018 1712
rect -5594 9428 -5560 9444
rect -5594 1696 -5560 1712
rect -5136 9428 -5102 9444
rect -5136 1696 -5102 1712
rect -4678 9428 -4644 9444
rect -4678 1696 -4644 1712
rect -4220 9428 -4186 9444
rect -4220 1696 -4186 1712
rect -3762 9428 -3728 9444
rect -2842 9428 -2808 9444
rect -3762 1696 -3728 1712
rect -3590 9102 -2990 9302
rect -3590 2102 -3390 9102
rect -3190 2102 -2990 9102
rect -8754 1619 -8738 1653
rect -8370 1619 -8354 1653
rect -8296 1619 -8280 1653
rect -7912 1619 -7896 1653
rect -7838 1619 -7822 1653
rect -7454 1619 -7438 1653
rect -7380 1619 -7364 1653
rect -6996 1619 -6980 1653
rect -6922 1619 -6906 1653
rect -6538 1619 -6522 1653
rect -6464 1619 -6448 1653
rect -6080 1619 -6064 1653
rect -6006 1619 -5990 1653
rect -5622 1619 -5606 1653
rect -5548 1619 -5532 1653
rect -5164 1619 -5148 1653
rect -5090 1619 -5074 1653
rect -4706 1619 -4690 1653
rect -4632 1619 -4616 1653
rect -4248 1619 -4232 1653
rect -4174 1619 -4158 1653
rect -3790 1619 -3774 1653
rect -9500 1102 -9400 1202
rect -9000 1102 -8900 1202
rect -9500 1002 -8900 1102
rect -3590 1202 -2990 2102
rect -2842 1696 -2808 1712
rect -2384 9428 -2350 9444
rect -2384 1696 -2350 1712
rect -1926 9428 -1892 9444
rect -1926 1696 -1892 1712
rect -1468 9428 -1434 9444
rect -1468 1696 -1434 1712
rect -1010 9428 -976 9444
rect -1010 1696 -976 1712
rect -552 9428 -518 9444
rect -552 1696 -518 1712
rect -94 9428 -60 9444
rect -94 1696 -60 1712
rect 364 9428 398 9444
rect 364 1696 398 1712
rect 822 9428 856 9444
rect 822 1696 856 1712
rect 1280 9428 1314 9444
rect 1280 1696 1314 1712
rect 1738 9428 1772 9444
rect 2658 9428 2692 9444
rect 1738 1696 1772 1712
rect 1910 9102 2510 9302
rect 1910 2102 2110 9102
rect 2310 2102 2510 9102
rect -2796 1619 -2780 1653
rect -2412 1619 -2396 1653
rect -2338 1619 -2322 1653
rect -1954 1619 -1938 1653
rect -1880 1619 -1864 1653
rect -1496 1619 -1480 1653
rect -1422 1619 -1406 1653
rect -1038 1619 -1022 1653
rect -964 1619 -948 1653
rect -580 1619 -564 1653
rect -506 1619 -490 1653
rect -122 1619 -106 1653
rect -48 1619 -32 1653
rect 336 1619 352 1653
rect 410 1619 426 1653
rect 794 1619 810 1653
rect 868 1619 884 1653
rect 1252 1619 1268 1653
rect 1326 1619 1342 1653
rect 1710 1619 1726 1653
rect -3590 1102 -3490 1202
rect -3090 1102 -2990 1202
rect -3590 1002 -2990 1102
rect 1910 1202 2510 2102
rect 2658 1696 2692 1712
rect 3116 9428 3150 9444
rect 3116 1696 3150 1712
rect 3574 9428 3608 9444
rect 3574 1696 3608 1712
rect 4032 9428 4066 9444
rect 4032 1696 4066 1712
rect 4490 9428 4524 9444
rect 4490 1696 4524 1712
rect 4948 9428 4982 9444
rect 4948 1696 4982 1712
rect 5406 9428 5440 9444
rect 5406 1696 5440 1712
rect 5864 9428 5898 9444
rect 5864 1696 5898 1712
rect 6322 9428 6356 9444
rect 6322 1696 6356 1712
rect 6780 9428 6814 9444
rect 6780 1696 6814 1712
rect 7238 9428 7272 9444
rect 7238 1696 7272 1712
rect 7696 9428 7730 9444
rect 12444 9418 12477 9452
rect 12511 9442 12718 9452
rect 12752 9442 12808 9476
rect 12842 9442 12898 9476
rect 12932 9442 12988 9476
rect 13022 9442 13078 9476
rect 13112 9442 13168 9476
rect 13202 9442 13258 9476
rect 13292 9442 13348 9476
rect 13382 9442 13438 9476
rect 13472 9452 14006 9476
rect 13472 9442 13664 9452
rect 12511 9423 13664 9442
rect 12511 9418 12684 9423
rect 12444 9382 12684 9418
rect 12444 9362 12626 9382
rect 12444 9328 12477 9362
rect 12511 9348 12626 9362
rect 12660 9348 12684 9382
rect 13484 9418 13664 9423
rect 13698 9418 13765 9452
rect 13799 9442 14006 9452
rect 14040 9442 14096 9476
rect 14130 9442 14186 9476
rect 14220 9442 14276 9476
rect 14310 9442 14366 9476
rect 14400 9442 14456 9476
rect 14490 9442 14546 9476
rect 14580 9442 14636 9476
rect 14670 9442 14726 9476
rect 14760 9452 15294 9476
rect 14760 9442 14952 9452
rect 13799 9423 14952 9442
rect 13799 9418 13984 9423
rect 13484 9382 13984 9418
rect 13484 9363 13914 9382
rect 12511 9328 12684 9348
rect 7696 1696 7730 1712
rect 7866 9100 8466 9300
rect 7866 2100 8066 9100
rect 8266 2100 8466 9100
rect 2704 1619 2720 1653
rect 3088 1619 3104 1653
rect 3162 1619 3178 1653
rect 3546 1619 3562 1653
rect 3620 1619 3636 1653
rect 4004 1619 4020 1653
rect 4078 1619 4094 1653
rect 4462 1619 4478 1653
rect 4536 1619 4552 1653
rect 4920 1619 4936 1653
rect 4994 1619 5010 1653
rect 5378 1619 5394 1653
rect 5452 1619 5468 1653
rect 5836 1619 5852 1653
rect 5910 1619 5926 1653
rect 6294 1619 6310 1653
rect 6368 1619 6384 1653
rect 6752 1619 6768 1653
rect 6826 1619 6842 1653
rect 7210 1619 7226 1653
rect 7284 1619 7300 1653
rect 7668 1619 7684 1653
rect 1910 1102 2010 1202
rect 2410 1102 2510 1202
rect 1910 1002 2510 1102
rect 7866 1200 8466 2100
rect 12444 9292 12684 9328
rect 12444 9272 12626 9292
rect 12444 9238 12477 9272
rect 12511 9258 12626 9272
rect 12660 9258 12684 9292
rect 12511 9238 12684 9258
rect 12444 9202 12684 9238
rect 12444 9182 12626 9202
rect 12444 9148 12477 9182
rect 12511 9168 12626 9182
rect 12660 9168 12684 9202
rect 12511 9148 12684 9168
rect 12444 9112 12684 9148
rect 12444 9092 12626 9112
rect 12444 9058 12477 9092
rect 12511 9078 12626 9092
rect 12660 9078 12684 9112
rect 12511 9058 12684 9078
rect 12444 9022 12684 9058
rect 12444 9002 12626 9022
rect 12444 8968 12477 9002
rect 12511 8988 12626 9002
rect 12660 8988 12684 9022
rect 12511 8968 12684 8988
rect 12444 8932 12684 8968
rect 12444 8912 12626 8932
rect 12444 8878 12477 8912
rect 12511 8898 12626 8912
rect 12660 8898 12684 8932
rect 12511 8878 12684 8898
rect 12444 8842 12684 8878
rect 12444 8822 12626 8842
rect 12444 8788 12477 8822
rect 12511 8808 12626 8822
rect 12660 8808 12684 8842
rect 12511 8788 12684 8808
rect 12444 8752 12684 8788
rect 12444 8732 12626 8752
rect 12444 8698 12477 8732
rect 12511 8718 12626 8732
rect 12660 8718 12684 8752
rect 12511 8698 12684 8718
rect 12444 8662 12684 8698
rect 12741 9300 13435 9361
rect 12741 9266 12800 9300
rect 12834 9288 12890 9300
rect 12862 9266 12890 9288
rect 12924 9288 12980 9300
rect 12924 9266 12928 9288
rect 12741 9254 12828 9266
rect 12862 9254 12928 9266
rect 12962 9266 12980 9288
rect 13014 9288 13070 9300
rect 13014 9266 13028 9288
rect 12962 9254 13028 9266
rect 13062 9266 13070 9288
rect 13104 9288 13160 9300
rect 13194 9288 13250 9300
rect 13284 9288 13340 9300
rect 13104 9266 13128 9288
rect 13194 9266 13228 9288
rect 13284 9266 13328 9288
rect 13374 9266 13435 9300
rect 13062 9254 13128 9266
rect 13162 9254 13228 9266
rect 13262 9254 13328 9266
rect 13362 9254 13435 9266
rect 12741 9210 13435 9254
rect 12741 9176 12800 9210
rect 12834 9188 12890 9210
rect 12862 9176 12890 9188
rect 12924 9188 12980 9210
rect 12924 9176 12928 9188
rect 12741 9154 12828 9176
rect 12862 9154 12928 9176
rect 12962 9176 12980 9188
rect 13014 9188 13070 9210
rect 13014 9176 13028 9188
rect 12962 9154 13028 9176
rect 13062 9176 13070 9188
rect 13104 9188 13160 9210
rect 13194 9188 13250 9210
rect 13284 9188 13340 9210
rect 13104 9176 13128 9188
rect 13194 9176 13228 9188
rect 13284 9176 13328 9188
rect 13374 9176 13435 9210
rect 13062 9154 13128 9176
rect 13162 9154 13228 9176
rect 13262 9154 13328 9176
rect 13362 9154 13435 9176
rect 12741 9120 13435 9154
rect 12741 9086 12800 9120
rect 12834 9088 12890 9120
rect 12862 9086 12890 9088
rect 12924 9088 12980 9120
rect 12924 9086 12928 9088
rect 12741 9054 12828 9086
rect 12862 9054 12928 9086
rect 12962 9086 12980 9088
rect 13014 9088 13070 9120
rect 13014 9086 13028 9088
rect 12962 9054 13028 9086
rect 13062 9086 13070 9088
rect 13104 9088 13160 9120
rect 13194 9088 13250 9120
rect 13284 9088 13340 9120
rect 13104 9086 13128 9088
rect 13194 9086 13228 9088
rect 13284 9086 13328 9088
rect 13374 9086 13435 9120
rect 13062 9054 13128 9086
rect 13162 9054 13228 9086
rect 13262 9054 13328 9086
rect 13362 9054 13435 9086
rect 12741 9030 13435 9054
rect 12741 8996 12800 9030
rect 12834 8996 12890 9030
rect 12924 8996 12980 9030
rect 13014 8996 13070 9030
rect 13104 8996 13160 9030
rect 13194 8996 13250 9030
rect 13284 8996 13340 9030
rect 13374 8996 13435 9030
rect 12741 8988 13435 8996
rect 12741 8954 12828 8988
rect 12862 8954 12928 8988
rect 12962 8954 13028 8988
rect 13062 8954 13128 8988
rect 13162 8954 13228 8988
rect 13262 8954 13328 8988
rect 13362 8954 13435 8988
rect 12741 8940 13435 8954
rect 12741 8906 12800 8940
rect 12834 8906 12890 8940
rect 12924 8906 12980 8940
rect 13014 8906 13070 8940
rect 13104 8906 13160 8940
rect 13194 8906 13250 8940
rect 13284 8906 13340 8940
rect 13374 8906 13435 8940
rect 12741 8888 13435 8906
rect 12741 8854 12828 8888
rect 12862 8854 12928 8888
rect 12962 8854 13028 8888
rect 13062 8854 13128 8888
rect 13162 8854 13228 8888
rect 13262 8854 13328 8888
rect 13362 8854 13435 8888
rect 12741 8850 13435 8854
rect 12741 8816 12800 8850
rect 12834 8816 12890 8850
rect 12924 8816 12980 8850
rect 13014 8816 13070 8850
rect 13104 8816 13160 8850
rect 13194 8816 13250 8850
rect 13284 8816 13340 8850
rect 13374 8816 13435 8850
rect 12741 8788 13435 8816
rect 12741 8760 12828 8788
rect 12862 8760 12928 8788
rect 12741 8726 12800 8760
rect 12862 8754 12890 8760
rect 12834 8726 12890 8754
rect 12924 8754 12928 8760
rect 12962 8760 13028 8788
rect 12962 8754 12980 8760
rect 12924 8726 12980 8754
rect 13014 8754 13028 8760
rect 13062 8760 13128 8788
rect 13162 8760 13228 8788
rect 13262 8760 13328 8788
rect 13362 8760 13435 8788
rect 13062 8754 13070 8760
rect 13014 8726 13070 8754
rect 13104 8754 13128 8760
rect 13194 8754 13228 8760
rect 13284 8754 13328 8760
rect 13104 8726 13160 8754
rect 13194 8726 13250 8754
rect 13284 8726 13340 8754
rect 13374 8726 13435 8760
rect 12741 8667 13435 8726
rect 13484 9329 13516 9363
rect 13550 9362 13914 9363
rect 13550 9329 13664 9362
rect 13484 9328 13664 9329
rect 13698 9328 13765 9362
rect 13799 9348 13914 9362
rect 13948 9348 13984 9382
rect 14784 9418 14952 9423
rect 14986 9418 15053 9452
rect 15087 9442 15294 9452
rect 15328 9442 15384 9476
rect 15418 9442 15474 9476
rect 15508 9442 15564 9476
rect 15598 9442 15654 9476
rect 15688 9442 15744 9476
rect 15778 9442 15834 9476
rect 15868 9442 15924 9476
rect 15958 9442 16014 9476
rect 16048 9452 16582 9476
rect 16048 9442 16240 9452
rect 15087 9423 16240 9442
rect 15087 9418 15255 9423
rect 14784 9382 15255 9418
rect 14784 9363 15202 9382
rect 13799 9328 13984 9348
rect 13484 9292 13984 9328
rect 13484 9273 13914 9292
rect 13484 9239 13516 9273
rect 13550 9272 13914 9273
rect 13550 9239 13664 9272
rect 13484 9238 13664 9239
rect 13698 9238 13765 9272
rect 13799 9258 13914 9272
rect 13948 9258 13984 9292
rect 13799 9238 13984 9258
rect 13484 9202 13984 9238
rect 13484 9183 13914 9202
rect 13484 9149 13516 9183
rect 13550 9182 13914 9183
rect 13550 9149 13664 9182
rect 13484 9148 13664 9149
rect 13698 9148 13765 9182
rect 13799 9168 13914 9182
rect 13948 9168 13984 9202
rect 13799 9148 13984 9168
rect 13484 9112 13984 9148
rect 13484 9093 13914 9112
rect 13484 9059 13516 9093
rect 13550 9092 13914 9093
rect 13550 9059 13664 9092
rect 13484 9058 13664 9059
rect 13698 9058 13765 9092
rect 13799 9078 13914 9092
rect 13948 9078 13984 9112
rect 13799 9058 13984 9078
rect 13484 9022 13984 9058
rect 13484 9003 13914 9022
rect 13484 8969 13516 9003
rect 13550 9002 13914 9003
rect 13550 8969 13664 9002
rect 13484 8968 13664 8969
rect 13698 8968 13765 9002
rect 13799 8988 13914 9002
rect 13948 8988 13984 9022
rect 13799 8968 13984 8988
rect 13484 8932 13984 8968
rect 13484 8913 13914 8932
rect 13484 8879 13516 8913
rect 13550 8912 13914 8913
rect 13550 8879 13664 8912
rect 13484 8878 13664 8879
rect 13698 8878 13765 8912
rect 13799 8898 13914 8912
rect 13948 8898 13984 8932
rect 13799 8878 13984 8898
rect 13484 8842 13984 8878
rect 13484 8823 13914 8842
rect 13484 8789 13516 8823
rect 13550 8822 13914 8823
rect 13550 8789 13664 8822
rect 13484 8788 13664 8789
rect 13698 8788 13765 8822
rect 13799 8808 13914 8822
rect 13948 8808 13984 8842
rect 13799 8788 13984 8808
rect 13484 8752 13984 8788
rect 13484 8733 13914 8752
rect 13484 8699 13516 8733
rect 13550 8732 13914 8733
rect 13550 8699 13664 8732
rect 13484 8698 13664 8699
rect 13698 8698 13765 8732
rect 13799 8718 13914 8732
rect 13948 8718 13984 8752
rect 13799 8698 13984 8718
rect 12444 8642 12626 8662
rect 12444 8608 12477 8642
rect 12511 8628 12626 8642
rect 12660 8628 12684 8662
rect 12511 8608 12684 8628
rect 12444 8605 12684 8608
rect 13484 8662 13984 8698
rect 14029 9300 14723 9361
rect 14029 9266 14088 9300
rect 14122 9288 14178 9300
rect 14150 9266 14178 9288
rect 14212 9288 14268 9300
rect 14212 9266 14216 9288
rect 14029 9254 14116 9266
rect 14150 9254 14216 9266
rect 14250 9266 14268 9288
rect 14302 9288 14358 9300
rect 14302 9266 14316 9288
rect 14250 9254 14316 9266
rect 14350 9266 14358 9288
rect 14392 9288 14448 9300
rect 14482 9288 14538 9300
rect 14572 9288 14628 9300
rect 14392 9266 14416 9288
rect 14482 9266 14516 9288
rect 14572 9266 14616 9288
rect 14662 9266 14723 9300
rect 14350 9254 14416 9266
rect 14450 9254 14516 9266
rect 14550 9254 14616 9266
rect 14650 9254 14723 9266
rect 14029 9210 14723 9254
rect 14029 9176 14088 9210
rect 14122 9188 14178 9210
rect 14150 9176 14178 9188
rect 14212 9188 14268 9210
rect 14212 9176 14216 9188
rect 14029 9154 14116 9176
rect 14150 9154 14216 9176
rect 14250 9176 14268 9188
rect 14302 9188 14358 9210
rect 14302 9176 14316 9188
rect 14250 9154 14316 9176
rect 14350 9176 14358 9188
rect 14392 9188 14448 9210
rect 14482 9188 14538 9210
rect 14572 9188 14628 9210
rect 14392 9176 14416 9188
rect 14482 9176 14516 9188
rect 14572 9176 14616 9188
rect 14662 9176 14723 9210
rect 14350 9154 14416 9176
rect 14450 9154 14516 9176
rect 14550 9154 14616 9176
rect 14650 9154 14723 9176
rect 14029 9120 14723 9154
rect 14029 9086 14088 9120
rect 14122 9088 14178 9120
rect 14150 9086 14178 9088
rect 14212 9088 14268 9120
rect 14212 9086 14216 9088
rect 14029 9054 14116 9086
rect 14150 9054 14216 9086
rect 14250 9086 14268 9088
rect 14302 9088 14358 9120
rect 14302 9086 14316 9088
rect 14250 9054 14316 9086
rect 14350 9086 14358 9088
rect 14392 9088 14448 9120
rect 14482 9088 14538 9120
rect 14572 9088 14628 9120
rect 14392 9086 14416 9088
rect 14482 9086 14516 9088
rect 14572 9086 14616 9088
rect 14662 9086 14723 9120
rect 14350 9054 14416 9086
rect 14450 9054 14516 9086
rect 14550 9054 14616 9086
rect 14650 9054 14723 9086
rect 14029 9030 14723 9054
rect 14029 8996 14088 9030
rect 14122 8996 14178 9030
rect 14212 8996 14268 9030
rect 14302 8996 14358 9030
rect 14392 8996 14448 9030
rect 14482 8996 14538 9030
rect 14572 8996 14628 9030
rect 14662 8996 14723 9030
rect 14029 8988 14723 8996
rect 14029 8954 14116 8988
rect 14150 8954 14216 8988
rect 14250 8954 14316 8988
rect 14350 8954 14416 8988
rect 14450 8954 14516 8988
rect 14550 8954 14616 8988
rect 14650 8954 14723 8988
rect 14029 8940 14723 8954
rect 14029 8906 14088 8940
rect 14122 8906 14178 8940
rect 14212 8906 14268 8940
rect 14302 8906 14358 8940
rect 14392 8906 14448 8940
rect 14482 8906 14538 8940
rect 14572 8906 14628 8940
rect 14662 8906 14723 8940
rect 14029 8888 14723 8906
rect 14029 8854 14116 8888
rect 14150 8854 14216 8888
rect 14250 8854 14316 8888
rect 14350 8854 14416 8888
rect 14450 8854 14516 8888
rect 14550 8854 14616 8888
rect 14650 8854 14723 8888
rect 14029 8850 14723 8854
rect 14029 8816 14088 8850
rect 14122 8816 14178 8850
rect 14212 8816 14268 8850
rect 14302 8816 14358 8850
rect 14392 8816 14448 8850
rect 14482 8816 14538 8850
rect 14572 8816 14628 8850
rect 14662 8816 14723 8850
rect 14029 8788 14723 8816
rect 14029 8760 14116 8788
rect 14150 8760 14216 8788
rect 14029 8726 14088 8760
rect 14150 8754 14178 8760
rect 14122 8726 14178 8754
rect 14212 8754 14216 8760
rect 14250 8760 14316 8788
rect 14250 8754 14268 8760
rect 14212 8726 14268 8754
rect 14302 8754 14316 8760
rect 14350 8760 14416 8788
rect 14450 8760 14516 8788
rect 14550 8760 14616 8788
rect 14650 8760 14723 8788
rect 14350 8754 14358 8760
rect 14302 8726 14358 8754
rect 14392 8754 14416 8760
rect 14482 8754 14516 8760
rect 14572 8754 14616 8760
rect 14392 8726 14448 8754
rect 14482 8726 14538 8754
rect 14572 8726 14628 8754
rect 14662 8726 14723 8760
rect 14029 8667 14723 8726
rect 14784 9329 14804 9363
rect 14838 9362 15202 9363
rect 14838 9329 14952 9362
rect 14784 9328 14952 9329
rect 14986 9328 15053 9362
rect 15087 9348 15202 9362
rect 15236 9348 15255 9382
rect 16073 9418 16240 9423
rect 16274 9418 16341 9452
rect 16375 9442 16582 9452
rect 16616 9442 16672 9476
rect 16706 9442 16762 9476
rect 16796 9442 16852 9476
rect 16886 9442 16942 9476
rect 16976 9442 17032 9476
rect 17066 9442 17122 9476
rect 17156 9442 17212 9476
rect 17246 9442 17302 9476
rect 17336 9452 17870 9476
rect 17336 9442 17528 9452
rect 16375 9423 17528 9442
rect 16375 9418 16543 9423
rect 16073 9382 16543 9418
rect 16073 9363 16490 9382
rect 15087 9328 15255 9348
rect 14784 9292 15255 9328
rect 14784 9273 15202 9292
rect 14784 9239 14804 9273
rect 14838 9272 15202 9273
rect 14838 9239 14952 9272
rect 14784 9238 14952 9239
rect 14986 9238 15053 9272
rect 15087 9258 15202 9272
rect 15236 9258 15255 9292
rect 15087 9238 15255 9258
rect 14784 9202 15255 9238
rect 14784 9183 15202 9202
rect 14784 9149 14804 9183
rect 14838 9182 15202 9183
rect 14838 9149 14952 9182
rect 14784 9148 14952 9149
rect 14986 9148 15053 9182
rect 15087 9168 15202 9182
rect 15236 9168 15255 9202
rect 15087 9148 15255 9168
rect 14784 9112 15255 9148
rect 14784 9093 15202 9112
rect 14784 9059 14804 9093
rect 14838 9092 15202 9093
rect 14838 9059 14952 9092
rect 14784 9058 14952 9059
rect 14986 9058 15053 9092
rect 15087 9078 15202 9092
rect 15236 9078 15255 9112
rect 15087 9058 15255 9078
rect 14784 9022 15255 9058
rect 14784 9003 15202 9022
rect 14784 8969 14804 9003
rect 14838 9002 15202 9003
rect 14838 8969 14952 9002
rect 14784 8968 14952 8969
rect 14986 8968 15053 9002
rect 15087 8988 15202 9002
rect 15236 8988 15255 9022
rect 15087 8968 15255 8988
rect 14784 8932 15255 8968
rect 14784 8913 15202 8932
rect 14784 8879 14804 8913
rect 14838 8912 15202 8913
rect 14838 8879 14952 8912
rect 14784 8878 14952 8879
rect 14986 8878 15053 8912
rect 15087 8898 15202 8912
rect 15236 8898 15255 8932
rect 15087 8878 15255 8898
rect 14784 8842 15255 8878
rect 14784 8823 15202 8842
rect 14784 8789 14804 8823
rect 14838 8822 15202 8823
rect 14838 8789 14952 8822
rect 14784 8788 14952 8789
rect 14986 8788 15053 8822
rect 15087 8808 15202 8822
rect 15236 8808 15255 8842
rect 15087 8788 15255 8808
rect 14784 8752 15255 8788
rect 14784 8733 15202 8752
rect 14784 8699 14804 8733
rect 14838 8732 15202 8733
rect 14838 8699 14952 8732
rect 14784 8698 14952 8699
rect 14986 8698 15053 8732
rect 15087 8718 15202 8732
rect 15236 8718 15255 8752
rect 15087 8698 15255 8718
rect 13484 8643 13914 8662
rect 13484 8609 13516 8643
rect 13550 8642 13914 8643
rect 13550 8609 13664 8642
rect 13484 8608 13664 8609
rect 13698 8608 13765 8642
rect 13799 8628 13914 8642
rect 13948 8628 13984 8662
rect 13799 8608 13984 8628
rect 13484 8605 13984 8608
rect 14784 8662 15255 8698
rect 15317 9300 16011 9361
rect 15317 9266 15376 9300
rect 15410 9288 15466 9300
rect 15438 9266 15466 9288
rect 15500 9288 15556 9300
rect 15500 9266 15504 9288
rect 15317 9254 15404 9266
rect 15438 9254 15504 9266
rect 15538 9266 15556 9288
rect 15590 9288 15646 9300
rect 15590 9266 15604 9288
rect 15538 9254 15604 9266
rect 15638 9266 15646 9288
rect 15680 9288 15736 9300
rect 15770 9288 15826 9300
rect 15860 9288 15916 9300
rect 15680 9266 15704 9288
rect 15770 9266 15804 9288
rect 15860 9266 15904 9288
rect 15950 9266 16011 9300
rect 15638 9254 15704 9266
rect 15738 9254 15804 9266
rect 15838 9254 15904 9266
rect 15938 9254 16011 9266
rect 15317 9210 16011 9254
rect 15317 9176 15376 9210
rect 15410 9188 15466 9210
rect 15438 9176 15466 9188
rect 15500 9188 15556 9210
rect 15500 9176 15504 9188
rect 15317 9154 15404 9176
rect 15438 9154 15504 9176
rect 15538 9176 15556 9188
rect 15590 9188 15646 9210
rect 15590 9176 15604 9188
rect 15538 9154 15604 9176
rect 15638 9176 15646 9188
rect 15680 9188 15736 9210
rect 15770 9188 15826 9210
rect 15860 9188 15916 9210
rect 15680 9176 15704 9188
rect 15770 9176 15804 9188
rect 15860 9176 15904 9188
rect 15950 9176 16011 9210
rect 15638 9154 15704 9176
rect 15738 9154 15804 9176
rect 15838 9154 15904 9176
rect 15938 9154 16011 9176
rect 15317 9120 16011 9154
rect 15317 9086 15376 9120
rect 15410 9088 15466 9120
rect 15438 9086 15466 9088
rect 15500 9088 15556 9120
rect 15500 9086 15504 9088
rect 15317 9054 15404 9086
rect 15438 9054 15504 9086
rect 15538 9086 15556 9088
rect 15590 9088 15646 9120
rect 15590 9086 15604 9088
rect 15538 9054 15604 9086
rect 15638 9086 15646 9088
rect 15680 9088 15736 9120
rect 15770 9088 15826 9120
rect 15860 9088 15916 9120
rect 15680 9086 15704 9088
rect 15770 9086 15804 9088
rect 15860 9086 15904 9088
rect 15950 9086 16011 9120
rect 15638 9054 15704 9086
rect 15738 9054 15804 9086
rect 15838 9054 15904 9086
rect 15938 9054 16011 9086
rect 15317 9030 16011 9054
rect 15317 8996 15376 9030
rect 15410 8996 15466 9030
rect 15500 8996 15556 9030
rect 15590 8996 15646 9030
rect 15680 8996 15736 9030
rect 15770 8996 15826 9030
rect 15860 8996 15916 9030
rect 15950 8996 16011 9030
rect 15317 8988 16011 8996
rect 15317 8954 15404 8988
rect 15438 8954 15504 8988
rect 15538 8954 15604 8988
rect 15638 8954 15704 8988
rect 15738 8954 15804 8988
rect 15838 8954 15904 8988
rect 15938 8954 16011 8988
rect 15317 8940 16011 8954
rect 15317 8906 15376 8940
rect 15410 8906 15466 8940
rect 15500 8906 15556 8940
rect 15590 8906 15646 8940
rect 15680 8906 15736 8940
rect 15770 8906 15826 8940
rect 15860 8906 15916 8940
rect 15950 8906 16011 8940
rect 15317 8888 16011 8906
rect 15317 8854 15404 8888
rect 15438 8854 15504 8888
rect 15538 8854 15604 8888
rect 15638 8854 15704 8888
rect 15738 8854 15804 8888
rect 15838 8854 15904 8888
rect 15938 8854 16011 8888
rect 15317 8850 16011 8854
rect 15317 8816 15376 8850
rect 15410 8816 15466 8850
rect 15500 8816 15556 8850
rect 15590 8816 15646 8850
rect 15680 8816 15736 8850
rect 15770 8816 15826 8850
rect 15860 8816 15916 8850
rect 15950 8816 16011 8850
rect 15317 8788 16011 8816
rect 15317 8760 15404 8788
rect 15438 8760 15504 8788
rect 15317 8726 15376 8760
rect 15438 8754 15466 8760
rect 15410 8726 15466 8754
rect 15500 8754 15504 8760
rect 15538 8760 15604 8788
rect 15538 8754 15556 8760
rect 15500 8726 15556 8754
rect 15590 8754 15604 8760
rect 15638 8760 15704 8788
rect 15738 8760 15804 8788
rect 15838 8760 15904 8788
rect 15938 8760 16011 8788
rect 15638 8754 15646 8760
rect 15590 8726 15646 8754
rect 15680 8754 15704 8760
rect 15770 8754 15804 8760
rect 15860 8754 15904 8760
rect 15680 8726 15736 8754
rect 15770 8726 15826 8754
rect 15860 8726 15916 8754
rect 15950 8726 16011 8760
rect 15317 8667 16011 8726
rect 16073 9329 16092 9363
rect 16126 9362 16490 9363
rect 16126 9329 16240 9362
rect 16073 9328 16240 9329
rect 16274 9328 16341 9362
rect 16375 9348 16490 9362
rect 16524 9348 16543 9382
rect 17361 9418 17528 9423
rect 17562 9418 17629 9452
rect 17663 9442 17870 9452
rect 17904 9442 17960 9476
rect 17994 9442 18050 9476
rect 18084 9442 18140 9476
rect 18174 9442 18230 9476
rect 18264 9442 18320 9476
rect 18354 9442 18410 9476
rect 18444 9442 18500 9476
rect 18534 9442 18590 9476
rect 18624 9452 18884 9476
rect 18624 9442 18816 9452
rect 17663 9423 18816 9442
rect 17663 9418 17831 9423
rect 17361 9382 17831 9418
rect 17361 9363 17778 9382
rect 16375 9328 16543 9348
rect 16073 9292 16543 9328
rect 16073 9273 16490 9292
rect 16073 9239 16092 9273
rect 16126 9272 16490 9273
rect 16126 9239 16240 9272
rect 16073 9238 16240 9239
rect 16274 9238 16341 9272
rect 16375 9258 16490 9272
rect 16524 9258 16543 9292
rect 16375 9238 16543 9258
rect 16073 9202 16543 9238
rect 16073 9183 16490 9202
rect 16073 9149 16092 9183
rect 16126 9182 16490 9183
rect 16126 9149 16240 9182
rect 16073 9148 16240 9149
rect 16274 9148 16341 9182
rect 16375 9168 16490 9182
rect 16524 9168 16543 9202
rect 16375 9148 16543 9168
rect 16073 9112 16543 9148
rect 16073 9093 16490 9112
rect 16073 9059 16092 9093
rect 16126 9092 16490 9093
rect 16126 9059 16240 9092
rect 16073 9058 16240 9059
rect 16274 9058 16341 9092
rect 16375 9078 16490 9092
rect 16524 9078 16543 9112
rect 16375 9058 16543 9078
rect 16073 9022 16543 9058
rect 16073 9003 16490 9022
rect 16073 8969 16092 9003
rect 16126 9002 16490 9003
rect 16126 8969 16240 9002
rect 16073 8968 16240 8969
rect 16274 8968 16341 9002
rect 16375 8988 16490 9002
rect 16524 8988 16543 9022
rect 16375 8968 16543 8988
rect 16073 8932 16543 8968
rect 16073 8913 16490 8932
rect 16073 8879 16092 8913
rect 16126 8912 16490 8913
rect 16126 8879 16240 8912
rect 16073 8878 16240 8879
rect 16274 8878 16341 8912
rect 16375 8898 16490 8912
rect 16524 8898 16543 8932
rect 16375 8878 16543 8898
rect 16073 8842 16543 8878
rect 16073 8823 16490 8842
rect 16073 8789 16092 8823
rect 16126 8822 16490 8823
rect 16126 8789 16240 8822
rect 16073 8788 16240 8789
rect 16274 8788 16341 8822
rect 16375 8808 16490 8822
rect 16524 8808 16543 8842
rect 16375 8788 16543 8808
rect 16073 8752 16543 8788
rect 16073 8733 16490 8752
rect 16073 8699 16092 8733
rect 16126 8732 16490 8733
rect 16126 8699 16240 8732
rect 16073 8698 16240 8699
rect 16274 8698 16341 8732
rect 16375 8718 16490 8732
rect 16524 8718 16543 8752
rect 16375 8698 16543 8718
rect 14784 8643 15202 8662
rect 14784 8609 14804 8643
rect 14838 8642 15202 8643
rect 14838 8609 14952 8642
rect 14784 8608 14952 8609
rect 14986 8608 15053 8642
rect 15087 8628 15202 8642
rect 15236 8628 15255 8662
rect 15087 8608 15255 8628
rect 14784 8605 15255 8608
rect 16073 8662 16543 8698
rect 16605 9300 17299 9361
rect 16605 9266 16664 9300
rect 16698 9288 16754 9300
rect 16726 9266 16754 9288
rect 16788 9288 16844 9300
rect 16788 9266 16792 9288
rect 16605 9254 16692 9266
rect 16726 9254 16792 9266
rect 16826 9266 16844 9288
rect 16878 9288 16934 9300
rect 16878 9266 16892 9288
rect 16826 9254 16892 9266
rect 16926 9266 16934 9288
rect 16968 9288 17024 9300
rect 17058 9288 17114 9300
rect 17148 9288 17204 9300
rect 16968 9266 16992 9288
rect 17058 9266 17092 9288
rect 17148 9266 17192 9288
rect 17238 9266 17299 9300
rect 16926 9254 16992 9266
rect 17026 9254 17092 9266
rect 17126 9254 17192 9266
rect 17226 9254 17299 9266
rect 16605 9210 17299 9254
rect 16605 9176 16664 9210
rect 16698 9188 16754 9210
rect 16726 9176 16754 9188
rect 16788 9188 16844 9210
rect 16788 9176 16792 9188
rect 16605 9154 16692 9176
rect 16726 9154 16792 9176
rect 16826 9176 16844 9188
rect 16878 9188 16934 9210
rect 16878 9176 16892 9188
rect 16826 9154 16892 9176
rect 16926 9176 16934 9188
rect 16968 9188 17024 9210
rect 17058 9188 17114 9210
rect 17148 9188 17204 9210
rect 16968 9176 16992 9188
rect 17058 9176 17092 9188
rect 17148 9176 17192 9188
rect 17238 9176 17299 9210
rect 16926 9154 16992 9176
rect 17026 9154 17092 9176
rect 17126 9154 17192 9176
rect 17226 9154 17299 9176
rect 16605 9120 17299 9154
rect 16605 9086 16664 9120
rect 16698 9088 16754 9120
rect 16726 9086 16754 9088
rect 16788 9088 16844 9120
rect 16788 9086 16792 9088
rect 16605 9054 16692 9086
rect 16726 9054 16792 9086
rect 16826 9086 16844 9088
rect 16878 9088 16934 9120
rect 16878 9086 16892 9088
rect 16826 9054 16892 9086
rect 16926 9086 16934 9088
rect 16968 9088 17024 9120
rect 17058 9088 17114 9120
rect 17148 9088 17204 9120
rect 16968 9086 16992 9088
rect 17058 9086 17092 9088
rect 17148 9086 17192 9088
rect 17238 9086 17299 9120
rect 16926 9054 16992 9086
rect 17026 9054 17092 9086
rect 17126 9054 17192 9086
rect 17226 9054 17299 9086
rect 16605 9030 17299 9054
rect 16605 8996 16664 9030
rect 16698 8996 16754 9030
rect 16788 8996 16844 9030
rect 16878 8996 16934 9030
rect 16968 8996 17024 9030
rect 17058 8996 17114 9030
rect 17148 8996 17204 9030
rect 17238 8996 17299 9030
rect 16605 8988 17299 8996
rect 16605 8954 16692 8988
rect 16726 8954 16792 8988
rect 16826 8954 16892 8988
rect 16926 8954 16992 8988
rect 17026 8954 17092 8988
rect 17126 8954 17192 8988
rect 17226 8954 17299 8988
rect 16605 8940 17299 8954
rect 16605 8906 16664 8940
rect 16698 8906 16754 8940
rect 16788 8906 16844 8940
rect 16878 8906 16934 8940
rect 16968 8906 17024 8940
rect 17058 8906 17114 8940
rect 17148 8906 17204 8940
rect 17238 8906 17299 8940
rect 16605 8888 17299 8906
rect 16605 8854 16692 8888
rect 16726 8854 16792 8888
rect 16826 8854 16892 8888
rect 16926 8854 16992 8888
rect 17026 8854 17092 8888
rect 17126 8854 17192 8888
rect 17226 8854 17299 8888
rect 16605 8850 17299 8854
rect 16605 8816 16664 8850
rect 16698 8816 16754 8850
rect 16788 8816 16844 8850
rect 16878 8816 16934 8850
rect 16968 8816 17024 8850
rect 17058 8816 17114 8850
rect 17148 8816 17204 8850
rect 17238 8816 17299 8850
rect 16605 8788 17299 8816
rect 16605 8760 16692 8788
rect 16726 8760 16792 8788
rect 16605 8726 16664 8760
rect 16726 8754 16754 8760
rect 16698 8726 16754 8754
rect 16788 8754 16792 8760
rect 16826 8760 16892 8788
rect 16826 8754 16844 8760
rect 16788 8726 16844 8754
rect 16878 8754 16892 8760
rect 16926 8760 16992 8788
rect 17026 8760 17092 8788
rect 17126 8760 17192 8788
rect 17226 8760 17299 8788
rect 16926 8754 16934 8760
rect 16878 8726 16934 8754
rect 16968 8754 16992 8760
rect 17058 8754 17092 8760
rect 17148 8754 17192 8760
rect 16968 8726 17024 8754
rect 17058 8726 17114 8754
rect 17148 8726 17204 8754
rect 17238 8726 17299 8760
rect 16605 8667 17299 8726
rect 17361 9329 17380 9363
rect 17414 9362 17778 9363
rect 17414 9329 17528 9362
rect 17361 9328 17528 9329
rect 17562 9328 17629 9362
rect 17663 9348 17778 9362
rect 17812 9348 17831 9382
rect 18649 9418 18816 9423
rect 18850 9418 18884 9452
rect 18649 9363 18884 9418
rect 17663 9328 17831 9348
rect 17361 9292 17831 9328
rect 17361 9273 17778 9292
rect 17361 9239 17380 9273
rect 17414 9272 17778 9273
rect 17414 9239 17528 9272
rect 17361 9238 17528 9239
rect 17562 9238 17629 9272
rect 17663 9258 17778 9272
rect 17812 9258 17831 9292
rect 17663 9238 17831 9258
rect 17361 9202 17831 9238
rect 17361 9183 17778 9202
rect 17361 9149 17380 9183
rect 17414 9182 17778 9183
rect 17414 9149 17528 9182
rect 17361 9148 17528 9149
rect 17562 9148 17629 9182
rect 17663 9168 17778 9182
rect 17812 9168 17831 9202
rect 17663 9148 17831 9168
rect 17361 9112 17831 9148
rect 17361 9093 17778 9112
rect 17361 9059 17380 9093
rect 17414 9092 17778 9093
rect 17414 9059 17528 9092
rect 17361 9058 17528 9059
rect 17562 9058 17629 9092
rect 17663 9078 17778 9092
rect 17812 9078 17831 9112
rect 17663 9058 17831 9078
rect 17361 9022 17831 9058
rect 17361 9003 17778 9022
rect 17361 8969 17380 9003
rect 17414 9002 17778 9003
rect 17414 8969 17528 9002
rect 17361 8968 17528 8969
rect 17562 8968 17629 9002
rect 17663 8988 17778 9002
rect 17812 8988 17831 9022
rect 17663 8968 17831 8988
rect 17361 8932 17831 8968
rect 17361 8913 17778 8932
rect 17361 8879 17380 8913
rect 17414 8912 17778 8913
rect 17414 8879 17528 8912
rect 17361 8878 17528 8879
rect 17562 8878 17629 8912
rect 17663 8898 17778 8912
rect 17812 8898 17831 8932
rect 17663 8878 17831 8898
rect 17361 8842 17831 8878
rect 17361 8823 17778 8842
rect 17361 8789 17380 8823
rect 17414 8822 17778 8823
rect 17414 8789 17528 8822
rect 17361 8788 17528 8789
rect 17562 8788 17629 8822
rect 17663 8808 17778 8822
rect 17812 8808 17831 8842
rect 17663 8788 17831 8808
rect 17361 8752 17831 8788
rect 17361 8733 17778 8752
rect 17361 8699 17380 8733
rect 17414 8732 17778 8733
rect 17414 8699 17528 8732
rect 17361 8698 17528 8699
rect 17562 8698 17629 8732
rect 17663 8718 17778 8732
rect 17812 8718 17831 8752
rect 17663 8698 17831 8718
rect 16073 8643 16490 8662
rect 16073 8609 16092 8643
rect 16126 8642 16490 8643
rect 16126 8609 16240 8642
rect 16073 8608 16240 8609
rect 16274 8608 16341 8642
rect 16375 8628 16490 8642
rect 16524 8628 16543 8662
rect 16375 8608 16543 8628
rect 16073 8605 16543 8608
rect 17361 8662 17831 8698
rect 17893 9300 18587 9361
rect 17893 9266 17952 9300
rect 17986 9288 18042 9300
rect 18014 9266 18042 9288
rect 18076 9288 18132 9300
rect 18076 9266 18080 9288
rect 17893 9254 17980 9266
rect 18014 9254 18080 9266
rect 18114 9266 18132 9288
rect 18166 9288 18222 9300
rect 18166 9266 18180 9288
rect 18114 9254 18180 9266
rect 18214 9266 18222 9288
rect 18256 9288 18312 9300
rect 18346 9288 18402 9300
rect 18436 9288 18492 9300
rect 18256 9266 18280 9288
rect 18346 9266 18380 9288
rect 18436 9266 18480 9288
rect 18526 9266 18587 9300
rect 18214 9254 18280 9266
rect 18314 9254 18380 9266
rect 18414 9254 18480 9266
rect 18514 9254 18587 9266
rect 17893 9210 18587 9254
rect 17893 9176 17952 9210
rect 17986 9188 18042 9210
rect 18014 9176 18042 9188
rect 18076 9188 18132 9210
rect 18076 9176 18080 9188
rect 17893 9154 17980 9176
rect 18014 9154 18080 9176
rect 18114 9176 18132 9188
rect 18166 9188 18222 9210
rect 18166 9176 18180 9188
rect 18114 9154 18180 9176
rect 18214 9176 18222 9188
rect 18256 9188 18312 9210
rect 18346 9188 18402 9210
rect 18436 9188 18492 9210
rect 18256 9176 18280 9188
rect 18346 9176 18380 9188
rect 18436 9176 18480 9188
rect 18526 9176 18587 9210
rect 18214 9154 18280 9176
rect 18314 9154 18380 9176
rect 18414 9154 18480 9176
rect 18514 9154 18587 9176
rect 17893 9120 18587 9154
rect 17893 9086 17952 9120
rect 17986 9088 18042 9120
rect 18014 9086 18042 9088
rect 18076 9088 18132 9120
rect 18076 9086 18080 9088
rect 17893 9054 17980 9086
rect 18014 9054 18080 9086
rect 18114 9086 18132 9088
rect 18166 9088 18222 9120
rect 18166 9086 18180 9088
rect 18114 9054 18180 9086
rect 18214 9086 18222 9088
rect 18256 9088 18312 9120
rect 18346 9088 18402 9120
rect 18436 9088 18492 9120
rect 18256 9086 18280 9088
rect 18346 9086 18380 9088
rect 18436 9086 18480 9088
rect 18526 9086 18587 9120
rect 18214 9054 18280 9086
rect 18314 9054 18380 9086
rect 18414 9054 18480 9086
rect 18514 9054 18587 9086
rect 17893 9030 18587 9054
rect 17893 8996 17952 9030
rect 17986 8996 18042 9030
rect 18076 8996 18132 9030
rect 18166 8996 18222 9030
rect 18256 8996 18312 9030
rect 18346 8996 18402 9030
rect 18436 8996 18492 9030
rect 18526 8996 18587 9030
rect 17893 8988 18587 8996
rect 17893 8954 17980 8988
rect 18014 8954 18080 8988
rect 18114 8954 18180 8988
rect 18214 8954 18280 8988
rect 18314 8954 18380 8988
rect 18414 8954 18480 8988
rect 18514 8954 18587 8988
rect 17893 8940 18587 8954
rect 17893 8906 17952 8940
rect 17986 8906 18042 8940
rect 18076 8906 18132 8940
rect 18166 8906 18222 8940
rect 18256 8906 18312 8940
rect 18346 8906 18402 8940
rect 18436 8906 18492 8940
rect 18526 8906 18587 8940
rect 17893 8888 18587 8906
rect 17893 8854 17980 8888
rect 18014 8854 18080 8888
rect 18114 8854 18180 8888
rect 18214 8854 18280 8888
rect 18314 8854 18380 8888
rect 18414 8854 18480 8888
rect 18514 8854 18587 8888
rect 17893 8850 18587 8854
rect 17893 8816 17952 8850
rect 17986 8816 18042 8850
rect 18076 8816 18132 8850
rect 18166 8816 18222 8850
rect 18256 8816 18312 8850
rect 18346 8816 18402 8850
rect 18436 8816 18492 8850
rect 18526 8816 18587 8850
rect 17893 8788 18587 8816
rect 17893 8760 17980 8788
rect 18014 8760 18080 8788
rect 17893 8726 17952 8760
rect 18014 8754 18042 8760
rect 17986 8726 18042 8754
rect 18076 8754 18080 8760
rect 18114 8760 18180 8788
rect 18114 8754 18132 8760
rect 18076 8726 18132 8754
rect 18166 8754 18180 8760
rect 18214 8760 18280 8788
rect 18314 8760 18380 8788
rect 18414 8760 18480 8788
rect 18514 8760 18587 8788
rect 18214 8754 18222 8760
rect 18166 8726 18222 8754
rect 18256 8754 18280 8760
rect 18346 8754 18380 8760
rect 18436 8754 18480 8760
rect 18256 8726 18312 8754
rect 18346 8726 18402 8754
rect 18436 8726 18492 8754
rect 18526 8726 18587 8760
rect 17893 8667 18587 8726
rect 18649 9329 18668 9363
rect 18702 9362 18884 9363
rect 18702 9329 18816 9362
rect 18649 9328 18816 9329
rect 18850 9328 18884 9362
rect 18649 9273 18884 9328
rect 18649 9239 18668 9273
rect 18702 9272 18884 9273
rect 18702 9239 18816 9272
rect 18649 9238 18816 9239
rect 18850 9238 18884 9272
rect 18649 9183 18884 9238
rect 18649 9149 18668 9183
rect 18702 9182 18884 9183
rect 18702 9149 18816 9182
rect 18649 9148 18816 9149
rect 18850 9148 18884 9182
rect 18649 9093 18884 9148
rect 18649 9059 18668 9093
rect 18702 9092 18884 9093
rect 18702 9059 18816 9092
rect 18649 9058 18816 9059
rect 18850 9058 18884 9092
rect 18649 9003 18884 9058
rect 18649 8969 18668 9003
rect 18702 9002 18884 9003
rect 18702 8969 18816 9002
rect 18649 8968 18816 8969
rect 18850 8968 18884 9002
rect 18649 8913 18884 8968
rect 18649 8879 18668 8913
rect 18702 8912 18884 8913
rect 18702 8879 18816 8912
rect 18649 8878 18816 8879
rect 18850 8878 18884 8912
rect 18649 8823 18884 8878
rect 18649 8789 18668 8823
rect 18702 8822 18884 8823
rect 18702 8789 18816 8822
rect 18649 8788 18816 8789
rect 18850 8788 18884 8822
rect 18649 8733 18884 8788
rect 18649 8699 18668 8733
rect 18702 8732 18884 8733
rect 18702 8699 18816 8732
rect 18649 8698 18816 8699
rect 18850 8698 18884 8732
rect 17361 8643 17778 8662
rect 17361 8609 17380 8643
rect 17414 8642 17778 8643
rect 17414 8609 17528 8642
rect 17361 8608 17528 8609
rect 17562 8608 17629 8642
rect 17663 8628 17778 8642
rect 17812 8628 17831 8662
rect 17663 8608 17831 8628
rect 17361 8605 17831 8608
rect 18649 8643 18884 8698
rect 18649 8609 18668 8643
rect 18702 8642 18884 8643
rect 18702 8609 18816 8642
rect 18649 8608 18816 8609
rect 18850 8608 18884 8642
rect 18649 8605 18884 8608
rect 12444 8586 18884 8605
rect 12444 8552 12684 8586
rect 12718 8552 12774 8586
rect 12808 8552 12864 8586
rect 12898 8552 12954 8586
rect 12988 8552 13044 8586
rect 13078 8552 13134 8586
rect 13168 8552 13224 8586
rect 13258 8552 13314 8586
rect 13348 8552 13404 8586
rect 13438 8552 13972 8586
rect 14006 8552 14062 8586
rect 14096 8552 14152 8586
rect 14186 8552 14242 8586
rect 14276 8552 14332 8586
rect 14366 8552 14422 8586
rect 14456 8552 14512 8586
rect 14546 8552 14602 8586
rect 14636 8552 14692 8586
rect 14726 8552 15260 8586
rect 15294 8552 15350 8586
rect 15384 8552 15440 8586
rect 15474 8552 15530 8586
rect 15564 8552 15620 8586
rect 15654 8552 15710 8586
rect 15744 8552 15800 8586
rect 15834 8552 15890 8586
rect 15924 8552 15980 8586
rect 16014 8552 16548 8586
rect 16582 8552 16638 8586
rect 16672 8552 16728 8586
rect 16762 8552 16818 8586
rect 16852 8552 16908 8586
rect 16942 8552 16998 8586
rect 17032 8552 17088 8586
rect 17122 8552 17178 8586
rect 17212 8552 17268 8586
rect 17302 8552 17836 8586
rect 17870 8552 17926 8586
rect 17960 8552 18016 8586
rect 18050 8552 18106 8586
rect 18140 8552 18196 8586
rect 18230 8552 18286 8586
rect 18320 8552 18376 8586
rect 18410 8552 18466 8586
rect 18500 8552 18556 8586
rect 18590 8552 18884 8586
rect 12444 8518 12477 8552
rect 12511 8533 13664 8552
rect 12511 8518 12684 8533
rect 12444 8469 12684 8518
rect 13484 8518 13664 8533
rect 13698 8518 13765 8552
rect 13799 8533 14952 8552
rect 13799 8518 13984 8533
rect 13484 8469 13984 8518
rect 14784 8518 14952 8533
rect 14986 8518 15053 8552
rect 15087 8533 16240 8552
rect 15087 8518 15184 8533
rect 14784 8469 15184 8518
rect 16084 8518 16240 8533
rect 16274 8518 16341 8552
rect 16375 8533 17528 8552
rect 16375 8518 16484 8533
rect 16084 8469 16484 8518
rect 17384 8518 17528 8533
rect 17562 8518 17629 8552
rect 17663 8533 18816 8552
rect 17663 8518 17784 8533
rect 17384 8469 17784 8518
rect 18684 8518 18816 8533
rect 18850 8518 18884 8552
rect 18684 8469 18884 8518
rect 12444 8462 18884 8469
rect 12444 8428 12477 8462
rect 12511 8439 13664 8462
rect 12511 8428 12578 8439
rect 12444 8405 12578 8428
rect 12612 8405 12668 8439
rect 12702 8405 12758 8439
rect 12792 8405 12848 8439
rect 12882 8405 12938 8439
rect 12972 8405 13028 8439
rect 13062 8405 13118 8439
rect 13152 8405 13208 8439
rect 13242 8405 13298 8439
rect 13332 8405 13388 8439
rect 13422 8405 13478 8439
rect 13512 8405 13568 8439
rect 13602 8428 13664 8439
rect 13698 8428 13765 8462
rect 13799 8439 14952 8462
rect 13799 8428 13866 8439
rect 13602 8405 13866 8428
rect 13900 8405 13956 8439
rect 13990 8405 14046 8439
rect 14080 8405 14136 8439
rect 14170 8405 14226 8439
rect 14260 8405 14316 8439
rect 14350 8405 14406 8439
rect 14440 8405 14496 8439
rect 14530 8405 14586 8439
rect 14620 8405 14676 8439
rect 14710 8405 14766 8439
rect 14800 8405 14856 8439
rect 14890 8428 14952 8439
rect 14986 8428 15053 8462
rect 15087 8439 16240 8462
rect 15087 8428 15154 8439
rect 14890 8405 15154 8428
rect 15188 8405 15244 8439
rect 15278 8405 15334 8439
rect 15368 8405 15424 8439
rect 15458 8405 15514 8439
rect 15548 8405 15604 8439
rect 15638 8405 15694 8439
rect 15728 8405 15784 8439
rect 15818 8405 15874 8439
rect 15908 8405 15964 8439
rect 15998 8405 16054 8439
rect 16088 8405 16144 8439
rect 16178 8428 16240 8439
rect 16274 8428 16341 8462
rect 16375 8439 17528 8462
rect 16375 8428 16442 8439
rect 16178 8405 16442 8428
rect 16476 8405 16532 8439
rect 16566 8405 16622 8439
rect 16656 8405 16712 8439
rect 16746 8405 16802 8439
rect 16836 8405 16892 8439
rect 16926 8405 16982 8439
rect 17016 8405 17072 8439
rect 17106 8405 17162 8439
rect 17196 8405 17252 8439
rect 17286 8405 17342 8439
rect 17376 8405 17432 8439
rect 17466 8428 17528 8439
rect 17562 8428 17629 8462
rect 17663 8439 18816 8462
rect 17663 8428 17730 8439
rect 17466 8405 17730 8428
rect 17764 8405 17820 8439
rect 17854 8405 17910 8439
rect 17944 8405 18000 8439
rect 18034 8405 18090 8439
rect 18124 8405 18180 8439
rect 18214 8405 18270 8439
rect 18304 8405 18360 8439
rect 18394 8405 18450 8439
rect 18484 8405 18540 8439
rect 18574 8405 18630 8439
rect 18664 8405 18720 8439
rect 18754 8428 18816 8439
rect 18850 8428 18884 8462
rect 18754 8405 18884 8428
rect 12444 8338 18884 8405
rect 12444 8304 12578 8338
rect 12612 8304 12668 8338
rect 12702 8304 12758 8338
rect 12792 8304 12848 8338
rect 12882 8304 12938 8338
rect 12972 8304 13028 8338
rect 13062 8304 13118 8338
rect 13152 8304 13208 8338
rect 13242 8304 13298 8338
rect 13332 8304 13388 8338
rect 13422 8304 13478 8338
rect 13512 8304 13568 8338
rect 13602 8304 13866 8338
rect 13900 8304 13956 8338
rect 13990 8304 14046 8338
rect 14080 8304 14136 8338
rect 14170 8304 14226 8338
rect 14260 8304 14316 8338
rect 14350 8304 14406 8338
rect 14440 8304 14496 8338
rect 14530 8304 14586 8338
rect 14620 8304 14676 8338
rect 14710 8304 14766 8338
rect 14800 8304 14856 8338
rect 14890 8304 15154 8338
rect 15188 8304 15244 8338
rect 15278 8304 15334 8338
rect 15368 8304 15424 8338
rect 15458 8304 15514 8338
rect 15548 8304 15604 8338
rect 15638 8304 15694 8338
rect 15728 8304 15784 8338
rect 15818 8304 15874 8338
rect 15908 8304 15964 8338
rect 15998 8304 16054 8338
rect 16088 8304 16144 8338
rect 16178 8304 16442 8338
rect 16476 8304 16532 8338
rect 16566 8304 16622 8338
rect 16656 8304 16712 8338
rect 16746 8304 16802 8338
rect 16836 8304 16892 8338
rect 16926 8304 16982 8338
rect 17016 8304 17072 8338
rect 17106 8304 17162 8338
rect 17196 8304 17252 8338
rect 17286 8304 17342 8338
rect 17376 8304 17432 8338
rect 17466 8304 17730 8338
rect 17764 8304 17820 8338
rect 17854 8304 17910 8338
rect 17944 8304 18000 8338
rect 18034 8304 18090 8338
rect 18124 8304 18180 8338
rect 18214 8304 18270 8338
rect 18304 8304 18360 8338
rect 18394 8304 18450 8338
rect 18484 8304 18540 8338
rect 18574 8304 18630 8338
rect 18664 8304 18720 8338
rect 18754 8304 18884 8338
rect 12444 8271 18884 8304
rect 12444 8254 12684 8271
rect 12444 8220 12477 8254
rect 12511 8220 12684 8254
rect 12444 8207 12684 8220
rect 13484 8254 13984 8271
rect 13484 8220 13664 8254
rect 13698 8220 13765 8254
rect 13799 8220 13984 8254
rect 13484 8207 13984 8220
rect 14784 8254 15184 8271
rect 14784 8220 14952 8254
rect 14986 8220 15053 8254
rect 15087 8220 15184 8254
rect 14784 8207 15184 8220
rect 16084 8254 16484 8271
rect 16084 8220 16240 8254
rect 16274 8220 16341 8254
rect 16375 8220 16484 8254
rect 16084 8207 16484 8220
rect 17384 8254 17784 8271
rect 17384 8220 17528 8254
rect 17562 8220 17629 8254
rect 17663 8220 17784 8254
rect 17384 8207 17784 8220
rect 18684 8254 18884 8271
rect 18684 8220 18816 8254
rect 18850 8220 18884 8254
rect 18684 8207 18884 8220
rect 12444 8188 18884 8207
rect 12444 8164 12718 8188
rect 12444 8130 12477 8164
rect 12511 8154 12718 8164
rect 12752 8154 12808 8188
rect 12842 8154 12898 8188
rect 12932 8154 12988 8188
rect 13022 8154 13078 8188
rect 13112 8154 13168 8188
rect 13202 8154 13258 8188
rect 13292 8154 13348 8188
rect 13382 8154 13438 8188
rect 13472 8164 14006 8188
rect 13472 8154 13664 8164
rect 12511 8135 13664 8154
rect 12511 8130 12684 8135
rect 12444 8094 12684 8130
rect 12444 8074 12626 8094
rect 12444 8040 12477 8074
rect 12511 8060 12626 8074
rect 12660 8060 12684 8094
rect 13484 8130 13664 8135
rect 13698 8130 13765 8164
rect 13799 8154 14006 8164
rect 14040 8154 14096 8188
rect 14130 8154 14186 8188
rect 14220 8154 14276 8188
rect 14310 8154 14366 8188
rect 14400 8154 14456 8188
rect 14490 8154 14546 8188
rect 14580 8154 14636 8188
rect 14670 8154 14726 8188
rect 14760 8164 15294 8188
rect 14760 8154 14952 8164
rect 13799 8135 14952 8154
rect 13799 8130 13984 8135
rect 13484 8094 13984 8130
rect 13484 8075 13914 8094
rect 12511 8040 12684 8060
rect 12444 8004 12684 8040
rect 12444 7984 12626 8004
rect 12444 7950 12477 7984
rect 12511 7970 12626 7984
rect 12660 7970 12684 8004
rect 12511 7950 12684 7970
rect 12444 7914 12684 7950
rect 12444 7894 12626 7914
rect 12444 7860 12477 7894
rect 12511 7880 12626 7894
rect 12660 7880 12684 7914
rect 12511 7860 12684 7880
rect 12444 7824 12684 7860
rect 12444 7804 12626 7824
rect 12444 7770 12477 7804
rect 12511 7790 12626 7804
rect 12660 7790 12684 7824
rect 12511 7770 12684 7790
rect 12444 7734 12684 7770
rect 12444 7714 12626 7734
rect 12444 7680 12477 7714
rect 12511 7700 12626 7714
rect 12660 7700 12684 7734
rect 12511 7680 12684 7700
rect 12444 7644 12684 7680
rect 12444 7624 12626 7644
rect 12444 7590 12477 7624
rect 12511 7610 12626 7624
rect 12660 7610 12684 7644
rect 12511 7590 12684 7610
rect 12444 7554 12684 7590
rect 12444 7534 12626 7554
rect 12444 7500 12477 7534
rect 12511 7520 12626 7534
rect 12660 7520 12684 7554
rect 12511 7500 12684 7520
rect 12444 7464 12684 7500
rect 12444 7444 12626 7464
rect 12444 7410 12477 7444
rect 12511 7430 12626 7444
rect 12660 7430 12684 7464
rect 12511 7410 12684 7430
rect 12444 7374 12684 7410
rect 12741 8012 13435 8073
rect 12741 7978 12800 8012
rect 12834 8000 12890 8012
rect 12862 7978 12890 8000
rect 12924 8000 12980 8012
rect 12924 7978 12928 8000
rect 12741 7966 12828 7978
rect 12862 7966 12928 7978
rect 12962 7978 12980 8000
rect 13014 8000 13070 8012
rect 13014 7978 13028 8000
rect 12962 7966 13028 7978
rect 13062 7978 13070 8000
rect 13104 8000 13160 8012
rect 13194 8000 13250 8012
rect 13284 8000 13340 8012
rect 13104 7978 13128 8000
rect 13194 7978 13228 8000
rect 13284 7978 13328 8000
rect 13374 7978 13435 8012
rect 13062 7966 13128 7978
rect 13162 7966 13228 7978
rect 13262 7966 13328 7978
rect 13362 7966 13435 7978
rect 12741 7922 13435 7966
rect 12741 7888 12800 7922
rect 12834 7900 12890 7922
rect 12862 7888 12890 7900
rect 12924 7900 12980 7922
rect 12924 7888 12928 7900
rect 12741 7866 12828 7888
rect 12862 7866 12928 7888
rect 12962 7888 12980 7900
rect 13014 7900 13070 7922
rect 13014 7888 13028 7900
rect 12962 7866 13028 7888
rect 13062 7888 13070 7900
rect 13104 7900 13160 7922
rect 13194 7900 13250 7922
rect 13284 7900 13340 7922
rect 13104 7888 13128 7900
rect 13194 7888 13228 7900
rect 13284 7888 13328 7900
rect 13374 7888 13435 7922
rect 13062 7866 13128 7888
rect 13162 7866 13228 7888
rect 13262 7866 13328 7888
rect 13362 7866 13435 7888
rect 12741 7832 13435 7866
rect 12741 7798 12800 7832
rect 12834 7800 12890 7832
rect 12862 7798 12890 7800
rect 12924 7800 12980 7832
rect 12924 7798 12928 7800
rect 12741 7766 12828 7798
rect 12862 7766 12928 7798
rect 12962 7798 12980 7800
rect 13014 7800 13070 7832
rect 13014 7798 13028 7800
rect 12962 7766 13028 7798
rect 13062 7798 13070 7800
rect 13104 7800 13160 7832
rect 13194 7800 13250 7832
rect 13284 7800 13340 7832
rect 13104 7798 13128 7800
rect 13194 7798 13228 7800
rect 13284 7798 13328 7800
rect 13374 7798 13435 7832
rect 13062 7766 13128 7798
rect 13162 7766 13228 7798
rect 13262 7766 13328 7798
rect 13362 7766 13435 7798
rect 12741 7742 13435 7766
rect 12741 7708 12800 7742
rect 12834 7708 12890 7742
rect 12924 7708 12980 7742
rect 13014 7708 13070 7742
rect 13104 7708 13160 7742
rect 13194 7708 13250 7742
rect 13284 7708 13340 7742
rect 13374 7708 13435 7742
rect 12741 7700 13435 7708
rect 12741 7666 12828 7700
rect 12862 7666 12928 7700
rect 12962 7666 13028 7700
rect 13062 7666 13128 7700
rect 13162 7666 13228 7700
rect 13262 7666 13328 7700
rect 13362 7666 13435 7700
rect 12741 7652 13435 7666
rect 12741 7618 12800 7652
rect 12834 7618 12890 7652
rect 12924 7618 12980 7652
rect 13014 7618 13070 7652
rect 13104 7618 13160 7652
rect 13194 7618 13250 7652
rect 13284 7618 13340 7652
rect 13374 7618 13435 7652
rect 12741 7600 13435 7618
rect 12741 7566 12828 7600
rect 12862 7566 12928 7600
rect 12962 7566 13028 7600
rect 13062 7566 13128 7600
rect 13162 7566 13228 7600
rect 13262 7566 13328 7600
rect 13362 7566 13435 7600
rect 12741 7562 13435 7566
rect 12741 7528 12800 7562
rect 12834 7528 12890 7562
rect 12924 7528 12980 7562
rect 13014 7528 13070 7562
rect 13104 7528 13160 7562
rect 13194 7528 13250 7562
rect 13284 7528 13340 7562
rect 13374 7528 13435 7562
rect 12741 7500 13435 7528
rect 12741 7472 12828 7500
rect 12862 7472 12928 7500
rect 12741 7438 12800 7472
rect 12862 7466 12890 7472
rect 12834 7438 12890 7466
rect 12924 7466 12928 7472
rect 12962 7472 13028 7500
rect 12962 7466 12980 7472
rect 12924 7438 12980 7466
rect 13014 7466 13028 7472
rect 13062 7472 13128 7500
rect 13162 7472 13228 7500
rect 13262 7472 13328 7500
rect 13362 7472 13435 7500
rect 13062 7466 13070 7472
rect 13014 7438 13070 7466
rect 13104 7466 13128 7472
rect 13194 7466 13228 7472
rect 13284 7466 13328 7472
rect 13104 7438 13160 7466
rect 13194 7438 13250 7466
rect 13284 7438 13340 7466
rect 13374 7438 13435 7472
rect 12741 7379 13435 7438
rect 13484 8041 13516 8075
rect 13550 8074 13914 8075
rect 13550 8041 13664 8074
rect 13484 8040 13664 8041
rect 13698 8040 13765 8074
rect 13799 8060 13914 8074
rect 13948 8060 13984 8094
rect 14784 8130 14952 8135
rect 14986 8130 15053 8164
rect 15087 8154 15294 8164
rect 15328 8154 15384 8188
rect 15418 8154 15474 8188
rect 15508 8154 15564 8188
rect 15598 8154 15654 8188
rect 15688 8154 15744 8188
rect 15778 8154 15834 8188
rect 15868 8154 15924 8188
rect 15958 8154 16014 8188
rect 16048 8164 16582 8188
rect 16048 8154 16240 8164
rect 15087 8135 16240 8154
rect 15087 8130 15255 8135
rect 14784 8094 15255 8130
rect 14784 8075 15202 8094
rect 13799 8040 13984 8060
rect 13484 8004 13984 8040
rect 13484 7985 13914 8004
rect 13484 7951 13516 7985
rect 13550 7984 13914 7985
rect 13550 7951 13664 7984
rect 13484 7950 13664 7951
rect 13698 7950 13765 7984
rect 13799 7970 13914 7984
rect 13948 7970 13984 8004
rect 13799 7950 13984 7970
rect 13484 7914 13984 7950
rect 13484 7895 13914 7914
rect 13484 7861 13516 7895
rect 13550 7894 13914 7895
rect 13550 7861 13664 7894
rect 13484 7860 13664 7861
rect 13698 7860 13765 7894
rect 13799 7880 13914 7894
rect 13948 7880 13984 7914
rect 13799 7860 13984 7880
rect 13484 7824 13984 7860
rect 13484 7805 13914 7824
rect 13484 7771 13516 7805
rect 13550 7804 13914 7805
rect 13550 7771 13664 7804
rect 13484 7770 13664 7771
rect 13698 7770 13765 7804
rect 13799 7790 13914 7804
rect 13948 7790 13984 7824
rect 13799 7770 13984 7790
rect 13484 7734 13984 7770
rect 13484 7715 13914 7734
rect 13484 7681 13516 7715
rect 13550 7714 13914 7715
rect 13550 7681 13664 7714
rect 13484 7680 13664 7681
rect 13698 7680 13765 7714
rect 13799 7700 13914 7714
rect 13948 7700 13984 7734
rect 13799 7680 13984 7700
rect 13484 7644 13984 7680
rect 13484 7625 13914 7644
rect 13484 7591 13516 7625
rect 13550 7624 13914 7625
rect 13550 7591 13664 7624
rect 13484 7590 13664 7591
rect 13698 7590 13765 7624
rect 13799 7610 13914 7624
rect 13948 7610 13984 7644
rect 13799 7590 13984 7610
rect 13484 7554 13984 7590
rect 13484 7535 13914 7554
rect 13484 7501 13516 7535
rect 13550 7534 13914 7535
rect 13550 7501 13664 7534
rect 13484 7500 13664 7501
rect 13698 7500 13765 7534
rect 13799 7520 13914 7534
rect 13948 7520 13984 7554
rect 13799 7500 13984 7520
rect 13484 7464 13984 7500
rect 13484 7445 13914 7464
rect 13484 7411 13516 7445
rect 13550 7444 13914 7445
rect 13550 7411 13664 7444
rect 13484 7410 13664 7411
rect 13698 7410 13765 7444
rect 13799 7430 13914 7444
rect 13948 7430 13984 7464
rect 13799 7410 13984 7430
rect 12444 7354 12626 7374
rect 12444 7320 12477 7354
rect 12511 7340 12626 7354
rect 12660 7340 12684 7374
rect 12511 7320 12684 7340
rect 12444 7317 12684 7320
rect 13484 7374 13984 7410
rect 14029 8012 14723 8073
rect 14029 7978 14088 8012
rect 14122 8000 14178 8012
rect 14150 7978 14178 8000
rect 14212 8000 14268 8012
rect 14212 7978 14216 8000
rect 14029 7966 14116 7978
rect 14150 7966 14216 7978
rect 14250 7978 14268 8000
rect 14302 8000 14358 8012
rect 14302 7978 14316 8000
rect 14250 7966 14316 7978
rect 14350 7978 14358 8000
rect 14392 8000 14448 8012
rect 14482 8000 14538 8012
rect 14572 8000 14628 8012
rect 14392 7978 14416 8000
rect 14482 7978 14516 8000
rect 14572 7978 14616 8000
rect 14662 7978 14723 8012
rect 14350 7966 14416 7978
rect 14450 7966 14516 7978
rect 14550 7966 14616 7978
rect 14650 7966 14723 7978
rect 14029 7922 14723 7966
rect 14029 7888 14088 7922
rect 14122 7900 14178 7922
rect 14150 7888 14178 7900
rect 14212 7900 14268 7922
rect 14212 7888 14216 7900
rect 14029 7866 14116 7888
rect 14150 7866 14216 7888
rect 14250 7888 14268 7900
rect 14302 7900 14358 7922
rect 14302 7888 14316 7900
rect 14250 7866 14316 7888
rect 14350 7888 14358 7900
rect 14392 7900 14448 7922
rect 14482 7900 14538 7922
rect 14572 7900 14628 7922
rect 14392 7888 14416 7900
rect 14482 7888 14516 7900
rect 14572 7888 14616 7900
rect 14662 7888 14723 7922
rect 14350 7866 14416 7888
rect 14450 7866 14516 7888
rect 14550 7866 14616 7888
rect 14650 7866 14723 7888
rect 14029 7832 14723 7866
rect 14029 7798 14088 7832
rect 14122 7800 14178 7832
rect 14150 7798 14178 7800
rect 14212 7800 14268 7832
rect 14212 7798 14216 7800
rect 14029 7766 14116 7798
rect 14150 7766 14216 7798
rect 14250 7798 14268 7800
rect 14302 7800 14358 7832
rect 14302 7798 14316 7800
rect 14250 7766 14316 7798
rect 14350 7798 14358 7800
rect 14392 7800 14448 7832
rect 14482 7800 14538 7832
rect 14572 7800 14628 7832
rect 14392 7798 14416 7800
rect 14482 7798 14516 7800
rect 14572 7798 14616 7800
rect 14662 7798 14723 7832
rect 14350 7766 14416 7798
rect 14450 7766 14516 7798
rect 14550 7766 14616 7798
rect 14650 7766 14723 7798
rect 14029 7742 14723 7766
rect 14029 7708 14088 7742
rect 14122 7708 14178 7742
rect 14212 7708 14268 7742
rect 14302 7708 14358 7742
rect 14392 7708 14448 7742
rect 14482 7708 14538 7742
rect 14572 7708 14628 7742
rect 14662 7708 14723 7742
rect 14029 7700 14723 7708
rect 14029 7666 14116 7700
rect 14150 7666 14216 7700
rect 14250 7666 14316 7700
rect 14350 7666 14416 7700
rect 14450 7666 14516 7700
rect 14550 7666 14616 7700
rect 14650 7666 14723 7700
rect 14029 7652 14723 7666
rect 14029 7618 14088 7652
rect 14122 7618 14178 7652
rect 14212 7618 14268 7652
rect 14302 7618 14358 7652
rect 14392 7618 14448 7652
rect 14482 7618 14538 7652
rect 14572 7618 14628 7652
rect 14662 7618 14723 7652
rect 14029 7600 14723 7618
rect 14029 7566 14116 7600
rect 14150 7566 14216 7600
rect 14250 7566 14316 7600
rect 14350 7566 14416 7600
rect 14450 7566 14516 7600
rect 14550 7566 14616 7600
rect 14650 7566 14723 7600
rect 14029 7562 14723 7566
rect 14029 7528 14088 7562
rect 14122 7528 14178 7562
rect 14212 7528 14268 7562
rect 14302 7528 14358 7562
rect 14392 7528 14448 7562
rect 14482 7528 14538 7562
rect 14572 7528 14628 7562
rect 14662 7528 14723 7562
rect 14029 7500 14723 7528
rect 14029 7472 14116 7500
rect 14150 7472 14216 7500
rect 14029 7438 14088 7472
rect 14150 7466 14178 7472
rect 14122 7438 14178 7466
rect 14212 7466 14216 7472
rect 14250 7472 14316 7500
rect 14250 7466 14268 7472
rect 14212 7438 14268 7466
rect 14302 7466 14316 7472
rect 14350 7472 14416 7500
rect 14450 7472 14516 7500
rect 14550 7472 14616 7500
rect 14650 7472 14723 7500
rect 14350 7466 14358 7472
rect 14302 7438 14358 7466
rect 14392 7466 14416 7472
rect 14482 7466 14516 7472
rect 14572 7466 14616 7472
rect 14392 7438 14448 7466
rect 14482 7438 14538 7466
rect 14572 7438 14628 7466
rect 14662 7438 14723 7472
rect 14029 7379 14723 7438
rect 14784 8041 14804 8075
rect 14838 8074 15202 8075
rect 14838 8041 14952 8074
rect 14784 8040 14952 8041
rect 14986 8040 15053 8074
rect 15087 8060 15202 8074
rect 15236 8060 15255 8094
rect 16073 8130 16240 8135
rect 16274 8130 16341 8164
rect 16375 8154 16582 8164
rect 16616 8154 16672 8188
rect 16706 8154 16762 8188
rect 16796 8154 16852 8188
rect 16886 8154 16942 8188
rect 16976 8154 17032 8188
rect 17066 8154 17122 8188
rect 17156 8154 17212 8188
rect 17246 8154 17302 8188
rect 17336 8164 17870 8188
rect 17336 8154 17528 8164
rect 16375 8135 17528 8154
rect 16375 8130 16543 8135
rect 16073 8094 16543 8130
rect 16073 8075 16490 8094
rect 15087 8040 15255 8060
rect 14784 8004 15255 8040
rect 14784 7985 15202 8004
rect 14784 7951 14804 7985
rect 14838 7984 15202 7985
rect 14838 7951 14952 7984
rect 14784 7950 14952 7951
rect 14986 7950 15053 7984
rect 15087 7970 15202 7984
rect 15236 7970 15255 8004
rect 15087 7950 15255 7970
rect 14784 7914 15255 7950
rect 14784 7895 15202 7914
rect 14784 7861 14804 7895
rect 14838 7894 15202 7895
rect 14838 7861 14952 7894
rect 14784 7860 14952 7861
rect 14986 7860 15053 7894
rect 15087 7880 15202 7894
rect 15236 7880 15255 7914
rect 15087 7860 15255 7880
rect 14784 7824 15255 7860
rect 14784 7805 15202 7824
rect 14784 7771 14804 7805
rect 14838 7804 15202 7805
rect 14838 7771 14952 7804
rect 14784 7770 14952 7771
rect 14986 7770 15053 7804
rect 15087 7790 15202 7804
rect 15236 7790 15255 7824
rect 15087 7770 15255 7790
rect 14784 7734 15255 7770
rect 14784 7715 15202 7734
rect 14784 7681 14804 7715
rect 14838 7714 15202 7715
rect 14838 7681 14952 7714
rect 14784 7680 14952 7681
rect 14986 7680 15053 7714
rect 15087 7700 15202 7714
rect 15236 7700 15255 7734
rect 15087 7680 15255 7700
rect 14784 7644 15255 7680
rect 14784 7625 15202 7644
rect 14784 7591 14804 7625
rect 14838 7624 15202 7625
rect 14838 7591 14952 7624
rect 14784 7590 14952 7591
rect 14986 7590 15053 7624
rect 15087 7610 15202 7624
rect 15236 7610 15255 7644
rect 15087 7590 15255 7610
rect 14784 7554 15255 7590
rect 14784 7535 15202 7554
rect 14784 7501 14804 7535
rect 14838 7534 15202 7535
rect 14838 7501 14952 7534
rect 14784 7500 14952 7501
rect 14986 7500 15053 7534
rect 15087 7520 15202 7534
rect 15236 7520 15255 7554
rect 15087 7500 15255 7520
rect 14784 7464 15255 7500
rect 14784 7445 15202 7464
rect 14784 7411 14804 7445
rect 14838 7444 15202 7445
rect 14838 7411 14952 7444
rect 14784 7410 14952 7411
rect 14986 7410 15053 7444
rect 15087 7430 15202 7444
rect 15236 7430 15255 7464
rect 15087 7410 15255 7430
rect 13484 7355 13914 7374
rect 13484 7321 13516 7355
rect 13550 7354 13914 7355
rect 13550 7321 13664 7354
rect 13484 7320 13664 7321
rect 13698 7320 13765 7354
rect 13799 7340 13914 7354
rect 13948 7340 13984 7374
rect 13799 7320 13984 7340
rect 13484 7317 13984 7320
rect 14784 7374 15255 7410
rect 15317 8012 16011 8073
rect 15317 7978 15376 8012
rect 15410 8000 15466 8012
rect 15438 7978 15466 8000
rect 15500 8000 15556 8012
rect 15500 7978 15504 8000
rect 15317 7966 15404 7978
rect 15438 7966 15504 7978
rect 15538 7978 15556 8000
rect 15590 8000 15646 8012
rect 15590 7978 15604 8000
rect 15538 7966 15604 7978
rect 15638 7978 15646 8000
rect 15680 8000 15736 8012
rect 15770 8000 15826 8012
rect 15860 8000 15916 8012
rect 15680 7978 15704 8000
rect 15770 7978 15804 8000
rect 15860 7978 15904 8000
rect 15950 7978 16011 8012
rect 15638 7966 15704 7978
rect 15738 7966 15804 7978
rect 15838 7966 15904 7978
rect 15938 7966 16011 7978
rect 15317 7922 16011 7966
rect 15317 7888 15376 7922
rect 15410 7900 15466 7922
rect 15438 7888 15466 7900
rect 15500 7900 15556 7922
rect 15500 7888 15504 7900
rect 15317 7866 15404 7888
rect 15438 7866 15504 7888
rect 15538 7888 15556 7900
rect 15590 7900 15646 7922
rect 15590 7888 15604 7900
rect 15538 7866 15604 7888
rect 15638 7888 15646 7900
rect 15680 7900 15736 7922
rect 15770 7900 15826 7922
rect 15860 7900 15916 7922
rect 15680 7888 15704 7900
rect 15770 7888 15804 7900
rect 15860 7888 15904 7900
rect 15950 7888 16011 7922
rect 15638 7866 15704 7888
rect 15738 7866 15804 7888
rect 15838 7866 15904 7888
rect 15938 7866 16011 7888
rect 15317 7832 16011 7866
rect 15317 7798 15376 7832
rect 15410 7800 15466 7832
rect 15438 7798 15466 7800
rect 15500 7800 15556 7832
rect 15500 7798 15504 7800
rect 15317 7766 15404 7798
rect 15438 7766 15504 7798
rect 15538 7798 15556 7800
rect 15590 7800 15646 7832
rect 15590 7798 15604 7800
rect 15538 7766 15604 7798
rect 15638 7798 15646 7800
rect 15680 7800 15736 7832
rect 15770 7800 15826 7832
rect 15860 7800 15916 7832
rect 15680 7798 15704 7800
rect 15770 7798 15804 7800
rect 15860 7798 15904 7800
rect 15950 7798 16011 7832
rect 15638 7766 15704 7798
rect 15738 7766 15804 7798
rect 15838 7766 15904 7798
rect 15938 7766 16011 7798
rect 15317 7742 16011 7766
rect 15317 7708 15376 7742
rect 15410 7708 15466 7742
rect 15500 7708 15556 7742
rect 15590 7708 15646 7742
rect 15680 7708 15736 7742
rect 15770 7708 15826 7742
rect 15860 7708 15916 7742
rect 15950 7708 16011 7742
rect 15317 7700 16011 7708
rect 15317 7666 15404 7700
rect 15438 7666 15504 7700
rect 15538 7666 15604 7700
rect 15638 7666 15704 7700
rect 15738 7666 15804 7700
rect 15838 7666 15904 7700
rect 15938 7666 16011 7700
rect 15317 7652 16011 7666
rect 15317 7618 15376 7652
rect 15410 7618 15466 7652
rect 15500 7618 15556 7652
rect 15590 7618 15646 7652
rect 15680 7618 15736 7652
rect 15770 7618 15826 7652
rect 15860 7618 15916 7652
rect 15950 7618 16011 7652
rect 15317 7600 16011 7618
rect 15317 7566 15404 7600
rect 15438 7566 15504 7600
rect 15538 7566 15604 7600
rect 15638 7566 15704 7600
rect 15738 7566 15804 7600
rect 15838 7566 15904 7600
rect 15938 7566 16011 7600
rect 15317 7562 16011 7566
rect 15317 7528 15376 7562
rect 15410 7528 15466 7562
rect 15500 7528 15556 7562
rect 15590 7528 15646 7562
rect 15680 7528 15736 7562
rect 15770 7528 15826 7562
rect 15860 7528 15916 7562
rect 15950 7528 16011 7562
rect 15317 7500 16011 7528
rect 15317 7472 15404 7500
rect 15438 7472 15504 7500
rect 15317 7438 15376 7472
rect 15438 7466 15466 7472
rect 15410 7438 15466 7466
rect 15500 7466 15504 7472
rect 15538 7472 15604 7500
rect 15538 7466 15556 7472
rect 15500 7438 15556 7466
rect 15590 7466 15604 7472
rect 15638 7472 15704 7500
rect 15738 7472 15804 7500
rect 15838 7472 15904 7500
rect 15938 7472 16011 7500
rect 15638 7466 15646 7472
rect 15590 7438 15646 7466
rect 15680 7466 15704 7472
rect 15770 7466 15804 7472
rect 15860 7466 15904 7472
rect 15680 7438 15736 7466
rect 15770 7438 15826 7466
rect 15860 7438 15916 7466
rect 15950 7438 16011 7472
rect 15317 7379 16011 7438
rect 16073 8041 16092 8075
rect 16126 8074 16490 8075
rect 16126 8041 16240 8074
rect 16073 8040 16240 8041
rect 16274 8040 16341 8074
rect 16375 8060 16490 8074
rect 16524 8060 16543 8094
rect 17361 8130 17528 8135
rect 17562 8130 17629 8164
rect 17663 8154 17870 8164
rect 17904 8154 17960 8188
rect 17994 8154 18050 8188
rect 18084 8154 18140 8188
rect 18174 8154 18230 8188
rect 18264 8154 18320 8188
rect 18354 8154 18410 8188
rect 18444 8154 18500 8188
rect 18534 8154 18590 8188
rect 18624 8164 18884 8188
rect 18624 8154 18816 8164
rect 17663 8135 18816 8154
rect 17663 8130 17831 8135
rect 17361 8094 17831 8130
rect 17361 8075 17778 8094
rect 16375 8040 16543 8060
rect 16073 8004 16543 8040
rect 16073 7985 16490 8004
rect 16073 7951 16092 7985
rect 16126 7984 16490 7985
rect 16126 7951 16240 7984
rect 16073 7950 16240 7951
rect 16274 7950 16341 7984
rect 16375 7970 16490 7984
rect 16524 7970 16543 8004
rect 16375 7950 16543 7970
rect 16073 7914 16543 7950
rect 16073 7895 16490 7914
rect 16073 7861 16092 7895
rect 16126 7894 16490 7895
rect 16126 7861 16240 7894
rect 16073 7860 16240 7861
rect 16274 7860 16341 7894
rect 16375 7880 16490 7894
rect 16524 7880 16543 7914
rect 16375 7860 16543 7880
rect 16073 7824 16543 7860
rect 16073 7805 16490 7824
rect 16073 7771 16092 7805
rect 16126 7804 16490 7805
rect 16126 7771 16240 7804
rect 16073 7770 16240 7771
rect 16274 7770 16341 7804
rect 16375 7790 16490 7804
rect 16524 7790 16543 7824
rect 16375 7770 16543 7790
rect 16073 7734 16543 7770
rect 16073 7715 16490 7734
rect 16073 7681 16092 7715
rect 16126 7714 16490 7715
rect 16126 7681 16240 7714
rect 16073 7680 16240 7681
rect 16274 7680 16341 7714
rect 16375 7700 16490 7714
rect 16524 7700 16543 7734
rect 16375 7680 16543 7700
rect 16073 7644 16543 7680
rect 16073 7625 16490 7644
rect 16073 7591 16092 7625
rect 16126 7624 16490 7625
rect 16126 7591 16240 7624
rect 16073 7590 16240 7591
rect 16274 7590 16341 7624
rect 16375 7610 16490 7624
rect 16524 7610 16543 7644
rect 16375 7590 16543 7610
rect 16073 7554 16543 7590
rect 16073 7535 16490 7554
rect 16073 7501 16092 7535
rect 16126 7534 16490 7535
rect 16126 7501 16240 7534
rect 16073 7500 16240 7501
rect 16274 7500 16341 7534
rect 16375 7520 16490 7534
rect 16524 7520 16543 7554
rect 16375 7500 16543 7520
rect 16073 7464 16543 7500
rect 16073 7445 16490 7464
rect 16073 7411 16092 7445
rect 16126 7444 16490 7445
rect 16126 7411 16240 7444
rect 16073 7410 16240 7411
rect 16274 7410 16341 7444
rect 16375 7430 16490 7444
rect 16524 7430 16543 7464
rect 16375 7410 16543 7430
rect 14784 7355 15202 7374
rect 14784 7321 14804 7355
rect 14838 7354 15202 7355
rect 14838 7321 14952 7354
rect 14784 7320 14952 7321
rect 14986 7320 15053 7354
rect 15087 7340 15202 7354
rect 15236 7340 15255 7374
rect 15087 7320 15255 7340
rect 14784 7317 15255 7320
rect 16073 7374 16543 7410
rect 16605 8012 17299 8073
rect 16605 7978 16664 8012
rect 16698 8000 16754 8012
rect 16726 7978 16754 8000
rect 16788 8000 16844 8012
rect 16788 7978 16792 8000
rect 16605 7966 16692 7978
rect 16726 7966 16792 7978
rect 16826 7978 16844 8000
rect 16878 8000 16934 8012
rect 16878 7978 16892 8000
rect 16826 7966 16892 7978
rect 16926 7978 16934 8000
rect 16968 8000 17024 8012
rect 17058 8000 17114 8012
rect 17148 8000 17204 8012
rect 16968 7978 16992 8000
rect 17058 7978 17092 8000
rect 17148 7978 17192 8000
rect 17238 7978 17299 8012
rect 16926 7966 16992 7978
rect 17026 7966 17092 7978
rect 17126 7966 17192 7978
rect 17226 7966 17299 7978
rect 16605 7922 17299 7966
rect 16605 7888 16664 7922
rect 16698 7900 16754 7922
rect 16726 7888 16754 7900
rect 16788 7900 16844 7922
rect 16788 7888 16792 7900
rect 16605 7866 16692 7888
rect 16726 7866 16792 7888
rect 16826 7888 16844 7900
rect 16878 7900 16934 7922
rect 16878 7888 16892 7900
rect 16826 7866 16892 7888
rect 16926 7888 16934 7900
rect 16968 7900 17024 7922
rect 17058 7900 17114 7922
rect 17148 7900 17204 7922
rect 16968 7888 16992 7900
rect 17058 7888 17092 7900
rect 17148 7888 17192 7900
rect 17238 7888 17299 7922
rect 16926 7866 16992 7888
rect 17026 7866 17092 7888
rect 17126 7866 17192 7888
rect 17226 7866 17299 7888
rect 16605 7832 17299 7866
rect 16605 7798 16664 7832
rect 16698 7800 16754 7832
rect 16726 7798 16754 7800
rect 16788 7800 16844 7832
rect 16788 7798 16792 7800
rect 16605 7766 16692 7798
rect 16726 7766 16792 7798
rect 16826 7798 16844 7800
rect 16878 7800 16934 7832
rect 16878 7798 16892 7800
rect 16826 7766 16892 7798
rect 16926 7798 16934 7800
rect 16968 7800 17024 7832
rect 17058 7800 17114 7832
rect 17148 7800 17204 7832
rect 16968 7798 16992 7800
rect 17058 7798 17092 7800
rect 17148 7798 17192 7800
rect 17238 7798 17299 7832
rect 16926 7766 16992 7798
rect 17026 7766 17092 7798
rect 17126 7766 17192 7798
rect 17226 7766 17299 7798
rect 16605 7742 17299 7766
rect 16605 7708 16664 7742
rect 16698 7708 16754 7742
rect 16788 7708 16844 7742
rect 16878 7708 16934 7742
rect 16968 7708 17024 7742
rect 17058 7708 17114 7742
rect 17148 7708 17204 7742
rect 17238 7708 17299 7742
rect 16605 7700 17299 7708
rect 16605 7666 16692 7700
rect 16726 7666 16792 7700
rect 16826 7666 16892 7700
rect 16926 7666 16992 7700
rect 17026 7666 17092 7700
rect 17126 7666 17192 7700
rect 17226 7666 17299 7700
rect 16605 7652 17299 7666
rect 16605 7618 16664 7652
rect 16698 7618 16754 7652
rect 16788 7618 16844 7652
rect 16878 7618 16934 7652
rect 16968 7618 17024 7652
rect 17058 7618 17114 7652
rect 17148 7618 17204 7652
rect 17238 7618 17299 7652
rect 16605 7600 17299 7618
rect 16605 7566 16692 7600
rect 16726 7566 16792 7600
rect 16826 7566 16892 7600
rect 16926 7566 16992 7600
rect 17026 7566 17092 7600
rect 17126 7566 17192 7600
rect 17226 7566 17299 7600
rect 16605 7562 17299 7566
rect 16605 7528 16664 7562
rect 16698 7528 16754 7562
rect 16788 7528 16844 7562
rect 16878 7528 16934 7562
rect 16968 7528 17024 7562
rect 17058 7528 17114 7562
rect 17148 7528 17204 7562
rect 17238 7528 17299 7562
rect 16605 7500 17299 7528
rect 16605 7472 16692 7500
rect 16726 7472 16792 7500
rect 16605 7438 16664 7472
rect 16726 7466 16754 7472
rect 16698 7438 16754 7466
rect 16788 7466 16792 7472
rect 16826 7472 16892 7500
rect 16826 7466 16844 7472
rect 16788 7438 16844 7466
rect 16878 7466 16892 7472
rect 16926 7472 16992 7500
rect 17026 7472 17092 7500
rect 17126 7472 17192 7500
rect 17226 7472 17299 7500
rect 16926 7466 16934 7472
rect 16878 7438 16934 7466
rect 16968 7466 16992 7472
rect 17058 7466 17092 7472
rect 17148 7466 17192 7472
rect 16968 7438 17024 7466
rect 17058 7438 17114 7466
rect 17148 7438 17204 7466
rect 17238 7438 17299 7472
rect 16605 7379 17299 7438
rect 17361 8041 17380 8075
rect 17414 8074 17778 8075
rect 17414 8041 17528 8074
rect 17361 8040 17528 8041
rect 17562 8040 17629 8074
rect 17663 8060 17778 8074
rect 17812 8060 17831 8094
rect 18649 8130 18816 8135
rect 18850 8130 18884 8164
rect 18649 8075 18884 8130
rect 17663 8040 17831 8060
rect 17361 8004 17831 8040
rect 17361 7985 17778 8004
rect 17361 7951 17380 7985
rect 17414 7984 17778 7985
rect 17414 7951 17528 7984
rect 17361 7950 17528 7951
rect 17562 7950 17629 7984
rect 17663 7970 17778 7984
rect 17812 7970 17831 8004
rect 17663 7950 17831 7970
rect 17361 7914 17831 7950
rect 17361 7895 17778 7914
rect 17361 7861 17380 7895
rect 17414 7894 17778 7895
rect 17414 7861 17528 7894
rect 17361 7860 17528 7861
rect 17562 7860 17629 7894
rect 17663 7880 17778 7894
rect 17812 7880 17831 7914
rect 17663 7860 17831 7880
rect 17361 7824 17831 7860
rect 17361 7805 17778 7824
rect 17361 7771 17380 7805
rect 17414 7804 17778 7805
rect 17414 7771 17528 7804
rect 17361 7770 17528 7771
rect 17562 7770 17629 7804
rect 17663 7790 17778 7804
rect 17812 7790 17831 7824
rect 17663 7770 17831 7790
rect 17361 7734 17831 7770
rect 17361 7715 17778 7734
rect 17361 7681 17380 7715
rect 17414 7714 17778 7715
rect 17414 7681 17528 7714
rect 17361 7680 17528 7681
rect 17562 7680 17629 7714
rect 17663 7700 17778 7714
rect 17812 7700 17831 7734
rect 17663 7680 17831 7700
rect 17361 7644 17831 7680
rect 17361 7625 17778 7644
rect 17361 7591 17380 7625
rect 17414 7624 17778 7625
rect 17414 7591 17528 7624
rect 17361 7590 17528 7591
rect 17562 7590 17629 7624
rect 17663 7610 17778 7624
rect 17812 7610 17831 7644
rect 17663 7590 17831 7610
rect 17361 7554 17831 7590
rect 17361 7535 17778 7554
rect 17361 7501 17380 7535
rect 17414 7534 17778 7535
rect 17414 7501 17528 7534
rect 17361 7500 17528 7501
rect 17562 7500 17629 7534
rect 17663 7520 17778 7534
rect 17812 7520 17831 7554
rect 17663 7500 17831 7520
rect 17361 7464 17831 7500
rect 17361 7445 17778 7464
rect 17361 7411 17380 7445
rect 17414 7444 17778 7445
rect 17414 7411 17528 7444
rect 17361 7410 17528 7411
rect 17562 7410 17629 7444
rect 17663 7430 17778 7444
rect 17812 7430 17831 7464
rect 17663 7410 17831 7430
rect 16073 7355 16490 7374
rect 16073 7321 16092 7355
rect 16126 7354 16490 7355
rect 16126 7321 16240 7354
rect 16073 7320 16240 7321
rect 16274 7320 16341 7354
rect 16375 7340 16490 7354
rect 16524 7340 16543 7374
rect 16375 7320 16543 7340
rect 16073 7317 16543 7320
rect 17361 7374 17831 7410
rect 17893 8012 18587 8073
rect 17893 7978 17952 8012
rect 17986 8000 18042 8012
rect 18014 7978 18042 8000
rect 18076 8000 18132 8012
rect 18076 7978 18080 8000
rect 17893 7966 17980 7978
rect 18014 7966 18080 7978
rect 18114 7978 18132 8000
rect 18166 8000 18222 8012
rect 18166 7978 18180 8000
rect 18114 7966 18180 7978
rect 18214 7978 18222 8000
rect 18256 8000 18312 8012
rect 18346 8000 18402 8012
rect 18436 8000 18492 8012
rect 18256 7978 18280 8000
rect 18346 7978 18380 8000
rect 18436 7978 18480 8000
rect 18526 7978 18587 8012
rect 18214 7966 18280 7978
rect 18314 7966 18380 7978
rect 18414 7966 18480 7978
rect 18514 7966 18587 7978
rect 17893 7922 18587 7966
rect 17893 7888 17952 7922
rect 17986 7900 18042 7922
rect 18014 7888 18042 7900
rect 18076 7900 18132 7922
rect 18076 7888 18080 7900
rect 17893 7866 17980 7888
rect 18014 7866 18080 7888
rect 18114 7888 18132 7900
rect 18166 7900 18222 7922
rect 18166 7888 18180 7900
rect 18114 7866 18180 7888
rect 18214 7888 18222 7900
rect 18256 7900 18312 7922
rect 18346 7900 18402 7922
rect 18436 7900 18492 7922
rect 18256 7888 18280 7900
rect 18346 7888 18380 7900
rect 18436 7888 18480 7900
rect 18526 7888 18587 7922
rect 18214 7866 18280 7888
rect 18314 7866 18380 7888
rect 18414 7866 18480 7888
rect 18514 7866 18587 7888
rect 17893 7832 18587 7866
rect 17893 7798 17952 7832
rect 17986 7800 18042 7832
rect 18014 7798 18042 7800
rect 18076 7800 18132 7832
rect 18076 7798 18080 7800
rect 17893 7766 17980 7798
rect 18014 7766 18080 7798
rect 18114 7798 18132 7800
rect 18166 7800 18222 7832
rect 18166 7798 18180 7800
rect 18114 7766 18180 7798
rect 18214 7798 18222 7800
rect 18256 7800 18312 7832
rect 18346 7800 18402 7832
rect 18436 7800 18492 7832
rect 18256 7798 18280 7800
rect 18346 7798 18380 7800
rect 18436 7798 18480 7800
rect 18526 7798 18587 7832
rect 18214 7766 18280 7798
rect 18314 7766 18380 7798
rect 18414 7766 18480 7798
rect 18514 7766 18587 7798
rect 17893 7742 18587 7766
rect 17893 7708 17952 7742
rect 17986 7708 18042 7742
rect 18076 7708 18132 7742
rect 18166 7708 18222 7742
rect 18256 7708 18312 7742
rect 18346 7708 18402 7742
rect 18436 7708 18492 7742
rect 18526 7708 18587 7742
rect 17893 7700 18587 7708
rect 17893 7666 17980 7700
rect 18014 7666 18080 7700
rect 18114 7666 18180 7700
rect 18214 7666 18280 7700
rect 18314 7666 18380 7700
rect 18414 7666 18480 7700
rect 18514 7666 18587 7700
rect 17893 7652 18587 7666
rect 17893 7618 17952 7652
rect 17986 7618 18042 7652
rect 18076 7618 18132 7652
rect 18166 7618 18222 7652
rect 18256 7618 18312 7652
rect 18346 7618 18402 7652
rect 18436 7618 18492 7652
rect 18526 7618 18587 7652
rect 17893 7600 18587 7618
rect 17893 7566 17980 7600
rect 18014 7566 18080 7600
rect 18114 7566 18180 7600
rect 18214 7566 18280 7600
rect 18314 7566 18380 7600
rect 18414 7566 18480 7600
rect 18514 7566 18587 7600
rect 17893 7562 18587 7566
rect 17893 7528 17952 7562
rect 17986 7528 18042 7562
rect 18076 7528 18132 7562
rect 18166 7528 18222 7562
rect 18256 7528 18312 7562
rect 18346 7528 18402 7562
rect 18436 7528 18492 7562
rect 18526 7528 18587 7562
rect 17893 7500 18587 7528
rect 17893 7472 17980 7500
rect 18014 7472 18080 7500
rect 17893 7438 17952 7472
rect 18014 7466 18042 7472
rect 17986 7438 18042 7466
rect 18076 7466 18080 7472
rect 18114 7472 18180 7500
rect 18114 7466 18132 7472
rect 18076 7438 18132 7466
rect 18166 7466 18180 7472
rect 18214 7472 18280 7500
rect 18314 7472 18380 7500
rect 18414 7472 18480 7500
rect 18514 7472 18587 7500
rect 18214 7466 18222 7472
rect 18166 7438 18222 7466
rect 18256 7466 18280 7472
rect 18346 7466 18380 7472
rect 18436 7466 18480 7472
rect 18256 7438 18312 7466
rect 18346 7438 18402 7466
rect 18436 7438 18492 7466
rect 18526 7438 18587 7472
rect 17893 7379 18587 7438
rect 18649 8041 18668 8075
rect 18702 8074 18884 8075
rect 18702 8041 18816 8074
rect 18649 8040 18816 8041
rect 18850 8040 18884 8074
rect 18649 7985 18884 8040
rect 18649 7951 18668 7985
rect 18702 7984 18884 7985
rect 18702 7951 18816 7984
rect 18649 7950 18816 7951
rect 18850 7950 18884 7984
rect 18649 7895 18884 7950
rect 18649 7861 18668 7895
rect 18702 7894 18884 7895
rect 18702 7861 18816 7894
rect 18649 7860 18816 7861
rect 18850 7860 18884 7894
rect 18649 7805 18884 7860
rect 18649 7771 18668 7805
rect 18702 7804 18884 7805
rect 18702 7771 18816 7804
rect 18649 7770 18816 7771
rect 18850 7770 18884 7804
rect 18649 7715 18884 7770
rect 18649 7681 18668 7715
rect 18702 7714 18884 7715
rect 18702 7681 18816 7714
rect 18649 7680 18816 7681
rect 18850 7680 18884 7714
rect 18649 7625 18884 7680
rect 18649 7591 18668 7625
rect 18702 7624 18884 7625
rect 18702 7591 18816 7624
rect 18649 7590 18816 7591
rect 18850 7590 18884 7624
rect 18649 7535 18884 7590
rect 18649 7501 18668 7535
rect 18702 7534 18884 7535
rect 18702 7501 18816 7534
rect 18649 7500 18816 7501
rect 18850 7500 18884 7534
rect 18649 7445 18884 7500
rect 18649 7411 18668 7445
rect 18702 7444 18884 7445
rect 18702 7411 18816 7444
rect 18649 7410 18816 7411
rect 18850 7410 18884 7444
rect 17361 7355 17778 7374
rect 17361 7321 17380 7355
rect 17414 7354 17778 7355
rect 17414 7321 17528 7354
rect 17361 7320 17528 7321
rect 17562 7320 17629 7354
rect 17663 7340 17778 7354
rect 17812 7340 17831 7374
rect 17663 7320 17831 7340
rect 17361 7317 17831 7320
rect 18649 7355 18884 7410
rect 18649 7321 18668 7355
rect 18702 7354 18884 7355
rect 18702 7321 18816 7354
rect 18649 7320 18816 7321
rect 18850 7320 18884 7354
rect 18649 7317 18884 7320
rect 12444 7298 18884 7317
rect 12444 7264 12684 7298
rect 12718 7264 12774 7298
rect 12808 7264 12864 7298
rect 12898 7264 12954 7298
rect 12988 7264 13044 7298
rect 13078 7264 13134 7298
rect 13168 7264 13224 7298
rect 13258 7264 13314 7298
rect 13348 7264 13404 7298
rect 13438 7264 13972 7298
rect 14006 7264 14062 7298
rect 14096 7264 14152 7298
rect 14186 7264 14242 7298
rect 14276 7264 14332 7298
rect 14366 7264 14422 7298
rect 14456 7264 14512 7298
rect 14546 7264 14602 7298
rect 14636 7264 14692 7298
rect 14726 7264 15260 7298
rect 15294 7264 15350 7298
rect 15384 7264 15440 7298
rect 15474 7264 15530 7298
rect 15564 7264 15620 7298
rect 15654 7264 15710 7298
rect 15744 7264 15800 7298
rect 15834 7264 15890 7298
rect 15924 7264 15980 7298
rect 16014 7264 16548 7298
rect 16582 7264 16638 7298
rect 16672 7264 16728 7298
rect 16762 7264 16818 7298
rect 16852 7264 16908 7298
rect 16942 7264 16998 7298
rect 17032 7264 17088 7298
rect 17122 7264 17178 7298
rect 17212 7264 17268 7298
rect 17302 7264 17836 7298
rect 17870 7264 17926 7298
rect 17960 7264 18016 7298
rect 18050 7264 18106 7298
rect 18140 7264 18196 7298
rect 18230 7264 18286 7298
rect 18320 7264 18376 7298
rect 18410 7264 18466 7298
rect 18500 7264 18556 7298
rect 18590 7264 18884 7298
rect 12444 7230 12477 7264
rect 12511 7245 13664 7264
rect 12511 7230 12684 7245
rect 12444 7181 12684 7230
rect 13484 7230 13664 7245
rect 13698 7230 13765 7264
rect 13799 7245 14952 7264
rect 13799 7230 13984 7245
rect 13484 7181 13984 7230
rect 14784 7230 14952 7245
rect 14986 7230 15053 7264
rect 15087 7245 16240 7264
rect 15087 7230 15184 7245
rect 14784 7181 15184 7230
rect 16084 7230 16240 7245
rect 16274 7230 16341 7264
rect 16375 7245 17528 7264
rect 16375 7230 16484 7245
rect 16084 7181 16484 7230
rect 17384 7230 17528 7245
rect 17562 7230 17629 7264
rect 17663 7245 18816 7264
rect 17663 7230 17784 7245
rect 17384 7181 17784 7230
rect 18684 7230 18816 7245
rect 18850 7230 18884 7264
rect 18684 7181 18884 7230
rect 12444 7174 18884 7181
rect 12444 7140 12477 7174
rect 12511 7151 13664 7174
rect 12511 7140 12578 7151
rect 12444 7117 12578 7140
rect 12612 7117 12668 7151
rect 12702 7117 12758 7151
rect 12792 7117 12848 7151
rect 12882 7117 12938 7151
rect 12972 7117 13028 7151
rect 13062 7117 13118 7151
rect 13152 7117 13208 7151
rect 13242 7117 13298 7151
rect 13332 7117 13388 7151
rect 13422 7117 13478 7151
rect 13512 7117 13568 7151
rect 13602 7140 13664 7151
rect 13698 7140 13765 7174
rect 13799 7151 14952 7174
rect 13799 7140 13866 7151
rect 13602 7117 13866 7140
rect 13900 7117 13956 7151
rect 13990 7117 14046 7151
rect 14080 7117 14136 7151
rect 14170 7117 14226 7151
rect 14260 7117 14316 7151
rect 14350 7117 14406 7151
rect 14440 7117 14496 7151
rect 14530 7117 14586 7151
rect 14620 7117 14676 7151
rect 14710 7117 14766 7151
rect 14800 7117 14856 7151
rect 14890 7140 14952 7151
rect 14986 7140 15053 7174
rect 15087 7151 16240 7174
rect 15087 7140 15154 7151
rect 14890 7117 15154 7140
rect 15188 7117 15244 7151
rect 15278 7117 15334 7151
rect 15368 7117 15424 7151
rect 15458 7117 15514 7151
rect 15548 7117 15604 7151
rect 15638 7117 15694 7151
rect 15728 7117 15784 7151
rect 15818 7117 15874 7151
rect 15908 7117 15964 7151
rect 15998 7117 16054 7151
rect 16088 7117 16144 7151
rect 16178 7140 16240 7151
rect 16274 7140 16341 7174
rect 16375 7151 17528 7174
rect 16375 7140 16442 7151
rect 16178 7117 16442 7140
rect 16476 7117 16532 7151
rect 16566 7117 16622 7151
rect 16656 7117 16712 7151
rect 16746 7117 16802 7151
rect 16836 7117 16892 7151
rect 16926 7117 16982 7151
rect 17016 7117 17072 7151
rect 17106 7117 17162 7151
rect 17196 7117 17252 7151
rect 17286 7117 17342 7151
rect 17376 7117 17432 7151
rect 17466 7140 17528 7151
rect 17562 7140 17629 7174
rect 17663 7151 18816 7174
rect 17663 7140 17730 7151
rect 17466 7117 17730 7140
rect 17764 7117 17820 7151
rect 17854 7117 17910 7151
rect 17944 7117 18000 7151
rect 18034 7117 18090 7151
rect 18124 7117 18180 7151
rect 18214 7117 18270 7151
rect 18304 7117 18360 7151
rect 18394 7117 18450 7151
rect 18484 7117 18540 7151
rect 18574 7117 18630 7151
rect 18664 7117 18720 7151
rect 18754 7140 18816 7151
rect 18850 7140 18884 7174
rect 18754 7117 18884 7140
rect 12444 7050 18884 7117
rect 12444 7016 12578 7050
rect 12612 7016 12668 7050
rect 12702 7016 12758 7050
rect 12792 7016 12848 7050
rect 12882 7016 12938 7050
rect 12972 7016 13028 7050
rect 13062 7016 13118 7050
rect 13152 7016 13208 7050
rect 13242 7016 13298 7050
rect 13332 7016 13388 7050
rect 13422 7016 13478 7050
rect 13512 7016 13568 7050
rect 13602 7016 13866 7050
rect 13900 7016 13956 7050
rect 13990 7016 14046 7050
rect 14080 7016 14136 7050
rect 14170 7016 14226 7050
rect 14260 7016 14316 7050
rect 14350 7016 14406 7050
rect 14440 7016 14496 7050
rect 14530 7016 14586 7050
rect 14620 7016 14676 7050
rect 14710 7016 14766 7050
rect 14800 7016 14856 7050
rect 14890 7016 15154 7050
rect 15188 7016 15244 7050
rect 15278 7016 15334 7050
rect 15368 7016 15424 7050
rect 15458 7016 15514 7050
rect 15548 7016 15604 7050
rect 15638 7016 15694 7050
rect 15728 7016 15784 7050
rect 15818 7016 15874 7050
rect 15908 7016 15964 7050
rect 15998 7016 16054 7050
rect 16088 7016 16144 7050
rect 16178 7016 16442 7050
rect 16476 7016 16532 7050
rect 16566 7016 16622 7050
rect 16656 7016 16712 7050
rect 16746 7016 16802 7050
rect 16836 7016 16892 7050
rect 16926 7016 16982 7050
rect 17016 7016 17072 7050
rect 17106 7016 17162 7050
rect 17196 7016 17252 7050
rect 17286 7016 17342 7050
rect 17376 7016 17432 7050
rect 17466 7016 17730 7050
rect 17764 7016 17820 7050
rect 17854 7016 17910 7050
rect 17944 7016 18000 7050
rect 18034 7016 18090 7050
rect 18124 7016 18180 7050
rect 18214 7016 18270 7050
rect 18304 7016 18360 7050
rect 18394 7016 18450 7050
rect 18484 7016 18540 7050
rect 18574 7016 18630 7050
rect 18664 7016 18720 7050
rect 18754 7016 18884 7050
rect 12444 6983 18884 7016
rect 12444 6966 12684 6983
rect 12444 6932 12477 6966
rect 12511 6932 12684 6966
rect 12444 6919 12684 6932
rect 13484 6966 13984 6983
rect 13484 6932 13664 6966
rect 13698 6932 13765 6966
rect 13799 6932 13984 6966
rect 13484 6919 13984 6932
rect 14784 6966 15184 6983
rect 14784 6932 14952 6966
rect 14986 6932 15053 6966
rect 15087 6932 15184 6966
rect 14784 6919 15184 6932
rect 16084 6966 16484 6983
rect 16084 6932 16240 6966
rect 16274 6932 16341 6966
rect 16375 6932 16484 6966
rect 16084 6919 16484 6932
rect 17384 6966 17784 6983
rect 17384 6932 17528 6966
rect 17562 6932 17629 6966
rect 17663 6932 17784 6966
rect 17384 6919 17784 6932
rect 18684 6966 18884 6983
rect 18684 6932 18816 6966
rect 18850 6932 18884 6966
rect 18684 6919 18884 6932
rect 12444 6900 18884 6919
rect 12444 6876 12718 6900
rect 12444 6842 12477 6876
rect 12511 6866 12718 6876
rect 12752 6866 12808 6900
rect 12842 6866 12898 6900
rect 12932 6866 12988 6900
rect 13022 6866 13078 6900
rect 13112 6866 13168 6900
rect 13202 6866 13258 6900
rect 13292 6866 13348 6900
rect 13382 6866 13438 6900
rect 13472 6876 14006 6900
rect 13472 6866 13664 6876
rect 12511 6847 13664 6866
rect 12511 6842 12684 6847
rect 12444 6806 12684 6842
rect 12444 6786 12626 6806
rect 12444 6752 12477 6786
rect 12511 6772 12626 6786
rect 12660 6772 12684 6806
rect 13484 6842 13664 6847
rect 13698 6842 13765 6876
rect 13799 6866 14006 6876
rect 14040 6866 14096 6900
rect 14130 6866 14186 6900
rect 14220 6866 14276 6900
rect 14310 6866 14366 6900
rect 14400 6866 14456 6900
rect 14490 6866 14546 6900
rect 14580 6866 14636 6900
rect 14670 6866 14726 6900
rect 14760 6876 15294 6900
rect 14760 6866 14952 6876
rect 13799 6847 14952 6866
rect 13799 6842 13984 6847
rect 13484 6806 13984 6842
rect 13484 6787 13914 6806
rect 12511 6752 12684 6772
rect 12444 6716 12684 6752
rect 12444 6696 12626 6716
rect 12444 6662 12477 6696
rect 12511 6682 12626 6696
rect 12660 6682 12684 6716
rect 12511 6662 12684 6682
rect 12444 6626 12684 6662
rect 12444 6606 12626 6626
rect 12444 6572 12477 6606
rect 12511 6592 12626 6606
rect 12660 6592 12684 6626
rect 12511 6572 12684 6592
rect 12444 6536 12684 6572
rect 12444 6516 12626 6536
rect 12444 6482 12477 6516
rect 12511 6502 12626 6516
rect 12660 6502 12684 6536
rect 12511 6482 12684 6502
rect 12444 6446 12684 6482
rect 12444 6426 12626 6446
rect 12444 6392 12477 6426
rect 12511 6412 12626 6426
rect 12660 6412 12684 6446
rect 12511 6392 12684 6412
rect 12444 6356 12684 6392
rect 12444 6336 12626 6356
rect 12444 6302 12477 6336
rect 12511 6322 12626 6336
rect 12660 6322 12684 6356
rect 12511 6302 12684 6322
rect 12444 6266 12684 6302
rect 12444 6246 12626 6266
rect 12444 6212 12477 6246
rect 12511 6232 12626 6246
rect 12660 6232 12684 6266
rect 12511 6212 12684 6232
rect 12444 6176 12684 6212
rect 12444 6156 12626 6176
rect 12444 6122 12477 6156
rect 12511 6142 12626 6156
rect 12660 6142 12684 6176
rect 12511 6122 12684 6142
rect 12444 6086 12684 6122
rect 12741 6724 13435 6785
rect 12741 6690 12800 6724
rect 12834 6712 12890 6724
rect 12862 6690 12890 6712
rect 12924 6712 12980 6724
rect 12924 6690 12928 6712
rect 12741 6678 12828 6690
rect 12862 6678 12928 6690
rect 12962 6690 12980 6712
rect 13014 6712 13070 6724
rect 13014 6690 13028 6712
rect 12962 6678 13028 6690
rect 13062 6690 13070 6712
rect 13104 6712 13160 6724
rect 13194 6712 13250 6724
rect 13284 6712 13340 6724
rect 13104 6690 13128 6712
rect 13194 6690 13228 6712
rect 13284 6690 13328 6712
rect 13374 6690 13435 6724
rect 13062 6678 13128 6690
rect 13162 6678 13228 6690
rect 13262 6678 13328 6690
rect 13362 6678 13435 6690
rect 12741 6634 13435 6678
rect 12741 6600 12800 6634
rect 12834 6612 12890 6634
rect 12862 6600 12890 6612
rect 12924 6612 12980 6634
rect 12924 6600 12928 6612
rect 12741 6578 12828 6600
rect 12862 6578 12928 6600
rect 12962 6600 12980 6612
rect 13014 6612 13070 6634
rect 13014 6600 13028 6612
rect 12962 6578 13028 6600
rect 13062 6600 13070 6612
rect 13104 6612 13160 6634
rect 13194 6612 13250 6634
rect 13284 6612 13340 6634
rect 13104 6600 13128 6612
rect 13194 6600 13228 6612
rect 13284 6600 13328 6612
rect 13374 6600 13435 6634
rect 13062 6578 13128 6600
rect 13162 6578 13228 6600
rect 13262 6578 13328 6600
rect 13362 6578 13435 6600
rect 12741 6544 13435 6578
rect 12741 6510 12800 6544
rect 12834 6512 12890 6544
rect 12862 6510 12890 6512
rect 12924 6512 12980 6544
rect 12924 6510 12928 6512
rect 12741 6478 12828 6510
rect 12862 6478 12928 6510
rect 12962 6510 12980 6512
rect 13014 6512 13070 6544
rect 13014 6510 13028 6512
rect 12962 6478 13028 6510
rect 13062 6510 13070 6512
rect 13104 6512 13160 6544
rect 13194 6512 13250 6544
rect 13284 6512 13340 6544
rect 13104 6510 13128 6512
rect 13194 6510 13228 6512
rect 13284 6510 13328 6512
rect 13374 6510 13435 6544
rect 13062 6478 13128 6510
rect 13162 6478 13228 6510
rect 13262 6478 13328 6510
rect 13362 6478 13435 6510
rect 12741 6454 13435 6478
rect 12741 6420 12800 6454
rect 12834 6420 12890 6454
rect 12924 6420 12980 6454
rect 13014 6420 13070 6454
rect 13104 6420 13160 6454
rect 13194 6420 13250 6454
rect 13284 6420 13340 6454
rect 13374 6420 13435 6454
rect 12741 6412 13435 6420
rect 12741 6378 12828 6412
rect 12862 6378 12928 6412
rect 12962 6378 13028 6412
rect 13062 6378 13128 6412
rect 13162 6378 13228 6412
rect 13262 6378 13328 6412
rect 13362 6378 13435 6412
rect 12741 6364 13435 6378
rect 12741 6330 12800 6364
rect 12834 6330 12890 6364
rect 12924 6330 12980 6364
rect 13014 6330 13070 6364
rect 13104 6330 13160 6364
rect 13194 6330 13250 6364
rect 13284 6330 13340 6364
rect 13374 6330 13435 6364
rect 12741 6312 13435 6330
rect 12741 6278 12828 6312
rect 12862 6278 12928 6312
rect 12962 6278 13028 6312
rect 13062 6278 13128 6312
rect 13162 6278 13228 6312
rect 13262 6278 13328 6312
rect 13362 6278 13435 6312
rect 12741 6274 13435 6278
rect 12741 6240 12800 6274
rect 12834 6240 12890 6274
rect 12924 6240 12980 6274
rect 13014 6240 13070 6274
rect 13104 6240 13160 6274
rect 13194 6240 13250 6274
rect 13284 6240 13340 6274
rect 13374 6240 13435 6274
rect 12741 6212 13435 6240
rect 12741 6184 12828 6212
rect 12862 6184 12928 6212
rect 12741 6150 12800 6184
rect 12862 6178 12890 6184
rect 12834 6150 12890 6178
rect 12924 6178 12928 6184
rect 12962 6184 13028 6212
rect 12962 6178 12980 6184
rect 12924 6150 12980 6178
rect 13014 6178 13028 6184
rect 13062 6184 13128 6212
rect 13162 6184 13228 6212
rect 13262 6184 13328 6212
rect 13362 6184 13435 6212
rect 13062 6178 13070 6184
rect 13014 6150 13070 6178
rect 13104 6178 13128 6184
rect 13194 6178 13228 6184
rect 13284 6178 13328 6184
rect 13104 6150 13160 6178
rect 13194 6150 13250 6178
rect 13284 6150 13340 6178
rect 13374 6150 13435 6184
rect 12741 6091 13435 6150
rect 13484 6753 13516 6787
rect 13550 6786 13914 6787
rect 13550 6753 13664 6786
rect 13484 6752 13664 6753
rect 13698 6752 13765 6786
rect 13799 6772 13914 6786
rect 13948 6772 13984 6806
rect 14784 6842 14952 6847
rect 14986 6842 15053 6876
rect 15087 6866 15294 6876
rect 15328 6866 15384 6900
rect 15418 6866 15474 6900
rect 15508 6866 15564 6900
rect 15598 6866 15654 6900
rect 15688 6866 15744 6900
rect 15778 6866 15834 6900
rect 15868 6866 15924 6900
rect 15958 6866 16014 6900
rect 16048 6876 16582 6900
rect 16048 6866 16240 6876
rect 15087 6847 16240 6866
rect 15087 6842 15255 6847
rect 14784 6806 15255 6842
rect 14784 6787 15202 6806
rect 13799 6752 13984 6772
rect 13484 6716 13984 6752
rect 13484 6697 13914 6716
rect 13484 6663 13516 6697
rect 13550 6696 13914 6697
rect 13550 6663 13664 6696
rect 13484 6662 13664 6663
rect 13698 6662 13765 6696
rect 13799 6682 13914 6696
rect 13948 6682 13984 6716
rect 13799 6662 13984 6682
rect 13484 6626 13984 6662
rect 13484 6607 13914 6626
rect 13484 6573 13516 6607
rect 13550 6606 13914 6607
rect 13550 6573 13664 6606
rect 13484 6572 13664 6573
rect 13698 6572 13765 6606
rect 13799 6592 13914 6606
rect 13948 6592 13984 6626
rect 13799 6572 13984 6592
rect 13484 6536 13984 6572
rect 13484 6517 13914 6536
rect 13484 6483 13516 6517
rect 13550 6516 13914 6517
rect 13550 6483 13664 6516
rect 13484 6482 13664 6483
rect 13698 6482 13765 6516
rect 13799 6502 13914 6516
rect 13948 6502 13984 6536
rect 13799 6482 13984 6502
rect 13484 6446 13984 6482
rect 13484 6427 13914 6446
rect 13484 6393 13516 6427
rect 13550 6426 13914 6427
rect 13550 6393 13664 6426
rect 13484 6392 13664 6393
rect 13698 6392 13765 6426
rect 13799 6412 13914 6426
rect 13948 6412 13984 6446
rect 13799 6392 13984 6412
rect 13484 6356 13984 6392
rect 13484 6337 13914 6356
rect 13484 6303 13516 6337
rect 13550 6336 13914 6337
rect 13550 6303 13664 6336
rect 13484 6302 13664 6303
rect 13698 6302 13765 6336
rect 13799 6322 13914 6336
rect 13948 6322 13984 6356
rect 13799 6302 13984 6322
rect 13484 6266 13984 6302
rect 13484 6247 13914 6266
rect 13484 6213 13516 6247
rect 13550 6246 13914 6247
rect 13550 6213 13664 6246
rect 13484 6212 13664 6213
rect 13698 6212 13765 6246
rect 13799 6232 13914 6246
rect 13948 6232 13984 6266
rect 13799 6212 13984 6232
rect 13484 6176 13984 6212
rect 13484 6157 13914 6176
rect 13484 6123 13516 6157
rect 13550 6156 13914 6157
rect 13550 6123 13664 6156
rect 13484 6122 13664 6123
rect 13698 6122 13765 6156
rect 13799 6142 13914 6156
rect 13948 6142 13984 6176
rect 13799 6122 13984 6142
rect 12444 6066 12626 6086
rect 12444 6032 12477 6066
rect 12511 6052 12626 6066
rect 12660 6052 12684 6086
rect 12511 6032 12684 6052
rect 12444 6029 12684 6032
rect 13484 6086 13984 6122
rect 14029 6724 14723 6785
rect 14029 6690 14088 6724
rect 14122 6712 14178 6724
rect 14150 6690 14178 6712
rect 14212 6712 14268 6724
rect 14212 6690 14216 6712
rect 14029 6678 14116 6690
rect 14150 6678 14216 6690
rect 14250 6690 14268 6712
rect 14302 6712 14358 6724
rect 14302 6690 14316 6712
rect 14250 6678 14316 6690
rect 14350 6690 14358 6712
rect 14392 6712 14448 6724
rect 14482 6712 14538 6724
rect 14572 6712 14628 6724
rect 14392 6690 14416 6712
rect 14482 6690 14516 6712
rect 14572 6690 14616 6712
rect 14662 6690 14723 6724
rect 14350 6678 14416 6690
rect 14450 6678 14516 6690
rect 14550 6678 14616 6690
rect 14650 6678 14723 6690
rect 14029 6634 14723 6678
rect 14029 6600 14088 6634
rect 14122 6612 14178 6634
rect 14150 6600 14178 6612
rect 14212 6612 14268 6634
rect 14212 6600 14216 6612
rect 14029 6578 14116 6600
rect 14150 6578 14216 6600
rect 14250 6600 14268 6612
rect 14302 6612 14358 6634
rect 14302 6600 14316 6612
rect 14250 6578 14316 6600
rect 14350 6600 14358 6612
rect 14392 6612 14448 6634
rect 14482 6612 14538 6634
rect 14572 6612 14628 6634
rect 14392 6600 14416 6612
rect 14482 6600 14516 6612
rect 14572 6600 14616 6612
rect 14662 6600 14723 6634
rect 14350 6578 14416 6600
rect 14450 6578 14516 6600
rect 14550 6578 14616 6600
rect 14650 6578 14723 6600
rect 14029 6544 14723 6578
rect 14029 6510 14088 6544
rect 14122 6512 14178 6544
rect 14150 6510 14178 6512
rect 14212 6512 14268 6544
rect 14212 6510 14216 6512
rect 14029 6478 14116 6510
rect 14150 6478 14216 6510
rect 14250 6510 14268 6512
rect 14302 6512 14358 6544
rect 14302 6510 14316 6512
rect 14250 6478 14316 6510
rect 14350 6510 14358 6512
rect 14392 6512 14448 6544
rect 14482 6512 14538 6544
rect 14572 6512 14628 6544
rect 14392 6510 14416 6512
rect 14482 6510 14516 6512
rect 14572 6510 14616 6512
rect 14662 6510 14723 6544
rect 14350 6478 14416 6510
rect 14450 6478 14516 6510
rect 14550 6478 14616 6510
rect 14650 6478 14723 6510
rect 14029 6454 14723 6478
rect 14029 6420 14088 6454
rect 14122 6420 14178 6454
rect 14212 6420 14268 6454
rect 14302 6420 14358 6454
rect 14392 6420 14448 6454
rect 14482 6420 14538 6454
rect 14572 6420 14628 6454
rect 14662 6420 14723 6454
rect 14029 6412 14723 6420
rect 14029 6378 14116 6412
rect 14150 6378 14216 6412
rect 14250 6378 14316 6412
rect 14350 6378 14416 6412
rect 14450 6378 14516 6412
rect 14550 6378 14616 6412
rect 14650 6378 14723 6412
rect 14029 6364 14723 6378
rect 14029 6330 14088 6364
rect 14122 6330 14178 6364
rect 14212 6330 14268 6364
rect 14302 6330 14358 6364
rect 14392 6330 14448 6364
rect 14482 6330 14538 6364
rect 14572 6330 14628 6364
rect 14662 6330 14723 6364
rect 14029 6312 14723 6330
rect 14029 6278 14116 6312
rect 14150 6278 14216 6312
rect 14250 6278 14316 6312
rect 14350 6278 14416 6312
rect 14450 6278 14516 6312
rect 14550 6278 14616 6312
rect 14650 6278 14723 6312
rect 14029 6274 14723 6278
rect 14029 6240 14088 6274
rect 14122 6240 14178 6274
rect 14212 6240 14268 6274
rect 14302 6240 14358 6274
rect 14392 6240 14448 6274
rect 14482 6240 14538 6274
rect 14572 6240 14628 6274
rect 14662 6240 14723 6274
rect 14029 6212 14723 6240
rect 14029 6184 14116 6212
rect 14150 6184 14216 6212
rect 14029 6150 14088 6184
rect 14150 6178 14178 6184
rect 14122 6150 14178 6178
rect 14212 6178 14216 6184
rect 14250 6184 14316 6212
rect 14250 6178 14268 6184
rect 14212 6150 14268 6178
rect 14302 6178 14316 6184
rect 14350 6184 14416 6212
rect 14450 6184 14516 6212
rect 14550 6184 14616 6212
rect 14650 6184 14723 6212
rect 14350 6178 14358 6184
rect 14302 6150 14358 6178
rect 14392 6178 14416 6184
rect 14482 6178 14516 6184
rect 14572 6178 14616 6184
rect 14392 6150 14448 6178
rect 14482 6150 14538 6178
rect 14572 6150 14628 6178
rect 14662 6150 14723 6184
rect 14029 6091 14723 6150
rect 14784 6753 14804 6787
rect 14838 6786 15202 6787
rect 14838 6753 14952 6786
rect 14784 6752 14952 6753
rect 14986 6752 15053 6786
rect 15087 6772 15202 6786
rect 15236 6772 15255 6806
rect 16073 6842 16240 6847
rect 16274 6842 16341 6876
rect 16375 6866 16582 6876
rect 16616 6866 16672 6900
rect 16706 6866 16762 6900
rect 16796 6866 16852 6900
rect 16886 6866 16942 6900
rect 16976 6866 17032 6900
rect 17066 6866 17122 6900
rect 17156 6866 17212 6900
rect 17246 6866 17302 6900
rect 17336 6876 17870 6900
rect 17336 6866 17528 6876
rect 16375 6847 17528 6866
rect 16375 6842 16543 6847
rect 16073 6806 16543 6842
rect 16073 6787 16490 6806
rect 15087 6752 15255 6772
rect 14784 6716 15255 6752
rect 14784 6697 15202 6716
rect 14784 6663 14804 6697
rect 14838 6696 15202 6697
rect 14838 6663 14952 6696
rect 14784 6662 14952 6663
rect 14986 6662 15053 6696
rect 15087 6682 15202 6696
rect 15236 6682 15255 6716
rect 15087 6662 15255 6682
rect 14784 6626 15255 6662
rect 14784 6607 15202 6626
rect 14784 6573 14804 6607
rect 14838 6606 15202 6607
rect 14838 6573 14952 6606
rect 14784 6572 14952 6573
rect 14986 6572 15053 6606
rect 15087 6592 15202 6606
rect 15236 6592 15255 6626
rect 15087 6572 15255 6592
rect 14784 6536 15255 6572
rect 14784 6517 15202 6536
rect 14784 6483 14804 6517
rect 14838 6516 15202 6517
rect 14838 6483 14952 6516
rect 14784 6482 14952 6483
rect 14986 6482 15053 6516
rect 15087 6502 15202 6516
rect 15236 6502 15255 6536
rect 15087 6482 15255 6502
rect 14784 6446 15255 6482
rect 14784 6427 15202 6446
rect 14784 6393 14804 6427
rect 14838 6426 15202 6427
rect 14838 6393 14952 6426
rect 14784 6392 14952 6393
rect 14986 6392 15053 6426
rect 15087 6412 15202 6426
rect 15236 6412 15255 6446
rect 15087 6392 15255 6412
rect 14784 6356 15255 6392
rect 14784 6337 15202 6356
rect 14784 6303 14804 6337
rect 14838 6336 15202 6337
rect 14838 6303 14952 6336
rect 14784 6302 14952 6303
rect 14986 6302 15053 6336
rect 15087 6322 15202 6336
rect 15236 6322 15255 6356
rect 15087 6302 15255 6322
rect 14784 6266 15255 6302
rect 14784 6247 15202 6266
rect 14784 6213 14804 6247
rect 14838 6246 15202 6247
rect 14838 6213 14952 6246
rect 14784 6212 14952 6213
rect 14986 6212 15053 6246
rect 15087 6232 15202 6246
rect 15236 6232 15255 6266
rect 15087 6212 15255 6232
rect 14784 6176 15255 6212
rect 14784 6157 15202 6176
rect 14784 6123 14804 6157
rect 14838 6156 15202 6157
rect 14838 6123 14952 6156
rect 14784 6122 14952 6123
rect 14986 6122 15053 6156
rect 15087 6142 15202 6156
rect 15236 6142 15255 6176
rect 15087 6122 15255 6142
rect 13484 6067 13914 6086
rect 13484 6033 13516 6067
rect 13550 6066 13914 6067
rect 13550 6033 13664 6066
rect 13484 6032 13664 6033
rect 13698 6032 13765 6066
rect 13799 6052 13914 6066
rect 13948 6052 13984 6086
rect 13799 6032 13984 6052
rect 13484 6029 13984 6032
rect 14784 6086 15255 6122
rect 15317 6724 16011 6785
rect 15317 6690 15376 6724
rect 15410 6712 15466 6724
rect 15438 6690 15466 6712
rect 15500 6712 15556 6724
rect 15500 6690 15504 6712
rect 15317 6678 15404 6690
rect 15438 6678 15504 6690
rect 15538 6690 15556 6712
rect 15590 6712 15646 6724
rect 15590 6690 15604 6712
rect 15538 6678 15604 6690
rect 15638 6690 15646 6712
rect 15680 6712 15736 6724
rect 15770 6712 15826 6724
rect 15860 6712 15916 6724
rect 15680 6690 15704 6712
rect 15770 6690 15804 6712
rect 15860 6690 15904 6712
rect 15950 6690 16011 6724
rect 15638 6678 15704 6690
rect 15738 6678 15804 6690
rect 15838 6678 15904 6690
rect 15938 6678 16011 6690
rect 15317 6634 16011 6678
rect 15317 6600 15376 6634
rect 15410 6612 15466 6634
rect 15438 6600 15466 6612
rect 15500 6612 15556 6634
rect 15500 6600 15504 6612
rect 15317 6578 15404 6600
rect 15438 6578 15504 6600
rect 15538 6600 15556 6612
rect 15590 6612 15646 6634
rect 15590 6600 15604 6612
rect 15538 6578 15604 6600
rect 15638 6600 15646 6612
rect 15680 6612 15736 6634
rect 15770 6612 15826 6634
rect 15860 6612 15916 6634
rect 15680 6600 15704 6612
rect 15770 6600 15804 6612
rect 15860 6600 15904 6612
rect 15950 6600 16011 6634
rect 15638 6578 15704 6600
rect 15738 6578 15804 6600
rect 15838 6578 15904 6600
rect 15938 6578 16011 6600
rect 15317 6544 16011 6578
rect 15317 6510 15376 6544
rect 15410 6512 15466 6544
rect 15438 6510 15466 6512
rect 15500 6512 15556 6544
rect 15500 6510 15504 6512
rect 15317 6478 15404 6510
rect 15438 6478 15504 6510
rect 15538 6510 15556 6512
rect 15590 6512 15646 6544
rect 15590 6510 15604 6512
rect 15538 6478 15604 6510
rect 15638 6510 15646 6512
rect 15680 6512 15736 6544
rect 15770 6512 15826 6544
rect 15860 6512 15916 6544
rect 15680 6510 15704 6512
rect 15770 6510 15804 6512
rect 15860 6510 15904 6512
rect 15950 6510 16011 6544
rect 15638 6478 15704 6510
rect 15738 6478 15804 6510
rect 15838 6478 15904 6510
rect 15938 6478 16011 6510
rect 15317 6454 16011 6478
rect 15317 6420 15376 6454
rect 15410 6420 15466 6454
rect 15500 6420 15556 6454
rect 15590 6420 15646 6454
rect 15680 6420 15736 6454
rect 15770 6420 15826 6454
rect 15860 6420 15916 6454
rect 15950 6420 16011 6454
rect 15317 6412 16011 6420
rect 15317 6378 15404 6412
rect 15438 6378 15504 6412
rect 15538 6378 15604 6412
rect 15638 6378 15704 6412
rect 15738 6378 15804 6412
rect 15838 6378 15904 6412
rect 15938 6378 16011 6412
rect 15317 6364 16011 6378
rect 15317 6330 15376 6364
rect 15410 6330 15466 6364
rect 15500 6330 15556 6364
rect 15590 6330 15646 6364
rect 15680 6330 15736 6364
rect 15770 6330 15826 6364
rect 15860 6330 15916 6364
rect 15950 6330 16011 6364
rect 15317 6312 16011 6330
rect 15317 6278 15404 6312
rect 15438 6278 15504 6312
rect 15538 6278 15604 6312
rect 15638 6278 15704 6312
rect 15738 6278 15804 6312
rect 15838 6278 15904 6312
rect 15938 6278 16011 6312
rect 15317 6274 16011 6278
rect 15317 6240 15376 6274
rect 15410 6240 15466 6274
rect 15500 6240 15556 6274
rect 15590 6240 15646 6274
rect 15680 6240 15736 6274
rect 15770 6240 15826 6274
rect 15860 6240 15916 6274
rect 15950 6240 16011 6274
rect 15317 6212 16011 6240
rect 15317 6184 15404 6212
rect 15438 6184 15504 6212
rect 15317 6150 15376 6184
rect 15438 6178 15466 6184
rect 15410 6150 15466 6178
rect 15500 6178 15504 6184
rect 15538 6184 15604 6212
rect 15538 6178 15556 6184
rect 15500 6150 15556 6178
rect 15590 6178 15604 6184
rect 15638 6184 15704 6212
rect 15738 6184 15804 6212
rect 15838 6184 15904 6212
rect 15938 6184 16011 6212
rect 15638 6178 15646 6184
rect 15590 6150 15646 6178
rect 15680 6178 15704 6184
rect 15770 6178 15804 6184
rect 15860 6178 15904 6184
rect 15680 6150 15736 6178
rect 15770 6150 15826 6178
rect 15860 6150 15916 6178
rect 15950 6150 16011 6184
rect 15317 6091 16011 6150
rect 16073 6753 16092 6787
rect 16126 6786 16490 6787
rect 16126 6753 16240 6786
rect 16073 6752 16240 6753
rect 16274 6752 16341 6786
rect 16375 6772 16490 6786
rect 16524 6772 16543 6806
rect 17361 6842 17528 6847
rect 17562 6842 17629 6876
rect 17663 6866 17870 6876
rect 17904 6866 17960 6900
rect 17994 6866 18050 6900
rect 18084 6866 18140 6900
rect 18174 6866 18230 6900
rect 18264 6866 18320 6900
rect 18354 6866 18410 6900
rect 18444 6866 18500 6900
rect 18534 6866 18590 6900
rect 18624 6876 18884 6900
rect 18624 6866 18816 6876
rect 17663 6847 18816 6866
rect 17663 6842 17831 6847
rect 17361 6806 17831 6842
rect 17361 6787 17778 6806
rect 16375 6752 16543 6772
rect 16073 6716 16543 6752
rect 16073 6697 16490 6716
rect 16073 6663 16092 6697
rect 16126 6696 16490 6697
rect 16126 6663 16240 6696
rect 16073 6662 16240 6663
rect 16274 6662 16341 6696
rect 16375 6682 16490 6696
rect 16524 6682 16543 6716
rect 16375 6662 16543 6682
rect 16073 6626 16543 6662
rect 16073 6607 16490 6626
rect 16073 6573 16092 6607
rect 16126 6606 16490 6607
rect 16126 6573 16240 6606
rect 16073 6572 16240 6573
rect 16274 6572 16341 6606
rect 16375 6592 16490 6606
rect 16524 6592 16543 6626
rect 16375 6572 16543 6592
rect 16073 6536 16543 6572
rect 16073 6517 16490 6536
rect 16073 6483 16092 6517
rect 16126 6516 16490 6517
rect 16126 6483 16240 6516
rect 16073 6482 16240 6483
rect 16274 6482 16341 6516
rect 16375 6502 16490 6516
rect 16524 6502 16543 6536
rect 16375 6482 16543 6502
rect 16073 6446 16543 6482
rect 16073 6427 16490 6446
rect 16073 6393 16092 6427
rect 16126 6426 16490 6427
rect 16126 6393 16240 6426
rect 16073 6392 16240 6393
rect 16274 6392 16341 6426
rect 16375 6412 16490 6426
rect 16524 6412 16543 6446
rect 16375 6392 16543 6412
rect 16073 6356 16543 6392
rect 16073 6337 16490 6356
rect 16073 6303 16092 6337
rect 16126 6336 16490 6337
rect 16126 6303 16240 6336
rect 16073 6302 16240 6303
rect 16274 6302 16341 6336
rect 16375 6322 16490 6336
rect 16524 6322 16543 6356
rect 16375 6302 16543 6322
rect 16073 6266 16543 6302
rect 16073 6247 16490 6266
rect 16073 6213 16092 6247
rect 16126 6246 16490 6247
rect 16126 6213 16240 6246
rect 16073 6212 16240 6213
rect 16274 6212 16341 6246
rect 16375 6232 16490 6246
rect 16524 6232 16543 6266
rect 16375 6212 16543 6232
rect 16073 6176 16543 6212
rect 16073 6157 16490 6176
rect 16073 6123 16092 6157
rect 16126 6156 16490 6157
rect 16126 6123 16240 6156
rect 16073 6122 16240 6123
rect 16274 6122 16341 6156
rect 16375 6142 16490 6156
rect 16524 6142 16543 6176
rect 16375 6122 16543 6142
rect 14784 6067 15202 6086
rect 14784 6033 14804 6067
rect 14838 6066 15202 6067
rect 14838 6033 14952 6066
rect 14784 6032 14952 6033
rect 14986 6032 15053 6066
rect 15087 6052 15202 6066
rect 15236 6052 15255 6086
rect 15087 6032 15255 6052
rect 14784 6029 15255 6032
rect 16073 6086 16543 6122
rect 16605 6724 17299 6785
rect 16605 6690 16664 6724
rect 16698 6712 16754 6724
rect 16726 6690 16754 6712
rect 16788 6712 16844 6724
rect 16788 6690 16792 6712
rect 16605 6678 16692 6690
rect 16726 6678 16792 6690
rect 16826 6690 16844 6712
rect 16878 6712 16934 6724
rect 16878 6690 16892 6712
rect 16826 6678 16892 6690
rect 16926 6690 16934 6712
rect 16968 6712 17024 6724
rect 17058 6712 17114 6724
rect 17148 6712 17204 6724
rect 16968 6690 16992 6712
rect 17058 6690 17092 6712
rect 17148 6690 17192 6712
rect 17238 6690 17299 6724
rect 16926 6678 16992 6690
rect 17026 6678 17092 6690
rect 17126 6678 17192 6690
rect 17226 6678 17299 6690
rect 16605 6634 17299 6678
rect 16605 6600 16664 6634
rect 16698 6612 16754 6634
rect 16726 6600 16754 6612
rect 16788 6612 16844 6634
rect 16788 6600 16792 6612
rect 16605 6578 16692 6600
rect 16726 6578 16792 6600
rect 16826 6600 16844 6612
rect 16878 6612 16934 6634
rect 16878 6600 16892 6612
rect 16826 6578 16892 6600
rect 16926 6600 16934 6612
rect 16968 6612 17024 6634
rect 17058 6612 17114 6634
rect 17148 6612 17204 6634
rect 16968 6600 16992 6612
rect 17058 6600 17092 6612
rect 17148 6600 17192 6612
rect 17238 6600 17299 6634
rect 16926 6578 16992 6600
rect 17026 6578 17092 6600
rect 17126 6578 17192 6600
rect 17226 6578 17299 6600
rect 16605 6544 17299 6578
rect 16605 6510 16664 6544
rect 16698 6512 16754 6544
rect 16726 6510 16754 6512
rect 16788 6512 16844 6544
rect 16788 6510 16792 6512
rect 16605 6478 16692 6510
rect 16726 6478 16792 6510
rect 16826 6510 16844 6512
rect 16878 6512 16934 6544
rect 16878 6510 16892 6512
rect 16826 6478 16892 6510
rect 16926 6510 16934 6512
rect 16968 6512 17024 6544
rect 17058 6512 17114 6544
rect 17148 6512 17204 6544
rect 16968 6510 16992 6512
rect 17058 6510 17092 6512
rect 17148 6510 17192 6512
rect 17238 6510 17299 6544
rect 16926 6478 16992 6510
rect 17026 6478 17092 6510
rect 17126 6478 17192 6510
rect 17226 6478 17299 6510
rect 16605 6454 17299 6478
rect 16605 6420 16664 6454
rect 16698 6420 16754 6454
rect 16788 6420 16844 6454
rect 16878 6420 16934 6454
rect 16968 6420 17024 6454
rect 17058 6420 17114 6454
rect 17148 6420 17204 6454
rect 17238 6420 17299 6454
rect 16605 6412 17299 6420
rect 16605 6378 16692 6412
rect 16726 6378 16792 6412
rect 16826 6378 16892 6412
rect 16926 6378 16992 6412
rect 17026 6378 17092 6412
rect 17126 6378 17192 6412
rect 17226 6378 17299 6412
rect 16605 6364 17299 6378
rect 16605 6330 16664 6364
rect 16698 6330 16754 6364
rect 16788 6330 16844 6364
rect 16878 6330 16934 6364
rect 16968 6330 17024 6364
rect 17058 6330 17114 6364
rect 17148 6330 17204 6364
rect 17238 6330 17299 6364
rect 16605 6312 17299 6330
rect 16605 6278 16692 6312
rect 16726 6278 16792 6312
rect 16826 6278 16892 6312
rect 16926 6278 16992 6312
rect 17026 6278 17092 6312
rect 17126 6278 17192 6312
rect 17226 6278 17299 6312
rect 16605 6274 17299 6278
rect 16605 6240 16664 6274
rect 16698 6240 16754 6274
rect 16788 6240 16844 6274
rect 16878 6240 16934 6274
rect 16968 6240 17024 6274
rect 17058 6240 17114 6274
rect 17148 6240 17204 6274
rect 17238 6240 17299 6274
rect 16605 6212 17299 6240
rect 16605 6184 16692 6212
rect 16726 6184 16792 6212
rect 16605 6150 16664 6184
rect 16726 6178 16754 6184
rect 16698 6150 16754 6178
rect 16788 6178 16792 6184
rect 16826 6184 16892 6212
rect 16826 6178 16844 6184
rect 16788 6150 16844 6178
rect 16878 6178 16892 6184
rect 16926 6184 16992 6212
rect 17026 6184 17092 6212
rect 17126 6184 17192 6212
rect 17226 6184 17299 6212
rect 16926 6178 16934 6184
rect 16878 6150 16934 6178
rect 16968 6178 16992 6184
rect 17058 6178 17092 6184
rect 17148 6178 17192 6184
rect 16968 6150 17024 6178
rect 17058 6150 17114 6178
rect 17148 6150 17204 6178
rect 17238 6150 17299 6184
rect 16605 6091 17299 6150
rect 17361 6753 17380 6787
rect 17414 6786 17778 6787
rect 17414 6753 17528 6786
rect 17361 6752 17528 6753
rect 17562 6752 17629 6786
rect 17663 6772 17778 6786
rect 17812 6772 17831 6806
rect 18649 6842 18816 6847
rect 18850 6842 18884 6876
rect 18649 6787 18884 6842
rect 17663 6752 17831 6772
rect 17361 6716 17831 6752
rect 17361 6697 17778 6716
rect 17361 6663 17380 6697
rect 17414 6696 17778 6697
rect 17414 6663 17528 6696
rect 17361 6662 17528 6663
rect 17562 6662 17629 6696
rect 17663 6682 17778 6696
rect 17812 6682 17831 6716
rect 17663 6662 17831 6682
rect 17361 6626 17831 6662
rect 17361 6607 17778 6626
rect 17361 6573 17380 6607
rect 17414 6606 17778 6607
rect 17414 6573 17528 6606
rect 17361 6572 17528 6573
rect 17562 6572 17629 6606
rect 17663 6592 17778 6606
rect 17812 6592 17831 6626
rect 17663 6572 17831 6592
rect 17361 6536 17831 6572
rect 17361 6517 17778 6536
rect 17361 6483 17380 6517
rect 17414 6516 17778 6517
rect 17414 6483 17528 6516
rect 17361 6482 17528 6483
rect 17562 6482 17629 6516
rect 17663 6502 17778 6516
rect 17812 6502 17831 6536
rect 17663 6482 17831 6502
rect 17361 6446 17831 6482
rect 17361 6427 17778 6446
rect 17361 6393 17380 6427
rect 17414 6426 17778 6427
rect 17414 6393 17528 6426
rect 17361 6392 17528 6393
rect 17562 6392 17629 6426
rect 17663 6412 17778 6426
rect 17812 6412 17831 6446
rect 17663 6392 17831 6412
rect 17361 6356 17831 6392
rect 17361 6337 17778 6356
rect 17361 6303 17380 6337
rect 17414 6336 17778 6337
rect 17414 6303 17528 6336
rect 17361 6302 17528 6303
rect 17562 6302 17629 6336
rect 17663 6322 17778 6336
rect 17812 6322 17831 6356
rect 17663 6302 17831 6322
rect 17361 6266 17831 6302
rect 17361 6247 17778 6266
rect 17361 6213 17380 6247
rect 17414 6246 17778 6247
rect 17414 6213 17528 6246
rect 17361 6212 17528 6213
rect 17562 6212 17629 6246
rect 17663 6232 17778 6246
rect 17812 6232 17831 6266
rect 17663 6212 17831 6232
rect 17361 6176 17831 6212
rect 17361 6157 17778 6176
rect 17361 6123 17380 6157
rect 17414 6156 17778 6157
rect 17414 6123 17528 6156
rect 17361 6122 17528 6123
rect 17562 6122 17629 6156
rect 17663 6142 17778 6156
rect 17812 6142 17831 6176
rect 17663 6122 17831 6142
rect 16073 6067 16490 6086
rect 16073 6033 16092 6067
rect 16126 6066 16490 6067
rect 16126 6033 16240 6066
rect 16073 6032 16240 6033
rect 16274 6032 16341 6066
rect 16375 6052 16490 6066
rect 16524 6052 16543 6086
rect 16375 6032 16543 6052
rect 16073 6029 16543 6032
rect 17361 6086 17831 6122
rect 17893 6724 18587 6785
rect 17893 6690 17952 6724
rect 17986 6712 18042 6724
rect 18014 6690 18042 6712
rect 18076 6712 18132 6724
rect 18076 6690 18080 6712
rect 17893 6678 17980 6690
rect 18014 6678 18080 6690
rect 18114 6690 18132 6712
rect 18166 6712 18222 6724
rect 18166 6690 18180 6712
rect 18114 6678 18180 6690
rect 18214 6690 18222 6712
rect 18256 6712 18312 6724
rect 18346 6712 18402 6724
rect 18436 6712 18492 6724
rect 18256 6690 18280 6712
rect 18346 6690 18380 6712
rect 18436 6690 18480 6712
rect 18526 6690 18587 6724
rect 18214 6678 18280 6690
rect 18314 6678 18380 6690
rect 18414 6678 18480 6690
rect 18514 6678 18587 6690
rect 17893 6634 18587 6678
rect 17893 6600 17952 6634
rect 17986 6612 18042 6634
rect 18014 6600 18042 6612
rect 18076 6612 18132 6634
rect 18076 6600 18080 6612
rect 17893 6578 17980 6600
rect 18014 6578 18080 6600
rect 18114 6600 18132 6612
rect 18166 6612 18222 6634
rect 18166 6600 18180 6612
rect 18114 6578 18180 6600
rect 18214 6600 18222 6612
rect 18256 6612 18312 6634
rect 18346 6612 18402 6634
rect 18436 6612 18492 6634
rect 18256 6600 18280 6612
rect 18346 6600 18380 6612
rect 18436 6600 18480 6612
rect 18526 6600 18587 6634
rect 18214 6578 18280 6600
rect 18314 6578 18380 6600
rect 18414 6578 18480 6600
rect 18514 6578 18587 6600
rect 17893 6544 18587 6578
rect 17893 6510 17952 6544
rect 17986 6512 18042 6544
rect 18014 6510 18042 6512
rect 18076 6512 18132 6544
rect 18076 6510 18080 6512
rect 17893 6478 17980 6510
rect 18014 6478 18080 6510
rect 18114 6510 18132 6512
rect 18166 6512 18222 6544
rect 18166 6510 18180 6512
rect 18114 6478 18180 6510
rect 18214 6510 18222 6512
rect 18256 6512 18312 6544
rect 18346 6512 18402 6544
rect 18436 6512 18492 6544
rect 18256 6510 18280 6512
rect 18346 6510 18380 6512
rect 18436 6510 18480 6512
rect 18526 6510 18587 6544
rect 18214 6478 18280 6510
rect 18314 6478 18380 6510
rect 18414 6478 18480 6510
rect 18514 6478 18587 6510
rect 17893 6454 18587 6478
rect 17893 6420 17952 6454
rect 17986 6420 18042 6454
rect 18076 6420 18132 6454
rect 18166 6420 18222 6454
rect 18256 6420 18312 6454
rect 18346 6420 18402 6454
rect 18436 6420 18492 6454
rect 18526 6420 18587 6454
rect 17893 6412 18587 6420
rect 17893 6378 17980 6412
rect 18014 6378 18080 6412
rect 18114 6378 18180 6412
rect 18214 6378 18280 6412
rect 18314 6378 18380 6412
rect 18414 6378 18480 6412
rect 18514 6378 18587 6412
rect 17893 6364 18587 6378
rect 17893 6330 17952 6364
rect 17986 6330 18042 6364
rect 18076 6330 18132 6364
rect 18166 6330 18222 6364
rect 18256 6330 18312 6364
rect 18346 6330 18402 6364
rect 18436 6330 18492 6364
rect 18526 6330 18587 6364
rect 17893 6312 18587 6330
rect 17893 6278 17980 6312
rect 18014 6278 18080 6312
rect 18114 6278 18180 6312
rect 18214 6278 18280 6312
rect 18314 6278 18380 6312
rect 18414 6278 18480 6312
rect 18514 6278 18587 6312
rect 17893 6274 18587 6278
rect 17893 6240 17952 6274
rect 17986 6240 18042 6274
rect 18076 6240 18132 6274
rect 18166 6240 18222 6274
rect 18256 6240 18312 6274
rect 18346 6240 18402 6274
rect 18436 6240 18492 6274
rect 18526 6240 18587 6274
rect 17893 6212 18587 6240
rect 17893 6184 17980 6212
rect 18014 6184 18080 6212
rect 17893 6150 17952 6184
rect 18014 6178 18042 6184
rect 17986 6150 18042 6178
rect 18076 6178 18080 6184
rect 18114 6184 18180 6212
rect 18114 6178 18132 6184
rect 18076 6150 18132 6178
rect 18166 6178 18180 6184
rect 18214 6184 18280 6212
rect 18314 6184 18380 6212
rect 18414 6184 18480 6212
rect 18514 6184 18587 6212
rect 18214 6178 18222 6184
rect 18166 6150 18222 6178
rect 18256 6178 18280 6184
rect 18346 6178 18380 6184
rect 18436 6178 18480 6184
rect 18256 6150 18312 6178
rect 18346 6150 18402 6178
rect 18436 6150 18492 6178
rect 18526 6150 18587 6184
rect 17893 6091 18587 6150
rect 18649 6753 18668 6787
rect 18702 6786 18884 6787
rect 18702 6753 18816 6786
rect 18649 6752 18816 6753
rect 18850 6752 18884 6786
rect 18649 6697 18884 6752
rect 18649 6663 18668 6697
rect 18702 6696 18884 6697
rect 18702 6663 18816 6696
rect 18649 6662 18816 6663
rect 18850 6662 18884 6696
rect 18649 6607 18884 6662
rect 18649 6573 18668 6607
rect 18702 6606 18884 6607
rect 18702 6573 18816 6606
rect 18649 6572 18816 6573
rect 18850 6572 18884 6606
rect 18649 6517 18884 6572
rect 18649 6483 18668 6517
rect 18702 6516 18884 6517
rect 18702 6483 18816 6516
rect 18649 6482 18816 6483
rect 18850 6482 18884 6516
rect 18649 6427 18884 6482
rect 18649 6393 18668 6427
rect 18702 6426 18884 6427
rect 18702 6393 18816 6426
rect 18649 6392 18816 6393
rect 18850 6392 18884 6426
rect 18649 6337 18884 6392
rect 18649 6303 18668 6337
rect 18702 6336 18884 6337
rect 18702 6303 18816 6336
rect 18649 6302 18816 6303
rect 18850 6302 18884 6336
rect 18649 6247 18884 6302
rect 18649 6213 18668 6247
rect 18702 6246 18884 6247
rect 18702 6213 18816 6246
rect 18649 6212 18816 6213
rect 18850 6212 18884 6246
rect 18649 6157 18884 6212
rect 18649 6123 18668 6157
rect 18702 6156 18884 6157
rect 18702 6123 18816 6156
rect 18649 6122 18816 6123
rect 18850 6122 18884 6156
rect 17361 6067 17778 6086
rect 17361 6033 17380 6067
rect 17414 6066 17778 6067
rect 17414 6033 17528 6066
rect 17361 6032 17528 6033
rect 17562 6032 17629 6066
rect 17663 6052 17778 6066
rect 17812 6052 17831 6086
rect 17663 6032 17831 6052
rect 17361 6029 17831 6032
rect 18649 6067 18884 6122
rect 18649 6033 18668 6067
rect 18702 6066 18884 6067
rect 18702 6033 18816 6066
rect 18649 6032 18816 6033
rect 18850 6032 18884 6066
rect 18649 6029 18884 6032
rect 12444 6010 18884 6029
rect 12444 5976 12684 6010
rect 12718 5976 12774 6010
rect 12808 5976 12864 6010
rect 12898 5976 12954 6010
rect 12988 5976 13044 6010
rect 13078 5976 13134 6010
rect 13168 5976 13224 6010
rect 13258 5976 13314 6010
rect 13348 5976 13404 6010
rect 13438 5976 13972 6010
rect 14006 5976 14062 6010
rect 14096 5976 14152 6010
rect 14186 5976 14242 6010
rect 14276 5976 14332 6010
rect 14366 5976 14422 6010
rect 14456 5976 14512 6010
rect 14546 5976 14602 6010
rect 14636 5976 14692 6010
rect 14726 5976 15260 6010
rect 15294 5976 15350 6010
rect 15384 5976 15440 6010
rect 15474 5976 15530 6010
rect 15564 5976 15620 6010
rect 15654 5976 15710 6010
rect 15744 5976 15800 6010
rect 15834 5976 15890 6010
rect 15924 5976 15980 6010
rect 16014 5976 16548 6010
rect 16582 5976 16638 6010
rect 16672 5976 16728 6010
rect 16762 5976 16818 6010
rect 16852 5976 16908 6010
rect 16942 5976 16998 6010
rect 17032 5976 17088 6010
rect 17122 5976 17178 6010
rect 17212 5976 17268 6010
rect 17302 5976 17836 6010
rect 17870 5976 17926 6010
rect 17960 5976 18016 6010
rect 18050 5976 18106 6010
rect 18140 5976 18196 6010
rect 18230 5976 18286 6010
rect 18320 5976 18376 6010
rect 18410 5976 18466 6010
rect 18500 5976 18556 6010
rect 18590 5976 18884 6010
rect 12444 5942 12477 5976
rect 12511 5957 13664 5976
rect 12511 5942 12684 5957
rect 12444 5893 12684 5942
rect 13484 5942 13664 5957
rect 13698 5942 13765 5976
rect 13799 5957 14952 5976
rect 13799 5942 13984 5957
rect 13484 5893 13984 5942
rect 14784 5942 14952 5957
rect 14986 5942 15053 5976
rect 15087 5957 16240 5976
rect 15087 5942 15184 5957
rect 14784 5893 15184 5942
rect 16084 5942 16240 5957
rect 16274 5942 16341 5976
rect 16375 5957 17528 5976
rect 16375 5942 16484 5957
rect 16084 5893 16484 5942
rect 17384 5942 17528 5957
rect 17562 5942 17629 5976
rect 17663 5957 18816 5976
rect 17663 5942 17784 5957
rect 17384 5893 17784 5942
rect 18684 5942 18816 5957
rect 18850 5942 18884 5976
rect 18684 5893 18884 5942
rect 12444 5886 18884 5893
rect 12444 5852 12477 5886
rect 12511 5863 13664 5886
rect 12511 5852 12578 5863
rect 12444 5829 12578 5852
rect 12612 5829 12668 5863
rect 12702 5829 12758 5863
rect 12792 5829 12848 5863
rect 12882 5829 12938 5863
rect 12972 5829 13028 5863
rect 13062 5829 13118 5863
rect 13152 5829 13208 5863
rect 13242 5829 13298 5863
rect 13332 5829 13388 5863
rect 13422 5829 13478 5863
rect 13512 5829 13568 5863
rect 13602 5852 13664 5863
rect 13698 5852 13765 5886
rect 13799 5863 14952 5886
rect 13799 5852 13866 5863
rect 13602 5829 13866 5852
rect 13900 5829 13956 5863
rect 13990 5829 14046 5863
rect 14080 5829 14136 5863
rect 14170 5829 14226 5863
rect 14260 5829 14316 5863
rect 14350 5829 14406 5863
rect 14440 5829 14496 5863
rect 14530 5829 14586 5863
rect 14620 5829 14676 5863
rect 14710 5829 14766 5863
rect 14800 5829 14856 5863
rect 14890 5852 14952 5863
rect 14986 5852 15053 5886
rect 15087 5863 16240 5886
rect 15087 5852 15154 5863
rect 14890 5829 15154 5852
rect 15188 5829 15244 5863
rect 15278 5829 15334 5863
rect 15368 5829 15424 5863
rect 15458 5829 15514 5863
rect 15548 5829 15604 5863
rect 15638 5829 15694 5863
rect 15728 5829 15784 5863
rect 15818 5829 15874 5863
rect 15908 5829 15964 5863
rect 15998 5829 16054 5863
rect 16088 5829 16144 5863
rect 16178 5852 16240 5863
rect 16274 5852 16341 5886
rect 16375 5863 17528 5886
rect 16375 5852 16442 5863
rect 16178 5829 16442 5852
rect 16476 5829 16532 5863
rect 16566 5829 16622 5863
rect 16656 5829 16712 5863
rect 16746 5829 16802 5863
rect 16836 5829 16892 5863
rect 16926 5829 16982 5863
rect 17016 5829 17072 5863
rect 17106 5829 17162 5863
rect 17196 5829 17252 5863
rect 17286 5829 17342 5863
rect 17376 5829 17432 5863
rect 17466 5852 17528 5863
rect 17562 5852 17629 5886
rect 17663 5863 18816 5886
rect 17663 5852 17730 5863
rect 17466 5829 17730 5852
rect 17764 5829 17820 5863
rect 17854 5829 17910 5863
rect 17944 5829 18000 5863
rect 18034 5829 18090 5863
rect 18124 5829 18180 5863
rect 18214 5829 18270 5863
rect 18304 5829 18360 5863
rect 18394 5829 18450 5863
rect 18484 5829 18540 5863
rect 18574 5829 18630 5863
rect 18664 5829 18720 5863
rect 18754 5852 18816 5863
rect 18850 5852 18884 5886
rect 18754 5829 18884 5852
rect 12444 5762 18884 5829
rect 12444 5728 12578 5762
rect 12612 5728 12668 5762
rect 12702 5728 12758 5762
rect 12792 5728 12848 5762
rect 12882 5728 12938 5762
rect 12972 5728 13028 5762
rect 13062 5728 13118 5762
rect 13152 5728 13208 5762
rect 13242 5728 13298 5762
rect 13332 5728 13388 5762
rect 13422 5728 13478 5762
rect 13512 5728 13568 5762
rect 13602 5728 13866 5762
rect 13900 5728 13956 5762
rect 13990 5728 14046 5762
rect 14080 5728 14136 5762
rect 14170 5728 14226 5762
rect 14260 5728 14316 5762
rect 14350 5728 14406 5762
rect 14440 5728 14496 5762
rect 14530 5728 14586 5762
rect 14620 5728 14676 5762
rect 14710 5728 14766 5762
rect 14800 5728 14856 5762
rect 14890 5728 15154 5762
rect 15188 5728 15244 5762
rect 15278 5728 15334 5762
rect 15368 5728 15424 5762
rect 15458 5728 15514 5762
rect 15548 5728 15604 5762
rect 15638 5728 15694 5762
rect 15728 5728 15784 5762
rect 15818 5728 15874 5762
rect 15908 5728 15964 5762
rect 15998 5728 16054 5762
rect 16088 5728 16144 5762
rect 16178 5728 16442 5762
rect 16476 5728 16532 5762
rect 16566 5728 16622 5762
rect 16656 5728 16712 5762
rect 16746 5728 16802 5762
rect 16836 5728 16892 5762
rect 16926 5728 16982 5762
rect 17016 5728 17072 5762
rect 17106 5728 17162 5762
rect 17196 5728 17252 5762
rect 17286 5728 17342 5762
rect 17376 5728 17432 5762
rect 17466 5728 17730 5762
rect 17764 5728 17820 5762
rect 17854 5728 17910 5762
rect 17944 5728 18000 5762
rect 18034 5728 18090 5762
rect 18124 5728 18180 5762
rect 18214 5728 18270 5762
rect 18304 5728 18360 5762
rect 18394 5728 18450 5762
rect 18484 5728 18540 5762
rect 18574 5728 18630 5762
rect 18664 5728 18720 5762
rect 18754 5728 18884 5762
rect 12444 5695 18884 5728
rect 12444 5678 12684 5695
rect 12444 5644 12477 5678
rect 12511 5644 12684 5678
rect 12444 5631 12684 5644
rect 13484 5678 13984 5695
rect 13484 5644 13664 5678
rect 13698 5644 13765 5678
rect 13799 5644 13984 5678
rect 13484 5631 13984 5644
rect 14784 5678 15184 5695
rect 14784 5644 14952 5678
rect 14986 5644 15053 5678
rect 15087 5644 15184 5678
rect 14784 5631 15184 5644
rect 16084 5678 16484 5695
rect 16084 5644 16240 5678
rect 16274 5644 16341 5678
rect 16375 5644 16484 5678
rect 16084 5631 16484 5644
rect 17384 5678 17784 5695
rect 17384 5644 17528 5678
rect 17562 5644 17629 5678
rect 17663 5644 17784 5678
rect 17384 5631 17784 5644
rect 18684 5678 18884 5695
rect 18684 5644 18816 5678
rect 18850 5644 18884 5678
rect 18684 5631 18884 5644
rect 12444 5612 18884 5631
rect 12444 5588 12718 5612
rect 12444 5554 12477 5588
rect 12511 5578 12718 5588
rect 12752 5578 12808 5612
rect 12842 5578 12898 5612
rect 12932 5578 12988 5612
rect 13022 5578 13078 5612
rect 13112 5578 13168 5612
rect 13202 5578 13258 5612
rect 13292 5578 13348 5612
rect 13382 5578 13438 5612
rect 13472 5588 14006 5612
rect 13472 5578 13664 5588
rect 12511 5559 13664 5578
rect 12511 5554 12684 5559
rect 12444 5518 12684 5554
rect 12444 5498 12626 5518
rect 12444 5464 12477 5498
rect 12511 5484 12626 5498
rect 12660 5484 12684 5518
rect 13484 5554 13664 5559
rect 13698 5554 13765 5588
rect 13799 5578 14006 5588
rect 14040 5578 14096 5612
rect 14130 5578 14186 5612
rect 14220 5578 14276 5612
rect 14310 5578 14366 5612
rect 14400 5578 14456 5612
rect 14490 5578 14546 5612
rect 14580 5578 14636 5612
rect 14670 5578 14726 5612
rect 14760 5588 15294 5612
rect 14760 5578 14952 5588
rect 13799 5559 14952 5578
rect 13799 5554 13984 5559
rect 13484 5518 13984 5554
rect 13484 5499 13914 5518
rect 12511 5464 12684 5484
rect 12444 5428 12684 5464
rect 12444 5408 12626 5428
rect 12444 5374 12477 5408
rect 12511 5394 12626 5408
rect 12660 5394 12684 5428
rect 12511 5374 12684 5394
rect 12444 5338 12684 5374
rect 12444 5318 12626 5338
rect 12444 5284 12477 5318
rect 12511 5304 12626 5318
rect 12660 5304 12684 5338
rect 12511 5284 12684 5304
rect 12444 5248 12684 5284
rect 12444 5228 12626 5248
rect 12444 5194 12477 5228
rect 12511 5214 12626 5228
rect 12660 5214 12684 5248
rect 12511 5194 12684 5214
rect 12444 5158 12684 5194
rect 12444 5138 12626 5158
rect 12444 5104 12477 5138
rect 12511 5124 12626 5138
rect 12660 5124 12684 5158
rect 12511 5104 12684 5124
rect 12444 5068 12684 5104
rect 12444 5048 12626 5068
rect 12444 5014 12477 5048
rect 12511 5034 12626 5048
rect 12660 5034 12684 5068
rect 12511 5014 12684 5034
rect 12444 4978 12684 5014
rect 12444 4958 12626 4978
rect 12444 4924 12477 4958
rect 12511 4944 12626 4958
rect 12660 4944 12684 4978
rect 12511 4924 12684 4944
rect 12444 4888 12684 4924
rect 12444 4868 12626 4888
rect 12444 4834 12477 4868
rect 12511 4854 12626 4868
rect 12660 4854 12684 4888
rect 12511 4834 12684 4854
rect 12444 4798 12684 4834
rect 12741 5436 13435 5497
rect 12741 5402 12800 5436
rect 12834 5424 12890 5436
rect 12862 5402 12890 5424
rect 12924 5424 12980 5436
rect 12924 5402 12928 5424
rect 12741 5390 12828 5402
rect 12862 5390 12928 5402
rect 12962 5402 12980 5424
rect 13014 5424 13070 5436
rect 13014 5402 13028 5424
rect 12962 5390 13028 5402
rect 13062 5402 13070 5424
rect 13104 5424 13160 5436
rect 13194 5424 13250 5436
rect 13284 5424 13340 5436
rect 13104 5402 13128 5424
rect 13194 5402 13228 5424
rect 13284 5402 13328 5424
rect 13374 5402 13435 5436
rect 13062 5390 13128 5402
rect 13162 5390 13228 5402
rect 13262 5390 13328 5402
rect 13362 5390 13435 5402
rect 12741 5346 13435 5390
rect 12741 5312 12800 5346
rect 12834 5324 12890 5346
rect 12862 5312 12890 5324
rect 12924 5324 12980 5346
rect 12924 5312 12928 5324
rect 12741 5290 12828 5312
rect 12862 5290 12928 5312
rect 12962 5312 12980 5324
rect 13014 5324 13070 5346
rect 13014 5312 13028 5324
rect 12962 5290 13028 5312
rect 13062 5312 13070 5324
rect 13104 5324 13160 5346
rect 13194 5324 13250 5346
rect 13284 5324 13340 5346
rect 13104 5312 13128 5324
rect 13194 5312 13228 5324
rect 13284 5312 13328 5324
rect 13374 5312 13435 5346
rect 13062 5290 13128 5312
rect 13162 5290 13228 5312
rect 13262 5290 13328 5312
rect 13362 5290 13435 5312
rect 12741 5256 13435 5290
rect 12741 5222 12800 5256
rect 12834 5224 12890 5256
rect 12862 5222 12890 5224
rect 12924 5224 12980 5256
rect 12924 5222 12928 5224
rect 12741 5190 12828 5222
rect 12862 5190 12928 5222
rect 12962 5222 12980 5224
rect 13014 5224 13070 5256
rect 13014 5222 13028 5224
rect 12962 5190 13028 5222
rect 13062 5222 13070 5224
rect 13104 5224 13160 5256
rect 13194 5224 13250 5256
rect 13284 5224 13340 5256
rect 13104 5222 13128 5224
rect 13194 5222 13228 5224
rect 13284 5222 13328 5224
rect 13374 5222 13435 5256
rect 13062 5190 13128 5222
rect 13162 5190 13228 5222
rect 13262 5190 13328 5222
rect 13362 5190 13435 5222
rect 12741 5166 13435 5190
rect 12741 5132 12800 5166
rect 12834 5132 12890 5166
rect 12924 5132 12980 5166
rect 13014 5132 13070 5166
rect 13104 5132 13160 5166
rect 13194 5132 13250 5166
rect 13284 5132 13340 5166
rect 13374 5132 13435 5166
rect 12741 5124 13435 5132
rect 12741 5090 12828 5124
rect 12862 5090 12928 5124
rect 12962 5090 13028 5124
rect 13062 5090 13128 5124
rect 13162 5090 13228 5124
rect 13262 5090 13328 5124
rect 13362 5090 13435 5124
rect 12741 5076 13435 5090
rect 12741 5042 12800 5076
rect 12834 5042 12890 5076
rect 12924 5042 12980 5076
rect 13014 5042 13070 5076
rect 13104 5042 13160 5076
rect 13194 5042 13250 5076
rect 13284 5042 13340 5076
rect 13374 5042 13435 5076
rect 12741 5024 13435 5042
rect 12741 4990 12828 5024
rect 12862 4990 12928 5024
rect 12962 4990 13028 5024
rect 13062 4990 13128 5024
rect 13162 4990 13228 5024
rect 13262 4990 13328 5024
rect 13362 4990 13435 5024
rect 12741 4986 13435 4990
rect 12741 4952 12800 4986
rect 12834 4952 12890 4986
rect 12924 4952 12980 4986
rect 13014 4952 13070 4986
rect 13104 4952 13160 4986
rect 13194 4952 13250 4986
rect 13284 4952 13340 4986
rect 13374 4952 13435 4986
rect 12741 4924 13435 4952
rect 12741 4896 12828 4924
rect 12862 4896 12928 4924
rect 12741 4862 12800 4896
rect 12862 4890 12890 4896
rect 12834 4862 12890 4890
rect 12924 4890 12928 4896
rect 12962 4896 13028 4924
rect 12962 4890 12980 4896
rect 12924 4862 12980 4890
rect 13014 4890 13028 4896
rect 13062 4896 13128 4924
rect 13162 4896 13228 4924
rect 13262 4896 13328 4924
rect 13362 4896 13435 4924
rect 13062 4890 13070 4896
rect 13014 4862 13070 4890
rect 13104 4890 13128 4896
rect 13194 4890 13228 4896
rect 13284 4890 13328 4896
rect 13104 4862 13160 4890
rect 13194 4862 13250 4890
rect 13284 4862 13340 4890
rect 13374 4862 13435 4896
rect 12741 4803 13435 4862
rect 13484 5465 13516 5499
rect 13550 5498 13914 5499
rect 13550 5465 13664 5498
rect 13484 5464 13664 5465
rect 13698 5464 13765 5498
rect 13799 5484 13914 5498
rect 13948 5484 13984 5518
rect 14784 5554 14952 5559
rect 14986 5554 15053 5588
rect 15087 5578 15294 5588
rect 15328 5578 15384 5612
rect 15418 5578 15474 5612
rect 15508 5578 15564 5612
rect 15598 5578 15654 5612
rect 15688 5578 15744 5612
rect 15778 5578 15834 5612
rect 15868 5578 15924 5612
rect 15958 5578 16014 5612
rect 16048 5588 16582 5612
rect 16048 5578 16240 5588
rect 15087 5559 16240 5578
rect 15087 5554 15255 5559
rect 14784 5518 15255 5554
rect 14784 5499 15202 5518
rect 13799 5464 13984 5484
rect 13484 5428 13984 5464
rect 13484 5409 13914 5428
rect 13484 5375 13516 5409
rect 13550 5408 13914 5409
rect 13550 5375 13664 5408
rect 13484 5374 13664 5375
rect 13698 5374 13765 5408
rect 13799 5394 13914 5408
rect 13948 5394 13984 5428
rect 13799 5374 13984 5394
rect 13484 5338 13984 5374
rect 13484 5319 13914 5338
rect 13484 5285 13516 5319
rect 13550 5318 13914 5319
rect 13550 5285 13664 5318
rect 13484 5284 13664 5285
rect 13698 5284 13765 5318
rect 13799 5304 13914 5318
rect 13948 5304 13984 5338
rect 13799 5284 13984 5304
rect 13484 5248 13984 5284
rect 13484 5229 13914 5248
rect 13484 5195 13516 5229
rect 13550 5228 13914 5229
rect 13550 5195 13664 5228
rect 13484 5194 13664 5195
rect 13698 5194 13765 5228
rect 13799 5214 13914 5228
rect 13948 5214 13984 5248
rect 13799 5194 13984 5214
rect 13484 5158 13984 5194
rect 13484 5139 13914 5158
rect 13484 5105 13516 5139
rect 13550 5138 13914 5139
rect 13550 5105 13664 5138
rect 13484 5104 13664 5105
rect 13698 5104 13765 5138
rect 13799 5124 13914 5138
rect 13948 5124 13984 5158
rect 13799 5104 13984 5124
rect 13484 5068 13984 5104
rect 13484 5049 13914 5068
rect 13484 5015 13516 5049
rect 13550 5048 13914 5049
rect 13550 5015 13664 5048
rect 13484 5014 13664 5015
rect 13698 5014 13765 5048
rect 13799 5034 13914 5048
rect 13948 5034 13984 5068
rect 13799 5014 13984 5034
rect 13484 4978 13984 5014
rect 13484 4959 13914 4978
rect 13484 4925 13516 4959
rect 13550 4958 13914 4959
rect 13550 4925 13664 4958
rect 13484 4924 13664 4925
rect 13698 4924 13765 4958
rect 13799 4944 13914 4958
rect 13948 4944 13984 4978
rect 13799 4924 13984 4944
rect 13484 4888 13984 4924
rect 13484 4869 13914 4888
rect 13484 4835 13516 4869
rect 13550 4868 13914 4869
rect 13550 4835 13664 4868
rect 13484 4834 13664 4835
rect 13698 4834 13765 4868
rect 13799 4854 13914 4868
rect 13948 4854 13984 4888
rect 13799 4834 13984 4854
rect 12444 4778 12626 4798
rect 12444 4744 12477 4778
rect 12511 4764 12626 4778
rect 12660 4764 12684 4798
rect 12511 4744 12684 4764
rect 12444 4741 12684 4744
rect 13484 4798 13984 4834
rect 14029 5436 14723 5497
rect 14029 5402 14088 5436
rect 14122 5424 14178 5436
rect 14150 5402 14178 5424
rect 14212 5424 14268 5436
rect 14212 5402 14216 5424
rect 14029 5390 14116 5402
rect 14150 5390 14216 5402
rect 14250 5402 14268 5424
rect 14302 5424 14358 5436
rect 14302 5402 14316 5424
rect 14250 5390 14316 5402
rect 14350 5402 14358 5424
rect 14392 5424 14448 5436
rect 14482 5424 14538 5436
rect 14572 5424 14628 5436
rect 14392 5402 14416 5424
rect 14482 5402 14516 5424
rect 14572 5402 14616 5424
rect 14662 5402 14723 5436
rect 14350 5390 14416 5402
rect 14450 5390 14516 5402
rect 14550 5390 14616 5402
rect 14650 5390 14723 5402
rect 14029 5346 14723 5390
rect 14029 5312 14088 5346
rect 14122 5324 14178 5346
rect 14150 5312 14178 5324
rect 14212 5324 14268 5346
rect 14212 5312 14216 5324
rect 14029 5290 14116 5312
rect 14150 5290 14216 5312
rect 14250 5312 14268 5324
rect 14302 5324 14358 5346
rect 14302 5312 14316 5324
rect 14250 5290 14316 5312
rect 14350 5312 14358 5324
rect 14392 5324 14448 5346
rect 14482 5324 14538 5346
rect 14572 5324 14628 5346
rect 14392 5312 14416 5324
rect 14482 5312 14516 5324
rect 14572 5312 14616 5324
rect 14662 5312 14723 5346
rect 14350 5290 14416 5312
rect 14450 5290 14516 5312
rect 14550 5290 14616 5312
rect 14650 5290 14723 5312
rect 14029 5256 14723 5290
rect 14029 5222 14088 5256
rect 14122 5224 14178 5256
rect 14150 5222 14178 5224
rect 14212 5224 14268 5256
rect 14212 5222 14216 5224
rect 14029 5190 14116 5222
rect 14150 5190 14216 5222
rect 14250 5222 14268 5224
rect 14302 5224 14358 5256
rect 14302 5222 14316 5224
rect 14250 5190 14316 5222
rect 14350 5222 14358 5224
rect 14392 5224 14448 5256
rect 14482 5224 14538 5256
rect 14572 5224 14628 5256
rect 14392 5222 14416 5224
rect 14482 5222 14516 5224
rect 14572 5222 14616 5224
rect 14662 5222 14723 5256
rect 14350 5190 14416 5222
rect 14450 5190 14516 5222
rect 14550 5190 14616 5222
rect 14650 5190 14723 5222
rect 14029 5166 14723 5190
rect 14029 5132 14088 5166
rect 14122 5132 14178 5166
rect 14212 5132 14268 5166
rect 14302 5132 14358 5166
rect 14392 5132 14448 5166
rect 14482 5132 14538 5166
rect 14572 5132 14628 5166
rect 14662 5132 14723 5166
rect 14029 5124 14723 5132
rect 14029 5090 14116 5124
rect 14150 5090 14216 5124
rect 14250 5090 14316 5124
rect 14350 5090 14416 5124
rect 14450 5090 14516 5124
rect 14550 5090 14616 5124
rect 14650 5090 14723 5124
rect 14029 5076 14723 5090
rect 14029 5042 14088 5076
rect 14122 5042 14178 5076
rect 14212 5042 14268 5076
rect 14302 5042 14358 5076
rect 14392 5042 14448 5076
rect 14482 5042 14538 5076
rect 14572 5042 14628 5076
rect 14662 5042 14723 5076
rect 14029 5024 14723 5042
rect 14029 4990 14116 5024
rect 14150 4990 14216 5024
rect 14250 4990 14316 5024
rect 14350 4990 14416 5024
rect 14450 4990 14516 5024
rect 14550 4990 14616 5024
rect 14650 4990 14723 5024
rect 14029 4986 14723 4990
rect 14029 4952 14088 4986
rect 14122 4952 14178 4986
rect 14212 4952 14268 4986
rect 14302 4952 14358 4986
rect 14392 4952 14448 4986
rect 14482 4952 14538 4986
rect 14572 4952 14628 4986
rect 14662 4952 14723 4986
rect 14029 4924 14723 4952
rect 14029 4896 14116 4924
rect 14150 4896 14216 4924
rect 14029 4862 14088 4896
rect 14150 4890 14178 4896
rect 14122 4862 14178 4890
rect 14212 4890 14216 4896
rect 14250 4896 14316 4924
rect 14250 4890 14268 4896
rect 14212 4862 14268 4890
rect 14302 4890 14316 4896
rect 14350 4896 14416 4924
rect 14450 4896 14516 4924
rect 14550 4896 14616 4924
rect 14650 4896 14723 4924
rect 14350 4890 14358 4896
rect 14302 4862 14358 4890
rect 14392 4890 14416 4896
rect 14482 4890 14516 4896
rect 14572 4890 14616 4896
rect 14392 4862 14448 4890
rect 14482 4862 14538 4890
rect 14572 4862 14628 4890
rect 14662 4862 14723 4896
rect 14029 4803 14723 4862
rect 14784 5465 14804 5499
rect 14838 5498 15202 5499
rect 14838 5465 14952 5498
rect 14784 5464 14952 5465
rect 14986 5464 15053 5498
rect 15087 5484 15202 5498
rect 15236 5484 15255 5518
rect 16073 5554 16240 5559
rect 16274 5554 16341 5588
rect 16375 5578 16582 5588
rect 16616 5578 16672 5612
rect 16706 5578 16762 5612
rect 16796 5578 16852 5612
rect 16886 5578 16942 5612
rect 16976 5578 17032 5612
rect 17066 5578 17122 5612
rect 17156 5578 17212 5612
rect 17246 5578 17302 5612
rect 17336 5588 17870 5612
rect 17336 5578 17528 5588
rect 16375 5559 17528 5578
rect 16375 5554 16543 5559
rect 16073 5518 16543 5554
rect 16073 5499 16490 5518
rect 15087 5464 15255 5484
rect 14784 5428 15255 5464
rect 14784 5409 15202 5428
rect 14784 5375 14804 5409
rect 14838 5408 15202 5409
rect 14838 5375 14952 5408
rect 14784 5374 14952 5375
rect 14986 5374 15053 5408
rect 15087 5394 15202 5408
rect 15236 5394 15255 5428
rect 15087 5374 15255 5394
rect 14784 5338 15255 5374
rect 14784 5319 15202 5338
rect 14784 5285 14804 5319
rect 14838 5318 15202 5319
rect 14838 5285 14952 5318
rect 14784 5284 14952 5285
rect 14986 5284 15053 5318
rect 15087 5304 15202 5318
rect 15236 5304 15255 5338
rect 15087 5284 15255 5304
rect 14784 5248 15255 5284
rect 14784 5229 15202 5248
rect 14784 5195 14804 5229
rect 14838 5228 15202 5229
rect 14838 5195 14952 5228
rect 14784 5194 14952 5195
rect 14986 5194 15053 5228
rect 15087 5214 15202 5228
rect 15236 5214 15255 5248
rect 15087 5194 15255 5214
rect 14784 5158 15255 5194
rect 14784 5139 15202 5158
rect 14784 5105 14804 5139
rect 14838 5138 15202 5139
rect 14838 5105 14952 5138
rect 14784 5104 14952 5105
rect 14986 5104 15053 5138
rect 15087 5124 15202 5138
rect 15236 5124 15255 5158
rect 15087 5104 15255 5124
rect 14784 5068 15255 5104
rect 14784 5049 15202 5068
rect 14784 5015 14804 5049
rect 14838 5048 15202 5049
rect 14838 5015 14952 5048
rect 14784 5014 14952 5015
rect 14986 5014 15053 5048
rect 15087 5034 15202 5048
rect 15236 5034 15255 5068
rect 15087 5014 15255 5034
rect 14784 4978 15255 5014
rect 14784 4959 15202 4978
rect 14784 4925 14804 4959
rect 14838 4958 15202 4959
rect 14838 4925 14952 4958
rect 14784 4924 14952 4925
rect 14986 4924 15053 4958
rect 15087 4944 15202 4958
rect 15236 4944 15255 4978
rect 15087 4924 15255 4944
rect 14784 4888 15255 4924
rect 14784 4869 15202 4888
rect 14784 4835 14804 4869
rect 14838 4868 15202 4869
rect 14838 4835 14952 4868
rect 14784 4834 14952 4835
rect 14986 4834 15053 4868
rect 15087 4854 15202 4868
rect 15236 4854 15255 4888
rect 15087 4834 15255 4854
rect 13484 4779 13914 4798
rect 13484 4745 13516 4779
rect 13550 4778 13914 4779
rect 13550 4745 13664 4778
rect 13484 4744 13664 4745
rect 13698 4744 13765 4778
rect 13799 4764 13914 4778
rect 13948 4764 13984 4798
rect 13799 4744 13984 4764
rect 13484 4741 13984 4744
rect 14784 4798 15255 4834
rect 15317 5436 16011 5497
rect 15317 5402 15376 5436
rect 15410 5424 15466 5436
rect 15438 5402 15466 5424
rect 15500 5424 15556 5436
rect 15500 5402 15504 5424
rect 15317 5390 15404 5402
rect 15438 5390 15504 5402
rect 15538 5402 15556 5424
rect 15590 5424 15646 5436
rect 15590 5402 15604 5424
rect 15538 5390 15604 5402
rect 15638 5402 15646 5424
rect 15680 5424 15736 5436
rect 15770 5424 15826 5436
rect 15860 5424 15916 5436
rect 15680 5402 15704 5424
rect 15770 5402 15804 5424
rect 15860 5402 15904 5424
rect 15950 5402 16011 5436
rect 15638 5390 15704 5402
rect 15738 5390 15804 5402
rect 15838 5390 15904 5402
rect 15938 5390 16011 5402
rect 15317 5346 16011 5390
rect 15317 5312 15376 5346
rect 15410 5324 15466 5346
rect 15438 5312 15466 5324
rect 15500 5324 15556 5346
rect 15500 5312 15504 5324
rect 15317 5290 15404 5312
rect 15438 5290 15504 5312
rect 15538 5312 15556 5324
rect 15590 5324 15646 5346
rect 15590 5312 15604 5324
rect 15538 5290 15604 5312
rect 15638 5312 15646 5324
rect 15680 5324 15736 5346
rect 15770 5324 15826 5346
rect 15860 5324 15916 5346
rect 15680 5312 15704 5324
rect 15770 5312 15804 5324
rect 15860 5312 15904 5324
rect 15950 5312 16011 5346
rect 15638 5290 15704 5312
rect 15738 5290 15804 5312
rect 15838 5290 15904 5312
rect 15938 5290 16011 5312
rect 15317 5256 16011 5290
rect 15317 5222 15376 5256
rect 15410 5224 15466 5256
rect 15438 5222 15466 5224
rect 15500 5224 15556 5256
rect 15500 5222 15504 5224
rect 15317 5190 15404 5222
rect 15438 5190 15504 5222
rect 15538 5222 15556 5224
rect 15590 5224 15646 5256
rect 15590 5222 15604 5224
rect 15538 5190 15604 5222
rect 15638 5222 15646 5224
rect 15680 5224 15736 5256
rect 15770 5224 15826 5256
rect 15860 5224 15916 5256
rect 15680 5222 15704 5224
rect 15770 5222 15804 5224
rect 15860 5222 15904 5224
rect 15950 5222 16011 5256
rect 15638 5190 15704 5222
rect 15738 5190 15804 5222
rect 15838 5190 15904 5222
rect 15938 5190 16011 5222
rect 15317 5166 16011 5190
rect 15317 5132 15376 5166
rect 15410 5132 15466 5166
rect 15500 5132 15556 5166
rect 15590 5132 15646 5166
rect 15680 5132 15736 5166
rect 15770 5132 15826 5166
rect 15860 5132 15916 5166
rect 15950 5132 16011 5166
rect 15317 5124 16011 5132
rect 15317 5090 15404 5124
rect 15438 5090 15504 5124
rect 15538 5090 15604 5124
rect 15638 5090 15704 5124
rect 15738 5090 15804 5124
rect 15838 5090 15904 5124
rect 15938 5090 16011 5124
rect 15317 5076 16011 5090
rect 15317 5042 15376 5076
rect 15410 5042 15466 5076
rect 15500 5042 15556 5076
rect 15590 5042 15646 5076
rect 15680 5042 15736 5076
rect 15770 5042 15826 5076
rect 15860 5042 15916 5076
rect 15950 5042 16011 5076
rect 15317 5024 16011 5042
rect 15317 4990 15404 5024
rect 15438 4990 15504 5024
rect 15538 4990 15604 5024
rect 15638 4990 15704 5024
rect 15738 4990 15804 5024
rect 15838 4990 15904 5024
rect 15938 4990 16011 5024
rect 15317 4986 16011 4990
rect 15317 4952 15376 4986
rect 15410 4952 15466 4986
rect 15500 4952 15556 4986
rect 15590 4952 15646 4986
rect 15680 4952 15736 4986
rect 15770 4952 15826 4986
rect 15860 4952 15916 4986
rect 15950 4952 16011 4986
rect 15317 4924 16011 4952
rect 15317 4896 15404 4924
rect 15438 4896 15504 4924
rect 15317 4862 15376 4896
rect 15438 4890 15466 4896
rect 15410 4862 15466 4890
rect 15500 4890 15504 4896
rect 15538 4896 15604 4924
rect 15538 4890 15556 4896
rect 15500 4862 15556 4890
rect 15590 4890 15604 4896
rect 15638 4896 15704 4924
rect 15738 4896 15804 4924
rect 15838 4896 15904 4924
rect 15938 4896 16011 4924
rect 15638 4890 15646 4896
rect 15590 4862 15646 4890
rect 15680 4890 15704 4896
rect 15770 4890 15804 4896
rect 15860 4890 15904 4896
rect 15680 4862 15736 4890
rect 15770 4862 15826 4890
rect 15860 4862 15916 4890
rect 15950 4862 16011 4896
rect 15317 4803 16011 4862
rect 16073 5465 16092 5499
rect 16126 5498 16490 5499
rect 16126 5465 16240 5498
rect 16073 5464 16240 5465
rect 16274 5464 16341 5498
rect 16375 5484 16490 5498
rect 16524 5484 16543 5518
rect 17361 5554 17528 5559
rect 17562 5554 17629 5588
rect 17663 5578 17870 5588
rect 17904 5578 17960 5612
rect 17994 5578 18050 5612
rect 18084 5578 18140 5612
rect 18174 5578 18230 5612
rect 18264 5578 18320 5612
rect 18354 5578 18410 5612
rect 18444 5578 18500 5612
rect 18534 5578 18590 5612
rect 18624 5588 18884 5612
rect 18624 5578 18816 5588
rect 17663 5559 18816 5578
rect 17663 5554 17831 5559
rect 17361 5518 17831 5554
rect 17361 5499 17778 5518
rect 16375 5464 16543 5484
rect 16073 5428 16543 5464
rect 16073 5409 16490 5428
rect 16073 5375 16092 5409
rect 16126 5408 16490 5409
rect 16126 5375 16240 5408
rect 16073 5374 16240 5375
rect 16274 5374 16341 5408
rect 16375 5394 16490 5408
rect 16524 5394 16543 5428
rect 16375 5374 16543 5394
rect 16073 5338 16543 5374
rect 16073 5319 16490 5338
rect 16073 5285 16092 5319
rect 16126 5318 16490 5319
rect 16126 5285 16240 5318
rect 16073 5284 16240 5285
rect 16274 5284 16341 5318
rect 16375 5304 16490 5318
rect 16524 5304 16543 5338
rect 16375 5284 16543 5304
rect 16073 5248 16543 5284
rect 16073 5229 16490 5248
rect 16073 5195 16092 5229
rect 16126 5228 16490 5229
rect 16126 5195 16240 5228
rect 16073 5194 16240 5195
rect 16274 5194 16341 5228
rect 16375 5214 16490 5228
rect 16524 5214 16543 5248
rect 16375 5194 16543 5214
rect 16073 5158 16543 5194
rect 16073 5139 16490 5158
rect 16073 5105 16092 5139
rect 16126 5138 16490 5139
rect 16126 5105 16240 5138
rect 16073 5104 16240 5105
rect 16274 5104 16341 5138
rect 16375 5124 16490 5138
rect 16524 5124 16543 5158
rect 16375 5104 16543 5124
rect 16073 5068 16543 5104
rect 16073 5049 16490 5068
rect 16073 5015 16092 5049
rect 16126 5048 16490 5049
rect 16126 5015 16240 5048
rect 16073 5014 16240 5015
rect 16274 5014 16341 5048
rect 16375 5034 16490 5048
rect 16524 5034 16543 5068
rect 16375 5014 16543 5034
rect 16073 4978 16543 5014
rect 16073 4959 16490 4978
rect 16073 4925 16092 4959
rect 16126 4958 16490 4959
rect 16126 4925 16240 4958
rect 16073 4924 16240 4925
rect 16274 4924 16341 4958
rect 16375 4944 16490 4958
rect 16524 4944 16543 4978
rect 16375 4924 16543 4944
rect 16073 4888 16543 4924
rect 16073 4869 16490 4888
rect 16073 4835 16092 4869
rect 16126 4868 16490 4869
rect 16126 4835 16240 4868
rect 16073 4834 16240 4835
rect 16274 4834 16341 4868
rect 16375 4854 16490 4868
rect 16524 4854 16543 4888
rect 16375 4834 16543 4854
rect 14784 4779 15202 4798
rect 14784 4745 14804 4779
rect 14838 4778 15202 4779
rect 14838 4745 14952 4778
rect 14784 4744 14952 4745
rect 14986 4744 15053 4778
rect 15087 4764 15202 4778
rect 15236 4764 15255 4798
rect 15087 4744 15255 4764
rect 14784 4741 15255 4744
rect 16073 4798 16543 4834
rect 16605 5436 17299 5497
rect 16605 5402 16664 5436
rect 16698 5424 16754 5436
rect 16726 5402 16754 5424
rect 16788 5424 16844 5436
rect 16788 5402 16792 5424
rect 16605 5390 16692 5402
rect 16726 5390 16792 5402
rect 16826 5402 16844 5424
rect 16878 5424 16934 5436
rect 16878 5402 16892 5424
rect 16826 5390 16892 5402
rect 16926 5402 16934 5424
rect 16968 5424 17024 5436
rect 17058 5424 17114 5436
rect 17148 5424 17204 5436
rect 16968 5402 16992 5424
rect 17058 5402 17092 5424
rect 17148 5402 17192 5424
rect 17238 5402 17299 5436
rect 16926 5390 16992 5402
rect 17026 5390 17092 5402
rect 17126 5390 17192 5402
rect 17226 5390 17299 5402
rect 16605 5346 17299 5390
rect 16605 5312 16664 5346
rect 16698 5324 16754 5346
rect 16726 5312 16754 5324
rect 16788 5324 16844 5346
rect 16788 5312 16792 5324
rect 16605 5290 16692 5312
rect 16726 5290 16792 5312
rect 16826 5312 16844 5324
rect 16878 5324 16934 5346
rect 16878 5312 16892 5324
rect 16826 5290 16892 5312
rect 16926 5312 16934 5324
rect 16968 5324 17024 5346
rect 17058 5324 17114 5346
rect 17148 5324 17204 5346
rect 16968 5312 16992 5324
rect 17058 5312 17092 5324
rect 17148 5312 17192 5324
rect 17238 5312 17299 5346
rect 16926 5290 16992 5312
rect 17026 5290 17092 5312
rect 17126 5290 17192 5312
rect 17226 5290 17299 5312
rect 16605 5256 17299 5290
rect 16605 5222 16664 5256
rect 16698 5224 16754 5256
rect 16726 5222 16754 5224
rect 16788 5224 16844 5256
rect 16788 5222 16792 5224
rect 16605 5190 16692 5222
rect 16726 5190 16792 5222
rect 16826 5222 16844 5224
rect 16878 5224 16934 5256
rect 16878 5222 16892 5224
rect 16826 5190 16892 5222
rect 16926 5222 16934 5224
rect 16968 5224 17024 5256
rect 17058 5224 17114 5256
rect 17148 5224 17204 5256
rect 16968 5222 16992 5224
rect 17058 5222 17092 5224
rect 17148 5222 17192 5224
rect 17238 5222 17299 5256
rect 16926 5190 16992 5222
rect 17026 5190 17092 5222
rect 17126 5190 17192 5222
rect 17226 5190 17299 5222
rect 16605 5166 17299 5190
rect 16605 5132 16664 5166
rect 16698 5132 16754 5166
rect 16788 5132 16844 5166
rect 16878 5132 16934 5166
rect 16968 5132 17024 5166
rect 17058 5132 17114 5166
rect 17148 5132 17204 5166
rect 17238 5132 17299 5166
rect 16605 5124 17299 5132
rect 16605 5090 16692 5124
rect 16726 5090 16792 5124
rect 16826 5090 16892 5124
rect 16926 5090 16992 5124
rect 17026 5090 17092 5124
rect 17126 5090 17192 5124
rect 17226 5090 17299 5124
rect 16605 5076 17299 5090
rect 16605 5042 16664 5076
rect 16698 5042 16754 5076
rect 16788 5042 16844 5076
rect 16878 5042 16934 5076
rect 16968 5042 17024 5076
rect 17058 5042 17114 5076
rect 17148 5042 17204 5076
rect 17238 5042 17299 5076
rect 16605 5024 17299 5042
rect 16605 4990 16692 5024
rect 16726 4990 16792 5024
rect 16826 4990 16892 5024
rect 16926 4990 16992 5024
rect 17026 4990 17092 5024
rect 17126 4990 17192 5024
rect 17226 4990 17299 5024
rect 16605 4986 17299 4990
rect 16605 4952 16664 4986
rect 16698 4952 16754 4986
rect 16788 4952 16844 4986
rect 16878 4952 16934 4986
rect 16968 4952 17024 4986
rect 17058 4952 17114 4986
rect 17148 4952 17204 4986
rect 17238 4952 17299 4986
rect 16605 4924 17299 4952
rect 16605 4896 16692 4924
rect 16726 4896 16792 4924
rect 16605 4862 16664 4896
rect 16726 4890 16754 4896
rect 16698 4862 16754 4890
rect 16788 4890 16792 4896
rect 16826 4896 16892 4924
rect 16826 4890 16844 4896
rect 16788 4862 16844 4890
rect 16878 4890 16892 4896
rect 16926 4896 16992 4924
rect 17026 4896 17092 4924
rect 17126 4896 17192 4924
rect 17226 4896 17299 4924
rect 16926 4890 16934 4896
rect 16878 4862 16934 4890
rect 16968 4890 16992 4896
rect 17058 4890 17092 4896
rect 17148 4890 17192 4896
rect 16968 4862 17024 4890
rect 17058 4862 17114 4890
rect 17148 4862 17204 4890
rect 17238 4862 17299 4896
rect 16605 4803 17299 4862
rect 17361 5465 17380 5499
rect 17414 5498 17778 5499
rect 17414 5465 17528 5498
rect 17361 5464 17528 5465
rect 17562 5464 17629 5498
rect 17663 5484 17778 5498
rect 17812 5484 17831 5518
rect 18649 5554 18816 5559
rect 18850 5554 18884 5588
rect 18649 5499 18884 5554
rect 17663 5464 17831 5484
rect 17361 5428 17831 5464
rect 17361 5409 17778 5428
rect 17361 5375 17380 5409
rect 17414 5408 17778 5409
rect 17414 5375 17528 5408
rect 17361 5374 17528 5375
rect 17562 5374 17629 5408
rect 17663 5394 17778 5408
rect 17812 5394 17831 5428
rect 17663 5374 17831 5394
rect 17361 5338 17831 5374
rect 17361 5319 17778 5338
rect 17361 5285 17380 5319
rect 17414 5318 17778 5319
rect 17414 5285 17528 5318
rect 17361 5284 17528 5285
rect 17562 5284 17629 5318
rect 17663 5304 17778 5318
rect 17812 5304 17831 5338
rect 17663 5284 17831 5304
rect 17361 5248 17831 5284
rect 17361 5229 17778 5248
rect 17361 5195 17380 5229
rect 17414 5228 17778 5229
rect 17414 5195 17528 5228
rect 17361 5194 17528 5195
rect 17562 5194 17629 5228
rect 17663 5214 17778 5228
rect 17812 5214 17831 5248
rect 17663 5194 17831 5214
rect 17361 5158 17831 5194
rect 17361 5139 17778 5158
rect 17361 5105 17380 5139
rect 17414 5138 17778 5139
rect 17414 5105 17528 5138
rect 17361 5104 17528 5105
rect 17562 5104 17629 5138
rect 17663 5124 17778 5138
rect 17812 5124 17831 5158
rect 17663 5104 17831 5124
rect 17361 5068 17831 5104
rect 17361 5049 17778 5068
rect 17361 5015 17380 5049
rect 17414 5048 17778 5049
rect 17414 5015 17528 5048
rect 17361 5014 17528 5015
rect 17562 5014 17629 5048
rect 17663 5034 17778 5048
rect 17812 5034 17831 5068
rect 17663 5014 17831 5034
rect 17361 4978 17831 5014
rect 17361 4959 17778 4978
rect 17361 4925 17380 4959
rect 17414 4958 17778 4959
rect 17414 4925 17528 4958
rect 17361 4924 17528 4925
rect 17562 4924 17629 4958
rect 17663 4944 17778 4958
rect 17812 4944 17831 4978
rect 17663 4924 17831 4944
rect 17361 4888 17831 4924
rect 17361 4869 17778 4888
rect 17361 4835 17380 4869
rect 17414 4868 17778 4869
rect 17414 4835 17528 4868
rect 17361 4834 17528 4835
rect 17562 4834 17629 4868
rect 17663 4854 17778 4868
rect 17812 4854 17831 4888
rect 17663 4834 17831 4854
rect 16073 4779 16490 4798
rect 16073 4745 16092 4779
rect 16126 4778 16490 4779
rect 16126 4745 16240 4778
rect 16073 4744 16240 4745
rect 16274 4744 16341 4778
rect 16375 4764 16490 4778
rect 16524 4764 16543 4798
rect 16375 4744 16543 4764
rect 16073 4741 16543 4744
rect 17361 4798 17831 4834
rect 17893 5436 18587 5497
rect 17893 5402 17952 5436
rect 17986 5424 18042 5436
rect 18014 5402 18042 5424
rect 18076 5424 18132 5436
rect 18076 5402 18080 5424
rect 17893 5390 17980 5402
rect 18014 5390 18080 5402
rect 18114 5402 18132 5424
rect 18166 5424 18222 5436
rect 18166 5402 18180 5424
rect 18114 5390 18180 5402
rect 18214 5402 18222 5424
rect 18256 5424 18312 5436
rect 18346 5424 18402 5436
rect 18436 5424 18492 5436
rect 18256 5402 18280 5424
rect 18346 5402 18380 5424
rect 18436 5402 18480 5424
rect 18526 5402 18587 5436
rect 18214 5390 18280 5402
rect 18314 5390 18380 5402
rect 18414 5390 18480 5402
rect 18514 5390 18587 5402
rect 17893 5346 18587 5390
rect 17893 5312 17952 5346
rect 17986 5324 18042 5346
rect 18014 5312 18042 5324
rect 18076 5324 18132 5346
rect 18076 5312 18080 5324
rect 17893 5290 17980 5312
rect 18014 5290 18080 5312
rect 18114 5312 18132 5324
rect 18166 5324 18222 5346
rect 18166 5312 18180 5324
rect 18114 5290 18180 5312
rect 18214 5312 18222 5324
rect 18256 5324 18312 5346
rect 18346 5324 18402 5346
rect 18436 5324 18492 5346
rect 18256 5312 18280 5324
rect 18346 5312 18380 5324
rect 18436 5312 18480 5324
rect 18526 5312 18587 5346
rect 18214 5290 18280 5312
rect 18314 5290 18380 5312
rect 18414 5290 18480 5312
rect 18514 5290 18587 5312
rect 17893 5256 18587 5290
rect 17893 5222 17952 5256
rect 17986 5224 18042 5256
rect 18014 5222 18042 5224
rect 18076 5224 18132 5256
rect 18076 5222 18080 5224
rect 17893 5190 17980 5222
rect 18014 5190 18080 5222
rect 18114 5222 18132 5224
rect 18166 5224 18222 5256
rect 18166 5222 18180 5224
rect 18114 5190 18180 5222
rect 18214 5222 18222 5224
rect 18256 5224 18312 5256
rect 18346 5224 18402 5256
rect 18436 5224 18492 5256
rect 18256 5222 18280 5224
rect 18346 5222 18380 5224
rect 18436 5222 18480 5224
rect 18526 5222 18587 5256
rect 18214 5190 18280 5222
rect 18314 5190 18380 5222
rect 18414 5190 18480 5222
rect 18514 5190 18587 5222
rect 17893 5166 18587 5190
rect 17893 5132 17952 5166
rect 17986 5132 18042 5166
rect 18076 5132 18132 5166
rect 18166 5132 18222 5166
rect 18256 5132 18312 5166
rect 18346 5132 18402 5166
rect 18436 5132 18492 5166
rect 18526 5132 18587 5166
rect 17893 5124 18587 5132
rect 17893 5090 17980 5124
rect 18014 5090 18080 5124
rect 18114 5090 18180 5124
rect 18214 5090 18280 5124
rect 18314 5090 18380 5124
rect 18414 5090 18480 5124
rect 18514 5090 18587 5124
rect 17893 5076 18587 5090
rect 17893 5042 17952 5076
rect 17986 5042 18042 5076
rect 18076 5042 18132 5076
rect 18166 5042 18222 5076
rect 18256 5042 18312 5076
rect 18346 5042 18402 5076
rect 18436 5042 18492 5076
rect 18526 5042 18587 5076
rect 17893 5024 18587 5042
rect 17893 4990 17980 5024
rect 18014 4990 18080 5024
rect 18114 4990 18180 5024
rect 18214 4990 18280 5024
rect 18314 4990 18380 5024
rect 18414 4990 18480 5024
rect 18514 4990 18587 5024
rect 17893 4986 18587 4990
rect 17893 4952 17952 4986
rect 17986 4952 18042 4986
rect 18076 4952 18132 4986
rect 18166 4952 18222 4986
rect 18256 4952 18312 4986
rect 18346 4952 18402 4986
rect 18436 4952 18492 4986
rect 18526 4952 18587 4986
rect 17893 4924 18587 4952
rect 17893 4896 17980 4924
rect 18014 4896 18080 4924
rect 17893 4862 17952 4896
rect 18014 4890 18042 4896
rect 17986 4862 18042 4890
rect 18076 4890 18080 4896
rect 18114 4896 18180 4924
rect 18114 4890 18132 4896
rect 18076 4862 18132 4890
rect 18166 4890 18180 4896
rect 18214 4896 18280 4924
rect 18314 4896 18380 4924
rect 18414 4896 18480 4924
rect 18514 4896 18587 4924
rect 18214 4890 18222 4896
rect 18166 4862 18222 4890
rect 18256 4890 18280 4896
rect 18346 4890 18380 4896
rect 18436 4890 18480 4896
rect 18256 4862 18312 4890
rect 18346 4862 18402 4890
rect 18436 4862 18492 4890
rect 18526 4862 18587 4896
rect 17893 4803 18587 4862
rect 18649 5465 18668 5499
rect 18702 5498 18884 5499
rect 18702 5465 18816 5498
rect 18649 5464 18816 5465
rect 18850 5464 18884 5498
rect 18649 5409 18884 5464
rect 18649 5375 18668 5409
rect 18702 5408 18884 5409
rect 18702 5375 18816 5408
rect 18649 5374 18816 5375
rect 18850 5374 18884 5408
rect 18649 5319 18884 5374
rect 18649 5285 18668 5319
rect 18702 5318 18884 5319
rect 18702 5285 18816 5318
rect 18649 5284 18816 5285
rect 18850 5284 18884 5318
rect 18649 5229 18884 5284
rect 18649 5195 18668 5229
rect 18702 5228 18884 5229
rect 18702 5195 18816 5228
rect 18649 5194 18816 5195
rect 18850 5194 18884 5228
rect 18649 5139 18884 5194
rect 18649 5105 18668 5139
rect 18702 5138 18884 5139
rect 18702 5105 18816 5138
rect 18649 5104 18816 5105
rect 18850 5104 18884 5138
rect 18649 5049 18884 5104
rect 18649 5015 18668 5049
rect 18702 5048 18884 5049
rect 18702 5015 18816 5048
rect 18649 5014 18816 5015
rect 18850 5014 18884 5048
rect 18649 4959 18884 5014
rect 18649 4925 18668 4959
rect 18702 4958 18884 4959
rect 18702 4925 18816 4958
rect 18649 4924 18816 4925
rect 18850 4924 18884 4958
rect 18649 4869 18884 4924
rect 18649 4835 18668 4869
rect 18702 4868 18884 4869
rect 18702 4835 18816 4868
rect 18649 4834 18816 4835
rect 18850 4834 18884 4868
rect 17361 4779 17778 4798
rect 17361 4745 17380 4779
rect 17414 4778 17778 4779
rect 17414 4745 17528 4778
rect 17361 4744 17528 4745
rect 17562 4744 17629 4778
rect 17663 4764 17778 4778
rect 17812 4764 17831 4798
rect 17663 4744 17831 4764
rect 17361 4741 17831 4744
rect 18649 4779 18884 4834
rect 18649 4745 18668 4779
rect 18702 4778 18884 4779
rect 18702 4745 18816 4778
rect 18649 4744 18816 4745
rect 18850 4744 18884 4778
rect 18649 4741 18884 4744
rect 12444 4722 18884 4741
rect 12444 4688 12684 4722
rect 12718 4688 12774 4722
rect 12808 4688 12864 4722
rect 12898 4688 12954 4722
rect 12988 4688 13044 4722
rect 13078 4688 13134 4722
rect 13168 4688 13224 4722
rect 13258 4688 13314 4722
rect 13348 4688 13404 4722
rect 13438 4688 13972 4722
rect 14006 4688 14062 4722
rect 14096 4688 14152 4722
rect 14186 4688 14242 4722
rect 14276 4688 14332 4722
rect 14366 4688 14422 4722
rect 14456 4688 14512 4722
rect 14546 4688 14602 4722
rect 14636 4688 14692 4722
rect 14726 4688 15260 4722
rect 15294 4688 15350 4722
rect 15384 4688 15440 4722
rect 15474 4688 15530 4722
rect 15564 4688 15620 4722
rect 15654 4688 15710 4722
rect 15744 4688 15800 4722
rect 15834 4688 15890 4722
rect 15924 4688 15980 4722
rect 16014 4688 16548 4722
rect 16582 4688 16638 4722
rect 16672 4688 16728 4722
rect 16762 4688 16818 4722
rect 16852 4688 16908 4722
rect 16942 4688 16998 4722
rect 17032 4688 17088 4722
rect 17122 4688 17178 4722
rect 17212 4688 17268 4722
rect 17302 4688 17836 4722
rect 17870 4688 17926 4722
rect 17960 4688 18016 4722
rect 18050 4688 18106 4722
rect 18140 4688 18196 4722
rect 18230 4688 18286 4722
rect 18320 4688 18376 4722
rect 18410 4688 18466 4722
rect 18500 4688 18556 4722
rect 18590 4688 18884 4722
rect 12444 4654 12477 4688
rect 12511 4669 13664 4688
rect 12511 4654 12684 4669
rect 12444 4605 12684 4654
rect 13484 4654 13664 4669
rect 13698 4654 13765 4688
rect 13799 4669 14952 4688
rect 13799 4654 13984 4669
rect 13484 4605 13984 4654
rect 14784 4654 14952 4669
rect 14986 4654 15053 4688
rect 15087 4669 16240 4688
rect 15087 4654 15184 4669
rect 14784 4605 15184 4654
rect 16084 4654 16240 4669
rect 16274 4654 16341 4688
rect 16375 4669 17528 4688
rect 16375 4654 16484 4669
rect 16084 4605 16484 4654
rect 17384 4654 17528 4669
rect 17562 4654 17629 4688
rect 17663 4669 18816 4688
rect 17663 4654 17784 4669
rect 17384 4605 17784 4654
rect 18684 4654 18816 4669
rect 18850 4654 18884 4688
rect 18684 4605 18884 4654
rect 12444 4598 18884 4605
rect 12444 4564 12477 4598
rect 12511 4575 13664 4598
rect 12511 4564 12578 4575
rect 12444 4541 12578 4564
rect 12612 4541 12668 4575
rect 12702 4541 12758 4575
rect 12792 4541 12848 4575
rect 12882 4541 12938 4575
rect 12972 4541 13028 4575
rect 13062 4541 13118 4575
rect 13152 4541 13208 4575
rect 13242 4541 13298 4575
rect 13332 4541 13388 4575
rect 13422 4541 13478 4575
rect 13512 4541 13568 4575
rect 13602 4564 13664 4575
rect 13698 4564 13765 4598
rect 13799 4575 14952 4598
rect 13799 4564 13866 4575
rect 13602 4541 13866 4564
rect 13900 4541 13956 4575
rect 13990 4541 14046 4575
rect 14080 4541 14136 4575
rect 14170 4541 14226 4575
rect 14260 4541 14316 4575
rect 14350 4541 14406 4575
rect 14440 4541 14496 4575
rect 14530 4541 14586 4575
rect 14620 4541 14676 4575
rect 14710 4541 14766 4575
rect 14800 4541 14856 4575
rect 14890 4564 14952 4575
rect 14986 4564 15053 4598
rect 15087 4575 16240 4598
rect 15087 4564 15154 4575
rect 14890 4541 15154 4564
rect 15188 4541 15244 4575
rect 15278 4541 15334 4575
rect 15368 4541 15424 4575
rect 15458 4541 15514 4575
rect 15548 4541 15604 4575
rect 15638 4541 15694 4575
rect 15728 4541 15784 4575
rect 15818 4541 15874 4575
rect 15908 4541 15964 4575
rect 15998 4541 16054 4575
rect 16088 4541 16144 4575
rect 16178 4564 16240 4575
rect 16274 4564 16341 4598
rect 16375 4575 17528 4598
rect 16375 4564 16442 4575
rect 16178 4541 16442 4564
rect 16476 4541 16532 4575
rect 16566 4541 16622 4575
rect 16656 4541 16712 4575
rect 16746 4541 16802 4575
rect 16836 4541 16892 4575
rect 16926 4541 16982 4575
rect 17016 4541 17072 4575
rect 17106 4541 17162 4575
rect 17196 4541 17252 4575
rect 17286 4541 17342 4575
rect 17376 4541 17432 4575
rect 17466 4564 17528 4575
rect 17562 4564 17629 4598
rect 17663 4575 18816 4598
rect 17663 4564 17730 4575
rect 17466 4541 17730 4564
rect 17764 4541 17820 4575
rect 17854 4541 17910 4575
rect 17944 4541 18000 4575
rect 18034 4541 18090 4575
rect 18124 4541 18180 4575
rect 18214 4541 18270 4575
rect 18304 4541 18360 4575
rect 18394 4541 18450 4575
rect 18484 4541 18540 4575
rect 18574 4541 18630 4575
rect 18664 4541 18720 4575
rect 18754 4564 18816 4575
rect 18850 4564 18884 4598
rect 18754 4541 18884 4564
rect 12444 4474 18884 4541
rect 12444 4440 12578 4474
rect 12612 4440 12668 4474
rect 12702 4440 12758 4474
rect 12792 4440 12848 4474
rect 12882 4440 12938 4474
rect 12972 4440 13028 4474
rect 13062 4440 13118 4474
rect 13152 4440 13208 4474
rect 13242 4440 13298 4474
rect 13332 4440 13388 4474
rect 13422 4440 13478 4474
rect 13512 4440 13568 4474
rect 13602 4440 13866 4474
rect 13900 4440 13956 4474
rect 13990 4440 14046 4474
rect 14080 4440 14136 4474
rect 14170 4440 14226 4474
rect 14260 4440 14316 4474
rect 14350 4440 14406 4474
rect 14440 4440 14496 4474
rect 14530 4440 14586 4474
rect 14620 4440 14676 4474
rect 14710 4440 14766 4474
rect 14800 4440 14856 4474
rect 14890 4440 15154 4474
rect 15188 4440 15244 4474
rect 15278 4440 15334 4474
rect 15368 4440 15424 4474
rect 15458 4440 15514 4474
rect 15548 4440 15604 4474
rect 15638 4440 15694 4474
rect 15728 4440 15784 4474
rect 15818 4440 15874 4474
rect 15908 4440 15964 4474
rect 15998 4440 16054 4474
rect 16088 4440 16144 4474
rect 16178 4440 16442 4474
rect 16476 4440 16532 4474
rect 16566 4440 16622 4474
rect 16656 4440 16712 4474
rect 16746 4440 16802 4474
rect 16836 4440 16892 4474
rect 16926 4440 16982 4474
rect 17016 4440 17072 4474
rect 17106 4440 17162 4474
rect 17196 4440 17252 4474
rect 17286 4440 17342 4474
rect 17376 4440 17432 4474
rect 17466 4440 17730 4474
rect 17764 4440 17820 4474
rect 17854 4440 17910 4474
rect 17944 4440 18000 4474
rect 18034 4440 18090 4474
rect 18124 4440 18180 4474
rect 18214 4440 18270 4474
rect 18304 4440 18360 4474
rect 18394 4440 18450 4474
rect 18484 4440 18540 4474
rect 18574 4440 18630 4474
rect 18664 4440 18720 4474
rect 18754 4440 18884 4474
rect 12444 4407 18884 4440
rect 12444 4390 12684 4407
rect 12444 4356 12477 4390
rect 12511 4356 12684 4390
rect 12444 4343 12684 4356
rect 13484 4390 13984 4407
rect 13484 4356 13664 4390
rect 13698 4356 13765 4390
rect 13799 4356 13984 4390
rect 13484 4343 13984 4356
rect 14784 4390 15184 4407
rect 14784 4356 14952 4390
rect 14986 4356 15053 4390
rect 15087 4356 15184 4390
rect 14784 4343 15184 4356
rect 16084 4390 16484 4407
rect 16084 4356 16240 4390
rect 16274 4356 16341 4390
rect 16375 4356 16484 4390
rect 16084 4343 16484 4356
rect 17384 4390 17784 4407
rect 17384 4356 17528 4390
rect 17562 4356 17629 4390
rect 17663 4356 17784 4390
rect 17384 4343 17784 4356
rect 18684 4390 18884 4407
rect 18684 4356 18816 4390
rect 18850 4356 18884 4390
rect 18684 4343 18884 4356
rect 12444 4324 18884 4343
rect 12444 4300 12718 4324
rect 12444 4266 12477 4300
rect 12511 4290 12718 4300
rect 12752 4290 12808 4324
rect 12842 4290 12898 4324
rect 12932 4290 12988 4324
rect 13022 4290 13078 4324
rect 13112 4290 13168 4324
rect 13202 4290 13258 4324
rect 13292 4290 13348 4324
rect 13382 4290 13438 4324
rect 13472 4300 14006 4324
rect 13472 4290 13664 4300
rect 12511 4271 13664 4290
rect 12511 4266 12684 4271
rect 12444 4230 12684 4266
rect 12444 4210 12626 4230
rect 12444 4176 12477 4210
rect 12511 4196 12626 4210
rect 12660 4196 12684 4230
rect 13484 4266 13664 4271
rect 13698 4266 13765 4300
rect 13799 4290 14006 4300
rect 14040 4290 14096 4324
rect 14130 4290 14186 4324
rect 14220 4290 14276 4324
rect 14310 4290 14366 4324
rect 14400 4290 14456 4324
rect 14490 4290 14546 4324
rect 14580 4290 14636 4324
rect 14670 4290 14726 4324
rect 14760 4300 15294 4324
rect 14760 4290 14952 4300
rect 13799 4271 14952 4290
rect 13799 4266 13984 4271
rect 13484 4230 13984 4266
rect 13484 4211 13914 4230
rect 12511 4176 12684 4196
rect 12444 4140 12684 4176
rect 12444 4120 12626 4140
rect 12444 4086 12477 4120
rect 12511 4106 12626 4120
rect 12660 4106 12684 4140
rect 12511 4086 12684 4106
rect 12444 4050 12684 4086
rect 12444 4030 12626 4050
rect 12444 3996 12477 4030
rect 12511 4016 12626 4030
rect 12660 4016 12684 4050
rect 12511 3996 12684 4016
rect 12444 3960 12684 3996
rect 12444 3940 12626 3960
rect 12444 3906 12477 3940
rect 12511 3926 12626 3940
rect 12660 3926 12684 3960
rect 12511 3906 12684 3926
rect 12444 3870 12684 3906
rect 12444 3850 12626 3870
rect 12444 3816 12477 3850
rect 12511 3836 12626 3850
rect 12660 3836 12684 3870
rect 12511 3816 12684 3836
rect 12444 3780 12684 3816
rect 12444 3760 12626 3780
rect 12444 3726 12477 3760
rect 12511 3746 12626 3760
rect 12660 3746 12684 3780
rect 12511 3726 12684 3746
rect 12444 3690 12684 3726
rect 12444 3670 12626 3690
rect 12444 3636 12477 3670
rect 12511 3656 12626 3670
rect 12660 3656 12684 3690
rect 12511 3636 12684 3656
rect 12444 3600 12684 3636
rect 12444 3580 12626 3600
rect 12444 3546 12477 3580
rect 12511 3566 12626 3580
rect 12660 3566 12684 3600
rect 12511 3546 12684 3566
rect 12444 3510 12684 3546
rect 12741 4148 13435 4209
rect 12741 4114 12800 4148
rect 12834 4136 12890 4148
rect 12862 4114 12890 4136
rect 12924 4136 12980 4148
rect 12924 4114 12928 4136
rect 12741 4102 12828 4114
rect 12862 4102 12928 4114
rect 12962 4114 12980 4136
rect 13014 4136 13070 4148
rect 13014 4114 13028 4136
rect 12962 4102 13028 4114
rect 13062 4114 13070 4136
rect 13104 4136 13160 4148
rect 13194 4136 13250 4148
rect 13284 4136 13340 4148
rect 13104 4114 13128 4136
rect 13194 4114 13228 4136
rect 13284 4114 13328 4136
rect 13374 4114 13435 4148
rect 13062 4102 13128 4114
rect 13162 4102 13228 4114
rect 13262 4102 13328 4114
rect 13362 4102 13435 4114
rect 12741 4058 13435 4102
rect 12741 4024 12800 4058
rect 12834 4036 12890 4058
rect 12862 4024 12890 4036
rect 12924 4036 12980 4058
rect 12924 4024 12928 4036
rect 12741 4002 12828 4024
rect 12862 4002 12928 4024
rect 12962 4024 12980 4036
rect 13014 4036 13070 4058
rect 13014 4024 13028 4036
rect 12962 4002 13028 4024
rect 13062 4024 13070 4036
rect 13104 4036 13160 4058
rect 13194 4036 13250 4058
rect 13284 4036 13340 4058
rect 13104 4024 13128 4036
rect 13194 4024 13228 4036
rect 13284 4024 13328 4036
rect 13374 4024 13435 4058
rect 13062 4002 13128 4024
rect 13162 4002 13228 4024
rect 13262 4002 13328 4024
rect 13362 4002 13435 4024
rect 12741 3968 13435 4002
rect 12741 3934 12800 3968
rect 12834 3936 12890 3968
rect 12862 3934 12890 3936
rect 12924 3936 12980 3968
rect 12924 3934 12928 3936
rect 12741 3902 12828 3934
rect 12862 3902 12928 3934
rect 12962 3934 12980 3936
rect 13014 3936 13070 3968
rect 13014 3934 13028 3936
rect 12962 3902 13028 3934
rect 13062 3934 13070 3936
rect 13104 3936 13160 3968
rect 13194 3936 13250 3968
rect 13284 3936 13340 3968
rect 13104 3934 13128 3936
rect 13194 3934 13228 3936
rect 13284 3934 13328 3936
rect 13374 3934 13435 3968
rect 13062 3902 13128 3934
rect 13162 3902 13228 3934
rect 13262 3902 13328 3934
rect 13362 3902 13435 3934
rect 12741 3878 13435 3902
rect 12741 3844 12800 3878
rect 12834 3844 12890 3878
rect 12924 3844 12980 3878
rect 13014 3844 13070 3878
rect 13104 3844 13160 3878
rect 13194 3844 13250 3878
rect 13284 3844 13340 3878
rect 13374 3844 13435 3878
rect 12741 3836 13435 3844
rect 12741 3802 12828 3836
rect 12862 3802 12928 3836
rect 12962 3802 13028 3836
rect 13062 3802 13128 3836
rect 13162 3802 13228 3836
rect 13262 3802 13328 3836
rect 13362 3802 13435 3836
rect 12741 3788 13435 3802
rect 12741 3754 12800 3788
rect 12834 3754 12890 3788
rect 12924 3754 12980 3788
rect 13014 3754 13070 3788
rect 13104 3754 13160 3788
rect 13194 3754 13250 3788
rect 13284 3754 13340 3788
rect 13374 3754 13435 3788
rect 12741 3736 13435 3754
rect 12741 3702 12828 3736
rect 12862 3702 12928 3736
rect 12962 3702 13028 3736
rect 13062 3702 13128 3736
rect 13162 3702 13228 3736
rect 13262 3702 13328 3736
rect 13362 3702 13435 3736
rect 12741 3698 13435 3702
rect 12741 3664 12800 3698
rect 12834 3664 12890 3698
rect 12924 3664 12980 3698
rect 13014 3664 13070 3698
rect 13104 3664 13160 3698
rect 13194 3664 13250 3698
rect 13284 3664 13340 3698
rect 13374 3664 13435 3698
rect 12741 3636 13435 3664
rect 12741 3608 12828 3636
rect 12862 3608 12928 3636
rect 12741 3574 12800 3608
rect 12862 3602 12890 3608
rect 12834 3574 12890 3602
rect 12924 3602 12928 3608
rect 12962 3608 13028 3636
rect 12962 3602 12980 3608
rect 12924 3574 12980 3602
rect 13014 3602 13028 3608
rect 13062 3608 13128 3636
rect 13162 3608 13228 3636
rect 13262 3608 13328 3636
rect 13362 3608 13435 3636
rect 13062 3602 13070 3608
rect 13014 3574 13070 3602
rect 13104 3602 13128 3608
rect 13194 3602 13228 3608
rect 13284 3602 13328 3608
rect 13104 3574 13160 3602
rect 13194 3574 13250 3602
rect 13284 3574 13340 3602
rect 13374 3574 13435 3608
rect 12741 3515 13435 3574
rect 13484 4177 13516 4211
rect 13550 4210 13914 4211
rect 13550 4177 13664 4210
rect 13484 4176 13664 4177
rect 13698 4176 13765 4210
rect 13799 4196 13914 4210
rect 13948 4196 13984 4230
rect 14784 4266 14952 4271
rect 14986 4266 15053 4300
rect 15087 4290 15294 4300
rect 15328 4290 15384 4324
rect 15418 4290 15474 4324
rect 15508 4290 15564 4324
rect 15598 4290 15654 4324
rect 15688 4290 15744 4324
rect 15778 4290 15834 4324
rect 15868 4290 15924 4324
rect 15958 4290 16014 4324
rect 16048 4300 16582 4324
rect 16048 4290 16240 4300
rect 15087 4271 16240 4290
rect 15087 4266 15255 4271
rect 14784 4230 15255 4266
rect 14784 4211 15202 4230
rect 13799 4176 13984 4196
rect 13484 4140 13984 4176
rect 13484 4121 13914 4140
rect 13484 4087 13516 4121
rect 13550 4120 13914 4121
rect 13550 4087 13664 4120
rect 13484 4086 13664 4087
rect 13698 4086 13765 4120
rect 13799 4106 13914 4120
rect 13948 4106 13984 4140
rect 13799 4086 13984 4106
rect 13484 4050 13984 4086
rect 13484 4031 13914 4050
rect 13484 3997 13516 4031
rect 13550 4030 13914 4031
rect 13550 3997 13664 4030
rect 13484 3996 13664 3997
rect 13698 3996 13765 4030
rect 13799 4016 13914 4030
rect 13948 4016 13984 4050
rect 13799 3996 13984 4016
rect 13484 3960 13984 3996
rect 13484 3941 13914 3960
rect 13484 3907 13516 3941
rect 13550 3940 13914 3941
rect 13550 3907 13664 3940
rect 13484 3906 13664 3907
rect 13698 3906 13765 3940
rect 13799 3926 13914 3940
rect 13948 3926 13984 3960
rect 13799 3906 13984 3926
rect 13484 3870 13984 3906
rect 13484 3851 13914 3870
rect 13484 3817 13516 3851
rect 13550 3850 13914 3851
rect 13550 3817 13664 3850
rect 13484 3816 13664 3817
rect 13698 3816 13765 3850
rect 13799 3836 13914 3850
rect 13948 3836 13984 3870
rect 13799 3816 13984 3836
rect 13484 3780 13984 3816
rect 13484 3761 13914 3780
rect 13484 3727 13516 3761
rect 13550 3760 13914 3761
rect 13550 3727 13664 3760
rect 13484 3726 13664 3727
rect 13698 3726 13765 3760
rect 13799 3746 13914 3760
rect 13948 3746 13984 3780
rect 13799 3726 13984 3746
rect 13484 3690 13984 3726
rect 13484 3671 13914 3690
rect 13484 3637 13516 3671
rect 13550 3670 13914 3671
rect 13550 3637 13664 3670
rect 13484 3636 13664 3637
rect 13698 3636 13765 3670
rect 13799 3656 13914 3670
rect 13948 3656 13984 3690
rect 13799 3636 13984 3656
rect 13484 3600 13984 3636
rect 13484 3581 13914 3600
rect 13484 3547 13516 3581
rect 13550 3580 13914 3581
rect 13550 3547 13664 3580
rect 13484 3546 13664 3547
rect 13698 3546 13765 3580
rect 13799 3566 13914 3580
rect 13948 3566 13984 3600
rect 13799 3546 13984 3566
rect 12444 3490 12626 3510
rect 12444 3456 12477 3490
rect 12511 3476 12626 3490
rect 12660 3476 12684 3510
rect 12511 3456 12684 3476
rect 12444 3453 12684 3456
rect 13484 3510 13984 3546
rect 14029 4148 14723 4209
rect 14029 4114 14088 4148
rect 14122 4136 14178 4148
rect 14150 4114 14178 4136
rect 14212 4136 14268 4148
rect 14212 4114 14216 4136
rect 14029 4102 14116 4114
rect 14150 4102 14216 4114
rect 14250 4114 14268 4136
rect 14302 4136 14358 4148
rect 14302 4114 14316 4136
rect 14250 4102 14316 4114
rect 14350 4114 14358 4136
rect 14392 4136 14448 4148
rect 14482 4136 14538 4148
rect 14572 4136 14628 4148
rect 14392 4114 14416 4136
rect 14482 4114 14516 4136
rect 14572 4114 14616 4136
rect 14662 4114 14723 4148
rect 14350 4102 14416 4114
rect 14450 4102 14516 4114
rect 14550 4102 14616 4114
rect 14650 4102 14723 4114
rect 14029 4058 14723 4102
rect 14029 4024 14088 4058
rect 14122 4036 14178 4058
rect 14150 4024 14178 4036
rect 14212 4036 14268 4058
rect 14212 4024 14216 4036
rect 14029 4002 14116 4024
rect 14150 4002 14216 4024
rect 14250 4024 14268 4036
rect 14302 4036 14358 4058
rect 14302 4024 14316 4036
rect 14250 4002 14316 4024
rect 14350 4024 14358 4036
rect 14392 4036 14448 4058
rect 14482 4036 14538 4058
rect 14572 4036 14628 4058
rect 14392 4024 14416 4036
rect 14482 4024 14516 4036
rect 14572 4024 14616 4036
rect 14662 4024 14723 4058
rect 14350 4002 14416 4024
rect 14450 4002 14516 4024
rect 14550 4002 14616 4024
rect 14650 4002 14723 4024
rect 14029 3968 14723 4002
rect 14029 3934 14088 3968
rect 14122 3936 14178 3968
rect 14150 3934 14178 3936
rect 14212 3936 14268 3968
rect 14212 3934 14216 3936
rect 14029 3902 14116 3934
rect 14150 3902 14216 3934
rect 14250 3934 14268 3936
rect 14302 3936 14358 3968
rect 14302 3934 14316 3936
rect 14250 3902 14316 3934
rect 14350 3934 14358 3936
rect 14392 3936 14448 3968
rect 14482 3936 14538 3968
rect 14572 3936 14628 3968
rect 14392 3934 14416 3936
rect 14482 3934 14516 3936
rect 14572 3934 14616 3936
rect 14662 3934 14723 3968
rect 14350 3902 14416 3934
rect 14450 3902 14516 3934
rect 14550 3902 14616 3934
rect 14650 3902 14723 3934
rect 14029 3878 14723 3902
rect 14029 3844 14088 3878
rect 14122 3844 14178 3878
rect 14212 3844 14268 3878
rect 14302 3844 14358 3878
rect 14392 3844 14448 3878
rect 14482 3844 14538 3878
rect 14572 3844 14628 3878
rect 14662 3844 14723 3878
rect 14029 3836 14723 3844
rect 14029 3802 14116 3836
rect 14150 3802 14216 3836
rect 14250 3802 14316 3836
rect 14350 3802 14416 3836
rect 14450 3802 14516 3836
rect 14550 3802 14616 3836
rect 14650 3802 14723 3836
rect 14029 3788 14723 3802
rect 14029 3754 14088 3788
rect 14122 3754 14178 3788
rect 14212 3754 14268 3788
rect 14302 3754 14358 3788
rect 14392 3754 14448 3788
rect 14482 3754 14538 3788
rect 14572 3754 14628 3788
rect 14662 3754 14723 3788
rect 14029 3736 14723 3754
rect 14029 3702 14116 3736
rect 14150 3702 14216 3736
rect 14250 3702 14316 3736
rect 14350 3702 14416 3736
rect 14450 3702 14516 3736
rect 14550 3702 14616 3736
rect 14650 3702 14723 3736
rect 14029 3698 14723 3702
rect 14029 3664 14088 3698
rect 14122 3664 14178 3698
rect 14212 3664 14268 3698
rect 14302 3664 14358 3698
rect 14392 3664 14448 3698
rect 14482 3664 14538 3698
rect 14572 3664 14628 3698
rect 14662 3664 14723 3698
rect 14029 3636 14723 3664
rect 14029 3608 14116 3636
rect 14150 3608 14216 3636
rect 14029 3574 14088 3608
rect 14150 3602 14178 3608
rect 14122 3574 14178 3602
rect 14212 3602 14216 3608
rect 14250 3608 14316 3636
rect 14250 3602 14268 3608
rect 14212 3574 14268 3602
rect 14302 3602 14316 3608
rect 14350 3608 14416 3636
rect 14450 3608 14516 3636
rect 14550 3608 14616 3636
rect 14650 3608 14723 3636
rect 14350 3602 14358 3608
rect 14302 3574 14358 3602
rect 14392 3602 14416 3608
rect 14482 3602 14516 3608
rect 14572 3602 14616 3608
rect 14392 3574 14448 3602
rect 14482 3574 14538 3602
rect 14572 3574 14628 3602
rect 14662 3574 14723 3608
rect 14029 3515 14723 3574
rect 14784 4177 14804 4211
rect 14838 4210 15202 4211
rect 14838 4177 14952 4210
rect 14784 4176 14952 4177
rect 14986 4176 15053 4210
rect 15087 4196 15202 4210
rect 15236 4196 15255 4230
rect 16073 4266 16240 4271
rect 16274 4266 16341 4300
rect 16375 4290 16582 4300
rect 16616 4290 16672 4324
rect 16706 4290 16762 4324
rect 16796 4290 16852 4324
rect 16886 4290 16942 4324
rect 16976 4290 17032 4324
rect 17066 4290 17122 4324
rect 17156 4290 17212 4324
rect 17246 4290 17302 4324
rect 17336 4300 17870 4324
rect 17336 4290 17528 4300
rect 16375 4271 17528 4290
rect 16375 4266 16543 4271
rect 16073 4230 16543 4266
rect 16073 4211 16490 4230
rect 15087 4176 15255 4196
rect 14784 4140 15255 4176
rect 14784 4121 15202 4140
rect 14784 4087 14804 4121
rect 14838 4120 15202 4121
rect 14838 4087 14952 4120
rect 14784 4086 14952 4087
rect 14986 4086 15053 4120
rect 15087 4106 15202 4120
rect 15236 4106 15255 4140
rect 15087 4086 15255 4106
rect 14784 4050 15255 4086
rect 14784 4031 15202 4050
rect 14784 3997 14804 4031
rect 14838 4030 15202 4031
rect 14838 3997 14952 4030
rect 14784 3996 14952 3997
rect 14986 3996 15053 4030
rect 15087 4016 15202 4030
rect 15236 4016 15255 4050
rect 15087 3996 15255 4016
rect 14784 3960 15255 3996
rect 14784 3941 15202 3960
rect 14784 3907 14804 3941
rect 14838 3940 15202 3941
rect 14838 3907 14952 3940
rect 14784 3906 14952 3907
rect 14986 3906 15053 3940
rect 15087 3926 15202 3940
rect 15236 3926 15255 3960
rect 15087 3906 15255 3926
rect 14784 3870 15255 3906
rect 14784 3851 15202 3870
rect 14784 3817 14804 3851
rect 14838 3850 15202 3851
rect 14838 3817 14952 3850
rect 14784 3816 14952 3817
rect 14986 3816 15053 3850
rect 15087 3836 15202 3850
rect 15236 3836 15255 3870
rect 15087 3816 15255 3836
rect 14784 3780 15255 3816
rect 14784 3761 15202 3780
rect 14784 3727 14804 3761
rect 14838 3760 15202 3761
rect 14838 3727 14952 3760
rect 14784 3726 14952 3727
rect 14986 3726 15053 3760
rect 15087 3746 15202 3760
rect 15236 3746 15255 3780
rect 15087 3726 15255 3746
rect 14784 3690 15255 3726
rect 14784 3671 15202 3690
rect 14784 3637 14804 3671
rect 14838 3670 15202 3671
rect 14838 3637 14952 3670
rect 14784 3636 14952 3637
rect 14986 3636 15053 3670
rect 15087 3656 15202 3670
rect 15236 3656 15255 3690
rect 15087 3636 15255 3656
rect 14784 3600 15255 3636
rect 14784 3581 15202 3600
rect 14784 3547 14804 3581
rect 14838 3580 15202 3581
rect 14838 3547 14952 3580
rect 14784 3546 14952 3547
rect 14986 3546 15053 3580
rect 15087 3566 15202 3580
rect 15236 3566 15255 3600
rect 15087 3546 15255 3566
rect 13484 3491 13914 3510
rect 13484 3457 13516 3491
rect 13550 3490 13914 3491
rect 13550 3457 13664 3490
rect 13484 3456 13664 3457
rect 13698 3456 13765 3490
rect 13799 3476 13914 3490
rect 13948 3476 13984 3510
rect 13799 3456 13984 3476
rect 13484 3453 13984 3456
rect 14784 3510 15255 3546
rect 15317 4148 16011 4209
rect 15317 4114 15376 4148
rect 15410 4136 15466 4148
rect 15438 4114 15466 4136
rect 15500 4136 15556 4148
rect 15500 4114 15504 4136
rect 15317 4102 15404 4114
rect 15438 4102 15504 4114
rect 15538 4114 15556 4136
rect 15590 4136 15646 4148
rect 15590 4114 15604 4136
rect 15538 4102 15604 4114
rect 15638 4114 15646 4136
rect 15680 4136 15736 4148
rect 15770 4136 15826 4148
rect 15860 4136 15916 4148
rect 15680 4114 15704 4136
rect 15770 4114 15804 4136
rect 15860 4114 15904 4136
rect 15950 4114 16011 4148
rect 15638 4102 15704 4114
rect 15738 4102 15804 4114
rect 15838 4102 15904 4114
rect 15938 4102 16011 4114
rect 15317 4058 16011 4102
rect 15317 4024 15376 4058
rect 15410 4036 15466 4058
rect 15438 4024 15466 4036
rect 15500 4036 15556 4058
rect 15500 4024 15504 4036
rect 15317 4002 15404 4024
rect 15438 4002 15504 4024
rect 15538 4024 15556 4036
rect 15590 4036 15646 4058
rect 15590 4024 15604 4036
rect 15538 4002 15604 4024
rect 15638 4024 15646 4036
rect 15680 4036 15736 4058
rect 15770 4036 15826 4058
rect 15860 4036 15916 4058
rect 15680 4024 15704 4036
rect 15770 4024 15804 4036
rect 15860 4024 15904 4036
rect 15950 4024 16011 4058
rect 15638 4002 15704 4024
rect 15738 4002 15804 4024
rect 15838 4002 15904 4024
rect 15938 4002 16011 4024
rect 15317 3968 16011 4002
rect 15317 3934 15376 3968
rect 15410 3936 15466 3968
rect 15438 3934 15466 3936
rect 15500 3936 15556 3968
rect 15500 3934 15504 3936
rect 15317 3902 15404 3934
rect 15438 3902 15504 3934
rect 15538 3934 15556 3936
rect 15590 3936 15646 3968
rect 15590 3934 15604 3936
rect 15538 3902 15604 3934
rect 15638 3934 15646 3936
rect 15680 3936 15736 3968
rect 15770 3936 15826 3968
rect 15860 3936 15916 3968
rect 15680 3934 15704 3936
rect 15770 3934 15804 3936
rect 15860 3934 15904 3936
rect 15950 3934 16011 3968
rect 15638 3902 15704 3934
rect 15738 3902 15804 3934
rect 15838 3902 15904 3934
rect 15938 3902 16011 3934
rect 15317 3878 16011 3902
rect 15317 3844 15376 3878
rect 15410 3844 15466 3878
rect 15500 3844 15556 3878
rect 15590 3844 15646 3878
rect 15680 3844 15736 3878
rect 15770 3844 15826 3878
rect 15860 3844 15916 3878
rect 15950 3844 16011 3878
rect 15317 3836 16011 3844
rect 15317 3802 15404 3836
rect 15438 3802 15504 3836
rect 15538 3802 15604 3836
rect 15638 3802 15704 3836
rect 15738 3802 15804 3836
rect 15838 3802 15904 3836
rect 15938 3802 16011 3836
rect 15317 3788 16011 3802
rect 15317 3754 15376 3788
rect 15410 3754 15466 3788
rect 15500 3754 15556 3788
rect 15590 3754 15646 3788
rect 15680 3754 15736 3788
rect 15770 3754 15826 3788
rect 15860 3754 15916 3788
rect 15950 3754 16011 3788
rect 15317 3736 16011 3754
rect 15317 3702 15404 3736
rect 15438 3702 15504 3736
rect 15538 3702 15604 3736
rect 15638 3702 15704 3736
rect 15738 3702 15804 3736
rect 15838 3702 15904 3736
rect 15938 3702 16011 3736
rect 15317 3698 16011 3702
rect 15317 3664 15376 3698
rect 15410 3664 15466 3698
rect 15500 3664 15556 3698
rect 15590 3664 15646 3698
rect 15680 3664 15736 3698
rect 15770 3664 15826 3698
rect 15860 3664 15916 3698
rect 15950 3664 16011 3698
rect 15317 3636 16011 3664
rect 15317 3608 15404 3636
rect 15438 3608 15504 3636
rect 15317 3574 15376 3608
rect 15438 3602 15466 3608
rect 15410 3574 15466 3602
rect 15500 3602 15504 3608
rect 15538 3608 15604 3636
rect 15538 3602 15556 3608
rect 15500 3574 15556 3602
rect 15590 3602 15604 3608
rect 15638 3608 15704 3636
rect 15738 3608 15804 3636
rect 15838 3608 15904 3636
rect 15938 3608 16011 3636
rect 15638 3602 15646 3608
rect 15590 3574 15646 3602
rect 15680 3602 15704 3608
rect 15770 3602 15804 3608
rect 15860 3602 15904 3608
rect 15680 3574 15736 3602
rect 15770 3574 15826 3602
rect 15860 3574 15916 3602
rect 15950 3574 16011 3608
rect 15317 3515 16011 3574
rect 16073 4177 16092 4211
rect 16126 4210 16490 4211
rect 16126 4177 16240 4210
rect 16073 4176 16240 4177
rect 16274 4176 16341 4210
rect 16375 4196 16490 4210
rect 16524 4196 16543 4230
rect 17361 4266 17528 4271
rect 17562 4266 17629 4300
rect 17663 4290 17870 4300
rect 17904 4290 17960 4324
rect 17994 4290 18050 4324
rect 18084 4290 18140 4324
rect 18174 4290 18230 4324
rect 18264 4290 18320 4324
rect 18354 4290 18410 4324
rect 18444 4290 18500 4324
rect 18534 4290 18590 4324
rect 18624 4300 18884 4324
rect 18624 4290 18816 4300
rect 17663 4271 18816 4290
rect 17663 4266 17831 4271
rect 17361 4230 17831 4266
rect 17361 4211 17778 4230
rect 16375 4176 16543 4196
rect 16073 4140 16543 4176
rect 16073 4121 16490 4140
rect 16073 4087 16092 4121
rect 16126 4120 16490 4121
rect 16126 4087 16240 4120
rect 16073 4086 16240 4087
rect 16274 4086 16341 4120
rect 16375 4106 16490 4120
rect 16524 4106 16543 4140
rect 16375 4086 16543 4106
rect 16073 4050 16543 4086
rect 16073 4031 16490 4050
rect 16073 3997 16092 4031
rect 16126 4030 16490 4031
rect 16126 3997 16240 4030
rect 16073 3996 16240 3997
rect 16274 3996 16341 4030
rect 16375 4016 16490 4030
rect 16524 4016 16543 4050
rect 16375 3996 16543 4016
rect 16073 3960 16543 3996
rect 16073 3941 16490 3960
rect 16073 3907 16092 3941
rect 16126 3940 16490 3941
rect 16126 3907 16240 3940
rect 16073 3906 16240 3907
rect 16274 3906 16341 3940
rect 16375 3926 16490 3940
rect 16524 3926 16543 3960
rect 16375 3906 16543 3926
rect 16073 3870 16543 3906
rect 16073 3851 16490 3870
rect 16073 3817 16092 3851
rect 16126 3850 16490 3851
rect 16126 3817 16240 3850
rect 16073 3816 16240 3817
rect 16274 3816 16341 3850
rect 16375 3836 16490 3850
rect 16524 3836 16543 3870
rect 16375 3816 16543 3836
rect 16073 3780 16543 3816
rect 16073 3761 16490 3780
rect 16073 3727 16092 3761
rect 16126 3760 16490 3761
rect 16126 3727 16240 3760
rect 16073 3726 16240 3727
rect 16274 3726 16341 3760
rect 16375 3746 16490 3760
rect 16524 3746 16543 3780
rect 16375 3726 16543 3746
rect 16073 3690 16543 3726
rect 16073 3671 16490 3690
rect 16073 3637 16092 3671
rect 16126 3670 16490 3671
rect 16126 3637 16240 3670
rect 16073 3636 16240 3637
rect 16274 3636 16341 3670
rect 16375 3656 16490 3670
rect 16524 3656 16543 3690
rect 16375 3636 16543 3656
rect 16073 3600 16543 3636
rect 16073 3581 16490 3600
rect 16073 3547 16092 3581
rect 16126 3580 16490 3581
rect 16126 3547 16240 3580
rect 16073 3546 16240 3547
rect 16274 3546 16341 3580
rect 16375 3566 16490 3580
rect 16524 3566 16543 3600
rect 16375 3546 16543 3566
rect 14784 3491 15202 3510
rect 14784 3457 14804 3491
rect 14838 3490 15202 3491
rect 14838 3457 14952 3490
rect 14784 3456 14952 3457
rect 14986 3456 15053 3490
rect 15087 3476 15202 3490
rect 15236 3476 15255 3510
rect 15087 3456 15255 3476
rect 14784 3453 15255 3456
rect 16073 3510 16543 3546
rect 16605 4148 17299 4209
rect 16605 4114 16664 4148
rect 16698 4136 16754 4148
rect 16726 4114 16754 4136
rect 16788 4136 16844 4148
rect 16788 4114 16792 4136
rect 16605 4102 16692 4114
rect 16726 4102 16792 4114
rect 16826 4114 16844 4136
rect 16878 4136 16934 4148
rect 16878 4114 16892 4136
rect 16826 4102 16892 4114
rect 16926 4114 16934 4136
rect 16968 4136 17024 4148
rect 17058 4136 17114 4148
rect 17148 4136 17204 4148
rect 16968 4114 16992 4136
rect 17058 4114 17092 4136
rect 17148 4114 17192 4136
rect 17238 4114 17299 4148
rect 16926 4102 16992 4114
rect 17026 4102 17092 4114
rect 17126 4102 17192 4114
rect 17226 4102 17299 4114
rect 16605 4058 17299 4102
rect 16605 4024 16664 4058
rect 16698 4036 16754 4058
rect 16726 4024 16754 4036
rect 16788 4036 16844 4058
rect 16788 4024 16792 4036
rect 16605 4002 16692 4024
rect 16726 4002 16792 4024
rect 16826 4024 16844 4036
rect 16878 4036 16934 4058
rect 16878 4024 16892 4036
rect 16826 4002 16892 4024
rect 16926 4024 16934 4036
rect 16968 4036 17024 4058
rect 17058 4036 17114 4058
rect 17148 4036 17204 4058
rect 16968 4024 16992 4036
rect 17058 4024 17092 4036
rect 17148 4024 17192 4036
rect 17238 4024 17299 4058
rect 16926 4002 16992 4024
rect 17026 4002 17092 4024
rect 17126 4002 17192 4024
rect 17226 4002 17299 4024
rect 16605 3968 17299 4002
rect 16605 3934 16664 3968
rect 16698 3936 16754 3968
rect 16726 3934 16754 3936
rect 16788 3936 16844 3968
rect 16788 3934 16792 3936
rect 16605 3902 16692 3934
rect 16726 3902 16792 3934
rect 16826 3934 16844 3936
rect 16878 3936 16934 3968
rect 16878 3934 16892 3936
rect 16826 3902 16892 3934
rect 16926 3934 16934 3936
rect 16968 3936 17024 3968
rect 17058 3936 17114 3968
rect 17148 3936 17204 3968
rect 16968 3934 16992 3936
rect 17058 3934 17092 3936
rect 17148 3934 17192 3936
rect 17238 3934 17299 3968
rect 16926 3902 16992 3934
rect 17026 3902 17092 3934
rect 17126 3902 17192 3934
rect 17226 3902 17299 3934
rect 16605 3878 17299 3902
rect 16605 3844 16664 3878
rect 16698 3844 16754 3878
rect 16788 3844 16844 3878
rect 16878 3844 16934 3878
rect 16968 3844 17024 3878
rect 17058 3844 17114 3878
rect 17148 3844 17204 3878
rect 17238 3844 17299 3878
rect 16605 3836 17299 3844
rect 16605 3802 16692 3836
rect 16726 3802 16792 3836
rect 16826 3802 16892 3836
rect 16926 3802 16992 3836
rect 17026 3802 17092 3836
rect 17126 3802 17192 3836
rect 17226 3802 17299 3836
rect 16605 3788 17299 3802
rect 16605 3754 16664 3788
rect 16698 3754 16754 3788
rect 16788 3754 16844 3788
rect 16878 3754 16934 3788
rect 16968 3754 17024 3788
rect 17058 3754 17114 3788
rect 17148 3754 17204 3788
rect 17238 3754 17299 3788
rect 16605 3736 17299 3754
rect 16605 3702 16692 3736
rect 16726 3702 16792 3736
rect 16826 3702 16892 3736
rect 16926 3702 16992 3736
rect 17026 3702 17092 3736
rect 17126 3702 17192 3736
rect 17226 3702 17299 3736
rect 16605 3698 17299 3702
rect 16605 3664 16664 3698
rect 16698 3664 16754 3698
rect 16788 3664 16844 3698
rect 16878 3664 16934 3698
rect 16968 3664 17024 3698
rect 17058 3664 17114 3698
rect 17148 3664 17204 3698
rect 17238 3664 17299 3698
rect 16605 3636 17299 3664
rect 16605 3608 16692 3636
rect 16726 3608 16792 3636
rect 16605 3574 16664 3608
rect 16726 3602 16754 3608
rect 16698 3574 16754 3602
rect 16788 3602 16792 3608
rect 16826 3608 16892 3636
rect 16826 3602 16844 3608
rect 16788 3574 16844 3602
rect 16878 3602 16892 3608
rect 16926 3608 16992 3636
rect 17026 3608 17092 3636
rect 17126 3608 17192 3636
rect 17226 3608 17299 3636
rect 16926 3602 16934 3608
rect 16878 3574 16934 3602
rect 16968 3602 16992 3608
rect 17058 3602 17092 3608
rect 17148 3602 17192 3608
rect 16968 3574 17024 3602
rect 17058 3574 17114 3602
rect 17148 3574 17204 3602
rect 17238 3574 17299 3608
rect 16605 3515 17299 3574
rect 17361 4177 17380 4211
rect 17414 4210 17778 4211
rect 17414 4177 17528 4210
rect 17361 4176 17528 4177
rect 17562 4176 17629 4210
rect 17663 4196 17778 4210
rect 17812 4196 17831 4230
rect 18649 4266 18816 4271
rect 18850 4266 18884 4300
rect 18649 4211 18884 4266
rect 17663 4176 17831 4196
rect 17361 4140 17831 4176
rect 17361 4121 17778 4140
rect 17361 4087 17380 4121
rect 17414 4120 17778 4121
rect 17414 4087 17528 4120
rect 17361 4086 17528 4087
rect 17562 4086 17629 4120
rect 17663 4106 17778 4120
rect 17812 4106 17831 4140
rect 17663 4086 17831 4106
rect 17361 4050 17831 4086
rect 17361 4031 17778 4050
rect 17361 3997 17380 4031
rect 17414 4030 17778 4031
rect 17414 3997 17528 4030
rect 17361 3996 17528 3997
rect 17562 3996 17629 4030
rect 17663 4016 17778 4030
rect 17812 4016 17831 4050
rect 17663 3996 17831 4016
rect 17361 3960 17831 3996
rect 17361 3941 17778 3960
rect 17361 3907 17380 3941
rect 17414 3940 17778 3941
rect 17414 3907 17528 3940
rect 17361 3906 17528 3907
rect 17562 3906 17629 3940
rect 17663 3926 17778 3940
rect 17812 3926 17831 3960
rect 17663 3906 17831 3926
rect 17361 3870 17831 3906
rect 17361 3851 17778 3870
rect 17361 3817 17380 3851
rect 17414 3850 17778 3851
rect 17414 3817 17528 3850
rect 17361 3816 17528 3817
rect 17562 3816 17629 3850
rect 17663 3836 17778 3850
rect 17812 3836 17831 3870
rect 17663 3816 17831 3836
rect 17361 3780 17831 3816
rect 17361 3761 17778 3780
rect 17361 3727 17380 3761
rect 17414 3760 17778 3761
rect 17414 3727 17528 3760
rect 17361 3726 17528 3727
rect 17562 3726 17629 3760
rect 17663 3746 17778 3760
rect 17812 3746 17831 3780
rect 17663 3726 17831 3746
rect 17361 3690 17831 3726
rect 17361 3671 17778 3690
rect 17361 3637 17380 3671
rect 17414 3670 17778 3671
rect 17414 3637 17528 3670
rect 17361 3636 17528 3637
rect 17562 3636 17629 3670
rect 17663 3656 17778 3670
rect 17812 3656 17831 3690
rect 17663 3636 17831 3656
rect 17361 3600 17831 3636
rect 17361 3581 17778 3600
rect 17361 3547 17380 3581
rect 17414 3580 17778 3581
rect 17414 3547 17528 3580
rect 17361 3546 17528 3547
rect 17562 3546 17629 3580
rect 17663 3566 17778 3580
rect 17812 3566 17831 3600
rect 17663 3546 17831 3566
rect 16073 3491 16490 3510
rect 16073 3457 16092 3491
rect 16126 3490 16490 3491
rect 16126 3457 16240 3490
rect 16073 3456 16240 3457
rect 16274 3456 16341 3490
rect 16375 3476 16490 3490
rect 16524 3476 16543 3510
rect 16375 3456 16543 3476
rect 16073 3453 16543 3456
rect 17361 3510 17831 3546
rect 17893 4148 18587 4209
rect 17893 4114 17952 4148
rect 17986 4136 18042 4148
rect 18014 4114 18042 4136
rect 18076 4136 18132 4148
rect 18076 4114 18080 4136
rect 17893 4102 17980 4114
rect 18014 4102 18080 4114
rect 18114 4114 18132 4136
rect 18166 4136 18222 4148
rect 18166 4114 18180 4136
rect 18114 4102 18180 4114
rect 18214 4114 18222 4136
rect 18256 4136 18312 4148
rect 18346 4136 18402 4148
rect 18436 4136 18492 4148
rect 18256 4114 18280 4136
rect 18346 4114 18380 4136
rect 18436 4114 18480 4136
rect 18526 4114 18587 4148
rect 18214 4102 18280 4114
rect 18314 4102 18380 4114
rect 18414 4102 18480 4114
rect 18514 4102 18587 4114
rect 17893 4058 18587 4102
rect 17893 4024 17952 4058
rect 17986 4036 18042 4058
rect 18014 4024 18042 4036
rect 18076 4036 18132 4058
rect 18076 4024 18080 4036
rect 17893 4002 17980 4024
rect 18014 4002 18080 4024
rect 18114 4024 18132 4036
rect 18166 4036 18222 4058
rect 18166 4024 18180 4036
rect 18114 4002 18180 4024
rect 18214 4024 18222 4036
rect 18256 4036 18312 4058
rect 18346 4036 18402 4058
rect 18436 4036 18492 4058
rect 18256 4024 18280 4036
rect 18346 4024 18380 4036
rect 18436 4024 18480 4036
rect 18526 4024 18587 4058
rect 18214 4002 18280 4024
rect 18314 4002 18380 4024
rect 18414 4002 18480 4024
rect 18514 4002 18587 4024
rect 17893 3968 18587 4002
rect 17893 3934 17952 3968
rect 17986 3936 18042 3968
rect 18014 3934 18042 3936
rect 18076 3936 18132 3968
rect 18076 3934 18080 3936
rect 17893 3902 17980 3934
rect 18014 3902 18080 3934
rect 18114 3934 18132 3936
rect 18166 3936 18222 3968
rect 18166 3934 18180 3936
rect 18114 3902 18180 3934
rect 18214 3934 18222 3936
rect 18256 3936 18312 3968
rect 18346 3936 18402 3968
rect 18436 3936 18492 3968
rect 18256 3934 18280 3936
rect 18346 3934 18380 3936
rect 18436 3934 18480 3936
rect 18526 3934 18587 3968
rect 18214 3902 18280 3934
rect 18314 3902 18380 3934
rect 18414 3902 18480 3934
rect 18514 3902 18587 3934
rect 17893 3878 18587 3902
rect 17893 3844 17952 3878
rect 17986 3844 18042 3878
rect 18076 3844 18132 3878
rect 18166 3844 18222 3878
rect 18256 3844 18312 3878
rect 18346 3844 18402 3878
rect 18436 3844 18492 3878
rect 18526 3844 18587 3878
rect 17893 3836 18587 3844
rect 17893 3802 17980 3836
rect 18014 3802 18080 3836
rect 18114 3802 18180 3836
rect 18214 3802 18280 3836
rect 18314 3802 18380 3836
rect 18414 3802 18480 3836
rect 18514 3802 18587 3836
rect 17893 3788 18587 3802
rect 17893 3754 17952 3788
rect 17986 3754 18042 3788
rect 18076 3754 18132 3788
rect 18166 3754 18222 3788
rect 18256 3754 18312 3788
rect 18346 3754 18402 3788
rect 18436 3754 18492 3788
rect 18526 3754 18587 3788
rect 17893 3736 18587 3754
rect 17893 3702 17980 3736
rect 18014 3702 18080 3736
rect 18114 3702 18180 3736
rect 18214 3702 18280 3736
rect 18314 3702 18380 3736
rect 18414 3702 18480 3736
rect 18514 3702 18587 3736
rect 17893 3698 18587 3702
rect 17893 3664 17952 3698
rect 17986 3664 18042 3698
rect 18076 3664 18132 3698
rect 18166 3664 18222 3698
rect 18256 3664 18312 3698
rect 18346 3664 18402 3698
rect 18436 3664 18492 3698
rect 18526 3664 18587 3698
rect 17893 3636 18587 3664
rect 17893 3608 17980 3636
rect 18014 3608 18080 3636
rect 17893 3574 17952 3608
rect 18014 3602 18042 3608
rect 17986 3574 18042 3602
rect 18076 3602 18080 3608
rect 18114 3608 18180 3636
rect 18114 3602 18132 3608
rect 18076 3574 18132 3602
rect 18166 3602 18180 3608
rect 18214 3608 18280 3636
rect 18314 3608 18380 3636
rect 18414 3608 18480 3636
rect 18514 3608 18587 3636
rect 18214 3602 18222 3608
rect 18166 3574 18222 3602
rect 18256 3602 18280 3608
rect 18346 3602 18380 3608
rect 18436 3602 18480 3608
rect 18256 3574 18312 3602
rect 18346 3574 18402 3602
rect 18436 3574 18492 3602
rect 18526 3574 18587 3608
rect 17893 3515 18587 3574
rect 18649 4177 18668 4211
rect 18702 4210 18884 4211
rect 18702 4177 18816 4210
rect 18649 4176 18816 4177
rect 18850 4176 18884 4210
rect 18649 4121 18884 4176
rect 18649 4087 18668 4121
rect 18702 4120 18884 4121
rect 18702 4087 18816 4120
rect 18649 4086 18816 4087
rect 18850 4086 18884 4120
rect 18649 4031 18884 4086
rect 18649 3997 18668 4031
rect 18702 4030 18884 4031
rect 18702 3997 18816 4030
rect 18649 3996 18816 3997
rect 18850 3996 18884 4030
rect 18649 3941 18884 3996
rect 18649 3907 18668 3941
rect 18702 3940 18884 3941
rect 18702 3907 18816 3940
rect 18649 3906 18816 3907
rect 18850 3906 18884 3940
rect 18649 3851 18884 3906
rect 18649 3817 18668 3851
rect 18702 3850 18884 3851
rect 18702 3817 18816 3850
rect 18649 3816 18816 3817
rect 18850 3816 18884 3850
rect 18649 3761 18884 3816
rect 18649 3727 18668 3761
rect 18702 3760 18884 3761
rect 18702 3727 18816 3760
rect 18649 3726 18816 3727
rect 18850 3726 18884 3760
rect 18649 3671 18884 3726
rect 18649 3637 18668 3671
rect 18702 3670 18884 3671
rect 18702 3637 18816 3670
rect 18649 3636 18816 3637
rect 18850 3636 18884 3670
rect 18649 3581 18884 3636
rect 18649 3547 18668 3581
rect 18702 3580 18884 3581
rect 18702 3547 18816 3580
rect 18649 3546 18816 3547
rect 18850 3546 18884 3580
rect 17361 3491 17778 3510
rect 17361 3457 17380 3491
rect 17414 3490 17778 3491
rect 17414 3457 17528 3490
rect 17361 3456 17528 3457
rect 17562 3456 17629 3490
rect 17663 3476 17778 3490
rect 17812 3476 17831 3510
rect 17663 3456 17831 3476
rect 17361 3453 17831 3456
rect 18649 3491 18884 3546
rect 18649 3457 18668 3491
rect 18702 3490 18884 3491
rect 18702 3457 18816 3490
rect 18649 3456 18816 3457
rect 18850 3456 18884 3490
rect 18649 3453 18884 3456
rect 12444 3434 18884 3453
rect 12444 3400 12684 3434
rect 12718 3400 12774 3434
rect 12808 3400 12864 3434
rect 12898 3400 12954 3434
rect 12988 3400 13044 3434
rect 13078 3400 13134 3434
rect 13168 3400 13224 3434
rect 13258 3400 13314 3434
rect 13348 3400 13404 3434
rect 13438 3400 13972 3434
rect 14006 3400 14062 3434
rect 14096 3400 14152 3434
rect 14186 3400 14242 3434
rect 14276 3400 14332 3434
rect 14366 3400 14422 3434
rect 14456 3400 14512 3434
rect 14546 3400 14602 3434
rect 14636 3400 14692 3434
rect 14726 3400 15260 3434
rect 15294 3400 15350 3434
rect 15384 3400 15440 3434
rect 15474 3400 15530 3434
rect 15564 3400 15620 3434
rect 15654 3400 15710 3434
rect 15744 3400 15800 3434
rect 15834 3400 15890 3434
rect 15924 3400 15980 3434
rect 16014 3400 16548 3434
rect 16582 3400 16638 3434
rect 16672 3400 16728 3434
rect 16762 3400 16818 3434
rect 16852 3400 16908 3434
rect 16942 3400 16998 3434
rect 17032 3400 17088 3434
rect 17122 3400 17178 3434
rect 17212 3400 17268 3434
rect 17302 3400 17836 3434
rect 17870 3400 17926 3434
rect 17960 3400 18016 3434
rect 18050 3400 18106 3434
rect 18140 3400 18196 3434
rect 18230 3400 18286 3434
rect 18320 3400 18376 3434
rect 18410 3400 18466 3434
rect 18500 3400 18556 3434
rect 18590 3400 18884 3434
rect 12444 3366 12477 3400
rect 12511 3381 13664 3400
rect 12511 3366 12684 3381
rect 12444 3317 12684 3366
rect 13484 3366 13664 3381
rect 13698 3366 13765 3400
rect 13799 3381 14952 3400
rect 13799 3366 13984 3381
rect 13484 3317 13984 3366
rect 14784 3366 14952 3381
rect 14986 3366 15053 3400
rect 15087 3381 16240 3400
rect 15087 3366 15184 3381
rect 14784 3317 15184 3366
rect 16084 3366 16240 3381
rect 16274 3366 16341 3400
rect 16375 3381 17528 3400
rect 16375 3366 16484 3381
rect 16084 3317 16484 3366
rect 17384 3366 17528 3381
rect 17562 3366 17629 3400
rect 17663 3381 18816 3400
rect 17663 3366 17784 3381
rect 17384 3317 17784 3366
rect 18684 3366 18816 3381
rect 18850 3366 18884 3400
rect 18684 3317 18884 3366
rect 12444 3310 18884 3317
rect 12444 3276 12477 3310
rect 12511 3287 13664 3310
rect 12511 3276 12578 3287
rect 12444 3253 12578 3276
rect 12612 3253 12668 3287
rect 12702 3253 12758 3287
rect 12792 3253 12848 3287
rect 12882 3253 12938 3287
rect 12972 3253 13028 3287
rect 13062 3253 13118 3287
rect 13152 3253 13208 3287
rect 13242 3253 13298 3287
rect 13332 3253 13388 3287
rect 13422 3253 13478 3287
rect 13512 3253 13568 3287
rect 13602 3276 13664 3287
rect 13698 3276 13765 3310
rect 13799 3287 14952 3310
rect 13799 3276 13866 3287
rect 13602 3253 13866 3276
rect 13900 3253 13956 3287
rect 13990 3253 14046 3287
rect 14080 3253 14136 3287
rect 14170 3253 14226 3287
rect 14260 3253 14316 3287
rect 14350 3253 14406 3287
rect 14440 3253 14496 3287
rect 14530 3253 14586 3287
rect 14620 3253 14676 3287
rect 14710 3253 14766 3287
rect 14800 3253 14856 3287
rect 14890 3276 14952 3287
rect 14986 3276 15053 3310
rect 15087 3287 16240 3310
rect 15087 3276 15154 3287
rect 14890 3253 15154 3276
rect 15188 3253 15244 3287
rect 15278 3253 15334 3287
rect 15368 3253 15424 3287
rect 15458 3253 15514 3287
rect 15548 3253 15604 3287
rect 15638 3253 15694 3287
rect 15728 3253 15784 3287
rect 15818 3253 15874 3287
rect 15908 3253 15964 3287
rect 15998 3253 16054 3287
rect 16088 3253 16144 3287
rect 16178 3276 16240 3287
rect 16274 3276 16341 3310
rect 16375 3287 17528 3310
rect 16375 3276 16442 3287
rect 16178 3253 16442 3276
rect 16476 3253 16532 3287
rect 16566 3253 16622 3287
rect 16656 3253 16712 3287
rect 16746 3253 16802 3287
rect 16836 3253 16892 3287
rect 16926 3253 16982 3287
rect 17016 3253 17072 3287
rect 17106 3253 17162 3287
rect 17196 3253 17252 3287
rect 17286 3253 17342 3287
rect 17376 3253 17432 3287
rect 17466 3276 17528 3287
rect 17562 3276 17629 3310
rect 17663 3287 18816 3310
rect 17663 3276 17730 3287
rect 17466 3253 17730 3276
rect 17764 3253 17820 3287
rect 17854 3253 17910 3287
rect 17944 3253 18000 3287
rect 18034 3253 18090 3287
rect 18124 3253 18180 3287
rect 18214 3253 18270 3287
rect 18304 3253 18360 3287
rect 18394 3253 18450 3287
rect 18484 3253 18540 3287
rect 18574 3253 18630 3287
rect 18664 3253 18720 3287
rect 18754 3276 18816 3287
rect 18850 3276 18884 3310
rect 18754 3253 18884 3276
rect 12444 3186 18884 3253
rect 12444 3152 12578 3186
rect 12612 3152 12668 3186
rect 12702 3152 12758 3186
rect 12792 3152 12848 3186
rect 12882 3152 12938 3186
rect 12972 3152 13028 3186
rect 13062 3152 13118 3186
rect 13152 3152 13208 3186
rect 13242 3152 13298 3186
rect 13332 3152 13388 3186
rect 13422 3152 13478 3186
rect 13512 3152 13568 3186
rect 13602 3152 13866 3186
rect 13900 3152 13956 3186
rect 13990 3152 14046 3186
rect 14080 3152 14136 3186
rect 14170 3152 14226 3186
rect 14260 3152 14316 3186
rect 14350 3152 14406 3186
rect 14440 3152 14496 3186
rect 14530 3152 14586 3186
rect 14620 3152 14676 3186
rect 14710 3152 14766 3186
rect 14800 3152 14856 3186
rect 14890 3152 15154 3186
rect 15188 3152 15244 3186
rect 15278 3152 15334 3186
rect 15368 3152 15424 3186
rect 15458 3152 15514 3186
rect 15548 3152 15604 3186
rect 15638 3152 15694 3186
rect 15728 3152 15784 3186
rect 15818 3152 15874 3186
rect 15908 3152 15964 3186
rect 15998 3152 16054 3186
rect 16088 3152 16144 3186
rect 16178 3152 16442 3186
rect 16476 3152 16532 3186
rect 16566 3152 16622 3186
rect 16656 3152 16712 3186
rect 16746 3152 16802 3186
rect 16836 3152 16892 3186
rect 16926 3152 16982 3186
rect 17016 3152 17072 3186
rect 17106 3152 17162 3186
rect 17196 3152 17252 3186
rect 17286 3152 17342 3186
rect 17376 3152 17432 3186
rect 17466 3152 17730 3186
rect 17764 3152 17820 3186
rect 17854 3152 17910 3186
rect 17944 3152 18000 3186
rect 18034 3152 18090 3186
rect 18124 3152 18180 3186
rect 18214 3152 18270 3186
rect 18304 3152 18360 3186
rect 18394 3152 18450 3186
rect 18484 3152 18540 3186
rect 18574 3152 18630 3186
rect 18664 3152 18720 3186
rect 18754 3152 18884 3186
rect 12444 3119 18884 3152
rect 12444 3102 12684 3119
rect 12444 3068 12477 3102
rect 12511 3068 12684 3102
rect 12444 3055 12684 3068
rect 13484 3102 13984 3119
rect 13484 3068 13664 3102
rect 13698 3068 13765 3102
rect 13799 3068 13984 3102
rect 13484 3055 13984 3068
rect 14784 3102 15184 3119
rect 14784 3068 14952 3102
rect 14986 3068 15053 3102
rect 15087 3068 15184 3102
rect 14784 3055 15184 3068
rect 16084 3102 16484 3119
rect 16084 3068 16240 3102
rect 16274 3068 16341 3102
rect 16375 3068 16484 3102
rect 16084 3055 16484 3068
rect 17384 3102 17784 3119
rect 17384 3068 17528 3102
rect 17562 3068 17629 3102
rect 17663 3068 17784 3102
rect 17384 3055 17784 3068
rect 18684 3102 18884 3119
rect 18684 3068 18816 3102
rect 18850 3068 18884 3102
rect 18684 3055 18884 3068
rect 12444 3036 18884 3055
rect 12444 3012 12718 3036
rect 12444 2978 12477 3012
rect 12511 3002 12718 3012
rect 12752 3002 12808 3036
rect 12842 3002 12898 3036
rect 12932 3002 12988 3036
rect 13022 3002 13078 3036
rect 13112 3002 13168 3036
rect 13202 3002 13258 3036
rect 13292 3002 13348 3036
rect 13382 3002 13438 3036
rect 13472 3012 14006 3036
rect 13472 3002 13664 3012
rect 12511 2983 13664 3002
rect 12511 2978 12684 2983
rect 12444 2942 12684 2978
rect 12444 2922 12626 2942
rect 12444 2888 12477 2922
rect 12511 2908 12626 2922
rect 12660 2908 12684 2942
rect 13484 2978 13664 2983
rect 13698 2978 13765 3012
rect 13799 3002 14006 3012
rect 14040 3002 14096 3036
rect 14130 3002 14186 3036
rect 14220 3002 14276 3036
rect 14310 3002 14366 3036
rect 14400 3002 14456 3036
rect 14490 3002 14546 3036
rect 14580 3002 14636 3036
rect 14670 3002 14726 3036
rect 14760 3012 15294 3036
rect 14760 3002 14952 3012
rect 13799 2983 14952 3002
rect 13799 2978 13984 2983
rect 13484 2942 13984 2978
rect 13484 2923 13914 2942
rect 12511 2888 12684 2908
rect 12444 2852 12684 2888
rect 12444 2832 12626 2852
rect 12444 2798 12477 2832
rect 12511 2818 12626 2832
rect 12660 2818 12684 2852
rect 12511 2798 12684 2818
rect 12444 2762 12684 2798
rect 12444 2742 12626 2762
rect 12444 2708 12477 2742
rect 12511 2728 12626 2742
rect 12660 2728 12684 2762
rect 12511 2708 12684 2728
rect 12444 2672 12684 2708
rect 12444 2652 12626 2672
rect 12444 2618 12477 2652
rect 12511 2638 12626 2652
rect 12660 2638 12684 2672
rect 12511 2618 12684 2638
rect 12444 2582 12684 2618
rect 12444 2562 12626 2582
rect 12444 2528 12477 2562
rect 12511 2548 12626 2562
rect 12660 2548 12684 2582
rect 12511 2528 12684 2548
rect 12444 2492 12684 2528
rect 12444 2472 12626 2492
rect 12444 2438 12477 2472
rect 12511 2458 12626 2472
rect 12660 2458 12684 2492
rect 12511 2438 12684 2458
rect 12444 2402 12684 2438
rect 12444 2382 12626 2402
rect 12444 2348 12477 2382
rect 12511 2368 12626 2382
rect 12660 2368 12684 2402
rect 12511 2348 12684 2368
rect 12444 2312 12684 2348
rect 12444 2292 12626 2312
rect 12444 2258 12477 2292
rect 12511 2278 12626 2292
rect 12660 2278 12684 2312
rect 12511 2258 12684 2278
rect 12444 2222 12684 2258
rect 12741 2860 13435 2921
rect 12741 2826 12800 2860
rect 12834 2848 12890 2860
rect 12862 2826 12890 2848
rect 12924 2848 12980 2860
rect 12924 2826 12928 2848
rect 12741 2814 12828 2826
rect 12862 2814 12928 2826
rect 12962 2826 12980 2848
rect 13014 2848 13070 2860
rect 13014 2826 13028 2848
rect 12962 2814 13028 2826
rect 13062 2826 13070 2848
rect 13104 2848 13160 2860
rect 13194 2848 13250 2860
rect 13284 2848 13340 2860
rect 13104 2826 13128 2848
rect 13194 2826 13228 2848
rect 13284 2826 13328 2848
rect 13374 2826 13435 2860
rect 13062 2814 13128 2826
rect 13162 2814 13228 2826
rect 13262 2814 13328 2826
rect 13362 2814 13435 2826
rect 12741 2770 13435 2814
rect 12741 2736 12800 2770
rect 12834 2748 12890 2770
rect 12862 2736 12890 2748
rect 12924 2748 12980 2770
rect 12924 2736 12928 2748
rect 12741 2714 12828 2736
rect 12862 2714 12928 2736
rect 12962 2736 12980 2748
rect 13014 2748 13070 2770
rect 13014 2736 13028 2748
rect 12962 2714 13028 2736
rect 13062 2736 13070 2748
rect 13104 2748 13160 2770
rect 13194 2748 13250 2770
rect 13284 2748 13340 2770
rect 13104 2736 13128 2748
rect 13194 2736 13228 2748
rect 13284 2736 13328 2748
rect 13374 2736 13435 2770
rect 13062 2714 13128 2736
rect 13162 2714 13228 2736
rect 13262 2714 13328 2736
rect 13362 2714 13435 2736
rect 12741 2680 13435 2714
rect 12741 2646 12800 2680
rect 12834 2648 12890 2680
rect 12862 2646 12890 2648
rect 12924 2648 12980 2680
rect 12924 2646 12928 2648
rect 12741 2614 12828 2646
rect 12862 2614 12928 2646
rect 12962 2646 12980 2648
rect 13014 2648 13070 2680
rect 13014 2646 13028 2648
rect 12962 2614 13028 2646
rect 13062 2646 13070 2648
rect 13104 2648 13160 2680
rect 13194 2648 13250 2680
rect 13284 2648 13340 2680
rect 13104 2646 13128 2648
rect 13194 2646 13228 2648
rect 13284 2646 13328 2648
rect 13374 2646 13435 2680
rect 13062 2614 13128 2646
rect 13162 2614 13228 2646
rect 13262 2614 13328 2646
rect 13362 2614 13435 2646
rect 12741 2590 13435 2614
rect 12741 2556 12800 2590
rect 12834 2556 12890 2590
rect 12924 2556 12980 2590
rect 13014 2556 13070 2590
rect 13104 2556 13160 2590
rect 13194 2556 13250 2590
rect 13284 2556 13340 2590
rect 13374 2556 13435 2590
rect 12741 2548 13435 2556
rect 12741 2514 12828 2548
rect 12862 2514 12928 2548
rect 12962 2514 13028 2548
rect 13062 2514 13128 2548
rect 13162 2514 13228 2548
rect 13262 2514 13328 2548
rect 13362 2514 13435 2548
rect 12741 2500 13435 2514
rect 12741 2466 12800 2500
rect 12834 2466 12890 2500
rect 12924 2466 12980 2500
rect 13014 2466 13070 2500
rect 13104 2466 13160 2500
rect 13194 2466 13250 2500
rect 13284 2466 13340 2500
rect 13374 2466 13435 2500
rect 12741 2448 13435 2466
rect 12741 2414 12828 2448
rect 12862 2414 12928 2448
rect 12962 2414 13028 2448
rect 13062 2414 13128 2448
rect 13162 2414 13228 2448
rect 13262 2414 13328 2448
rect 13362 2414 13435 2448
rect 12741 2410 13435 2414
rect 12741 2376 12800 2410
rect 12834 2376 12890 2410
rect 12924 2376 12980 2410
rect 13014 2376 13070 2410
rect 13104 2376 13160 2410
rect 13194 2376 13250 2410
rect 13284 2376 13340 2410
rect 13374 2376 13435 2410
rect 12741 2348 13435 2376
rect 12741 2320 12828 2348
rect 12862 2320 12928 2348
rect 12741 2286 12800 2320
rect 12862 2314 12890 2320
rect 12834 2286 12890 2314
rect 12924 2314 12928 2320
rect 12962 2320 13028 2348
rect 12962 2314 12980 2320
rect 12924 2286 12980 2314
rect 13014 2314 13028 2320
rect 13062 2320 13128 2348
rect 13162 2320 13228 2348
rect 13262 2320 13328 2348
rect 13362 2320 13435 2348
rect 13062 2314 13070 2320
rect 13014 2286 13070 2314
rect 13104 2314 13128 2320
rect 13194 2314 13228 2320
rect 13284 2314 13328 2320
rect 13104 2286 13160 2314
rect 13194 2286 13250 2314
rect 13284 2286 13340 2314
rect 13374 2286 13435 2320
rect 12741 2227 13435 2286
rect 13484 2889 13516 2923
rect 13550 2922 13914 2923
rect 13550 2889 13664 2922
rect 13484 2888 13664 2889
rect 13698 2888 13765 2922
rect 13799 2908 13914 2922
rect 13948 2908 13984 2942
rect 14784 2978 14952 2983
rect 14986 2978 15053 3012
rect 15087 3002 15294 3012
rect 15328 3002 15384 3036
rect 15418 3002 15474 3036
rect 15508 3002 15564 3036
rect 15598 3002 15654 3036
rect 15688 3002 15744 3036
rect 15778 3002 15834 3036
rect 15868 3002 15924 3036
rect 15958 3002 16014 3036
rect 16048 3012 16582 3036
rect 16048 3002 16240 3012
rect 15087 2983 16240 3002
rect 15087 2978 15255 2983
rect 14784 2942 15255 2978
rect 14784 2923 15202 2942
rect 13799 2888 13984 2908
rect 13484 2852 13984 2888
rect 13484 2833 13914 2852
rect 13484 2799 13516 2833
rect 13550 2832 13914 2833
rect 13550 2799 13664 2832
rect 13484 2798 13664 2799
rect 13698 2798 13765 2832
rect 13799 2818 13914 2832
rect 13948 2818 13984 2852
rect 13799 2798 13984 2818
rect 13484 2762 13984 2798
rect 13484 2743 13914 2762
rect 13484 2709 13516 2743
rect 13550 2742 13914 2743
rect 13550 2709 13664 2742
rect 13484 2708 13664 2709
rect 13698 2708 13765 2742
rect 13799 2728 13914 2742
rect 13948 2728 13984 2762
rect 13799 2708 13984 2728
rect 13484 2672 13984 2708
rect 13484 2653 13914 2672
rect 13484 2619 13516 2653
rect 13550 2652 13914 2653
rect 13550 2619 13664 2652
rect 13484 2618 13664 2619
rect 13698 2618 13765 2652
rect 13799 2638 13914 2652
rect 13948 2638 13984 2672
rect 13799 2618 13984 2638
rect 13484 2582 13984 2618
rect 13484 2563 13914 2582
rect 13484 2529 13516 2563
rect 13550 2562 13914 2563
rect 13550 2529 13664 2562
rect 13484 2528 13664 2529
rect 13698 2528 13765 2562
rect 13799 2548 13914 2562
rect 13948 2548 13984 2582
rect 13799 2528 13984 2548
rect 13484 2492 13984 2528
rect 13484 2473 13914 2492
rect 13484 2439 13516 2473
rect 13550 2472 13914 2473
rect 13550 2439 13664 2472
rect 13484 2438 13664 2439
rect 13698 2438 13765 2472
rect 13799 2458 13914 2472
rect 13948 2458 13984 2492
rect 13799 2438 13984 2458
rect 13484 2402 13984 2438
rect 13484 2383 13914 2402
rect 13484 2349 13516 2383
rect 13550 2382 13914 2383
rect 13550 2349 13664 2382
rect 13484 2348 13664 2349
rect 13698 2348 13765 2382
rect 13799 2368 13914 2382
rect 13948 2368 13984 2402
rect 13799 2348 13984 2368
rect 13484 2312 13984 2348
rect 13484 2293 13914 2312
rect 13484 2259 13516 2293
rect 13550 2292 13914 2293
rect 13550 2259 13664 2292
rect 13484 2258 13664 2259
rect 13698 2258 13765 2292
rect 13799 2278 13914 2292
rect 13948 2278 13984 2312
rect 13799 2258 13984 2278
rect 12444 2202 12626 2222
rect 12444 2168 12477 2202
rect 12511 2188 12626 2202
rect 12660 2188 12684 2222
rect 12511 2168 12684 2188
rect 12444 2165 12684 2168
rect 13484 2222 13984 2258
rect 14029 2860 14723 2921
rect 14029 2826 14088 2860
rect 14122 2848 14178 2860
rect 14150 2826 14178 2848
rect 14212 2848 14268 2860
rect 14212 2826 14216 2848
rect 14029 2814 14116 2826
rect 14150 2814 14216 2826
rect 14250 2826 14268 2848
rect 14302 2848 14358 2860
rect 14302 2826 14316 2848
rect 14250 2814 14316 2826
rect 14350 2826 14358 2848
rect 14392 2848 14448 2860
rect 14482 2848 14538 2860
rect 14572 2848 14628 2860
rect 14392 2826 14416 2848
rect 14482 2826 14516 2848
rect 14572 2826 14616 2848
rect 14662 2826 14723 2860
rect 14350 2814 14416 2826
rect 14450 2814 14516 2826
rect 14550 2814 14616 2826
rect 14650 2814 14723 2826
rect 14029 2770 14723 2814
rect 14029 2736 14088 2770
rect 14122 2748 14178 2770
rect 14150 2736 14178 2748
rect 14212 2748 14268 2770
rect 14212 2736 14216 2748
rect 14029 2714 14116 2736
rect 14150 2714 14216 2736
rect 14250 2736 14268 2748
rect 14302 2748 14358 2770
rect 14302 2736 14316 2748
rect 14250 2714 14316 2736
rect 14350 2736 14358 2748
rect 14392 2748 14448 2770
rect 14482 2748 14538 2770
rect 14572 2748 14628 2770
rect 14392 2736 14416 2748
rect 14482 2736 14516 2748
rect 14572 2736 14616 2748
rect 14662 2736 14723 2770
rect 14350 2714 14416 2736
rect 14450 2714 14516 2736
rect 14550 2714 14616 2736
rect 14650 2714 14723 2736
rect 14029 2680 14723 2714
rect 14029 2646 14088 2680
rect 14122 2648 14178 2680
rect 14150 2646 14178 2648
rect 14212 2648 14268 2680
rect 14212 2646 14216 2648
rect 14029 2614 14116 2646
rect 14150 2614 14216 2646
rect 14250 2646 14268 2648
rect 14302 2648 14358 2680
rect 14302 2646 14316 2648
rect 14250 2614 14316 2646
rect 14350 2646 14358 2648
rect 14392 2648 14448 2680
rect 14482 2648 14538 2680
rect 14572 2648 14628 2680
rect 14392 2646 14416 2648
rect 14482 2646 14516 2648
rect 14572 2646 14616 2648
rect 14662 2646 14723 2680
rect 14350 2614 14416 2646
rect 14450 2614 14516 2646
rect 14550 2614 14616 2646
rect 14650 2614 14723 2646
rect 14029 2590 14723 2614
rect 14029 2556 14088 2590
rect 14122 2556 14178 2590
rect 14212 2556 14268 2590
rect 14302 2556 14358 2590
rect 14392 2556 14448 2590
rect 14482 2556 14538 2590
rect 14572 2556 14628 2590
rect 14662 2556 14723 2590
rect 14029 2548 14723 2556
rect 14029 2514 14116 2548
rect 14150 2514 14216 2548
rect 14250 2514 14316 2548
rect 14350 2514 14416 2548
rect 14450 2514 14516 2548
rect 14550 2514 14616 2548
rect 14650 2514 14723 2548
rect 14029 2500 14723 2514
rect 14029 2466 14088 2500
rect 14122 2466 14178 2500
rect 14212 2466 14268 2500
rect 14302 2466 14358 2500
rect 14392 2466 14448 2500
rect 14482 2466 14538 2500
rect 14572 2466 14628 2500
rect 14662 2466 14723 2500
rect 14029 2448 14723 2466
rect 14029 2414 14116 2448
rect 14150 2414 14216 2448
rect 14250 2414 14316 2448
rect 14350 2414 14416 2448
rect 14450 2414 14516 2448
rect 14550 2414 14616 2448
rect 14650 2414 14723 2448
rect 14029 2410 14723 2414
rect 14029 2376 14088 2410
rect 14122 2376 14178 2410
rect 14212 2376 14268 2410
rect 14302 2376 14358 2410
rect 14392 2376 14448 2410
rect 14482 2376 14538 2410
rect 14572 2376 14628 2410
rect 14662 2376 14723 2410
rect 14029 2348 14723 2376
rect 14029 2320 14116 2348
rect 14150 2320 14216 2348
rect 14029 2286 14088 2320
rect 14150 2314 14178 2320
rect 14122 2286 14178 2314
rect 14212 2314 14216 2320
rect 14250 2320 14316 2348
rect 14250 2314 14268 2320
rect 14212 2286 14268 2314
rect 14302 2314 14316 2320
rect 14350 2320 14416 2348
rect 14450 2320 14516 2348
rect 14550 2320 14616 2348
rect 14650 2320 14723 2348
rect 14350 2314 14358 2320
rect 14302 2286 14358 2314
rect 14392 2314 14416 2320
rect 14482 2314 14516 2320
rect 14572 2314 14616 2320
rect 14392 2286 14448 2314
rect 14482 2286 14538 2314
rect 14572 2286 14628 2314
rect 14662 2286 14723 2320
rect 14029 2227 14723 2286
rect 14784 2889 14804 2923
rect 14838 2922 15202 2923
rect 14838 2889 14952 2922
rect 14784 2888 14952 2889
rect 14986 2888 15053 2922
rect 15087 2908 15202 2922
rect 15236 2908 15255 2942
rect 16073 2978 16240 2983
rect 16274 2978 16341 3012
rect 16375 3002 16582 3012
rect 16616 3002 16672 3036
rect 16706 3002 16762 3036
rect 16796 3002 16852 3036
rect 16886 3002 16942 3036
rect 16976 3002 17032 3036
rect 17066 3002 17122 3036
rect 17156 3002 17212 3036
rect 17246 3002 17302 3036
rect 17336 3012 17870 3036
rect 17336 3002 17528 3012
rect 16375 2983 17528 3002
rect 16375 2978 16543 2983
rect 16073 2942 16543 2978
rect 16073 2923 16490 2942
rect 15087 2888 15255 2908
rect 14784 2852 15255 2888
rect 14784 2833 15202 2852
rect 14784 2799 14804 2833
rect 14838 2832 15202 2833
rect 14838 2799 14952 2832
rect 14784 2798 14952 2799
rect 14986 2798 15053 2832
rect 15087 2818 15202 2832
rect 15236 2818 15255 2852
rect 15087 2798 15255 2818
rect 14784 2762 15255 2798
rect 14784 2743 15202 2762
rect 14784 2709 14804 2743
rect 14838 2742 15202 2743
rect 14838 2709 14952 2742
rect 14784 2708 14952 2709
rect 14986 2708 15053 2742
rect 15087 2728 15202 2742
rect 15236 2728 15255 2762
rect 15087 2708 15255 2728
rect 14784 2672 15255 2708
rect 14784 2653 15202 2672
rect 14784 2619 14804 2653
rect 14838 2652 15202 2653
rect 14838 2619 14952 2652
rect 14784 2618 14952 2619
rect 14986 2618 15053 2652
rect 15087 2638 15202 2652
rect 15236 2638 15255 2672
rect 15087 2618 15255 2638
rect 14784 2582 15255 2618
rect 14784 2563 15202 2582
rect 14784 2529 14804 2563
rect 14838 2562 15202 2563
rect 14838 2529 14952 2562
rect 14784 2528 14952 2529
rect 14986 2528 15053 2562
rect 15087 2548 15202 2562
rect 15236 2548 15255 2582
rect 15087 2528 15255 2548
rect 14784 2492 15255 2528
rect 14784 2473 15202 2492
rect 14784 2439 14804 2473
rect 14838 2472 15202 2473
rect 14838 2439 14952 2472
rect 14784 2438 14952 2439
rect 14986 2438 15053 2472
rect 15087 2458 15202 2472
rect 15236 2458 15255 2492
rect 15087 2438 15255 2458
rect 14784 2402 15255 2438
rect 14784 2383 15202 2402
rect 14784 2349 14804 2383
rect 14838 2382 15202 2383
rect 14838 2349 14952 2382
rect 14784 2348 14952 2349
rect 14986 2348 15053 2382
rect 15087 2368 15202 2382
rect 15236 2368 15255 2402
rect 15087 2348 15255 2368
rect 14784 2312 15255 2348
rect 14784 2293 15202 2312
rect 14784 2259 14804 2293
rect 14838 2292 15202 2293
rect 14838 2259 14952 2292
rect 14784 2258 14952 2259
rect 14986 2258 15053 2292
rect 15087 2278 15202 2292
rect 15236 2278 15255 2312
rect 15087 2258 15255 2278
rect 13484 2203 13914 2222
rect 13484 2169 13516 2203
rect 13550 2202 13914 2203
rect 13550 2169 13664 2202
rect 13484 2168 13664 2169
rect 13698 2168 13765 2202
rect 13799 2188 13914 2202
rect 13948 2188 13984 2222
rect 13799 2168 13984 2188
rect 13484 2165 13984 2168
rect 14784 2222 15255 2258
rect 15317 2860 16011 2921
rect 15317 2826 15376 2860
rect 15410 2848 15466 2860
rect 15438 2826 15466 2848
rect 15500 2848 15556 2860
rect 15500 2826 15504 2848
rect 15317 2814 15404 2826
rect 15438 2814 15504 2826
rect 15538 2826 15556 2848
rect 15590 2848 15646 2860
rect 15590 2826 15604 2848
rect 15538 2814 15604 2826
rect 15638 2826 15646 2848
rect 15680 2848 15736 2860
rect 15770 2848 15826 2860
rect 15860 2848 15916 2860
rect 15680 2826 15704 2848
rect 15770 2826 15804 2848
rect 15860 2826 15904 2848
rect 15950 2826 16011 2860
rect 15638 2814 15704 2826
rect 15738 2814 15804 2826
rect 15838 2814 15904 2826
rect 15938 2814 16011 2826
rect 15317 2770 16011 2814
rect 15317 2736 15376 2770
rect 15410 2748 15466 2770
rect 15438 2736 15466 2748
rect 15500 2748 15556 2770
rect 15500 2736 15504 2748
rect 15317 2714 15404 2736
rect 15438 2714 15504 2736
rect 15538 2736 15556 2748
rect 15590 2748 15646 2770
rect 15590 2736 15604 2748
rect 15538 2714 15604 2736
rect 15638 2736 15646 2748
rect 15680 2748 15736 2770
rect 15770 2748 15826 2770
rect 15860 2748 15916 2770
rect 15680 2736 15704 2748
rect 15770 2736 15804 2748
rect 15860 2736 15904 2748
rect 15950 2736 16011 2770
rect 15638 2714 15704 2736
rect 15738 2714 15804 2736
rect 15838 2714 15904 2736
rect 15938 2714 16011 2736
rect 15317 2680 16011 2714
rect 15317 2646 15376 2680
rect 15410 2648 15466 2680
rect 15438 2646 15466 2648
rect 15500 2648 15556 2680
rect 15500 2646 15504 2648
rect 15317 2614 15404 2646
rect 15438 2614 15504 2646
rect 15538 2646 15556 2648
rect 15590 2648 15646 2680
rect 15590 2646 15604 2648
rect 15538 2614 15604 2646
rect 15638 2646 15646 2648
rect 15680 2648 15736 2680
rect 15770 2648 15826 2680
rect 15860 2648 15916 2680
rect 15680 2646 15704 2648
rect 15770 2646 15804 2648
rect 15860 2646 15904 2648
rect 15950 2646 16011 2680
rect 15638 2614 15704 2646
rect 15738 2614 15804 2646
rect 15838 2614 15904 2646
rect 15938 2614 16011 2646
rect 15317 2590 16011 2614
rect 15317 2556 15376 2590
rect 15410 2556 15466 2590
rect 15500 2556 15556 2590
rect 15590 2556 15646 2590
rect 15680 2556 15736 2590
rect 15770 2556 15826 2590
rect 15860 2556 15916 2590
rect 15950 2556 16011 2590
rect 15317 2548 16011 2556
rect 15317 2514 15404 2548
rect 15438 2514 15504 2548
rect 15538 2514 15604 2548
rect 15638 2514 15704 2548
rect 15738 2514 15804 2548
rect 15838 2514 15904 2548
rect 15938 2514 16011 2548
rect 15317 2500 16011 2514
rect 15317 2466 15376 2500
rect 15410 2466 15466 2500
rect 15500 2466 15556 2500
rect 15590 2466 15646 2500
rect 15680 2466 15736 2500
rect 15770 2466 15826 2500
rect 15860 2466 15916 2500
rect 15950 2466 16011 2500
rect 15317 2448 16011 2466
rect 15317 2414 15404 2448
rect 15438 2414 15504 2448
rect 15538 2414 15604 2448
rect 15638 2414 15704 2448
rect 15738 2414 15804 2448
rect 15838 2414 15904 2448
rect 15938 2414 16011 2448
rect 15317 2410 16011 2414
rect 15317 2376 15376 2410
rect 15410 2376 15466 2410
rect 15500 2376 15556 2410
rect 15590 2376 15646 2410
rect 15680 2376 15736 2410
rect 15770 2376 15826 2410
rect 15860 2376 15916 2410
rect 15950 2376 16011 2410
rect 15317 2348 16011 2376
rect 15317 2320 15404 2348
rect 15438 2320 15504 2348
rect 15317 2286 15376 2320
rect 15438 2314 15466 2320
rect 15410 2286 15466 2314
rect 15500 2314 15504 2320
rect 15538 2320 15604 2348
rect 15538 2314 15556 2320
rect 15500 2286 15556 2314
rect 15590 2314 15604 2320
rect 15638 2320 15704 2348
rect 15738 2320 15804 2348
rect 15838 2320 15904 2348
rect 15938 2320 16011 2348
rect 15638 2314 15646 2320
rect 15590 2286 15646 2314
rect 15680 2314 15704 2320
rect 15770 2314 15804 2320
rect 15860 2314 15904 2320
rect 15680 2286 15736 2314
rect 15770 2286 15826 2314
rect 15860 2286 15916 2314
rect 15950 2286 16011 2320
rect 15317 2227 16011 2286
rect 16073 2889 16092 2923
rect 16126 2922 16490 2923
rect 16126 2889 16240 2922
rect 16073 2888 16240 2889
rect 16274 2888 16341 2922
rect 16375 2908 16490 2922
rect 16524 2908 16543 2942
rect 17361 2978 17528 2983
rect 17562 2978 17629 3012
rect 17663 3002 17870 3012
rect 17904 3002 17960 3036
rect 17994 3002 18050 3036
rect 18084 3002 18140 3036
rect 18174 3002 18230 3036
rect 18264 3002 18320 3036
rect 18354 3002 18410 3036
rect 18444 3002 18500 3036
rect 18534 3002 18590 3036
rect 18624 3012 18884 3036
rect 18624 3002 18816 3012
rect 17663 2983 18816 3002
rect 17663 2978 17831 2983
rect 17361 2942 17831 2978
rect 17361 2923 17778 2942
rect 16375 2888 16543 2908
rect 16073 2852 16543 2888
rect 16073 2833 16490 2852
rect 16073 2799 16092 2833
rect 16126 2832 16490 2833
rect 16126 2799 16240 2832
rect 16073 2798 16240 2799
rect 16274 2798 16341 2832
rect 16375 2818 16490 2832
rect 16524 2818 16543 2852
rect 16375 2798 16543 2818
rect 16073 2762 16543 2798
rect 16073 2743 16490 2762
rect 16073 2709 16092 2743
rect 16126 2742 16490 2743
rect 16126 2709 16240 2742
rect 16073 2708 16240 2709
rect 16274 2708 16341 2742
rect 16375 2728 16490 2742
rect 16524 2728 16543 2762
rect 16375 2708 16543 2728
rect 16073 2672 16543 2708
rect 16073 2653 16490 2672
rect 16073 2619 16092 2653
rect 16126 2652 16490 2653
rect 16126 2619 16240 2652
rect 16073 2618 16240 2619
rect 16274 2618 16341 2652
rect 16375 2638 16490 2652
rect 16524 2638 16543 2672
rect 16375 2618 16543 2638
rect 16073 2582 16543 2618
rect 16073 2563 16490 2582
rect 16073 2529 16092 2563
rect 16126 2562 16490 2563
rect 16126 2529 16240 2562
rect 16073 2528 16240 2529
rect 16274 2528 16341 2562
rect 16375 2548 16490 2562
rect 16524 2548 16543 2582
rect 16375 2528 16543 2548
rect 16073 2492 16543 2528
rect 16073 2473 16490 2492
rect 16073 2439 16092 2473
rect 16126 2472 16490 2473
rect 16126 2439 16240 2472
rect 16073 2438 16240 2439
rect 16274 2438 16341 2472
rect 16375 2458 16490 2472
rect 16524 2458 16543 2492
rect 16375 2438 16543 2458
rect 16073 2402 16543 2438
rect 16073 2383 16490 2402
rect 16073 2349 16092 2383
rect 16126 2382 16490 2383
rect 16126 2349 16240 2382
rect 16073 2348 16240 2349
rect 16274 2348 16341 2382
rect 16375 2368 16490 2382
rect 16524 2368 16543 2402
rect 16375 2348 16543 2368
rect 16073 2312 16543 2348
rect 16073 2293 16490 2312
rect 16073 2259 16092 2293
rect 16126 2292 16490 2293
rect 16126 2259 16240 2292
rect 16073 2258 16240 2259
rect 16274 2258 16341 2292
rect 16375 2278 16490 2292
rect 16524 2278 16543 2312
rect 16375 2258 16543 2278
rect 14784 2203 15202 2222
rect 14784 2169 14804 2203
rect 14838 2202 15202 2203
rect 14838 2169 14952 2202
rect 14784 2168 14952 2169
rect 14986 2168 15053 2202
rect 15087 2188 15202 2202
rect 15236 2188 15255 2222
rect 15087 2168 15255 2188
rect 14784 2165 15255 2168
rect 16073 2222 16543 2258
rect 16605 2860 17299 2921
rect 16605 2826 16664 2860
rect 16698 2848 16754 2860
rect 16726 2826 16754 2848
rect 16788 2848 16844 2860
rect 16788 2826 16792 2848
rect 16605 2814 16692 2826
rect 16726 2814 16792 2826
rect 16826 2826 16844 2848
rect 16878 2848 16934 2860
rect 16878 2826 16892 2848
rect 16826 2814 16892 2826
rect 16926 2826 16934 2848
rect 16968 2848 17024 2860
rect 17058 2848 17114 2860
rect 17148 2848 17204 2860
rect 16968 2826 16992 2848
rect 17058 2826 17092 2848
rect 17148 2826 17192 2848
rect 17238 2826 17299 2860
rect 16926 2814 16992 2826
rect 17026 2814 17092 2826
rect 17126 2814 17192 2826
rect 17226 2814 17299 2826
rect 16605 2770 17299 2814
rect 16605 2736 16664 2770
rect 16698 2748 16754 2770
rect 16726 2736 16754 2748
rect 16788 2748 16844 2770
rect 16788 2736 16792 2748
rect 16605 2714 16692 2736
rect 16726 2714 16792 2736
rect 16826 2736 16844 2748
rect 16878 2748 16934 2770
rect 16878 2736 16892 2748
rect 16826 2714 16892 2736
rect 16926 2736 16934 2748
rect 16968 2748 17024 2770
rect 17058 2748 17114 2770
rect 17148 2748 17204 2770
rect 16968 2736 16992 2748
rect 17058 2736 17092 2748
rect 17148 2736 17192 2748
rect 17238 2736 17299 2770
rect 16926 2714 16992 2736
rect 17026 2714 17092 2736
rect 17126 2714 17192 2736
rect 17226 2714 17299 2736
rect 16605 2680 17299 2714
rect 16605 2646 16664 2680
rect 16698 2648 16754 2680
rect 16726 2646 16754 2648
rect 16788 2648 16844 2680
rect 16788 2646 16792 2648
rect 16605 2614 16692 2646
rect 16726 2614 16792 2646
rect 16826 2646 16844 2648
rect 16878 2648 16934 2680
rect 16878 2646 16892 2648
rect 16826 2614 16892 2646
rect 16926 2646 16934 2648
rect 16968 2648 17024 2680
rect 17058 2648 17114 2680
rect 17148 2648 17204 2680
rect 16968 2646 16992 2648
rect 17058 2646 17092 2648
rect 17148 2646 17192 2648
rect 17238 2646 17299 2680
rect 16926 2614 16992 2646
rect 17026 2614 17092 2646
rect 17126 2614 17192 2646
rect 17226 2614 17299 2646
rect 16605 2590 17299 2614
rect 16605 2556 16664 2590
rect 16698 2556 16754 2590
rect 16788 2556 16844 2590
rect 16878 2556 16934 2590
rect 16968 2556 17024 2590
rect 17058 2556 17114 2590
rect 17148 2556 17204 2590
rect 17238 2556 17299 2590
rect 16605 2548 17299 2556
rect 16605 2514 16692 2548
rect 16726 2514 16792 2548
rect 16826 2514 16892 2548
rect 16926 2514 16992 2548
rect 17026 2514 17092 2548
rect 17126 2514 17192 2548
rect 17226 2514 17299 2548
rect 16605 2500 17299 2514
rect 16605 2466 16664 2500
rect 16698 2466 16754 2500
rect 16788 2466 16844 2500
rect 16878 2466 16934 2500
rect 16968 2466 17024 2500
rect 17058 2466 17114 2500
rect 17148 2466 17204 2500
rect 17238 2466 17299 2500
rect 16605 2448 17299 2466
rect 16605 2414 16692 2448
rect 16726 2414 16792 2448
rect 16826 2414 16892 2448
rect 16926 2414 16992 2448
rect 17026 2414 17092 2448
rect 17126 2414 17192 2448
rect 17226 2414 17299 2448
rect 16605 2410 17299 2414
rect 16605 2376 16664 2410
rect 16698 2376 16754 2410
rect 16788 2376 16844 2410
rect 16878 2376 16934 2410
rect 16968 2376 17024 2410
rect 17058 2376 17114 2410
rect 17148 2376 17204 2410
rect 17238 2376 17299 2410
rect 16605 2348 17299 2376
rect 16605 2320 16692 2348
rect 16726 2320 16792 2348
rect 16605 2286 16664 2320
rect 16726 2314 16754 2320
rect 16698 2286 16754 2314
rect 16788 2314 16792 2320
rect 16826 2320 16892 2348
rect 16826 2314 16844 2320
rect 16788 2286 16844 2314
rect 16878 2314 16892 2320
rect 16926 2320 16992 2348
rect 17026 2320 17092 2348
rect 17126 2320 17192 2348
rect 17226 2320 17299 2348
rect 16926 2314 16934 2320
rect 16878 2286 16934 2314
rect 16968 2314 16992 2320
rect 17058 2314 17092 2320
rect 17148 2314 17192 2320
rect 16968 2286 17024 2314
rect 17058 2286 17114 2314
rect 17148 2286 17204 2314
rect 17238 2286 17299 2320
rect 16605 2227 17299 2286
rect 17361 2889 17380 2923
rect 17414 2922 17778 2923
rect 17414 2889 17528 2922
rect 17361 2888 17528 2889
rect 17562 2888 17629 2922
rect 17663 2908 17778 2922
rect 17812 2908 17831 2942
rect 18649 2978 18816 2983
rect 18850 2978 18884 3012
rect 18649 2923 18884 2978
rect 17663 2888 17831 2908
rect 17361 2852 17831 2888
rect 17361 2833 17778 2852
rect 17361 2799 17380 2833
rect 17414 2832 17778 2833
rect 17414 2799 17528 2832
rect 17361 2798 17528 2799
rect 17562 2798 17629 2832
rect 17663 2818 17778 2832
rect 17812 2818 17831 2852
rect 17663 2798 17831 2818
rect 17361 2762 17831 2798
rect 17361 2743 17778 2762
rect 17361 2709 17380 2743
rect 17414 2742 17778 2743
rect 17414 2709 17528 2742
rect 17361 2708 17528 2709
rect 17562 2708 17629 2742
rect 17663 2728 17778 2742
rect 17812 2728 17831 2762
rect 17663 2708 17831 2728
rect 17361 2672 17831 2708
rect 17361 2653 17778 2672
rect 17361 2619 17380 2653
rect 17414 2652 17778 2653
rect 17414 2619 17528 2652
rect 17361 2618 17528 2619
rect 17562 2618 17629 2652
rect 17663 2638 17778 2652
rect 17812 2638 17831 2672
rect 17663 2618 17831 2638
rect 17361 2582 17831 2618
rect 17361 2563 17778 2582
rect 17361 2529 17380 2563
rect 17414 2562 17778 2563
rect 17414 2529 17528 2562
rect 17361 2528 17528 2529
rect 17562 2528 17629 2562
rect 17663 2548 17778 2562
rect 17812 2548 17831 2582
rect 17663 2528 17831 2548
rect 17361 2492 17831 2528
rect 17361 2473 17778 2492
rect 17361 2439 17380 2473
rect 17414 2472 17778 2473
rect 17414 2439 17528 2472
rect 17361 2438 17528 2439
rect 17562 2438 17629 2472
rect 17663 2458 17778 2472
rect 17812 2458 17831 2492
rect 17663 2438 17831 2458
rect 17361 2402 17831 2438
rect 17361 2383 17778 2402
rect 17361 2349 17380 2383
rect 17414 2382 17778 2383
rect 17414 2349 17528 2382
rect 17361 2348 17528 2349
rect 17562 2348 17629 2382
rect 17663 2368 17778 2382
rect 17812 2368 17831 2402
rect 17663 2348 17831 2368
rect 17361 2312 17831 2348
rect 17361 2293 17778 2312
rect 17361 2259 17380 2293
rect 17414 2292 17778 2293
rect 17414 2259 17528 2292
rect 17361 2258 17528 2259
rect 17562 2258 17629 2292
rect 17663 2278 17778 2292
rect 17812 2278 17831 2312
rect 17663 2258 17831 2278
rect 16073 2203 16490 2222
rect 16073 2169 16092 2203
rect 16126 2202 16490 2203
rect 16126 2169 16240 2202
rect 16073 2168 16240 2169
rect 16274 2168 16341 2202
rect 16375 2188 16490 2202
rect 16524 2188 16543 2222
rect 16375 2168 16543 2188
rect 16073 2165 16543 2168
rect 17361 2222 17831 2258
rect 17893 2860 18587 2921
rect 17893 2826 17952 2860
rect 17986 2848 18042 2860
rect 18014 2826 18042 2848
rect 18076 2848 18132 2860
rect 18076 2826 18080 2848
rect 17893 2814 17980 2826
rect 18014 2814 18080 2826
rect 18114 2826 18132 2848
rect 18166 2848 18222 2860
rect 18166 2826 18180 2848
rect 18114 2814 18180 2826
rect 18214 2826 18222 2848
rect 18256 2848 18312 2860
rect 18346 2848 18402 2860
rect 18436 2848 18492 2860
rect 18256 2826 18280 2848
rect 18346 2826 18380 2848
rect 18436 2826 18480 2848
rect 18526 2826 18587 2860
rect 18214 2814 18280 2826
rect 18314 2814 18380 2826
rect 18414 2814 18480 2826
rect 18514 2814 18587 2826
rect 17893 2770 18587 2814
rect 17893 2736 17952 2770
rect 17986 2748 18042 2770
rect 18014 2736 18042 2748
rect 18076 2748 18132 2770
rect 18076 2736 18080 2748
rect 17893 2714 17980 2736
rect 18014 2714 18080 2736
rect 18114 2736 18132 2748
rect 18166 2748 18222 2770
rect 18166 2736 18180 2748
rect 18114 2714 18180 2736
rect 18214 2736 18222 2748
rect 18256 2748 18312 2770
rect 18346 2748 18402 2770
rect 18436 2748 18492 2770
rect 18256 2736 18280 2748
rect 18346 2736 18380 2748
rect 18436 2736 18480 2748
rect 18526 2736 18587 2770
rect 18214 2714 18280 2736
rect 18314 2714 18380 2736
rect 18414 2714 18480 2736
rect 18514 2714 18587 2736
rect 17893 2680 18587 2714
rect 17893 2646 17952 2680
rect 17986 2648 18042 2680
rect 18014 2646 18042 2648
rect 18076 2648 18132 2680
rect 18076 2646 18080 2648
rect 17893 2614 17980 2646
rect 18014 2614 18080 2646
rect 18114 2646 18132 2648
rect 18166 2648 18222 2680
rect 18166 2646 18180 2648
rect 18114 2614 18180 2646
rect 18214 2646 18222 2648
rect 18256 2648 18312 2680
rect 18346 2648 18402 2680
rect 18436 2648 18492 2680
rect 18256 2646 18280 2648
rect 18346 2646 18380 2648
rect 18436 2646 18480 2648
rect 18526 2646 18587 2680
rect 18214 2614 18280 2646
rect 18314 2614 18380 2646
rect 18414 2614 18480 2646
rect 18514 2614 18587 2646
rect 17893 2590 18587 2614
rect 17893 2556 17952 2590
rect 17986 2556 18042 2590
rect 18076 2556 18132 2590
rect 18166 2556 18222 2590
rect 18256 2556 18312 2590
rect 18346 2556 18402 2590
rect 18436 2556 18492 2590
rect 18526 2556 18587 2590
rect 17893 2548 18587 2556
rect 17893 2514 17980 2548
rect 18014 2514 18080 2548
rect 18114 2514 18180 2548
rect 18214 2514 18280 2548
rect 18314 2514 18380 2548
rect 18414 2514 18480 2548
rect 18514 2514 18587 2548
rect 17893 2500 18587 2514
rect 17893 2466 17952 2500
rect 17986 2466 18042 2500
rect 18076 2466 18132 2500
rect 18166 2466 18222 2500
rect 18256 2466 18312 2500
rect 18346 2466 18402 2500
rect 18436 2466 18492 2500
rect 18526 2466 18587 2500
rect 17893 2448 18587 2466
rect 17893 2414 17980 2448
rect 18014 2414 18080 2448
rect 18114 2414 18180 2448
rect 18214 2414 18280 2448
rect 18314 2414 18380 2448
rect 18414 2414 18480 2448
rect 18514 2414 18587 2448
rect 17893 2410 18587 2414
rect 17893 2376 17952 2410
rect 17986 2376 18042 2410
rect 18076 2376 18132 2410
rect 18166 2376 18222 2410
rect 18256 2376 18312 2410
rect 18346 2376 18402 2410
rect 18436 2376 18492 2410
rect 18526 2376 18587 2410
rect 17893 2348 18587 2376
rect 17893 2320 17980 2348
rect 18014 2320 18080 2348
rect 17893 2286 17952 2320
rect 18014 2314 18042 2320
rect 17986 2286 18042 2314
rect 18076 2314 18080 2320
rect 18114 2320 18180 2348
rect 18114 2314 18132 2320
rect 18076 2286 18132 2314
rect 18166 2314 18180 2320
rect 18214 2320 18280 2348
rect 18314 2320 18380 2348
rect 18414 2320 18480 2348
rect 18514 2320 18587 2348
rect 18214 2314 18222 2320
rect 18166 2286 18222 2314
rect 18256 2314 18280 2320
rect 18346 2314 18380 2320
rect 18436 2314 18480 2320
rect 18256 2286 18312 2314
rect 18346 2286 18402 2314
rect 18436 2286 18492 2314
rect 18526 2286 18587 2320
rect 17893 2227 18587 2286
rect 18649 2889 18668 2923
rect 18702 2922 18884 2923
rect 18702 2889 18816 2922
rect 18649 2888 18816 2889
rect 18850 2888 18884 2922
rect 18649 2833 18884 2888
rect 18649 2799 18668 2833
rect 18702 2832 18884 2833
rect 18702 2799 18816 2832
rect 18649 2798 18816 2799
rect 18850 2798 18884 2832
rect 18649 2743 18884 2798
rect 18649 2709 18668 2743
rect 18702 2742 18884 2743
rect 18702 2709 18816 2742
rect 18649 2708 18816 2709
rect 18850 2708 18884 2742
rect 18649 2653 18884 2708
rect 18649 2619 18668 2653
rect 18702 2652 18884 2653
rect 18702 2619 18816 2652
rect 18649 2618 18816 2619
rect 18850 2618 18884 2652
rect 18649 2563 18884 2618
rect 18649 2529 18668 2563
rect 18702 2562 18884 2563
rect 18702 2529 18816 2562
rect 18649 2528 18816 2529
rect 18850 2528 18884 2562
rect 18649 2473 18884 2528
rect 18649 2439 18668 2473
rect 18702 2472 18884 2473
rect 18702 2439 18816 2472
rect 18649 2438 18816 2439
rect 18850 2438 18884 2472
rect 18649 2383 18884 2438
rect 18649 2349 18668 2383
rect 18702 2382 18884 2383
rect 18702 2349 18816 2382
rect 18649 2348 18816 2349
rect 18850 2348 18884 2382
rect 18649 2293 18884 2348
rect 18649 2259 18668 2293
rect 18702 2292 18884 2293
rect 18702 2259 18816 2292
rect 18649 2258 18816 2259
rect 18850 2258 18884 2292
rect 17361 2203 17778 2222
rect 17361 2169 17380 2203
rect 17414 2202 17778 2203
rect 17414 2169 17528 2202
rect 17361 2168 17528 2169
rect 17562 2168 17629 2202
rect 17663 2188 17778 2202
rect 17812 2188 17831 2222
rect 17663 2168 17831 2188
rect 17361 2165 17831 2168
rect 18649 2203 18884 2258
rect 18649 2169 18668 2203
rect 18702 2202 18884 2203
rect 18702 2169 18816 2202
rect 18649 2168 18816 2169
rect 18850 2168 18884 2202
rect 18649 2165 18884 2168
rect 12444 2146 18884 2165
rect 12444 2112 12684 2146
rect 12718 2112 12774 2146
rect 12808 2112 12864 2146
rect 12898 2112 12954 2146
rect 12988 2112 13044 2146
rect 13078 2112 13134 2146
rect 13168 2112 13224 2146
rect 13258 2112 13314 2146
rect 13348 2112 13404 2146
rect 13438 2112 13972 2146
rect 14006 2112 14062 2146
rect 14096 2112 14152 2146
rect 14186 2112 14242 2146
rect 14276 2112 14332 2146
rect 14366 2112 14422 2146
rect 14456 2112 14512 2146
rect 14546 2112 14602 2146
rect 14636 2112 14692 2146
rect 14726 2112 15260 2146
rect 15294 2112 15350 2146
rect 15384 2112 15440 2146
rect 15474 2112 15530 2146
rect 15564 2112 15620 2146
rect 15654 2112 15710 2146
rect 15744 2112 15800 2146
rect 15834 2112 15890 2146
rect 15924 2112 15980 2146
rect 16014 2112 16548 2146
rect 16582 2112 16638 2146
rect 16672 2112 16728 2146
rect 16762 2112 16818 2146
rect 16852 2112 16908 2146
rect 16942 2112 16998 2146
rect 17032 2112 17088 2146
rect 17122 2112 17178 2146
rect 17212 2112 17268 2146
rect 17302 2112 17836 2146
rect 17870 2112 17926 2146
rect 17960 2112 18016 2146
rect 18050 2112 18106 2146
rect 18140 2112 18196 2146
rect 18230 2112 18286 2146
rect 18320 2112 18376 2146
rect 18410 2112 18466 2146
rect 18500 2112 18556 2146
rect 18590 2112 18884 2146
rect 12444 2078 12477 2112
rect 12511 2093 13664 2112
rect 12511 2078 12684 2093
rect 12444 2029 12684 2078
rect 13484 2078 13664 2093
rect 13698 2078 13765 2112
rect 13799 2093 14952 2112
rect 13799 2078 13984 2093
rect 13484 2029 13984 2078
rect 14784 2078 14952 2093
rect 14986 2078 15053 2112
rect 15087 2093 16240 2112
rect 15087 2078 15184 2093
rect 14784 2029 15184 2078
rect 16084 2078 16240 2093
rect 16274 2078 16341 2112
rect 16375 2093 17528 2112
rect 16375 2078 16484 2093
rect 16084 2029 16484 2078
rect 17384 2078 17528 2093
rect 17562 2078 17629 2112
rect 17663 2093 18816 2112
rect 17663 2078 17784 2093
rect 17384 2029 17784 2078
rect 18684 2078 18816 2093
rect 18850 2078 18884 2112
rect 18684 2029 18884 2078
rect 12444 2022 18884 2029
rect 12444 1988 12477 2022
rect 12511 1999 13664 2022
rect 12511 1988 12578 1999
rect 12444 1965 12578 1988
rect 12612 1965 12668 1999
rect 12702 1965 12758 1999
rect 12792 1965 12848 1999
rect 12882 1965 12938 1999
rect 12972 1965 13028 1999
rect 13062 1965 13118 1999
rect 13152 1965 13208 1999
rect 13242 1965 13298 1999
rect 13332 1965 13388 1999
rect 13422 1965 13478 1999
rect 13512 1965 13568 1999
rect 13602 1988 13664 1999
rect 13698 1988 13765 2022
rect 13799 1999 14952 2022
rect 13799 1988 13866 1999
rect 13602 1965 13866 1988
rect 13900 1965 13956 1999
rect 13990 1965 14046 1999
rect 14080 1965 14136 1999
rect 14170 1965 14226 1999
rect 14260 1965 14316 1999
rect 14350 1965 14406 1999
rect 14440 1965 14496 1999
rect 14530 1965 14586 1999
rect 14620 1965 14676 1999
rect 14710 1965 14766 1999
rect 14800 1965 14856 1999
rect 14890 1988 14952 1999
rect 14986 1988 15053 2022
rect 15087 1999 16240 2022
rect 15087 1988 15154 1999
rect 14890 1965 15154 1988
rect 15188 1965 15244 1999
rect 15278 1965 15334 1999
rect 15368 1965 15424 1999
rect 15458 1965 15514 1999
rect 15548 1965 15604 1999
rect 15638 1965 15694 1999
rect 15728 1965 15784 1999
rect 15818 1965 15874 1999
rect 15908 1965 15964 1999
rect 15998 1965 16054 1999
rect 16088 1965 16144 1999
rect 16178 1988 16240 1999
rect 16274 1988 16341 2022
rect 16375 1999 17528 2022
rect 16375 1988 16442 1999
rect 16178 1965 16442 1988
rect 16476 1965 16532 1999
rect 16566 1965 16622 1999
rect 16656 1965 16712 1999
rect 16746 1965 16802 1999
rect 16836 1965 16892 1999
rect 16926 1965 16982 1999
rect 17016 1965 17072 1999
rect 17106 1965 17162 1999
rect 17196 1965 17252 1999
rect 17286 1965 17342 1999
rect 17376 1965 17432 1999
rect 17466 1988 17528 1999
rect 17562 1988 17629 2022
rect 17663 1999 18816 2022
rect 17663 1988 17730 1999
rect 17466 1965 17730 1988
rect 17764 1965 17820 1999
rect 17854 1965 17910 1999
rect 17944 1965 18000 1999
rect 18034 1965 18090 1999
rect 18124 1965 18180 1999
rect 18214 1965 18270 1999
rect 18304 1965 18360 1999
rect 18394 1965 18450 1999
rect 18484 1965 18540 1999
rect 18574 1965 18630 1999
rect 18664 1965 18720 1999
rect 18754 1988 18816 1999
rect 18850 1988 18884 2022
rect 18754 1965 18884 1988
rect 12444 1930 18884 1965
rect 12484 1918 12684 1930
rect 13484 1918 13984 1930
rect 18684 1918 18884 1930
rect 7866 1100 7966 1200
rect 8366 1100 8466 1200
rect 7866 1000 8466 1100
<< viali >>
rect -21532 25036 -10316 25052
rect -21532 24270 -21516 25036
rect -21516 24270 -10332 25036
rect -10332 24270 -10316 25036
rect -21532 24254 -10316 24270
rect -5644 21579 -5106 21976
rect -4826 21579 -4288 21976
rect -4008 21579 -3470 21976
rect -3190 21579 -2652 21976
rect -736 21517 -198 21914
rect 82 21517 620 21914
rect 900 21517 1438 21914
rect 1718 21517 2256 21914
rect 2536 21517 3074 21914
rect 3354 21517 3892 21914
rect 4172 21517 4710 21914
rect 4990 21517 5528 21914
rect 5808 21517 6346 21914
rect 6626 21517 7164 21914
rect 7444 21517 7982 21914
rect 8262 21517 8800 21914
rect 9080 21517 9618 21914
rect 9898 21517 10436 21914
rect 10716 21517 11254 21914
rect 11534 21517 12072 21914
rect 12352 21517 12890 21914
rect -8916 20193 -8378 20590
rect -8098 20193 -7560 20590
rect -7280 20193 -6742 20590
rect -8916 16438 -8378 16835
rect -8098 16438 -7560 16835
rect -7280 16438 -6742 16835
rect -5644 16848 -5106 17245
rect -4826 16848 -4288 17245
rect -4008 16848 -3470 17245
rect -3190 16848 -2652 17245
rect -736 14782 -198 15179
rect 82 14781 620 15179
rect 900 14782 1438 15179
rect 1718 14782 2256 15179
rect 2536 14781 3074 15179
rect 3354 14782 3892 15179
rect 4172 14782 4710 15179
rect 4990 14781 5528 15179
rect 5808 14782 6346 15179
rect 6626 14782 7164 15179
rect 7444 14782 7982 15179
rect 8262 14781 8800 15179
rect 9080 14782 9618 15179
rect 9898 14782 10436 15179
rect 10716 14782 11254 15179
rect 11534 14782 12072 15179
rect 12352 14782 12890 15179
rect 12828 11842 12834 11864
rect 12834 11842 12862 11864
rect 12828 11830 12862 11842
rect 12928 11830 12962 11864
rect 13028 11830 13062 11864
rect 13128 11842 13160 11864
rect 13160 11842 13162 11864
rect 13228 11842 13250 11864
rect 13250 11842 13262 11864
rect 13328 11842 13340 11864
rect 13340 11842 13362 11864
rect 13128 11830 13162 11842
rect 13228 11830 13262 11842
rect 13328 11830 13362 11842
rect 12828 11752 12834 11764
rect 12834 11752 12862 11764
rect 12828 11730 12862 11752
rect 12928 11730 12962 11764
rect 13028 11730 13062 11764
rect 13128 11752 13160 11764
rect 13160 11752 13162 11764
rect 13228 11752 13250 11764
rect 13250 11752 13262 11764
rect 13328 11752 13340 11764
rect 13340 11752 13362 11764
rect 13128 11730 13162 11752
rect 13228 11730 13262 11752
rect 13328 11730 13362 11752
rect 12828 11662 12834 11664
rect 12834 11662 12862 11664
rect 12828 11630 12862 11662
rect 12928 11630 12962 11664
rect 13028 11630 13062 11664
rect 13128 11662 13160 11664
rect 13160 11662 13162 11664
rect 13228 11662 13250 11664
rect 13250 11662 13262 11664
rect 13328 11662 13340 11664
rect 13340 11662 13362 11664
rect 13128 11630 13162 11662
rect 13228 11630 13262 11662
rect 13328 11630 13362 11662
rect 12828 11530 12862 11564
rect 12928 11530 12962 11564
rect 13028 11530 13062 11564
rect 13128 11530 13162 11564
rect 13228 11530 13262 11564
rect 13328 11530 13362 11564
rect 12828 11430 12862 11464
rect 12928 11430 12962 11464
rect 13028 11430 13062 11464
rect 13128 11430 13162 11464
rect 13228 11430 13262 11464
rect 13328 11430 13362 11464
rect 12828 11336 12862 11364
rect 12828 11330 12834 11336
rect 12834 11330 12862 11336
rect 12928 11330 12962 11364
rect 13028 11330 13062 11364
rect 13128 11336 13162 11364
rect 13228 11336 13262 11364
rect 13328 11336 13362 11364
rect 13128 11330 13160 11336
rect 13160 11330 13162 11336
rect 13228 11330 13250 11336
rect 13250 11330 13262 11336
rect 13328 11330 13340 11336
rect 13340 11330 13362 11336
rect 14116 11842 14122 11864
rect 14122 11842 14150 11864
rect 14116 11830 14150 11842
rect 14216 11830 14250 11864
rect 14316 11830 14350 11864
rect 14416 11842 14448 11864
rect 14448 11842 14450 11864
rect 14516 11842 14538 11864
rect 14538 11842 14550 11864
rect 14616 11842 14628 11864
rect 14628 11842 14650 11864
rect 14416 11830 14450 11842
rect 14516 11830 14550 11842
rect 14616 11830 14650 11842
rect 14116 11752 14122 11764
rect 14122 11752 14150 11764
rect 14116 11730 14150 11752
rect 14216 11730 14250 11764
rect 14316 11730 14350 11764
rect 14416 11752 14448 11764
rect 14448 11752 14450 11764
rect 14516 11752 14538 11764
rect 14538 11752 14550 11764
rect 14616 11752 14628 11764
rect 14628 11752 14650 11764
rect 14416 11730 14450 11752
rect 14516 11730 14550 11752
rect 14616 11730 14650 11752
rect 14116 11662 14122 11664
rect 14122 11662 14150 11664
rect 14116 11630 14150 11662
rect 14216 11630 14250 11664
rect 14316 11630 14350 11664
rect 14416 11662 14448 11664
rect 14448 11662 14450 11664
rect 14516 11662 14538 11664
rect 14538 11662 14550 11664
rect 14616 11662 14628 11664
rect 14628 11662 14650 11664
rect 14416 11630 14450 11662
rect 14516 11630 14550 11662
rect 14616 11630 14650 11662
rect 14116 11530 14150 11564
rect 14216 11530 14250 11564
rect 14316 11530 14350 11564
rect 14416 11530 14450 11564
rect 14516 11530 14550 11564
rect 14616 11530 14650 11564
rect 14116 11430 14150 11464
rect 14216 11430 14250 11464
rect 14316 11430 14350 11464
rect 14416 11430 14450 11464
rect 14516 11430 14550 11464
rect 14616 11430 14650 11464
rect 14116 11336 14150 11364
rect 14116 11330 14122 11336
rect 14122 11330 14150 11336
rect 14216 11330 14250 11364
rect 14316 11330 14350 11364
rect 14416 11336 14450 11364
rect 14516 11336 14550 11364
rect 14616 11336 14650 11364
rect 14416 11330 14448 11336
rect 14448 11330 14450 11336
rect 14516 11330 14538 11336
rect 14538 11330 14550 11336
rect 14616 11330 14628 11336
rect 14628 11330 14650 11336
rect 15404 11842 15410 11864
rect 15410 11842 15438 11864
rect 15404 11830 15438 11842
rect 15504 11830 15538 11864
rect 15604 11830 15638 11864
rect 15704 11842 15736 11864
rect 15736 11842 15738 11864
rect 15804 11842 15826 11864
rect 15826 11842 15838 11864
rect 15904 11842 15916 11864
rect 15916 11842 15938 11864
rect 15704 11830 15738 11842
rect 15804 11830 15838 11842
rect 15904 11830 15938 11842
rect 15404 11752 15410 11764
rect 15410 11752 15438 11764
rect 15404 11730 15438 11752
rect 15504 11730 15538 11764
rect 15604 11730 15638 11764
rect 15704 11752 15736 11764
rect 15736 11752 15738 11764
rect 15804 11752 15826 11764
rect 15826 11752 15838 11764
rect 15904 11752 15916 11764
rect 15916 11752 15938 11764
rect 15704 11730 15738 11752
rect 15804 11730 15838 11752
rect 15904 11730 15938 11752
rect 15404 11662 15410 11664
rect 15410 11662 15438 11664
rect 15404 11630 15438 11662
rect 15504 11630 15538 11664
rect 15604 11630 15638 11664
rect 15704 11662 15736 11664
rect 15736 11662 15738 11664
rect 15804 11662 15826 11664
rect 15826 11662 15838 11664
rect 15904 11662 15916 11664
rect 15916 11662 15938 11664
rect 15704 11630 15738 11662
rect 15804 11630 15838 11662
rect 15904 11630 15938 11662
rect 15404 11530 15438 11564
rect 15504 11530 15538 11564
rect 15604 11530 15638 11564
rect 15704 11530 15738 11564
rect 15804 11530 15838 11564
rect 15904 11530 15938 11564
rect 15404 11430 15438 11464
rect 15504 11430 15538 11464
rect 15604 11430 15638 11464
rect 15704 11430 15738 11464
rect 15804 11430 15838 11464
rect 15904 11430 15938 11464
rect 15404 11336 15438 11364
rect 15404 11330 15410 11336
rect 15410 11330 15438 11336
rect 15504 11330 15538 11364
rect 15604 11330 15638 11364
rect 15704 11336 15738 11364
rect 15804 11336 15838 11364
rect 15904 11336 15938 11364
rect 15704 11330 15736 11336
rect 15736 11330 15738 11336
rect 15804 11330 15826 11336
rect 15826 11330 15838 11336
rect 15904 11330 15916 11336
rect 15916 11330 15938 11336
rect 16692 11842 16698 11864
rect 16698 11842 16726 11864
rect 16692 11830 16726 11842
rect 16792 11830 16826 11864
rect 16892 11830 16926 11864
rect 16992 11842 17024 11864
rect 17024 11842 17026 11864
rect 17092 11842 17114 11864
rect 17114 11842 17126 11864
rect 17192 11842 17204 11864
rect 17204 11842 17226 11864
rect 16992 11830 17026 11842
rect 17092 11830 17126 11842
rect 17192 11830 17226 11842
rect 16692 11752 16698 11764
rect 16698 11752 16726 11764
rect 16692 11730 16726 11752
rect 16792 11730 16826 11764
rect 16892 11730 16926 11764
rect 16992 11752 17024 11764
rect 17024 11752 17026 11764
rect 17092 11752 17114 11764
rect 17114 11752 17126 11764
rect 17192 11752 17204 11764
rect 17204 11752 17226 11764
rect 16992 11730 17026 11752
rect 17092 11730 17126 11752
rect 17192 11730 17226 11752
rect 16692 11662 16698 11664
rect 16698 11662 16726 11664
rect 16692 11630 16726 11662
rect 16792 11630 16826 11664
rect 16892 11630 16926 11664
rect 16992 11662 17024 11664
rect 17024 11662 17026 11664
rect 17092 11662 17114 11664
rect 17114 11662 17126 11664
rect 17192 11662 17204 11664
rect 17204 11662 17226 11664
rect 16992 11630 17026 11662
rect 17092 11630 17126 11662
rect 17192 11630 17226 11662
rect 16692 11530 16726 11564
rect 16792 11530 16826 11564
rect 16892 11530 16926 11564
rect 16992 11530 17026 11564
rect 17092 11530 17126 11564
rect 17192 11530 17226 11564
rect 16692 11430 16726 11464
rect 16792 11430 16826 11464
rect 16892 11430 16926 11464
rect 16992 11430 17026 11464
rect 17092 11430 17126 11464
rect 17192 11430 17226 11464
rect 16692 11336 16726 11364
rect 16692 11330 16698 11336
rect 16698 11330 16726 11336
rect 16792 11330 16826 11364
rect 16892 11330 16926 11364
rect 16992 11336 17026 11364
rect 17092 11336 17126 11364
rect 17192 11336 17226 11364
rect 16992 11330 17024 11336
rect 17024 11330 17026 11336
rect 17092 11330 17114 11336
rect 17114 11330 17126 11336
rect 17192 11330 17204 11336
rect 17204 11330 17226 11336
rect 17980 11842 17986 11864
rect 17986 11842 18014 11864
rect 17980 11830 18014 11842
rect 18080 11830 18114 11864
rect 18180 11830 18214 11864
rect 18280 11842 18312 11864
rect 18312 11842 18314 11864
rect 18380 11842 18402 11864
rect 18402 11842 18414 11864
rect 18480 11842 18492 11864
rect 18492 11842 18514 11864
rect 18280 11830 18314 11842
rect 18380 11830 18414 11842
rect 18480 11830 18514 11842
rect 17980 11752 17986 11764
rect 17986 11752 18014 11764
rect 17980 11730 18014 11752
rect 18080 11730 18114 11764
rect 18180 11730 18214 11764
rect 18280 11752 18312 11764
rect 18312 11752 18314 11764
rect 18380 11752 18402 11764
rect 18402 11752 18414 11764
rect 18480 11752 18492 11764
rect 18492 11752 18514 11764
rect 18280 11730 18314 11752
rect 18380 11730 18414 11752
rect 18480 11730 18514 11752
rect 17980 11662 17986 11664
rect 17986 11662 18014 11664
rect 17980 11630 18014 11662
rect 18080 11630 18114 11664
rect 18180 11630 18214 11664
rect 18280 11662 18312 11664
rect 18312 11662 18314 11664
rect 18380 11662 18402 11664
rect 18402 11662 18414 11664
rect 18480 11662 18492 11664
rect 18492 11662 18514 11664
rect 18280 11630 18314 11662
rect 18380 11630 18414 11662
rect 18480 11630 18514 11662
rect 17980 11530 18014 11564
rect 18080 11530 18114 11564
rect 18180 11530 18214 11564
rect 18280 11530 18314 11564
rect 18380 11530 18414 11564
rect 18480 11530 18514 11564
rect 17980 11430 18014 11464
rect 18080 11430 18114 11464
rect 18180 11430 18214 11464
rect 18280 11430 18314 11464
rect 18380 11430 18414 11464
rect 18480 11430 18514 11464
rect 17980 11336 18014 11364
rect 17980 11330 17986 11336
rect 17986 11330 18014 11336
rect 18080 11330 18114 11364
rect 18180 11330 18214 11364
rect 18280 11336 18314 11364
rect 18380 11336 18414 11364
rect 18480 11336 18514 11364
rect 18280 11330 18312 11336
rect 18312 11330 18314 11336
rect 18380 11330 18402 11336
rect 18402 11330 18414 11336
rect 18480 11330 18492 11336
rect 18492 11330 18514 11336
rect 12828 10554 12834 10576
rect 12834 10554 12862 10576
rect 12828 10542 12862 10554
rect 12928 10542 12962 10576
rect 13028 10542 13062 10576
rect 13128 10554 13160 10576
rect 13160 10554 13162 10576
rect 13228 10554 13250 10576
rect 13250 10554 13262 10576
rect 13328 10554 13340 10576
rect 13340 10554 13362 10576
rect 13128 10542 13162 10554
rect 13228 10542 13262 10554
rect 13328 10542 13362 10554
rect 12828 10464 12834 10476
rect 12834 10464 12862 10476
rect 12828 10442 12862 10464
rect 12928 10442 12962 10476
rect 13028 10442 13062 10476
rect 13128 10464 13160 10476
rect 13160 10464 13162 10476
rect 13228 10464 13250 10476
rect 13250 10464 13262 10476
rect 13328 10464 13340 10476
rect 13340 10464 13362 10476
rect 13128 10442 13162 10464
rect 13228 10442 13262 10464
rect 13328 10442 13362 10464
rect 12828 10374 12834 10376
rect 12834 10374 12862 10376
rect 12828 10342 12862 10374
rect 12928 10342 12962 10376
rect 13028 10342 13062 10376
rect 13128 10374 13160 10376
rect 13160 10374 13162 10376
rect 13228 10374 13250 10376
rect 13250 10374 13262 10376
rect 13328 10374 13340 10376
rect 13340 10374 13362 10376
rect 13128 10342 13162 10374
rect 13228 10342 13262 10374
rect 13328 10342 13362 10374
rect 12828 10242 12862 10276
rect 12928 10242 12962 10276
rect 13028 10242 13062 10276
rect 13128 10242 13162 10276
rect 13228 10242 13262 10276
rect 13328 10242 13362 10276
rect 12828 10142 12862 10176
rect 12928 10142 12962 10176
rect 13028 10142 13062 10176
rect 13128 10142 13162 10176
rect 13228 10142 13262 10176
rect 13328 10142 13362 10176
rect 12828 10048 12862 10076
rect 12828 10042 12834 10048
rect 12834 10042 12862 10048
rect 12928 10042 12962 10076
rect 13028 10042 13062 10076
rect 13128 10048 13162 10076
rect 13228 10048 13262 10076
rect 13328 10048 13362 10076
rect 13128 10042 13160 10048
rect 13160 10042 13162 10048
rect 13228 10042 13250 10048
rect 13250 10042 13262 10048
rect 13328 10042 13340 10048
rect 13340 10042 13362 10048
rect 14116 10554 14122 10576
rect 14122 10554 14150 10576
rect 14116 10542 14150 10554
rect 14216 10542 14250 10576
rect 14316 10542 14350 10576
rect 14416 10554 14448 10576
rect 14448 10554 14450 10576
rect 14516 10554 14538 10576
rect 14538 10554 14550 10576
rect 14616 10554 14628 10576
rect 14628 10554 14650 10576
rect 14416 10542 14450 10554
rect 14516 10542 14550 10554
rect 14616 10542 14650 10554
rect 14116 10464 14122 10476
rect 14122 10464 14150 10476
rect 14116 10442 14150 10464
rect 14216 10442 14250 10476
rect 14316 10442 14350 10476
rect 14416 10464 14448 10476
rect 14448 10464 14450 10476
rect 14516 10464 14538 10476
rect 14538 10464 14550 10476
rect 14616 10464 14628 10476
rect 14628 10464 14650 10476
rect 14416 10442 14450 10464
rect 14516 10442 14550 10464
rect 14616 10442 14650 10464
rect 14116 10374 14122 10376
rect 14122 10374 14150 10376
rect 14116 10342 14150 10374
rect 14216 10342 14250 10376
rect 14316 10342 14350 10376
rect 14416 10374 14448 10376
rect 14448 10374 14450 10376
rect 14516 10374 14538 10376
rect 14538 10374 14550 10376
rect 14616 10374 14628 10376
rect 14628 10374 14650 10376
rect 14416 10342 14450 10374
rect 14516 10342 14550 10374
rect 14616 10342 14650 10374
rect 14116 10242 14150 10276
rect 14216 10242 14250 10276
rect 14316 10242 14350 10276
rect 14416 10242 14450 10276
rect 14516 10242 14550 10276
rect 14616 10242 14650 10276
rect 14116 10142 14150 10176
rect 14216 10142 14250 10176
rect 14316 10142 14350 10176
rect 14416 10142 14450 10176
rect 14516 10142 14550 10176
rect 14616 10142 14650 10176
rect 14116 10048 14150 10076
rect 14116 10042 14122 10048
rect 14122 10042 14150 10048
rect 14216 10042 14250 10076
rect 14316 10042 14350 10076
rect 14416 10048 14450 10076
rect 14516 10048 14550 10076
rect 14616 10048 14650 10076
rect 14416 10042 14448 10048
rect 14448 10042 14450 10048
rect 14516 10042 14538 10048
rect 14538 10042 14550 10048
rect 14616 10042 14628 10048
rect 14628 10042 14650 10048
rect 15404 10554 15410 10576
rect 15410 10554 15438 10576
rect 15404 10542 15438 10554
rect 15504 10542 15538 10576
rect 15604 10542 15638 10576
rect 15704 10554 15736 10576
rect 15736 10554 15738 10576
rect 15804 10554 15826 10576
rect 15826 10554 15838 10576
rect 15904 10554 15916 10576
rect 15916 10554 15938 10576
rect 15704 10542 15738 10554
rect 15804 10542 15838 10554
rect 15904 10542 15938 10554
rect 15404 10464 15410 10476
rect 15410 10464 15438 10476
rect 15404 10442 15438 10464
rect 15504 10442 15538 10476
rect 15604 10442 15638 10476
rect 15704 10464 15736 10476
rect 15736 10464 15738 10476
rect 15804 10464 15826 10476
rect 15826 10464 15838 10476
rect 15904 10464 15916 10476
rect 15916 10464 15938 10476
rect 15704 10442 15738 10464
rect 15804 10442 15838 10464
rect 15904 10442 15938 10464
rect 15404 10374 15410 10376
rect 15410 10374 15438 10376
rect 15404 10342 15438 10374
rect 15504 10342 15538 10376
rect 15604 10342 15638 10376
rect 15704 10374 15736 10376
rect 15736 10374 15738 10376
rect 15804 10374 15826 10376
rect 15826 10374 15838 10376
rect 15904 10374 15916 10376
rect 15916 10374 15938 10376
rect 15704 10342 15738 10374
rect 15804 10342 15838 10374
rect 15904 10342 15938 10374
rect 15404 10242 15438 10276
rect 15504 10242 15538 10276
rect 15604 10242 15638 10276
rect 15704 10242 15738 10276
rect 15804 10242 15838 10276
rect 15904 10242 15938 10276
rect 15404 10142 15438 10176
rect 15504 10142 15538 10176
rect 15604 10142 15638 10176
rect 15704 10142 15738 10176
rect 15804 10142 15838 10176
rect 15904 10142 15938 10176
rect 15404 10048 15438 10076
rect 15404 10042 15410 10048
rect 15410 10042 15438 10048
rect 15504 10042 15538 10076
rect 15604 10042 15638 10076
rect 15704 10048 15738 10076
rect 15804 10048 15838 10076
rect 15904 10048 15938 10076
rect 15704 10042 15736 10048
rect 15736 10042 15738 10048
rect 15804 10042 15826 10048
rect 15826 10042 15838 10048
rect 15904 10042 15916 10048
rect 15916 10042 15938 10048
rect 16692 10554 16698 10576
rect 16698 10554 16726 10576
rect 16692 10542 16726 10554
rect 16792 10542 16826 10576
rect 16892 10542 16926 10576
rect 16992 10554 17024 10576
rect 17024 10554 17026 10576
rect 17092 10554 17114 10576
rect 17114 10554 17126 10576
rect 17192 10554 17204 10576
rect 17204 10554 17226 10576
rect 16992 10542 17026 10554
rect 17092 10542 17126 10554
rect 17192 10542 17226 10554
rect 16692 10464 16698 10476
rect 16698 10464 16726 10476
rect 16692 10442 16726 10464
rect 16792 10442 16826 10476
rect 16892 10442 16926 10476
rect 16992 10464 17024 10476
rect 17024 10464 17026 10476
rect 17092 10464 17114 10476
rect 17114 10464 17126 10476
rect 17192 10464 17204 10476
rect 17204 10464 17226 10476
rect 16992 10442 17026 10464
rect 17092 10442 17126 10464
rect 17192 10442 17226 10464
rect 16692 10374 16698 10376
rect 16698 10374 16726 10376
rect 16692 10342 16726 10374
rect 16792 10342 16826 10376
rect 16892 10342 16926 10376
rect 16992 10374 17024 10376
rect 17024 10374 17026 10376
rect 17092 10374 17114 10376
rect 17114 10374 17126 10376
rect 17192 10374 17204 10376
rect 17204 10374 17226 10376
rect 16992 10342 17026 10374
rect 17092 10342 17126 10374
rect 17192 10342 17226 10374
rect 16692 10242 16726 10276
rect 16792 10242 16826 10276
rect 16892 10242 16926 10276
rect 16992 10242 17026 10276
rect 17092 10242 17126 10276
rect 17192 10242 17226 10276
rect 16692 10142 16726 10176
rect 16792 10142 16826 10176
rect 16892 10142 16926 10176
rect 16992 10142 17026 10176
rect 17092 10142 17126 10176
rect 17192 10142 17226 10176
rect 16692 10048 16726 10076
rect 16692 10042 16698 10048
rect 16698 10042 16726 10048
rect 16792 10042 16826 10076
rect 16892 10042 16926 10076
rect 16992 10048 17026 10076
rect 17092 10048 17126 10076
rect 17192 10048 17226 10076
rect 16992 10042 17024 10048
rect 17024 10042 17026 10048
rect 17092 10042 17114 10048
rect 17114 10042 17126 10048
rect 17192 10042 17204 10048
rect 17204 10042 17226 10048
rect 17980 10554 17986 10576
rect 17986 10554 18014 10576
rect 17980 10542 18014 10554
rect 18080 10542 18114 10576
rect 18180 10542 18214 10576
rect 18280 10554 18312 10576
rect 18312 10554 18314 10576
rect 18380 10554 18402 10576
rect 18402 10554 18414 10576
rect 18480 10554 18492 10576
rect 18492 10554 18514 10576
rect 18280 10542 18314 10554
rect 18380 10542 18414 10554
rect 18480 10542 18514 10554
rect 17980 10464 17986 10476
rect 17986 10464 18014 10476
rect 17980 10442 18014 10464
rect 18080 10442 18114 10476
rect 18180 10442 18214 10476
rect 18280 10464 18312 10476
rect 18312 10464 18314 10476
rect 18380 10464 18402 10476
rect 18402 10464 18414 10476
rect 18480 10464 18492 10476
rect 18492 10464 18514 10476
rect 18280 10442 18314 10464
rect 18380 10442 18414 10464
rect 18480 10442 18514 10464
rect 17980 10374 17986 10376
rect 17986 10374 18014 10376
rect 17980 10342 18014 10374
rect 18080 10342 18114 10376
rect 18180 10342 18214 10376
rect 18280 10374 18312 10376
rect 18312 10374 18314 10376
rect 18380 10374 18402 10376
rect 18402 10374 18414 10376
rect 18480 10374 18492 10376
rect 18492 10374 18514 10376
rect 18280 10342 18314 10374
rect 18380 10342 18414 10374
rect 18480 10342 18514 10374
rect 17980 10242 18014 10276
rect 18080 10242 18114 10276
rect 18180 10242 18214 10276
rect 18280 10242 18314 10276
rect 18380 10242 18414 10276
rect 18480 10242 18514 10276
rect 17980 10142 18014 10176
rect 18080 10142 18114 10176
rect 18180 10142 18214 10176
rect 18280 10142 18314 10176
rect 18380 10142 18414 10176
rect 18480 10142 18514 10176
rect 17980 10048 18014 10076
rect 17980 10042 17986 10048
rect 17986 10042 18014 10048
rect 18080 10042 18114 10076
rect 18180 10042 18214 10076
rect 18280 10048 18314 10076
rect 18380 10048 18414 10076
rect 18480 10048 18514 10076
rect 18280 10042 18312 10048
rect 18312 10042 18314 10048
rect 18380 10042 18402 10048
rect 18402 10042 18414 10048
rect 18480 10042 18492 10048
rect 18492 10042 18514 10048
rect -17888 9382 -11424 9388
rect -17888 9050 -17882 9382
rect -17882 9050 -11430 9382
rect -11430 9050 -11424 9382
rect -17888 9044 -11424 9050
rect -17164 8818 -11788 8852
rect -17248 8514 -17214 8698
rect -17164 8360 -11788 8394
rect -16728 6692 -16544 6726
rect -16156 6692 -15972 6726
rect -15584 6692 -15400 6726
rect -15012 6692 -14828 6726
rect -14440 6692 -14256 6726
rect -13868 6692 -13684 6726
rect -13296 6692 -13112 6726
rect -12724 6692 -12540 6726
rect -20906 5668 -20854 5720
rect -19990 5668 -19938 5720
rect -21658 5570 -21474 5604
rect -21200 5570 -21016 5604
rect -20742 5570 -20558 5604
rect -20284 5570 -20100 5604
rect -19826 5570 -19642 5604
rect -19368 5570 -19184 5604
rect -21812 5144 -21778 5520
rect -21354 5144 -21320 5520
rect -20896 5144 -20862 5520
rect -20438 5144 -20404 5520
rect -19980 5144 -19946 5520
rect -19522 5144 -19488 5520
rect -19064 5144 -19030 5520
rect -17434 5044 -17334 6642
rect -16882 4866 -16848 6642
rect -16424 4866 -16390 6642
rect -16310 4866 -16276 6642
rect -15852 4866 -15818 6642
rect -15738 4866 -15704 6642
rect -15280 4866 -15246 6642
rect -15166 4866 -15132 6642
rect -14708 4866 -14674 6642
rect -14594 4866 -14560 6642
rect -14136 4866 -14102 6642
rect -14022 4866 -13988 6642
rect -13564 4866 -13530 6642
rect -13450 4866 -13416 6642
rect -12992 4866 -12958 6642
rect -12878 4866 -12844 6642
rect -12420 4866 -12386 6642
rect -11934 5044 -11834 6642
rect -18454 4289 -18270 4323
rect -17882 4289 -17698 4323
rect -17310 4289 -17126 4323
rect -16738 4289 -16554 4323
rect -16166 4289 -15982 4323
rect -15594 4289 -15410 4323
rect -15022 4289 -14838 4323
rect -14450 4289 -14266 4323
rect -13878 4289 -13694 4323
rect -13306 4289 -13122 4323
rect -12734 4289 -12550 4323
rect -12162 4289 -11978 4323
rect -11590 4289 -11406 4323
rect -11018 4289 -10834 4323
rect -19250 1800 -19150 4142
rect -18608 1674 -18574 4230
rect -18150 1674 -18116 4230
rect -18036 1674 -18002 4230
rect -17578 1674 -17544 4230
rect -17464 1674 -17430 4230
rect -17006 1674 -16972 4230
rect -16892 1674 -16858 4230
rect -16434 1674 -16400 4230
rect -16320 1674 -16286 4230
rect -15862 1674 -15828 4230
rect -15748 1674 -15714 4230
rect -15290 1674 -15256 4230
rect -15176 1674 -15142 4230
rect -14718 1674 -14684 4230
rect -14604 1674 -14570 4230
rect -14146 1674 -14112 4230
rect -14032 1674 -13998 4230
rect -13574 1674 -13540 4230
rect -13460 1674 -13426 4230
rect -13002 1674 -12968 4230
rect -12888 1674 -12854 4230
rect -12430 1674 -12396 4230
rect -12316 1674 -12282 4230
rect -11858 1674 -11824 4230
rect -11744 1674 -11710 4230
rect -11286 1674 -11252 4230
rect -11172 1674 -11138 4230
rect -10714 1674 -10680 4230
rect -10122 1800 -10022 4142
rect -15668 1196 -13326 1296
rect -8800 1712 -8766 9428
rect -8342 1712 -8308 9428
rect -7884 1712 -7850 9428
rect -7426 1712 -7392 9428
rect -6968 1712 -6934 9428
rect -6510 1712 -6476 9428
rect -6052 1712 -6018 9428
rect -5594 1712 -5560 9428
rect -5136 1712 -5102 9428
rect -4678 1712 -4644 9428
rect -4220 1712 -4186 9428
rect -3762 1712 -3728 9428
rect -8646 1619 -8462 1653
rect -8188 1619 -8004 1653
rect -7730 1619 -7546 1653
rect -7272 1619 -7088 1653
rect -6814 1619 -6630 1653
rect -6356 1619 -6172 1653
rect -5898 1619 -5714 1653
rect -5440 1619 -5256 1653
rect -4982 1619 -4798 1653
rect -4524 1619 -4340 1653
rect -4066 1619 -3882 1653
rect -9400 1102 -9000 1202
rect -2842 1712 -2808 9428
rect -2384 1712 -2350 9428
rect -1926 1712 -1892 9428
rect -1468 1712 -1434 9428
rect -1010 1712 -976 9428
rect -552 1712 -518 9428
rect -94 1712 -60 9428
rect 364 1712 398 9428
rect 822 1712 856 9428
rect 1280 1712 1314 9428
rect 1738 1712 1772 9428
rect -2688 1619 -2504 1653
rect -2230 1619 -2046 1653
rect -1772 1619 -1588 1653
rect -1314 1619 -1130 1653
rect -856 1619 -672 1653
rect -398 1619 -214 1653
rect 60 1619 244 1653
rect 518 1619 702 1653
rect 976 1619 1160 1653
rect 1434 1619 1618 1653
rect -3490 1102 -3090 1202
rect 2658 1712 2692 9428
rect 3116 1712 3150 9428
rect 3574 1712 3608 9428
rect 4032 1712 4066 9428
rect 4490 1712 4524 9428
rect 4948 1712 4982 9428
rect 5406 1712 5440 9428
rect 5864 1712 5898 9428
rect 6322 1712 6356 9428
rect 6780 1712 6814 9428
rect 7238 1712 7272 9428
rect 7696 1712 7730 9428
rect 2812 1619 2996 1653
rect 3270 1619 3454 1653
rect 3728 1619 3912 1653
rect 4186 1619 4370 1653
rect 4644 1619 4828 1653
rect 5102 1619 5286 1653
rect 5560 1619 5744 1653
rect 6018 1619 6202 1653
rect 6476 1619 6660 1653
rect 6934 1619 7118 1653
rect 7392 1619 7576 1653
rect 2010 1102 2410 1202
rect 12828 9266 12834 9288
rect 12834 9266 12862 9288
rect 12828 9254 12862 9266
rect 12928 9254 12962 9288
rect 13028 9254 13062 9288
rect 13128 9266 13160 9288
rect 13160 9266 13162 9288
rect 13228 9266 13250 9288
rect 13250 9266 13262 9288
rect 13328 9266 13340 9288
rect 13340 9266 13362 9288
rect 13128 9254 13162 9266
rect 13228 9254 13262 9266
rect 13328 9254 13362 9266
rect 12828 9176 12834 9188
rect 12834 9176 12862 9188
rect 12828 9154 12862 9176
rect 12928 9154 12962 9188
rect 13028 9154 13062 9188
rect 13128 9176 13160 9188
rect 13160 9176 13162 9188
rect 13228 9176 13250 9188
rect 13250 9176 13262 9188
rect 13328 9176 13340 9188
rect 13340 9176 13362 9188
rect 13128 9154 13162 9176
rect 13228 9154 13262 9176
rect 13328 9154 13362 9176
rect 12828 9086 12834 9088
rect 12834 9086 12862 9088
rect 12828 9054 12862 9086
rect 12928 9054 12962 9088
rect 13028 9054 13062 9088
rect 13128 9086 13160 9088
rect 13160 9086 13162 9088
rect 13228 9086 13250 9088
rect 13250 9086 13262 9088
rect 13328 9086 13340 9088
rect 13340 9086 13362 9088
rect 13128 9054 13162 9086
rect 13228 9054 13262 9086
rect 13328 9054 13362 9086
rect 12828 8954 12862 8988
rect 12928 8954 12962 8988
rect 13028 8954 13062 8988
rect 13128 8954 13162 8988
rect 13228 8954 13262 8988
rect 13328 8954 13362 8988
rect 12828 8854 12862 8888
rect 12928 8854 12962 8888
rect 13028 8854 13062 8888
rect 13128 8854 13162 8888
rect 13228 8854 13262 8888
rect 13328 8854 13362 8888
rect 12828 8760 12862 8788
rect 12828 8754 12834 8760
rect 12834 8754 12862 8760
rect 12928 8754 12962 8788
rect 13028 8754 13062 8788
rect 13128 8760 13162 8788
rect 13228 8760 13262 8788
rect 13328 8760 13362 8788
rect 13128 8754 13160 8760
rect 13160 8754 13162 8760
rect 13228 8754 13250 8760
rect 13250 8754 13262 8760
rect 13328 8754 13340 8760
rect 13340 8754 13362 8760
rect 14116 9266 14122 9288
rect 14122 9266 14150 9288
rect 14116 9254 14150 9266
rect 14216 9254 14250 9288
rect 14316 9254 14350 9288
rect 14416 9266 14448 9288
rect 14448 9266 14450 9288
rect 14516 9266 14538 9288
rect 14538 9266 14550 9288
rect 14616 9266 14628 9288
rect 14628 9266 14650 9288
rect 14416 9254 14450 9266
rect 14516 9254 14550 9266
rect 14616 9254 14650 9266
rect 14116 9176 14122 9188
rect 14122 9176 14150 9188
rect 14116 9154 14150 9176
rect 14216 9154 14250 9188
rect 14316 9154 14350 9188
rect 14416 9176 14448 9188
rect 14448 9176 14450 9188
rect 14516 9176 14538 9188
rect 14538 9176 14550 9188
rect 14616 9176 14628 9188
rect 14628 9176 14650 9188
rect 14416 9154 14450 9176
rect 14516 9154 14550 9176
rect 14616 9154 14650 9176
rect 14116 9086 14122 9088
rect 14122 9086 14150 9088
rect 14116 9054 14150 9086
rect 14216 9054 14250 9088
rect 14316 9054 14350 9088
rect 14416 9086 14448 9088
rect 14448 9086 14450 9088
rect 14516 9086 14538 9088
rect 14538 9086 14550 9088
rect 14616 9086 14628 9088
rect 14628 9086 14650 9088
rect 14416 9054 14450 9086
rect 14516 9054 14550 9086
rect 14616 9054 14650 9086
rect 14116 8954 14150 8988
rect 14216 8954 14250 8988
rect 14316 8954 14350 8988
rect 14416 8954 14450 8988
rect 14516 8954 14550 8988
rect 14616 8954 14650 8988
rect 14116 8854 14150 8888
rect 14216 8854 14250 8888
rect 14316 8854 14350 8888
rect 14416 8854 14450 8888
rect 14516 8854 14550 8888
rect 14616 8854 14650 8888
rect 14116 8760 14150 8788
rect 14116 8754 14122 8760
rect 14122 8754 14150 8760
rect 14216 8754 14250 8788
rect 14316 8754 14350 8788
rect 14416 8760 14450 8788
rect 14516 8760 14550 8788
rect 14616 8760 14650 8788
rect 14416 8754 14448 8760
rect 14448 8754 14450 8760
rect 14516 8754 14538 8760
rect 14538 8754 14550 8760
rect 14616 8754 14628 8760
rect 14628 8754 14650 8760
rect 15404 9266 15410 9288
rect 15410 9266 15438 9288
rect 15404 9254 15438 9266
rect 15504 9254 15538 9288
rect 15604 9254 15638 9288
rect 15704 9266 15736 9288
rect 15736 9266 15738 9288
rect 15804 9266 15826 9288
rect 15826 9266 15838 9288
rect 15904 9266 15916 9288
rect 15916 9266 15938 9288
rect 15704 9254 15738 9266
rect 15804 9254 15838 9266
rect 15904 9254 15938 9266
rect 15404 9176 15410 9188
rect 15410 9176 15438 9188
rect 15404 9154 15438 9176
rect 15504 9154 15538 9188
rect 15604 9154 15638 9188
rect 15704 9176 15736 9188
rect 15736 9176 15738 9188
rect 15804 9176 15826 9188
rect 15826 9176 15838 9188
rect 15904 9176 15916 9188
rect 15916 9176 15938 9188
rect 15704 9154 15738 9176
rect 15804 9154 15838 9176
rect 15904 9154 15938 9176
rect 15404 9086 15410 9088
rect 15410 9086 15438 9088
rect 15404 9054 15438 9086
rect 15504 9054 15538 9088
rect 15604 9054 15638 9088
rect 15704 9086 15736 9088
rect 15736 9086 15738 9088
rect 15804 9086 15826 9088
rect 15826 9086 15838 9088
rect 15904 9086 15916 9088
rect 15916 9086 15938 9088
rect 15704 9054 15738 9086
rect 15804 9054 15838 9086
rect 15904 9054 15938 9086
rect 15404 8954 15438 8988
rect 15504 8954 15538 8988
rect 15604 8954 15638 8988
rect 15704 8954 15738 8988
rect 15804 8954 15838 8988
rect 15904 8954 15938 8988
rect 15404 8854 15438 8888
rect 15504 8854 15538 8888
rect 15604 8854 15638 8888
rect 15704 8854 15738 8888
rect 15804 8854 15838 8888
rect 15904 8854 15938 8888
rect 15404 8760 15438 8788
rect 15404 8754 15410 8760
rect 15410 8754 15438 8760
rect 15504 8754 15538 8788
rect 15604 8754 15638 8788
rect 15704 8760 15738 8788
rect 15804 8760 15838 8788
rect 15904 8760 15938 8788
rect 15704 8754 15736 8760
rect 15736 8754 15738 8760
rect 15804 8754 15826 8760
rect 15826 8754 15838 8760
rect 15904 8754 15916 8760
rect 15916 8754 15938 8760
rect 16692 9266 16698 9288
rect 16698 9266 16726 9288
rect 16692 9254 16726 9266
rect 16792 9254 16826 9288
rect 16892 9254 16926 9288
rect 16992 9266 17024 9288
rect 17024 9266 17026 9288
rect 17092 9266 17114 9288
rect 17114 9266 17126 9288
rect 17192 9266 17204 9288
rect 17204 9266 17226 9288
rect 16992 9254 17026 9266
rect 17092 9254 17126 9266
rect 17192 9254 17226 9266
rect 16692 9176 16698 9188
rect 16698 9176 16726 9188
rect 16692 9154 16726 9176
rect 16792 9154 16826 9188
rect 16892 9154 16926 9188
rect 16992 9176 17024 9188
rect 17024 9176 17026 9188
rect 17092 9176 17114 9188
rect 17114 9176 17126 9188
rect 17192 9176 17204 9188
rect 17204 9176 17226 9188
rect 16992 9154 17026 9176
rect 17092 9154 17126 9176
rect 17192 9154 17226 9176
rect 16692 9086 16698 9088
rect 16698 9086 16726 9088
rect 16692 9054 16726 9086
rect 16792 9054 16826 9088
rect 16892 9054 16926 9088
rect 16992 9086 17024 9088
rect 17024 9086 17026 9088
rect 17092 9086 17114 9088
rect 17114 9086 17126 9088
rect 17192 9086 17204 9088
rect 17204 9086 17226 9088
rect 16992 9054 17026 9086
rect 17092 9054 17126 9086
rect 17192 9054 17226 9086
rect 16692 8954 16726 8988
rect 16792 8954 16826 8988
rect 16892 8954 16926 8988
rect 16992 8954 17026 8988
rect 17092 8954 17126 8988
rect 17192 8954 17226 8988
rect 16692 8854 16726 8888
rect 16792 8854 16826 8888
rect 16892 8854 16926 8888
rect 16992 8854 17026 8888
rect 17092 8854 17126 8888
rect 17192 8854 17226 8888
rect 16692 8760 16726 8788
rect 16692 8754 16698 8760
rect 16698 8754 16726 8760
rect 16792 8754 16826 8788
rect 16892 8754 16926 8788
rect 16992 8760 17026 8788
rect 17092 8760 17126 8788
rect 17192 8760 17226 8788
rect 16992 8754 17024 8760
rect 17024 8754 17026 8760
rect 17092 8754 17114 8760
rect 17114 8754 17126 8760
rect 17192 8754 17204 8760
rect 17204 8754 17226 8760
rect 17980 9266 17986 9288
rect 17986 9266 18014 9288
rect 17980 9254 18014 9266
rect 18080 9254 18114 9288
rect 18180 9254 18214 9288
rect 18280 9266 18312 9288
rect 18312 9266 18314 9288
rect 18380 9266 18402 9288
rect 18402 9266 18414 9288
rect 18480 9266 18492 9288
rect 18492 9266 18514 9288
rect 18280 9254 18314 9266
rect 18380 9254 18414 9266
rect 18480 9254 18514 9266
rect 17980 9176 17986 9188
rect 17986 9176 18014 9188
rect 17980 9154 18014 9176
rect 18080 9154 18114 9188
rect 18180 9154 18214 9188
rect 18280 9176 18312 9188
rect 18312 9176 18314 9188
rect 18380 9176 18402 9188
rect 18402 9176 18414 9188
rect 18480 9176 18492 9188
rect 18492 9176 18514 9188
rect 18280 9154 18314 9176
rect 18380 9154 18414 9176
rect 18480 9154 18514 9176
rect 17980 9086 17986 9088
rect 17986 9086 18014 9088
rect 17980 9054 18014 9086
rect 18080 9054 18114 9088
rect 18180 9054 18214 9088
rect 18280 9086 18312 9088
rect 18312 9086 18314 9088
rect 18380 9086 18402 9088
rect 18402 9086 18414 9088
rect 18480 9086 18492 9088
rect 18492 9086 18514 9088
rect 18280 9054 18314 9086
rect 18380 9054 18414 9086
rect 18480 9054 18514 9086
rect 17980 8954 18014 8988
rect 18080 8954 18114 8988
rect 18180 8954 18214 8988
rect 18280 8954 18314 8988
rect 18380 8954 18414 8988
rect 18480 8954 18514 8988
rect 17980 8854 18014 8888
rect 18080 8854 18114 8888
rect 18180 8854 18214 8888
rect 18280 8854 18314 8888
rect 18380 8854 18414 8888
rect 18480 8854 18514 8888
rect 17980 8760 18014 8788
rect 17980 8754 17986 8760
rect 17986 8754 18014 8760
rect 18080 8754 18114 8788
rect 18180 8754 18214 8788
rect 18280 8760 18314 8788
rect 18380 8760 18414 8788
rect 18480 8760 18514 8788
rect 18280 8754 18312 8760
rect 18312 8754 18314 8760
rect 18380 8754 18402 8760
rect 18402 8754 18414 8760
rect 18480 8754 18492 8760
rect 18492 8754 18514 8760
rect 12828 7978 12834 8000
rect 12834 7978 12862 8000
rect 12828 7966 12862 7978
rect 12928 7966 12962 8000
rect 13028 7966 13062 8000
rect 13128 7978 13160 8000
rect 13160 7978 13162 8000
rect 13228 7978 13250 8000
rect 13250 7978 13262 8000
rect 13328 7978 13340 8000
rect 13340 7978 13362 8000
rect 13128 7966 13162 7978
rect 13228 7966 13262 7978
rect 13328 7966 13362 7978
rect 12828 7888 12834 7900
rect 12834 7888 12862 7900
rect 12828 7866 12862 7888
rect 12928 7866 12962 7900
rect 13028 7866 13062 7900
rect 13128 7888 13160 7900
rect 13160 7888 13162 7900
rect 13228 7888 13250 7900
rect 13250 7888 13262 7900
rect 13328 7888 13340 7900
rect 13340 7888 13362 7900
rect 13128 7866 13162 7888
rect 13228 7866 13262 7888
rect 13328 7866 13362 7888
rect 12828 7798 12834 7800
rect 12834 7798 12862 7800
rect 12828 7766 12862 7798
rect 12928 7766 12962 7800
rect 13028 7766 13062 7800
rect 13128 7798 13160 7800
rect 13160 7798 13162 7800
rect 13228 7798 13250 7800
rect 13250 7798 13262 7800
rect 13328 7798 13340 7800
rect 13340 7798 13362 7800
rect 13128 7766 13162 7798
rect 13228 7766 13262 7798
rect 13328 7766 13362 7798
rect 12828 7666 12862 7700
rect 12928 7666 12962 7700
rect 13028 7666 13062 7700
rect 13128 7666 13162 7700
rect 13228 7666 13262 7700
rect 13328 7666 13362 7700
rect 12828 7566 12862 7600
rect 12928 7566 12962 7600
rect 13028 7566 13062 7600
rect 13128 7566 13162 7600
rect 13228 7566 13262 7600
rect 13328 7566 13362 7600
rect 12828 7472 12862 7500
rect 12828 7466 12834 7472
rect 12834 7466 12862 7472
rect 12928 7466 12962 7500
rect 13028 7466 13062 7500
rect 13128 7472 13162 7500
rect 13228 7472 13262 7500
rect 13328 7472 13362 7500
rect 13128 7466 13160 7472
rect 13160 7466 13162 7472
rect 13228 7466 13250 7472
rect 13250 7466 13262 7472
rect 13328 7466 13340 7472
rect 13340 7466 13362 7472
rect 14116 7978 14122 8000
rect 14122 7978 14150 8000
rect 14116 7966 14150 7978
rect 14216 7966 14250 8000
rect 14316 7966 14350 8000
rect 14416 7978 14448 8000
rect 14448 7978 14450 8000
rect 14516 7978 14538 8000
rect 14538 7978 14550 8000
rect 14616 7978 14628 8000
rect 14628 7978 14650 8000
rect 14416 7966 14450 7978
rect 14516 7966 14550 7978
rect 14616 7966 14650 7978
rect 14116 7888 14122 7900
rect 14122 7888 14150 7900
rect 14116 7866 14150 7888
rect 14216 7866 14250 7900
rect 14316 7866 14350 7900
rect 14416 7888 14448 7900
rect 14448 7888 14450 7900
rect 14516 7888 14538 7900
rect 14538 7888 14550 7900
rect 14616 7888 14628 7900
rect 14628 7888 14650 7900
rect 14416 7866 14450 7888
rect 14516 7866 14550 7888
rect 14616 7866 14650 7888
rect 14116 7798 14122 7800
rect 14122 7798 14150 7800
rect 14116 7766 14150 7798
rect 14216 7766 14250 7800
rect 14316 7766 14350 7800
rect 14416 7798 14448 7800
rect 14448 7798 14450 7800
rect 14516 7798 14538 7800
rect 14538 7798 14550 7800
rect 14616 7798 14628 7800
rect 14628 7798 14650 7800
rect 14416 7766 14450 7798
rect 14516 7766 14550 7798
rect 14616 7766 14650 7798
rect 14116 7666 14150 7700
rect 14216 7666 14250 7700
rect 14316 7666 14350 7700
rect 14416 7666 14450 7700
rect 14516 7666 14550 7700
rect 14616 7666 14650 7700
rect 14116 7566 14150 7600
rect 14216 7566 14250 7600
rect 14316 7566 14350 7600
rect 14416 7566 14450 7600
rect 14516 7566 14550 7600
rect 14616 7566 14650 7600
rect 14116 7472 14150 7500
rect 14116 7466 14122 7472
rect 14122 7466 14150 7472
rect 14216 7466 14250 7500
rect 14316 7466 14350 7500
rect 14416 7472 14450 7500
rect 14516 7472 14550 7500
rect 14616 7472 14650 7500
rect 14416 7466 14448 7472
rect 14448 7466 14450 7472
rect 14516 7466 14538 7472
rect 14538 7466 14550 7472
rect 14616 7466 14628 7472
rect 14628 7466 14650 7472
rect 15404 7978 15410 8000
rect 15410 7978 15438 8000
rect 15404 7966 15438 7978
rect 15504 7966 15538 8000
rect 15604 7966 15638 8000
rect 15704 7978 15736 8000
rect 15736 7978 15738 8000
rect 15804 7978 15826 8000
rect 15826 7978 15838 8000
rect 15904 7978 15916 8000
rect 15916 7978 15938 8000
rect 15704 7966 15738 7978
rect 15804 7966 15838 7978
rect 15904 7966 15938 7978
rect 15404 7888 15410 7900
rect 15410 7888 15438 7900
rect 15404 7866 15438 7888
rect 15504 7866 15538 7900
rect 15604 7866 15638 7900
rect 15704 7888 15736 7900
rect 15736 7888 15738 7900
rect 15804 7888 15826 7900
rect 15826 7888 15838 7900
rect 15904 7888 15916 7900
rect 15916 7888 15938 7900
rect 15704 7866 15738 7888
rect 15804 7866 15838 7888
rect 15904 7866 15938 7888
rect 15404 7798 15410 7800
rect 15410 7798 15438 7800
rect 15404 7766 15438 7798
rect 15504 7766 15538 7800
rect 15604 7766 15638 7800
rect 15704 7798 15736 7800
rect 15736 7798 15738 7800
rect 15804 7798 15826 7800
rect 15826 7798 15838 7800
rect 15904 7798 15916 7800
rect 15916 7798 15938 7800
rect 15704 7766 15738 7798
rect 15804 7766 15838 7798
rect 15904 7766 15938 7798
rect 15404 7666 15438 7700
rect 15504 7666 15538 7700
rect 15604 7666 15638 7700
rect 15704 7666 15738 7700
rect 15804 7666 15838 7700
rect 15904 7666 15938 7700
rect 15404 7566 15438 7600
rect 15504 7566 15538 7600
rect 15604 7566 15638 7600
rect 15704 7566 15738 7600
rect 15804 7566 15838 7600
rect 15904 7566 15938 7600
rect 15404 7472 15438 7500
rect 15404 7466 15410 7472
rect 15410 7466 15438 7472
rect 15504 7466 15538 7500
rect 15604 7466 15638 7500
rect 15704 7472 15738 7500
rect 15804 7472 15838 7500
rect 15904 7472 15938 7500
rect 15704 7466 15736 7472
rect 15736 7466 15738 7472
rect 15804 7466 15826 7472
rect 15826 7466 15838 7472
rect 15904 7466 15916 7472
rect 15916 7466 15938 7472
rect 16692 7978 16698 8000
rect 16698 7978 16726 8000
rect 16692 7966 16726 7978
rect 16792 7966 16826 8000
rect 16892 7966 16926 8000
rect 16992 7978 17024 8000
rect 17024 7978 17026 8000
rect 17092 7978 17114 8000
rect 17114 7978 17126 8000
rect 17192 7978 17204 8000
rect 17204 7978 17226 8000
rect 16992 7966 17026 7978
rect 17092 7966 17126 7978
rect 17192 7966 17226 7978
rect 16692 7888 16698 7900
rect 16698 7888 16726 7900
rect 16692 7866 16726 7888
rect 16792 7866 16826 7900
rect 16892 7866 16926 7900
rect 16992 7888 17024 7900
rect 17024 7888 17026 7900
rect 17092 7888 17114 7900
rect 17114 7888 17126 7900
rect 17192 7888 17204 7900
rect 17204 7888 17226 7900
rect 16992 7866 17026 7888
rect 17092 7866 17126 7888
rect 17192 7866 17226 7888
rect 16692 7798 16698 7800
rect 16698 7798 16726 7800
rect 16692 7766 16726 7798
rect 16792 7766 16826 7800
rect 16892 7766 16926 7800
rect 16992 7798 17024 7800
rect 17024 7798 17026 7800
rect 17092 7798 17114 7800
rect 17114 7798 17126 7800
rect 17192 7798 17204 7800
rect 17204 7798 17226 7800
rect 16992 7766 17026 7798
rect 17092 7766 17126 7798
rect 17192 7766 17226 7798
rect 16692 7666 16726 7700
rect 16792 7666 16826 7700
rect 16892 7666 16926 7700
rect 16992 7666 17026 7700
rect 17092 7666 17126 7700
rect 17192 7666 17226 7700
rect 16692 7566 16726 7600
rect 16792 7566 16826 7600
rect 16892 7566 16926 7600
rect 16992 7566 17026 7600
rect 17092 7566 17126 7600
rect 17192 7566 17226 7600
rect 16692 7472 16726 7500
rect 16692 7466 16698 7472
rect 16698 7466 16726 7472
rect 16792 7466 16826 7500
rect 16892 7466 16926 7500
rect 16992 7472 17026 7500
rect 17092 7472 17126 7500
rect 17192 7472 17226 7500
rect 16992 7466 17024 7472
rect 17024 7466 17026 7472
rect 17092 7466 17114 7472
rect 17114 7466 17126 7472
rect 17192 7466 17204 7472
rect 17204 7466 17226 7472
rect 17980 7978 17986 8000
rect 17986 7978 18014 8000
rect 17980 7966 18014 7978
rect 18080 7966 18114 8000
rect 18180 7966 18214 8000
rect 18280 7978 18312 8000
rect 18312 7978 18314 8000
rect 18380 7978 18402 8000
rect 18402 7978 18414 8000
rect 18480 7978 18492 8000
rect 18492 7978 18514 8000
rect 18280 7966 18314 7978
rect 18380 7966 18414 7978
rect 18480 7966 18514 7978
rect 17980 7888 17986 7900
rect 17986 7888 18014 7900
rect 17980 7866 18014 7888
rect 18080 7866 18114 7900
rect 18180 7866 18214 7900
rect 18280 7888 18312 7900
rect 18312 7888 18314 7900
rect 18380 7888 18402 7900
rect 18402 7888 18414 7900
rect 18480 7888 18492 7900
rect 18492 7888 18514 7900
rect 18280 7866 18314 7888
rect 18380 7866 18414 7888
rect 18480 7866 18514 7888
rect 17980 7798 17986 7800
rect 17986 7798 18014 7800
rect 17980 7766 18014 7798
rect 18080 7766 18114 7800
rect 18180 7766 18214 7800
rect 18280 7798 18312 7800
rect 18312 7798 18314 7800
rect 18380 7798 18402 7800
rect 18402 7798 18414 7800
rect 18480 7798 18492 7800
rect 18492 7798 18514 7800
rect 18280 7766 18314 7798
rect 18380 7766 18414 7798
rect 18480 7766 18514 7798
rect 17980 7666 18014 7700
rect 18080 7666 18114 7700
rect 18180 7666 18214 7700
rect 18280 7666 18314 7700
rect 18380 7666 18414 7700
rect 18480 7666 18514 7700
rect 17980 7566 18014 7600
rect 18080 7566 18114 7600
rect 18180 7566 18214 7600
rect 18280 7566 18314 7600
rect 18380 7566 18414 7600
rect 18480 7566 18514 7600
rect 17980 7472 18014 7500
rect 17980 7466 17986 7472
rect 17986 7466 18014 7472
rect 18080 7466 18114 7500
rect 18180 7466 18214 7500
rect 18280 7472 18314 7500
rect 18380 7472 18414 7500
rect 18480 7472 18514 7500
rect 18280 7466 18312 7472
rect 18312 7466 18314 7472
rect 18380 7466 18402 7472
rect 18402 7466 18414 7472
rect 18480 7466 18492 7472
rect 18492 7466 18514 7472
rect 12828 6690 12834 6712
rect 12834 6690 12862 6712
rect 12828 6678 12862 6690
rect 12928 6678 12962 6712
rect 13028 6678 13062 6712
rect 13128 6690 13160 6712
rect 13160 6690 13162 6712
rect 13228 6690 13250 6712
rect 13250 6690 13262 6712
rect 13328 6690 13340 6712
rect 13340 6690 13362 6712
rect 13128 6678 13162 6690
rect 13228 6678 13262 6690
rect 13328 6678 13362 6690
rect 12828 6600 12834 6612
rect 12834 6600 12862 6612
rect 12828 6578 12862 6600
rect 12928 6578 12962 6612
rect 13028 6578 13062 6612
rect 13128 6600 13160 6612
rect 13160 6600 13162 6612
rect 13228 6600 13250 6612
rect 13250 6600 13262 6612
rect 13328 6600 13340 6612
rect 13340 6600 13362 6612
rect 13128 6578 13162 6600
rect 13228 6578 13262 6600
rect 13328 6578 13362 6600
rect 12828 6510 12834 6512
rect 12834 6510 12862 6512
rect 12828 6478 12862 6510
rect 12928 6478 12962 6512
rect 13028 6478 13062 6512
rect 13128 6510 13160 6512
rect 13160 6510 13162 6512
rect 13228 6510 13250 6512
rect 13250 6510 13262 6512
rect 13328 6510 13340 6512
rect 13340 6510 13362 6512
rect 13128 6478 13162 6510
rect 13228 6478 13262 6510
rect 13328 6478 13362 6510
rect 12828 6378 12862 6412
rect 12928 6378 12962 6412
rect 13028 6378 13062 6412
rect 13128 6378 13162 6412
rect 13228 6378 13262 6412
rect 13328 6378 13362 6412
rect 12828 6278 12862 6312
rect 12928 6278 12962 6312
rect 13028 6278 13062 6312
rect 13128 6278 13162 6312
rect 13228 6278 13262 6312
rect 13328 6278 13362 6312
rect 12828 6184 12862 6212
rect 12828 6178 12834 6184
rect 12834 6178 12862 6184
rect 12928 6178 12962 6212
rect 13028 6178 13062 6212
rect 13128 6184 13162 6212
rect 13228 6184 13262 6212
rect 13328 6184 13362 6212
rect 13128 6178 13160 6184
rect 13160 6178 13162 6184
rect 13228 6178 13250 6184
rect 13250 6178 13262 6184
rect 13328 6178 13340 6184
rect 13340 6178 13362 6184
rect 14116 6690 14122 6712
rect 14122 6690 14150 6712
rect 14116 6678 14150 6690
rect 14216 6678 14250 6712
rect 14316 6678 14350 6712
rect 14416 6690 14448 6712
rect 14448 6690 14450 6712
rect 14516 6690 14538 6712
rect 14538 6690 14550 6712
rect 14616 6690 14628 6712
rect 14628 6690 14650 6712
rect 14416 6678 14450 6690
rect 14516 6678 14550 6690
rect 14616 6678 14650 6690
rect 14116 6600 14122 6612
rect 14122 6600 14150 6612
rect 14116 6578 14150 6600
rect 14216 6578 14250 6612
rect 14316 6578 14350 6612
rect 14416 6600 14448 6612
rect 14448 6600 14450 6612
rect 14516 6600 14538 6612
rect 14538 6600 14550 6612
rect 14616 6600 14628 6612
rect 14628 6600 14650 6612
rect 14416 6578 14450 6600
rect 14516 6578 14550 6600
rect 14616 6578 14650 6600
rect 14116 6510 14122 6512
rect 14122 6510 14150 6512
rect 14116 6478 14150 6510
rect 14216 6478 14250 6512
rect 14316 6478 14350 6512
rect 14416 6510 14448 6512
rect 14448 6510 14450 6512
rect 14516 6510 14538 6512
rect 14538 6510 14550 6512
rect 14616 6510 14628 6512
rect 14628 6510 14650 6512
rect 14416 6478 14450 6510
rect 14516 6478 14550 6510
rect 14616 6478 14650 6510
rect 14116 6378 14150 6412
rect 14216 6378 14250 6412
rect 14316 6378 14350 6412
rect 14416 6378 14450 6412
rect 14516 6378 14550 6412
rect 14616 6378 14650 6412
rect 14116 6278 14150 6312
rect 14216 6278 14250 6312
rect 14316 6278 14350 6312
rect 14416 6278 14450 6312
rect 14516 6278 14550 6312
rect 14616 6278 14650 6312
rect 14116 6184 14150 6212
rect 14116 6178 14122 6184
rect 14122 6178 14150 6184
rect 14216 6178 14250 6212
rect 14316 6178 14350 6212
rect 14416 6184 14450 6212
rect 14516 6184 14550 6212
rect 14616 6184 14650 6212
rect 14416 6178 14448 6184
rect 14448 6178 14450 6184
rect 14516 6178 14538 6184
rect 14538 6178 14550 6184
rect 14616 6178 14628 6184
rect 14628 6178 14650 6184
rect 15404 6690 15410 6712
rect 15410 6690 15438 6712
rect 15404 6678 15438 6690
rect 15504 6678 15538 6712
rect 15604 6678 15638 6712
rect 15704 6690 15736 6712
rect 15736 6690 15738 6712
rect 15804 6690 15826 6712
rect 15826 6690 15838 6712
rect 15904 6690 15916 6712
rect 15916 6690 15938 6712
rect 15704 6678 15738 6690
rect 15804 6678 15838 6690
rect 15904 6678 15938 6690
rect 15404 6600 15410 6612
rect 15410 6600 15438 6612
rect 15404 6578 15438 6600
rect 15504 6578 15538 6612
rect 15604 6578 15638 6612
rect 15704 6600 15736 6612
rect 15736 6600 15738 6612
rect 15804 6600 15826 6612
rect 15826 6600 15838 6612
rect 15904 6600 15916 6612
rect 15916 6600 15938 6612
rect 15704 6578 15738 6600
rect 15804 6578 15838 6600
rect 15904 6578 15938 6600
rect 15404 6510 15410 6512
rect 15410 6510 15438 6512
rect 15404 6478 15438 6510
rect 15504 6478 15538 6512
rect 15604 6478 15638 6512
rect 15704 6510 15736 6512
rect 15736 6510 15738 6512
rect 15804 6510 15826 6512
rect 15826 6510 15838 6512
rect 15904 6510 15916 6512
rect 15916 6510 15938 6512
rect 15704 6478 15738 6510
rect 15804 6478 15838 6510
rect 15904 6478 15938 6510
rect 15404 6378 15438 6412
rect 15504 6378 15538 6412
rect 15604 6378 15638 6412
rect 15704 6378 15738 6412
rect 15804 6378 15838 6412
rect 15904 6378 15938 6412
rect 15404 6278 15438 6312
rect 15504 6278 15538 6312
rect 15604 6278 15638 6312
rect 15704 6278 15738 6312
rect 15804 6278 15838 6312
rect 15904 6278 15938 6312
rect 15404 6184 15438 6212
rect 15404 6178 15410 6184
rect 15410 6178 15438 6184
rect 15504 6178 15538 6212
rect 15604 6178 15638 6212
rect 15704 6184 15738 6212
rect 15804 6184 15838 6212
rect 15904 6184 15938 6212
rect 15704 6178 15736 6184
rect 15736 6178 15738 6184
rect 15804 6178 15826 6184
rect 15826 6178 15838 6184
rect 15904 6178 15916 6184
rect 15916 6178 15938 6184
rect 16692 6690 16698 6712
rect 16698 6690 16726 6712
rect 16692 6678 16726 6690
rect 16792 6678 16826 6712
rect 16892 6678 16926 6712
rect 16992 6690 17024 6712
rect 17024 6690 17026 6712
rect 17092 6690 17114 6712
rect 17114 6690 17126 6712
rect 17192 6690 17204 6712
rect 17204 6690 17226 6712
rect 16992 6678 17026 6690
rect 17092 6678 17126 6690
rect 17192 6678 17226 6690
rect 16692 6600 16698 6612
rect 16698 6600 16726 6612
rect 16692 6578 16726 6600
rect 16792 6578 16826 6612
rect 16892 6578 16926 6612
rect 16992 6600 17024 6612
rect 17024 6600 17026 6612
rect 17092 6600 17114 6612
rect 17114 6600 17126 6612
rect 17192 6600 17204 6612
rect 17204 6600 17226 6612
rect 16992 6578 17026 6600
rect 17092 6578 17126 6600
rect 17192 6578 17226 6600
rect 16692 6510 16698 6512
rect 16698 6510 16726 6512
rect 16692 6478 16726 6510
rect 16792 6478 16826 6512
rect 16892 6478 16926 6512
rect 16992 6510 17024 6512
rect 17024 6510 17026 6512
rect 17092 6510 17114 6512
rect 17114 6510 17126 6512
rect 17192 6510 17204 6512
rect 17204 6510 17226 6512
rect 16992 6478 17026 6510
rect 17092 6478 17126 6510
rect 17192 6478 17226 6510
rect 16692 6378 16726 6412
rect 16792 6378 16826 6412
rect 16892 6378 16926 6412
rect 16992 6378 17026 6412
rect 17092 6378 17126 6412
rect 17192 6378 17226 6412
rect 16692 6278 16726 6312
rect 16792 6278 16826 6312
rect 16892 6278 16926 6312
rect 16992 6278 17026 6312
rect 17092 6278 17126 6312
rect 17192 6278 17226 6312
rect 16692 6184 16726 6212
rect 16692 6178 16698 6184
rect 16698 6178 16726 6184
rect 16792 6178 16826 6212
rect 16892 6178 16926 6212
rect 16992 6184 17026 6212
rect 17092 6184 17126 6212
rect 17192 6184 17226 6212
rect 16992 6178 17024 6184
rect 17024 6178 17026 6184
rect 17092 6178 17114 6184
rect 17114 6178 17126 6184
rect 17192 6178 17204 6184
rect 17204 6178 17226 6184
rect 17980 6690 17986 6712
rect 17986 6690 18014 6712
rect 17980 6678 18014 6690
rect 18080 6678 18114 6712
rect 18180 6678 18214 6712
rect 18280 6690 18312 6712
rect 18312 6690 18314 6712
rect 18380 6690 18402 6712
rect 18402 6690 18414 6712
rect 18480 6690 18492 6712
rect 18492 6690 18514 6712
rect 18280 6678 18314 6690
rect 18380 6678 18414 6690
rect 18480 6678 18514 6690
rect 17980 6600 17986 6612
rect 17986 6600 18014 6612
rect 17980 6578 18014 6600
rect 18080 6578 18114 6612
rect 18180 6578 18214 6612
rect 18280 6600 18312 6612
rect 18312 6600 18314 6612
rect 18380 6600 18402 6612
rect 18402 6600 18414 6612
rect 18480 6600 18492 6612
rect 18492 6600 18514 6612
rect 18280 6578 18314 6600
rect 18380 6578 18414 6600
rect 18480 6578 18514 6600
rect 17980 6510 17986 6512
rect 17986 6510 18014 6512
rect 17980 6478 18014 6510
rect 18080 6478 18114 6512
rect 18180 6478 18214 6512
rect 18280 6510 18312 6512
rect 18312 6510 18314 6512
rect 18380 6510 18402 6512
rect 18402 6510 18414 6512
rect 18480 6510 18492 6512
rect 18492 6510 18514 6512
rect 18280 6478 18314 6510
rect 18380 6478 18414 6510
rect 18480 6478 18514 6510
rect 17980 6378 18014 6412
rect 18080 6378 18114 6412
rect 18180 6378 18214 6412
rect 18280 6378 18314 6412
rect 18380 6378 18414 6412
rect 18480 6378 18514 6412
rect 17980 6278 18014 6312
rect 18080 6278 18114 6312
rect 18180 6278 18214 6312
rect 18280 6278 18314 6312
rect 18380 6278 18414 6312
rect 18480 6278 18514 6312
rect 17980 6184 18014 6212
rect 17980 6178 17986 6184
rect 17986 6178 18014 6184
rect 18080 6178 18114 6212
rect 18180 6178 18214 6212
rect 18280 6184 18314 6212
rect 18380 6184 18414 6212
rect 18480 6184 18514 6212
rect 18280 6178 18312 6184
rect 18312 6178 18314 6184
rect 18380 6178 18402 6184
rect 18402 6178 18414 6184
rect 18480 6178 18492 6184
rect 18492 6178 18514 6184
rect 12828 5402 12834 5424
rect 12834 5402 12862 5424
rect 12828 5390 12862 5402
rect 12928 5390 12962 5424
rect 13028 5390 13062 5424
rect 13128 5402 13160 5424
rect 13160 5402 13162 5424
rect 13228 5402 13250 5424
rect 13250 5402 13262 5424
rect 13328 5402 13340 5424
rect 13340 5402 13362 5424
rect 13128 5390 13162 5402
rect 13228 5390 13262 5402
rect 13328 5390 13362 5402
rect 12828 5312 12834 5324
rect 12834 5312 12862 5324
rect 12828 5290 12862 5312
rect 12928 5290 12962 5324
rect 13028 5290 13062 5324
rect 13128 5312 13160 5324
rect 13160 5312 13162 5324
rect 13228 5312 13250 5324
rect 13250 5312 13262 5324
rect 13328 5312 13340 5324
rect 13340 5312 13362 5324
rect 13128 5290 13162 5312
rect 13228 5290 13262 5312
rect 13328 5290 13362 5312
rect 12828 5222 12834 5224
rect 12834 5222 12862 5224
rect 12828 5190 12862 5222
rect 12928 5190 12962 5224
rect 13028 5190 13062 5224
rect 13128 5222 13160 5224
rect 13160 5222 13162 5224
rect 13228 5222 13250 5224
rect 13250 5222 13262 5224
rect 13328 5222 13340 5224
rect 13340 5222 13362 5224
rect 13128 5190 13162 5222
rect 13228 5190 13262 5222
rect 13328 5190 13362 5222
rect 12828 5090 12862 5124
rect 12928 5090 12962 5124
rect 13028 5090 13062 5124
rect 13128 5090 13162 5124
rect 13228 5090 13262 5124
rect 13328 5090 13362 5124
rect 12828 4990 12862 5024
rect 12928 4990 12962 5024
rect 13028 4990 13062 5024
rect 13128 4990 13162 5024
rect 13228 4990 13262 5024
rect 13328 4990 13362 5024
rect 12828 4896 12862 4924
rect 12828 4890 12834 4896
rect 12834 4890 12862 4896
rect 12928 4890 12962 4924
rect 13028 4890 13062 4924
rect 13128 4896 13162 4924
rect 13228 4896 13262 4924
rect 13328 4896 13362 4924
rect 13128 4890 13160 4896
rect 13160 4890 13162 4896
rect 13228 4890 13250 4896
rect 13250 4890 13262 4896
rect 13328 4890 13340 4896
rect 13340 4890 13362 4896
rect 14116 5402 14122 5424
rect 14122 5402 14150 5424
rect 14116 5390 14150 5402
rect 14216 5390 14250 5424
rect 14316 5390 14350 5424
rect 14416 5402 14448 5424
rect 14448 5402 14450 5424
rect 14516 5402 14538 5424
rect 14538 5402 14550 5424
rect 14616 5402 14628 5424
rect 14628 5402 14650 5424
rect 14416 5390 14450 5402
rect 14516 5390 14550 5402
rect 14616 5390 14650 5402
rect 14116 5312 14122 5324
rect 14122 5312 14150 5324
rect 14116 5290 14150 5312
rect 14216 5290 14250 5324
rect 14316 5290 14350 5324
rect 14416 5312 14448 5324
rect 14448 5312 14450 5324
rect 14516 5312 14538 5324
rect 14538 5312 14550 5324
rect 14616 5312 14628 5324
rect 14628 5312 14650 5324
rect 14416 5290 14450 5312
rect 14516 5290 14550 5312
rect 14616 5290 14650 5312
rect 14116 5222 14122 5224
rect 14122 5222 14150 5224
rect 14116 5190 14150 5222
rect 14216 5190 14250 5224
rect 14316 5190 14350 5224
rect 14416 5222 14448 5224
rect 14448 5222 14450 5224
rect 14516 5222 14538 5224
rect 14538 5222 14550 5224
rect 14616 5222 14628 5224
rect 14628 5222 14650 5224
rect 14416 5190 14450 5222
rect 14516 5190 14550 5222
rect 14616 5190 14650 5222
rect 14116 5090 14150 5124
rect 14216 5090 14250 5124
rect 14316 5090 14350 5124
rect 14416 5090 14450 5124
rect 14516 5090 14550 5124
rect 14616 5090 14650 5124
rect 14116 4990 14150 5024
rect 14216 4990 14250 5024
rect 14316 4990 14350 5024
rect 14416 4990 14450 5024
rect 14516 4990 14550 5024
rect 14616 4990 14650 5024
rect 14116 4896 14150 4924
rect 14116 4890 14122 4896
rect 14122 4890 14150 4896
rect 14216 4890 14250 4924
rect 14316 4890 14350 4924
rect 14416 4896 14450 4924
rect 14516 4896 14550 4924
rect 14616 4896 14650 4924
rect 14416 4890 14448 4896
rect 14448 4890 14450 4896
rect 14516 4890 14538 4896
rect 14538 4890 14550 4896
rect 14616 4890 14628 4896
rect 14628 4890 14650 4896
rect 15404 5402 15410 5424
rect 15410 5402 15438 5424
rect 15404 5390 15438 5402
rect 15504 5390 15538 5424
rect 15604 5390 15638 5424
rect 15704 5402 15736 5424
rect 15736 5402 15738 5424
rect 15804 5402 15826 5424
rect 15826 5402 15838 5424
rect 15904 5402 15916 5424
rect 15916 5402 15938 5424
rect 15704 5390 15738 5402
rect 15804 5390 15838 5402
rect 15904 5390 15938 5402
rect 15404 5312 15410 5324
rect 15410 5312 15438 5324
rect 15404 5290 15438 5312
rect 15504 5290 15538 5324
rect 15604 5290 15638 5324
rect 15704 5312 15736 5324
rect 15736 5312 15738 5324
rect 15804 5312 15826 5324
rect 15826 5312 15838 5324
rect 15904 5312 15916 5324
rect 15916 5312 15938 5324
rect 15704 5290 15738 5312
rect 15804 5290 15838 5312
rect 15904 5290 15938 5312
rect 15404 5222 15410 5224
rect 15410 5222 15438 5224
rect 15404 5190 15438 5222
rect 15504 5190 15538 5224
rect 15604 5190 15638 5224
rect 15704 5222 15736 5224
rect 15736 5222 15738 5224
rect 15804 5222 15826 5224
rect 15826 5222 15838 5224
rect 15904 5222 15916 5224
rect 15916 5222 15938 5224
rect 15704 5190 15738 5222
rect 15804 5190 15838 5222
rect 15904 5190 15938 5222
rect 15404 5090 15438 5124
rect 15504 5090 15538 5124
rect 15604 5090 15638 5124
rect 15704 5090 15738 5124
rect 15804 5090 15838 5124
rect 15904 5090 15938 5124
rect 15404 4990 15438 5024
rect 15504 4990 15538 5024
rect 15604 4990 15638 5024
rect 15704 4990 15738 5024
rect 15804 4990 15838 5024
rect 15904 4990 15938 5024
rect 15404 4896 15438 4924
rect 15404 4890 15410 4896
rect 15410 4890 15438 4896
rect 15504 4890 15538 4924
rect 15604 4890 15638 4924
rect 15704 4896 15738 4924
rect 15804 4896 15838 4924
rect 15904 4896 15938 4924
rect 15704 4890 15736 4896
rect 15736 4890 15738 4896
rect 15804 4890 15826 4896
rect 15826 4890 15838 4896
rect 15904 4890 15916 4896
rect 15916 4890 15938 4896
rect 16692 5402 16698 5424
rect 16698 5402 16726 5424
rect 16692 5390 16726 5402
rect 16792 5390 16826 5424
rect 16892 5390 16926 5424
rect 16992 5402 17024 5424
rect 17024 5402 17026 5424
rect 17092 5402 17114 5424
rect 17114 5402 17126 5424
rect 17192 5402 17204 5424
rect 17204 5402 17226 5424
rect 16992 5390 17026 5402
rect 17092 5390 17126 5402
rect 17192 5390 17226 5402
rect 16692 5312 16698 5324
rect 16698 5312 16726 5324
rect 16692 5290 16726 5312
rect 16792 5290 16826 5324
rect 16892 5290 16926 5324
rect 16992 5312 17024 5324
rect 17024 5312 17026 5324
rect 17092 5312 17114 5324
rect 17114 5312 17126 5324
rect 17192 5312 17204 5324
rect 17204 5312 17226 5324
rect 16992 5290 17026 5312
rect 17092 5290 17126 5312
rect 17192 5290 17226 5312
rect 16692 5222 16698 5224
rect 16698 5222 16726 5224
rect 16692 5190 16726 5222
rect 16792 5190 16826 5224
rect 16892 5190 16926 5224
rect 16992 5222 17024 5224
rect 17024 5222 17026 5224
rect 17092 5222 17114 5224
rect 17114 5222 17126 5224
rect 17192 5222 17204 5224
rect 17204 5222 17226 5224
rect 16992 5190 17026 5222
rect 17092 5190 17126 5222
rect 17192 5190 17226 5222
rect 16692 5090 16726 5124
rect 16792 5090 16826 5124
rect 16892 5090 16926 5124
rect 16992 5090 17026 5124
rect 17092 5090 17126 5124
rect 17192 5090 17226 5124
rect 16692 4990 16726 5024
rect 16792 4990 16826 5024
rect 16892 4990 16926 5024
rect 16992 4990 17026 5024
rect 17092 4990 17126 5024
rect 17192 4990 17226 5024
rect 16692 4896 16726 4924
rect 16692 4890 16698 4896
rect 16698 4890 16726 4896
rect 16792 4890 16826 4924
rect 16892 4890 16926 4924
rect 16992 4896 17026 4924
rect 17092 4896 17126 4924
rect 17192 4896 17226 4924
rect 16992 4890 17024 4896
rect 17024 4890 17026 4896
rect 17092 4890 17114 4896
rect 17114 4890 17126 4896
rect 17192 4890 17204 4896
rect 17204 4890 17226 4896
rect 17980 5402 17986 5424
rect 17986 5402 18014 5424
rect 17980 5390 18014 5402
rect 18080 5390 18114 5424
rect 18180 5390 18214 5424
rect 18280 5402 18312 5424
rect 18312 5402 18314 5424
rect 18380 5402 18402 5424
rect 18402 5402 18414 5424
rect 18480 5402 18492 5424
rect 18492 5402 18514 5424
rect 18280 5390 18314 5402
rect 18380 5390 18414 5402
rect 18480 5390 18514 5402
rect 17980 5312 17986 5324
rect 17986 5312 18014 5324
rect 17980 5290 18014 5312
rect 18080 5290 18114 5324
rect 18180 5290 18214 5324
rect 18280 5312 18312 5324
rect 18312 5312 18314 5324
rect 18380 5312 18402 5324
rect 18402 5312 18414 5324
rect 18480 5312 18492 5324
rect 18492 5312 18514 5324
rect 18280 5290 18314 5312
rect 18380 5290 18414 5312
rect 18480 5290 18514 5312
rect 17980 5222 17986 5224
rect 17986 5222 18014 5224
rect 17980 5190 18014 5222
rect 18080 5190 18114 5224
rect 18180 5190 18214 5224
rect 18280 5222 18312 5224
rect 18312 5222 18314 5224
rect 18380 5222 18402 5224
rect 18402 5222 18414 5224
rect 18480 5222 18492 5224
rect 18492 5222 18514 5224
rect 18280 5190 18314 5222
rect 18380 5190 18414 5222
rect 18480 5190 18514 5222
rect 17980 5090 18014 5124
rect 18080 5090 18114 5124
rect 18180 5090 18214 5124
rect 18280 5090 18314 5124
rect 18380 5090 18414 5124
rect 18480 5090 18514 5124
rect 17980 4990 18014 5024
rect 18080 4990 18114 5024
rect 18180 4990 18214 5024
rect 18280 4990 18314 5024
rect 18380 4990 18414 5024
rect 18480 4990 18514 5024
rect 17980 4896 18014 4924
rect 17980 4890 17986 4896
rect 17986 4890 18014 4896
rect 18080 4890 18114 4924
rect 18180 4890 18214 4924
rect 18280 4896 18314 4924
rect 18380 4896 18414 4924
rect 18480 4896 18514 4924
rect 18280 4890 18312 4896
rect 18312 4890 18314 4896
rect 18380 4890 18402 4896
rect 18402 4890 18414 4896
rect 18480 4890 18492 4896
rect 18492 4890 18514 4896
rect 12828 4114 12834 4136
rect 12834 4114 12862 4136
rect 12828 4102 12862 4114
rect 12928 4102 12962 4136
rect 13028 4102 13062 4136
rect 13128 4114 13160 4136
rect 13160 4114 13162 4136
rect 13228 4114 13250 4136
rect 13250 4114 13262 4136
rect 13328 4114 13340 4136
rect 13340 4114 13362 4136
rect 13128 4102 13162 4114
rect 13228 4102 13262 4114
rect 13328 4102 13362 4114
rect 12828 4024 12834 4036
rect 12834 4024 12862 4036
rect 12828 4002 12862 4024
rect 12928 4002 12962 4036
rect 13028 4002 13062 4036
rect 13128 4024 13160 4036
rect 13160 4024 13162 4036
rect 13228 4024 13250 4036
rect 13250 4024 13262 4036
rect 13328 4024 13340 4036
rect 13340 4024 13362 4036
rect 13128 4002 13162 4024
rect 13228 4002 13262 4024
rect 13328 4002 13362 4024
rect 12828 3934 12834 3936
rect 12834 3934 12862 3936
rect 12828 3902 12862 3934
rect 12928 3902 12962 3936
rect 13028 3902 13062 3936
rect 13128 3934 13160 3936
rect 13160 3934 13162 3936
rect 13228 3934 13250 3936
rect 13250 3934 13262 3936
rect 13328 3934 13340 3936
rect 13340 3934 13362 3936
rect 13128 3902 13162 3934
rect 13228 3902 13262 3934
rect 13328 3902 13362 3934
rect 12828 3802 12862 3836
rect 12928 3802 12962 3836
rect 13028 3802 13062 3836
rect 13128 3802 13162 3836
rect 13228 3802 13262 3836
rect 13328 3802 13362 3836
rect 12828 3702 12862 3736
rect 12928 3702 12962 3736
rect 13028 3702 13062 3736
rect 13128 3702 13162 3736
rect 13228 3702 13262 3736
rect 13328 3702 13362 3736
rect 12828 3608 12862 3636
rect 12828 3602 12834 3608
rect 12834 3602 12862 3608
rect 12928 3602 12962 3636
rect 13028 3602 13062 3636
rect 13128 3608 13162 3636
rect 13228 3608 13262 3636
rect 13328 3608 13362 3636
rect 13128 3602 13160 3608
rect 13160 3602 13162 3608
rect 13228 3602 13250 3608
rect 13250 3602 13262 3608
rect 13328 3602 13340 3608
rect 13340 3602 13362 3608
rect 14116 4114 14122 4136
rect 14122 4114 14150 4136
rect 14116 4102 14150 4114
rect 14216 4102 14250 4136
rect 14316 4102 14350 4136
rect 14416 4114 14448 4136
rect 14448 4114 14450 4136
rect 14516 4114 14538 4136
rect 14538 4114 14550 4136
rect 14616 4114 14628 4136
rect 14628 4114 14650 4136
rect 14416 4102 14450 4114
rect 14516 4102 14550 4114
rect 14616 4102 14650 4114
rect 14116 4024 14122 4036
rect 14122 4024 14150 4036
rect 14116 4002 14150 4024
rect 14216 4002 14250 4036
rect 14316 4002 14350 4036
rect 14416 4024 14448 4036
rect 14448 4024 14450 4036
rect 14516 4024 14538 4036
rect 14538 4024 14550 4036
rect 14616 4024 14628 4036
rect 14628 4024 14650 4036
rect 14416 4002 14450 4024
rect 14516 4002 14550 4024
rect 14616 4002 14650 4024
rect 14116 3934 14122 3936
rect 14122 3934 14150 3936
rect 14116 3902 14150 3934
rect 14216 3902 14250 3936
rect 14316 3902 14350 3936
rect 14416 3934 14448 3936
rect 14448 3934 14450 3936
rect 14516 3934 14538 3936
rect 14538 3934 14550 3936
rect 14616 3934 14628 3936
rect 14628 3934 14650 3936
rect 14416 3902 14450 3934
rect 14516 3902 14550 3934
rect 14616 3902 14650 3934
rect 14116 3802 14150 3836
rect 14216 3802 14250 3836
rect 14316 3802 14350 3836
rect 14416 3802 14450 3836
rect 14516 3802 14550 3836
rect 14616 3802 14650 3836
rect 14116 3702 14150 3736
rect 14216 3702 14250 3736
rect 14316 3702 14350 3736
rect 14416 3702 14450 3736
rect 14516 3702 14550 3736
rect 14616 3702 14650 3736
rect 14116 3608 14150 3636
rect 14116 3602 14122 3608
rect 14122 3602 14150 3608
rect 14216 3602 14250 3636
rect 14316 3602 14350 3636
rect 14416 3608 14450 3636
rect 14516 3608 14550 3636
rect 14616 3608 14650 3636
rect 14416 3602 14448 3608
rect 14448 3602 14450 3608
rect 14516 3602 14538 3608
rect 14538 3602 14550 3608
rect 14616 3602 14628 3608
rect 14628 3602 14650 3608
rect 15404 4114 15410 4136
rect 15410 4114 15438 4136
rect 15404 4102 15438 4114
rect 15504 4102 15538 4136
rect 15604 4102 15638 4136
rect 15704 4114 15736 4136
rect 15736 4114 15738 4136
rect 15804 4114 15826 4136
rect 15826 4114 15838 4136
rect 15904 4114 15916 4136
rect 15916 4114 15938 4136
rect 15704 4102 15738 4114
rect 15804 4102 15838 4114
rect 15904 4102 15938 4114
rect 15404 4024 15410 4036
rect 15410 4024 15438 4036
rect 15404 4002 15438 4024
rect 15504 4002 15538 4036
rect 15604 4002 15638 4036
rect 15704 4024 15736 4036
rect 15736 4024 15738 4036
rect 15804 4024 15826 4036
rect 15826 4024 15838 4036
rect 15904 4024 15916 4036
rect 15916 4024 15938 4036
rect 15704 4002 15738 4024
rect 15804 4002 15838 4024
rect 15904 4002 15938 4024
rect 15404 3934 15410 3936
rect 15410 3934 15438 3936
rect 15404 3902 15438 3934
rect 15504 3902 15538 3936
rect 15604 3902 15638 3936
rect 15704 3934 15736 3936
rect 15736 3934 15738 3936
rect 15804 3934 15826 3936
rect 15826 3934 15838 3936
rect 15904 3934 15916 3936
rect 15916 3934 15938 3936
rect 15704 3902 15738 3934
rect 15804 3902 15838 3934
rect 15904 3902 15938 3934
rect 15404 3802 15438 3836
rect 15504 3802 15538 3836
rect 15604 3802 15638 3836
rect 15704 3802 15738 3836
rect 15804 3802 15838 3836
rect 15904 3802 15938 3836
rect 15404 3702 15438 3736
rect 15504 3702 15538 3736
rect 15604 3702 15638 3736
rect 15704 3702 15738 3736
rect 15804 3702 15838 3736
rect 15904 3702 15938 3736
rect 15404 3608 15438 3636
rect 15404 3602 15410 3608
rect 15410 3602 15438 3608
rect 15504 3602 15538 3636
rect 15604 3602 15638 3636
rect 15704 3608 15738 3636
rect 15804 3608 15838 3636
rect 15904 3608 15938 3636
rect 15704 3602 15736 3608
rect 15736 3602 15738 3608
rect 15804 3602 15826 3608
rect 15826 3602 15838 3608
rect 15904 3602 15916 3608
rect 15916 3602 15938 3608
rect 16692 4114 16698 4136
rect 16698 4114 16726 4136
rect 16692 4102 16726 4114
rect 16792 4102 16826 4136
rect 16892 4102 16926 4136
rect 16992 4114 17024 4136
rect 17024 4114 17026 4136
rect 17092 4114 17114 4136
rect 17114 4114 17126 4136
rect 17192 4114 17204 4136
rect 17204 4114 17226 4136
rect 16992 4102 17026 4114
rect 17092 4102 17126 4114
rect 17192 4102 17226 4114
rect 16692 4024 16698 4036
rect 16698 4024 16726 4036
rect 16692 4002 16726 4024
rect 16792 4002 16826 4036
rect 16892 4002 16926 4036
rect 16992 4024 17024 4036
rect 17024 4024 17026 4036
rect 17092 4024 17114 4036
rect 17114 4024 17126 4036
rect 17192 4024 17204 4036
rect 17204 4024 17226 4036
rect 16992 4002 17026 4024
rect 17092 4002 17126 4024
rect 17192 4002 17226 4024
rect 16692 3934 16698 3936
rect 16698 3934 16726 3936
rect 16692 3902 16726 3934
rect 16792 3902 16826 3936
rect 16892 3902 16926 3936
rect 16992 3934 17024 3936
rect 17024 3934 17026 3936
rect 17092 3934 17114 3936
rect 17114 3934 17126 3936
rect 17192 3934 17204 3936
rect 17204 3934 17226 3936
rect 16992 3902 17026 3934
rect 17092 3902 17126 3934
rect 17192 3902 17226 3934
rect 16692 3802 16726 3836
rect 16792 3802 16826 3836
rect 16892 3802 16926 3836
rect 16992 3802 17026 3836
rect 17092 3802 17126 3836
rect 17192 3802 17226 3836
rect 16692 3702 16726 3736
rect 16792 3702 16826 3736
rect 16892 3702 16926 3736
rect 16992 3702 17026 3736
rect 17092 3702 17126 3736
rect 17192 3702 17226 3736
rect 16692 3608 16726 3636
rect 16692 3602 16698 3608
rect 16698 3602 16726 3608
rect 16792 3602 16826 3636
rect 16892 3602 16926 3636
rect 16992 3608 17026 3636
rect 17092 3608 17126 3636
rect 17192 3608 17226 3636
rect 16992 3602 17024 3608
rect 17024 3602 17026 3608
rect 17092 3602 17114 3608
rect 17114 3602 17126 3608
rect 17192 3602 17204 3608
rect 17204 3602 17226 3608
rect 17980 4114 17986 4136
rect 17986 4114 18014 4136
rect 17980 4102 18014 4114
rect 18080 4102 18114 4136
rect 18180 4102 18214 4136
rect 18280 4114 18312 4136
rect 18312 4114 18314 4136
rect 18380 4114 18402 4136
rect 18402 4114 18414 4136
rect 18480 4114 18492 4136
rect 18492 4114 18514 4136
rect 18280 4102 18314 4114
rect 18380 4102 18414 4114
rect 18480 4102 18514 4114
rect 17980 4024 17986 4036
rect 17986 4024 18014 4036
rect 17980 4002 18014 4024
rect 18080 4002 18114 4036
rect 18180 4002 18214 4036
rect 18280 4024 18312 4036
rect 18312 4024 18314 4036
rect 18380 4024 18402 4036
rect 18402 4024 18414 4036
rect 18480 4024 18492 4036
rect 18492 4024 18514 4036
rect 18280 4002 18314 4024
rect 18380 4002 18414 4024
rect 18480 4002 18514 4024
rect 17980 3934 17986 3936
rect 17986 3934 18014 3936
rect 17980 3902 18014 3934
rect 18080 3902 18114 3936
rect 18180 3902 18214 3936
rect 18280 3934 18312 3936
rect 18312 3934 18314 3936
rect 18380 3934 18402 3936
rect 18402 3934 18414 3936
rect 18480 3934 18492 3936
rect 18492 3934 18514 3936
rect 18280 3902 18314 3934
rect 18380 3902 18414 3934
rect 18480 3902 18514 3934
rect 17980 3802 18014 3836
rect 18080 3802 18114 3836
rect 18180 3802 18214 3836
rect 18280 3802 18314 3836
rect 18380 3802 18414 3836
rect 18480 3802 18514 3836
rect 17980 3702 18014 3736
rect 18080 3702 18114 3736
rect 18180 3702 18214 3736
rect 18280 3702 18314 3736
rect 18380 3702 18414 3736
rect 18480 3702 18514 3736
rect 17980 3608 18014 3636
rect 17980 3602 17986 3608
rect 17986 3602 18014 3608
rect 18080 3602 18114 3636
rect 18180 3602 18214 3636
rect 18280 3608 18314 3636
rect 18380 3608 18414 3636
rect 18480 3608 18514 3636
rect 18280 3602 18312 3608
rect 18312 3602 18314 3608
rect 18380 3602 18402 3608
rect 18402 3602 18414 3608
rect 18480 3602 18492 3608
rect 18492 3602 18514 3608
rect 12828 2826 12834 2848
rect 12834 2826 12862 2848
rect 12828 2814 12862 2826
rect 12928 2814 12962 2848
rect 13028 2814 13062 2848
rect 13128 2826 13160 2848
rect 13160 2826 13162 2848
rect 13228 2826 13250 2848
rect 13250 2826 13262 2848
rect 13328 2826 13340 2848
rect 13340 2826 13362 2848
rect 13128 2814 13162 2826
rect 13228 2814 13262 2826
rect 13328 2814 13362 2826
rect 12828 2736 12834 2748
rect 12834 2736 12862 2748
rect 12828 2714 12862 2736
rect 12928 2714 12962 2748
rect 13028 2714 13062 2748
rect 13128 2736 13160 2748
rect 13160 2736 13162 2748
rect 13228 2736 13250 2748
rect 13250 2736 13262 2748
rect 13328 2736 13340 2748
rect 13340 2736 13362 2748
rect 13128 2714 13162 2736
rect 13228 2714 13262 2736
rect 13328 2714 13362 2736
rect 12828 2646 12834 2648
rect 12834 2646 12862 2648
rect 12828 2614 12862 2646
rect 12928 2614 12962 2648
rect 13028 2614 13062 2648
rect 13128 2646 13160 2648
rect 13160 2646 13162 2648
rect 13228 2646 13250 2648
rect 13250 2646 13262 2648
rect 13328 2646 13340 2648
rect 13340 2646 13362 2648
rect 13128 2614 13162 2646
rect 13228 2614 13262 2646
rect 13328 2614 13362 2646
rect 12828 2514 12862 2548
rect 12928 2514 12962 2548
rect 13028 2514 13062 2548
rect 13128 2514 13162 2548
rect 13228 2514 13262 2548
rect 13328 2514 13362 2548
rect 12828 2414 12862 2448
rect 12928 2414 12962 2448
rect 13028 2414 13062 2448
rect 13128 2414 13162 2448
rect 13228 2414 13262 2448
rect 13328 2414 13362 2448
rect 12828 2320 12862 2348
rect 12828 2314 12834 2320
rect 12834 2314 12862 2320
rect 12928 2314 12962 2348
rect 13028 2314 13062 2348
rect 13128 2320 13162 2348
rect 13228 2320 13262 2348
rect 13328 2320 13362 2348
rect 13128 2314 13160 2320
rect 13160 2314 13162 2320
rect 13228 2314 13250 2320
rect 13250 2314 13262 2320
rect 13328 2314 13340 2320
rect 13340 2314 13362 2320
rect 14116 2826 14122 2848
rect 14122 2826 14150 2848
rect 14116 2814 14150 2826
rect 14216 2814 14250 2848
rect 14316 2814 14350 2848
rect 14416 2826 14448 2848
rect 14448 2826 14450 2848
rect 14516 2826 14538 2848
rect 14538 2826 14550 2848
rect 14616 2826 14628 2848
rect 14628 2826 14650 2848
rect 14416 2814 14450 2826
rect 14516 2814 14550 2826
rect 14616 2814 14650 2826
rect 14116 2736 14122 2748
rect 14122 2736 14150 2748
rect 14116 2714 14150 2736
rect 14216 2714 14250 2748
rect 14316 2714 14350 2748
rect 14416 2736 14448 2748
rect 14448 2736 14450 2748
rect 14516 2736 14538 2748
rect 14538 2736 14550 2748
rect 14616 2736 14628 2748
rect 14628 2736 14650 2748
rect 14416 2714 14450 2736
rect 14516 2714 14550 2736
rect 14616 2714 14650 2736
rect 14116 2646 14122 2648
rect 14122 2646 14150 2648
rect 14116 2614 14150 2646
rect 14216 2614 14250 2648
rect 14316 2614 14350 2648
rect 14416 2646 14448 2648
rect 14448 2646 14450 2648
rect 14516 2646 14538 2648
rect 14538 2646 14550 2648
rect 14616 2646 14628 2648
rect 14628 2646 14650 2648
rect 14416 2614 14450 2646
rect 14516 2614 14550 2646
rect 14616 2614 14650 2646
rect 14116 2514 14150 2548
rect 14216 2514 14250 2548
rect 14316 2514 14350 2548
rect 14416 2514 14450 2548
rect 14516 2514 14550 2548
rect 14616 2514 14650 2548
rect 14116 2414 14150 2448
rect 14216 2414 14250 2448
rect 14316 2414 14350 2448
rect 14416 2414 14450 2448
rect 14516 2414 14550 2448
rect 14616 2414 14650 2448
rect 14116 2320 14150 2348
rect 14116 2314 14122 2320
rect 14122 2314 14150 2320
rect 14216 2314 14250 2348
rect 14316 2314 14350 2348
rect 14416 2320 14450 2348
rect 14516 2320 14550 2348
rect 14616 2320 14650 2348
rect 14416 2314 14448 2320
rect 14448 2314 14450 2320
rect 14516 2314 14538 2320
rect 14538 2314 14550 2320
rect 14616 2314 14628 2320
rect 14628 2314 14650 2320
rect 15404 2826 15410 2848
rect 15410 2826 15438 2848
rect 15404 2814 15438 2826
rect 15504 2814 15538 2848
rect 15604 2814 15638 2848
rect 15704 2826 15736 2848
rect 15736 2826 15738 2848
rect 15804 2826 15826 2848
rect 15826 2826 15838 2848
rect 15904 2826 15916 2848
rect 15916 2826 15938 2848
rect 15704 2814 15738 2826
rect 15804 2814 15838 2826
rect 15904 2814 15938 2826
rect 15404 2736 15410 2748
rect 15410 2736 15438 2748
rect 15404 2714 15438 2736
rect 15504 2714 15538 2748
rect 15604 2714 15638 2748
rect 15704 2736 15736 2748
rect 15736 2736 15738 2748
rect 15804 2736 15826 2748
rect 15826 2736 15838 2748
rect 15904 2736 15916 2748
rect 15916 2736 15938 2748
rect 15704 2714 15738 2736
rect 15804 2714 15838 2736
rect 15904 2714 15938 2736
rect 15404 2646 15410 2648
rect 15410 2646 15438 2648
rect 15404 2614 15438 2646
rect 15504 2614 15538 2648
rect 15604 2614 15638 2648
rect 15704 2646 15736 2648
rect 15736 2646 15738 2648
rect 15804 2646 15826 2648
rect 15826 2646 15838 2648
rect 15904 2646 15916 2648
rect 15916 2646 15938 2648
rect 15704 2614 15738 2646
rect 15804 2614 15838 2646
rect 15904 2614 15938 2646
rect 15404 2514 15438 2548
rect 15504 2514 15538 2548
rect 15604 2514 15638 2548
rect 15704 2514 15738 2548
rect 15804 2514 15838 2548
rect 15904 2514 15938 2548
rect 15404 2414 15438 2448
rect 15504 2414 15538 2448
rect 15604 2414 15638 2448
rect 15704 2414 15738 2448
rect 15804 2414 15838 2448
rect 15904 2414 15938 2448
rect 15404 2320 15438 2348
rect 15404 2314 15410 2320
rect 15410 2314 15438 2320
rect 15504 2314 15538 2348
rect 15604 2314 15638 2348
rect 15704 2320 15738 2348
rect 15804 2320 15838 2348
rect 15904 2320 15938 2348
rect 15704 2314 15736 2320
rect 15736 2314 15738 2320
rect 15804 2314 15826 2320
rect 15826 2314 15838 2320
rect 15904 2314 15916 2320
rect 15916 2314 15938 2320
rect 16692 2826 16698 2848
rect 16698 2826 16726 2848
rect 16692 2814 16726 2826
rect 16792 2814 16826 2848
rect 16892 2814 16926 2848
rect 16992 2826 17024 2848
rect 17024 2826 17026 2848
rect 17092 2826 17114 2848
rect 17114 2826 17126 2848
rect 17192 2826 17204 2848
rect 17204 2826 17226 2848
rect 16992 2814 17026 2826
rect 17092 2814 17126 2826
rect 17192 2814 17226 2826
rect 16692 2736 16698 2748
rect 16698 2736 16726 2748
rect 16692 2714 16726 2736
rect 16792 2714 16826 2748
rect 16892 2714 16926 2748
rect 16992 2736 17024 2748
rect 17024 2736 17026 2748
rect 17092 2736 17114 2748
rect 17114 2736 17126 2748
rect 17192 2736 17204 2748
rect 17204 2736 17226 2748
rect 16992 2714 17026 2736
rect 17092 2714 17126 2736
rect 17192 2714 17226 2736
rect 16692 2646 16698 2648
rect 16698 2646 16726 2648
rect 16692 2614 16726 2646
rect 16792 2614 16826 2648
rect 16892 2614 16926 2648
rect 16992 2646 17024 2648
rect 17024 2646 17026 2648
rect 17092 2646 17114 2648
rect 17114 2646 17126 2648
rect 17192 2646 17204 2648
rect 17204 2646 17226 2648
rect 16992 2614 17026 2646
rect 17092 2614 17126 2646
rect 17192 2614 17226 2646
rect 16692 2514 16726 2548
rect 16792 2514 16826 2548
rect 16892 2514 16926 2548
rect 16992 2514 17026 2548
rect 17092 2514 17126 2548
rect 17192 2514 17226 2548
rect 16692 2414 16726 2448
rect 16792 2414 16826 2448
rect 16892 2414 16926 2448
rect 16992 2414 17026 2448
rect 17092 2414 17126 2448
rect 17192 2414 17226 2448
rect 16692 2320 16726 2348
rect 16692 2314 16698 2320
rect 16698 2314 16726 2320
rect 16792 2314 16826 2348
rect 16892 2314 16926 2348
rect 16992 2320 17026 2348
rect 17092 2320 17126 2348
rect 17192 2320 17226 2348
rect 16992 2314 17024 2320
rect 17024 2314 17026 2320
rect 17092 2314 17114 2320
rect 17114 2314 17126 2320
rect 17192 2314 17204 2320
rect 17204 2314 17226 2320
rect 17980 2826 17986 2848
rect 17986 2826 18014 2848
rect 17980 2814 18014 2826
rect 18080 2814 18114 2848
rect 18180 2814 18214 2848
rect 18280 2826 18312 2848
rect 18312 2826 18314 2848
rect 18380 2826 18402 2848
rect 18402 2826 18414 2848
rect 18480 2826 18492 2848
rect 18492 2826 18514 2848
rect 18280 2814 18314 2826
rect 18380 2814 18414 2826
rect 18480 2814 18514 2826
rect 17980 2736 17986 2748
rect 17986 2736 18014 2748
rect 17980 2714 18014 2736
rect 18080 2714 18114 2748
rect 18180 2714 18214 2748
rect 18280 2736 18312 2748
rect 18312 2736 18314 2748
rect 18380 2736 18402 2748
rect 18402 2736 18414 2748
rect 18480 2736 18492 2748
rect 18492 2736 18514 2748
rect 18280 2714 18314 2736
rect 18380 2714 18414 2736
rect 18480 2714 18514 2736
rect 17980 2646 17986 2648
rect 17986 2646 18014 2648
rect 17980 2614 18014 2646
rect 18080 2614 18114 2648
rect 18180 2614 18214 2648
rect 18280 2646 18312 2648
rect 18312 2646 18314 2648
rect 18380 2646 18402 2648
rect 18402 2646 18414 2648
rect 18480 2646 18492 2648
rect 18492 2646 18514 2648
rect 18280 2614 18314 2646
rect 18380 2614 18414 2646
rect 18480 2614 18514 2646
rect 17980 2514 18014 2548
rect 18080 2514 18114 2548
rect 18180 2514 18214 2548
rect 18280 2514 18314 2548
rect 18380 2514 18414 2548
rect 18480 2514 18514 2548
rect 17980 2414 18014 2448
rect 18080 2414 18114 2448
rect 18180 2414 18214 2448
rect 18280 2414 18314 2448
rect 18380 2414 18414 2448
rect 18480 2414 18514 2448
rect 17980 2320 18014 2348
rect 17980 2314 17986 2320
rect 17986 2314 18014 2320
rect 18080 2314 18114 2348
rect 18180 2314 18214 2348
rect 18280 2320 18314 2348
rect 18380 2320 18414 2348
rect 18480 2320 18514 2348
rect 18280 2314 18312 2320
rect 18312 2314 18314 2320
rect 18380 2314 18402 2320
rect 18402 2314 18414 2320
rect 18480 2314 18492 2320
rect 18492 2314 18514 2320
rect 7966 1100 8366 1200
<< metal1 >>
rect -21552 25066 -10296 25072
rect -21552 24240 -21546 25066
rect -10302 24240 -10296 25066
rect -21552 24234 -10296 24240
rect 1714 23526 3908 23532
rect 1714 22968 1720 23526
rect 2278 22968 3344 23526
rect 3902 22968 3908 23526
rect 1714 22962 3908 22968
rect 7260 23526 10458 23532
rect 7260 22968 7434 23526
rect 7992 22968 9888 23526
rect 10446 22968 10458 23526
rect 7260 22962 10458 22968
rect -4842 22732 -4150 22734
rect -4842 22726 1454 22732
rect -4842 22168 890 22726
rect 1448 22168 1454 22726
rect -4842 22162 1454 22168
rect 4034 22726 7180 22732
rect 4034 22168 4162 22726
rect 4720 22168 6616 22726
rect 7174 22168 7180 22726
rect 4034 22162 7180 22168
rect 8950 22726 12088 22732
rect 8950 22168 9070 22726
rect 9628 22168 11524 22726
rect 12082 22168 12088 22726
rect 8950 22162 12088 22168
rect -5656 21976 -5094 21982
rect -5656 21579 -5644 21976
rect -5106 21579 -5094 21976
rect -5656 21573 -5094 21579
rect -4842 21976 -4272 22162
rect -4842 21579 -4826 21976
rect -4288 21579 -4272 21976
rect -4842 21562 -4272 21579
rect -4024 21976 -3452 21994
rect -4024 21579 -4008 21976
rect -3470 21579 -3452 21976
rect -4024 21270 -3452 21579
rect -3202 21976 -2640 21982
rect -3202 21579 -3190 21976
rect -2652 21579 -2640 21976
rect 66 21926 636 21932
rect -3202 21573 -2640 21579
rect -748 21914 -186 21920
rect -748 21517 -736 21914
rect -198 21517 -186 21914
rect -748 21511 -186 21517
rect 66 21506 72 21926
rect 630 21506 636 21926
rect 66 21500 636 21506
rect 884 21926 1454 21932
rect 884 21506 890 21926
rect 1448 21506 1454 21926
rect 884 21500 1454 21506
rect 1702 21926 2272 21932
rect 1702 21506 1708 21926
rect 2266 21506 2272 21926
rect 1702 21500 2272 21506
rect 2520 21926 3090 21932
rect 2520 21506 2526 21926
rect 3084 21506 3090 21926
rect 2520 21500 3090 21506
rect 3338 21926 3908 21932
rect 3338 21506 3344 21926
rect 3902 21506 3908 21926
rect 3338 21500 3908 21506
rect 4156 21926 4726 21932
rect 4156 21506 4162 21926
rect 4720 21506 4726 21926
rect 4156 21500 4726 21506
rect 4974 21926 5544 21932
rect 4974 21506 4980 21926
rect 5538 21506 5544 21926
rect 4974 21500 5544 21506
rect 5792 21926 6362 21932
rect 5792 21506 5798 21926
rect 6356 21506 6362 21926
rect 5792 21500 6362 21506
rect 6610 21926 7180 21932
rect 6610 21506 6616 21926
rect 7174 21506 7180 21926
rect 6610 21500 7180 21506
rect 7428 21926 7998 21932
rect 7428 21506 7434 21926
rect 7992 21506 7998 21926
rect 7428 21500 7998 21506
rect 8246 21926 8816 21932
rect 8246 21506 8252 21926
rect 8810 21506 8816 21926
rect 8246 21500 8816 21506
rect 9064 21926 9634 21932
rect 9064 21506 9070 21926
rect 9628 21506 9634 21926
rect 9064 21500 9634 21506
rect 9882 21926 10452 21932
rect 9882 21506 9888 21926
rect 10446 21506 10452 21926
rect 9882 21500 10452 21506
rect 10700 21926 11270 21932
rect 10700 21506 10706 21926
rect 11264 21506 11270 21926
rect 10700 21500 11270 21506
rect 11518 21926 12088 21932
rect 11518 21506 11524 21926
rect 12082 21506 12088 21926
rect 12340 21914 12902 21920
rect 12340 21517 12352 21914
rect 12890 21517 12902 21914
rect 12340 21511 12902 21517
rect 11518 21500 12088 21506
rect -4024 21264 636 21270
rect -4024 20706 72 21264
rect 630 20706 636 21264
rect -4024 20700 636 20706
rect 2520 21264 5544 21270
rect 2520 20706 2526 21264
rect 3084 20706 4980 21264
rect 5538 20706 5544 21264
rect 2520 20700 5544 20706
rect 8246 21264 11270 21270
rect 8246 20706 8252 21264
rect 8810 20706 10706 21264
rect 11264 20706 11270 21264
rect 8246 20700 11270 20706
rect -8928 20590 -8366 20596
rect -8928 20193 -8916 20590
rect -8378 20193 -8366 20590
rect -8928 20187 -8366 20193
rect -8110 20590 -7548 20596
rect -8110 20193 -8098 20590
rect -7560 20193 -7548 20590
rect -8110 20187 -7548 20193
rect -7292 20590 -6730 20596
rect -7292 20193 -7280 20590
rect -6742 20193 -6730 20590
rect -7292 20187 -6730 20193
rect -5656 17245 -5094 17251
rect -5656 16848 -5644 17245
rect -5106 16848 -5094 17245
rect -5656 16842 -5094 16848
rect -4838 17245 -4276 17251
rect -4838 16848 -4826 17245
rect -4288 16848 -4276 17245
rect -4838 16842 -4276 16848
rect -4020 17245 -3458 17251
rect -4020 16848 -4008 17245
rect -3470 16848 -3458 17245
rect -4020 16842 -3458 16848
rect -3202 17245 -2640 17251
rect -3202 16848 -3190 17245
rect -2652 16848 -2640 17245
rect -3202 16842 -2640 16848
rect -8928 16835 -8366 16841
rect -8928 16438 -8916 16835
rect -8378 16438 -8366 16835
rect -8928 16432 -8366 16438
rect -8110 16835 -7548 16841
rect -8110 16438 -8098 16835
rect -7560 16438 -7548 16835
rect -8110 16432 -7548 16438
rect -7292 16835 -6730 16841
rect -7292 16438 -7280 16835
rect -6742 16438 -6730 16835
rect -7292 16432 -6730 16438
rect 884 16790 4726 16796
rect -8104 15996 -7556 16432
rect 884 16232 890 16790
rect 1448 16232 4162 16790
rect 4720 16232 4726 16790
rect 884 16226 4726 16232
rect 6616 16790 9634 16796
rect 7174 16232 9070 16790
rect 9628 16232 9634 16790
rect 6616 16226 9634 16232
rect -8104 15990 2272 15996
rect -8104 15432 1708 15990
rect 2266 15432 2272 15990
rect -8104 15426 2272 15432
rect 3338 15990 7998 15996
rect 3338 15432 3344 15990
rect 3902 15432 7434 15990
rect 7992 15432 7998 15990
rect 3338 15426 7998 15432
rect 66 15190 636 15196
rect -748 15179 -186 15185
rect -748 14782 -736 15179
rect -198 14782 -186 15179
rect -748 14776 -186 14782
rect 66 14770 72 15190
rect 630 14770 636 15190
rect 66 14764 636 14770
rect 884 15190 1454 15196
rect 884 14770 890 15190
rect 1448 14770 1454 15190
rect 884 14764 1454 14770
rect 1702 15190 2272 15196
rect 1702 14770 1708 15190
rect 2266 14770 2272 15190
rect 1702 14764 2272 14770
rect 2520 15190 3090 15196
rect 2520 14770 2526 15190
rect 3084 14770 3090 15190
rect 2520 14764 3090 14770
rect 3338 15190 3908 15196
rect 3338 14770 3344 15190
rect 3902 14770 3908 15190
rect 3338 14764 3908 14770
rect 4156 15190 4726 15196
rect 4156 14770 4162 15190
rect 4720 14770 4726 15190
rect 4156 14764 4726 14770
rect 4974 15190 5544 15196
rect 4974 14770 4980 15190
rect 5538 14770 5544 15190
rect 4974 14764 5544 14770
rect 5714 15190 6418 15196
rect 5714 15158 5798 15190
rect 5714 14640 5720 15158
rect 6356 15158 6418 15190
rect 6412 14640 6418 15158
rect 6610 15190 7180 15196
rect 6610 14770 6616 15190
rect 7174 14770 7180 15190
rect 6610 14764 7180 14770
rect 7428 15190 7998 15196
rect 7428 14770 7434 15190
rect 7992 14770 7998 15190
rect 7428 14764 7998 14770
rect 8246 15190 8816 15196
rect 8246 14770 8252 15190
rect 8810 14770 8816 15190
rect 8246 14764 8816 14770
rect 9064 15190 9634 15196
rect 9064 14770 9070 15190
rect 9628 14770 9634 15190
rect 9064 14764 9634 14770
rect 9804 15190 10508 15196
rect 66 14528 3090 14534
rect 66 13970 72 14528
rect 630 13970 2526 14528
rect 3084 13970 3090 14528
rect 66 13964 3090 13970
rect 4974 14528 8816 14534
rect 4974 13970 4980 14528
rect 5538 13970 8252 14528
rect 8810 13970 8816 14528
rect 4974 13964 8816 13970
rect 9804 14498 9810 15190
rect 10502 14498 10508 15190
rect 9804 13500 10508 14498
rect -2890 12808 10508 13500
rect 10622 15190 11326 15196
rect 10622 14498 10628 15190
rect 11320 14498 11326 15190
rect -8390 11860 -6390 11902
rect -8390 11410 -8384 11860
rect -6396 11410 -6390 11860
rect -9908 11104 -9776 11110
rect -9908 10690 -9902 11104
rect -9782 10690 -9776 11104
rect -10364 10398 -10232 10684
rect -10364 10106 -10358 10398
rect -10238 10106 -10232 10398
rect -17900 9388 -11412 9400
rect -17900 9044 -17888 9388
rect -11424 9044 -11412 9388
rect -17900 8852 -11412 9044
rect -17900 8832 -17164 8852
rect -17176 8818 -17164 8832
rect -11788 8832 -11412 8852
rect -11788 8818 -11776 8832
rect -17176 8812 -11776 8818
rect -19254 8698 -17208 8710
rect -19254 8514 -17248 8698
rect -17214 8514 -17208 8698
rect -19254 8502 -17208 8514
rect -17176 8394 -11776 8400
rect -17894 8360 -17164 8394
rect -11788 8360 -11418 8394
rect -17894 8038 -11418 8360
rect -20918 5720 -20842 5732
rect -20918 5668 -20906 5720
rect -20854 5668 -20842 5720
rect -20918 5656 -20842 5668
rect -20002 5720 -19926 5732
rect -20002 5668 -19990 5720
rect -19938 5668 -19926 5720
rect -20002 5656 -19926 5668
rect -21670 5604 -21462 5610
rect -21224 5604 -20992 5616
rect -21670 5570 -21658 5604
rect -21474 5570 -21462 5604
rect -21670 5564 -21462 5570
rect -21360 5570 -21200 5604
rect -21016 5570 -20992 5604
rect -21360 5532 -21316 5570
rect -21224 5552 -20992 5570
rect -21818 5520 -21772 5532
rect -21818 5144 -21812 5520
rect -21778 5144 -21772 5520
rect -21818 5132 -21772 5144
rect -21360 5520 -21314 5532
rect -21360 5144 -21354 5520
rect -21320 5144 -21314 5520
rect -21360 5002 -21314 5144
rect -20902 5520 -20856 5656
rect -20754 5604 -20546 5610
rect -20754 5570 -20742 5604
rect -20558 5570 -20546 5604
rect -20754 5564 -20546 5570
rect -20296 5604 -20088 5610
rect -20296 5570 -20284 5604
rect -20100 5570 -20088 5604
rect -20296 5564 -20088 5570
rect -20902 5144 -20896 5520
rect -20862 5144 -20856 5520
rect -20902 5132 -20856 5144
rect -20444 5520 -20398 5532
rect -20444 5144 -20438 5520
rect -20404 5144 -20398 5520
rect -21370 4996 -21306 5002
rect -21370 4944 -21364 4996
rect -21312 4944 -21306 4996
rect -21370 4938 -21306 4944
rect -20444 4796 -20398 5144
rect -19986 5520 -19940 5656
rect -19860 5604 -19628 5616
rect -19380 5604 -19172 5610
rect -19860 5570 -19826 5604
rect -19642 5570 -19482 5604
rect -19860 5552 -19628 5570
rect -19986 5144 -19980 5520
rect -19946 5144 -19940 5520
rect -19986 5132 -19940 5144
rect -19528 5520 -19482 5570
rect -19380 5570 -19368 5604
rect -19184 5570 -19172 5604
rect -19380 5564 -19172 5570
rect -19528 5144 -19522 5520
rect -19488 5144 -19482 5520
rect -19528 5008 -19482 5144
rect -19070 5520 -19024 5532
rect -19070 5144 -19064 5520
rect -19030 5144 -19024 5520
rect -19070 5132 -19024 5144
rect -19536 5002 -19472 5008
rect -19536 4950 -19530 5002
rect -19478 4950 -19472 5002
rect -19536 4944 -19472 4950
rect -18930 5002 -18724 5008
rect -18930 4944 -18924 5002
rect -18730 4944 -18724 5002
rect -20452 4790 -20388 4796
rect -20452 4738 -20446 4790
rect -20394 4738 -20388 4790
rect -20452 4732 -20388 4738
rect -19266 4142 -19134 4154
rect -19266 1800 -19250 4142
rect -19150 1800 -19134 4142
rect -19266 1552 -19134 1800
rect -19266 1448 -19240 1552
rect -19188 1448 -19134 1552
rect -19266 1438 -19134 1448
rect -18930 1358 -18724 4944
rect -17894 4630 -17686 8038
rect -15584 6986 -15400 7006
rect -15584 6932 -15564 6986
rect -15420 6932 -15400 6986
rect -16156 6846 -15972 6866
rect -16156 6792 -16136 6846
rect -15992 6792 -15972 6846
rect -16156 6732 -15972 6792
rect -15584 6732 -15400 6932
rect -14440 6986 -14256 7006
rect -14440 6932 -14420 6986
rect -14276 6932 -14256 6986
rect -15012 6846 -14828 6866
rect -15012 6792 -14992 6846
rect -14848 6792 -14828 6846
rect -15012 6732 -14828 6792
rect -14440 6732 -14256 6932
rect -13296 6986 -13112 7006
rect -13296 6932 -13276 6986
rect -13132 6932 -13112 6986
rect -13868 6846 -13684 6866
rect -13868 6792 -13848 6846
rect -13704 6792 -13684 6846
rect -13868 6732 -13684 6792
rect -13296 6732 -13112 6932
rect -17440 6726 -16384 6732
rect -17440 6692 -16728 6726
rect -16544 6692 -16384 6726
rect -17440 6686 -16384 6692
rect -16168 6726 -15960 6732
rect -16168 6692 -16156 6726
rect -15972 6692 -15960 6726
rect -16168 6686 -15960 6692
rect -15596 6726 -15388 6732
rect -15596 6692 -15584 6726
rect -15400 6692 -15388 6726
rect -15596 6686 -15388 6692
rect -15024 6726 -14816 6732
rect -15024 6692 -15012 6726
rect -14828 6692 -14816 6726
rect -15024 6686 -14816 6692
rect -14452 6726 -14244 6732
rect -14452 6692 -14440 6726
rect -14256 6692 -14244 6726
rect -14452 6686 -14244 6692
rect -13880 6726 -13672 6732
rect -13880 6692 -13868 6726
rect -13684 6692 -13672 6726
rect -13880 6686 -13672 6692
rect -13308 6726 -13100 6732
rect -13308 6692 -13296 6726
rect -13112 6692 -13100 6726
rect -13308 6686 -13100 6692
rect -12884 6726 -11828 6732
rect -12884 6692 -12724 6726
rect -12540 6692 -11828 6726
rect -12884 6686 -11828 6692
rect -17440 6658 -17326 6686
rect -17450 6642 -17318 6658
rect -17450 5044 -17434 6642
rect -17334 5044 -17318 6642
rect -17450 5026 -17318 5044
rect -16888 6642 -16842 6686
rect -16888 4866 -16882 6642
rect -16848 4866 -16842 6642
rect -16888 4854 -16842 4866
rect -16430 6642 -16384 6686
rect -16430 4866 -16424 6642
rect -16390 4866 -16384 6642
rect -16430 4854 -16384 4866
rect -16316 6642 -16270 6654
rect -16316 4866 -16310 6642
rect -16276 4866 -16270 6642
rect -16316 4854 -16270 4866
rect -15858 6642 -15812 6654
rect -15858 4866 -15852 6642
rect -15818 4866 -15812 6642
rect -15858 4854 -15812 4866
rect -15744 6642 -15698 6654
rect -15744 4866 -15738 6642
rect -15704 4866 -15698 6642
rect -15744 4854 -15698 4866
rect -15286 6642 -15240 6654
rect -15286 4866 -15280 6642
rect -15246 4866 -15240 6642
rect -15286 4854 -15240 4866
rect -15172 6642 -15126 6654
rect -15172 4866 -15166 6642
rect -15132 4866 -15126 6642
rect -15172 4854 -15126 4866
rect -14714 6642 -14668 6654
rect -14714 4866 -14708 6642
rect -14674 4866 -14668 6642
rect -14714 4854 -14668 4866
rect -14600 6642 -14554 6654
rect -14600 4866 -14594 6642
rect -14560 4866 -14554 6642
rect -14600 4854 -14554 4866
rect -14142 6642 -14096 6654
rect -14142 4866 -14136 6642
rect -14102 4866 -14096 6642
rect -14142 4854 -14096 4866
rect -14028 6642 -13982 6654
rect -14028 4866 -14022 6642
rect -13988 4866 -13982 6642
rect -14028 4854 -13982 4866
rect -13570 6642 -13524 6654
rect -13570 4866 -13564 6642
rect -13530 4866 -13524 6642
rect -13570 4854 -13524 4866
rect -13456 6642 -13410 6654
rect -13456 4866 -13450 6642
rect -13416 4866 -13410 6642
rect -13456 4854 -13410 4866
rect -12998 6642 -12952 6654
rect -12998 4866 -12992 6642
rect -12958 4866 -12952 6642
rect -12998 4854 -12952 4866
rect -12884 6642 -12838 6686
rect -12884 4866 -12878 6642
rect -12844 4866 -12838 6642
rect -12884 4854 -12838 4866
rect -12426 6642 -12380 6686
rect -11942 6658 -11828 6686
rect -12426 4866 -12420 6642
rect -12386 4866 -12380 6642
rect -11950 6642 -11818 6658
rect -11950 5044 -11934 6642
rect -11834 5044 -11818 6642
rect -11950 5026 -11818 5044
rect -12426 4854 -12380 4866
rect -17894 4376 -17768 4630
rect -17716 4376 -17686 4630
rect -18614 4323 -18110 4330
rect -18614 4289 -18454 4323
rect -18270 4289 -18110 4323
rect -18614 4282 -18110 4289
rect -17894 4323 -17686 4376
rect -17894 4289 -17882 4323
rect -17698 4289 -17686 4323
rect -17894 4282 -17686 4289
rect -17334 4630 -17126 4636
rect -17334 4376 -17208 4630
rect -17156 4376 -17126 4630
rect -17334 4329 -17126 4376
rect -16774 4630 -16566 4636
rect -16774 4376 -16648 4630
rect -16596 4376 -16566 4630
rect -16774 4329 -16566 4376
rect -17334 4323 -17114 4329
rect -17334 4289 -17310 4323
rect -17126 4289 -17114 4323
rect -17334 4283 -17114 4289
rect -16774 4323 -16542 4329
rect -16774 4289 -16738 4323
rect -16554 4289 -16542 4323
rect -16774 4283 -16542 4289
rect -16312 4324 -16278 4854
rect -15852 4790 -15818 4854
rect -15878 4780 -15806 4790
rect -15878 4676 -15868 4780
rect -15816 4676 -15806 4780
rect -15878 4666 -15806 4676
rect -15740 4636 -15706 4854
rect -15280 4790 -15246 4854
rect -15306 4780 -15234 4790
rect -15306 4676 -15296 4780
rect -15244 4676 -15234 4780
rect -15306 4666 -15234 4676
rect -15754 4630 -15690 4636
rect -15754 4376 -15748 4630
rect -15696 4376 -15690 4630
rect -15754 4370 -15690 4376
rect -16176 4340 -15956 4342
rect -16176 4329 -16170 4340
rect -16178 4324 -16170 4329
rect -16312 4284 -16170 4324
rect -15962 4320 -15956 4340
rect -17334 4282 -17126 4283
rect -16774 4282 -16566 4283
rect -18614 4230 -18568 4282
rect -18614 1674 -18608 4230
rect -18574 1674 -18568 4230
rect -18614 1562 -18568 1674
rect -18156 4230 -18110 4282
rect -16312 4242 -16278 4284
rect -16178 4283 -16170 4284
rect -16176 4282 -16170 4283
rect -15962 4284 -15866 4320
rect -15962 4282 -15956 4284
rect -16176 4272 -15956 4282
rect -15740 4242 -15706 4370
rect -15604 4336 -15384 4342
rect -15604 4329 -15598 4336
rect -15606 4283 -15598 4329
rect -15604 4278 -15598 4283
rect -15390 4278 -15384 4336
rect -15604 4272 -15384 4278
rect -15168 4324 -15134 4854
rect -14708 4790 -14674 4854
rect -14734 4780 -14662 4790
rect -14734 4676 -14724 4780
rect -14672 4676 -14662 4780
rect -14734 4666 -14662 4676
rect -14596 4636 -14562 4854
rect -14136 4790 -14102 4854
rect -14162 4780 -14090 4790
rect -14162 4676 -14152 4780
rect -14100 4676 -14090 4780
rect -14162 4666 -14090 4676
rect -14610 4630 -14546 4636
rect -14610 4376 -14604 4630
rect -14552 4376 -14546 4630
rect -14610 4370 -14546 4376
rect -15032 4340 -14812 4346
rect -15032 4329 -15026 4340
rect -15034 4324 -15026 4329
rect -15168 4288 -15026 4324
rect -14818 4324 -14812 4340
rect -15168 4242 -15134 4288
rect -15034 4283 -15026 4288
rect -15032 4282 -15026 4283
rect -14818 4288 -14722 4324
rect -14818 4282 -14812 4288
rect -15032 4276 -14812 4282
rect -14596 4242 -14562 4370
rect -14460 4340 -14240 4346
rect -14460 4329 -14454 4340
rect -14462 4283 -14454 4329
rect -14460 4282 -14454 4283
rect -14246 4282 -14240 4340
rect -14460 4276 -14240 4282
rect -14024 4324 -13990 4854
rect -13564 4790 -13530 4854
rect -13590 4780 -13518 4790
rect -13590 4676 -13580 4780
rect -13528 4676 -13518 4780
rect -13590 4666 -13518 4676
rect -13452 4636 -13418 4854
rect -12992 4790 -12958 4854
rect -13018 4780 -12946 4790
rect -13018 4676 -13008 4780
rect -12956 4676 -12946 4780
rect -13018 4666 -12946 4676
rect -13466 4630 -13402 4636
rect -13466 4376 -13460 4630
rect -13408 4376 -13402 4630
rect -13466 4370 -13402 4376
rect -12746 4630 -12538 4636
rect -12746 4376 -12660 4630
rect -12608 4376 -12538 4630
rect -13888 4340 -13668 4346
rect -13888 4329 -13882 4340
rect -13890 4324 -13882 4329
rect -14024 4288 -13882 4324
rect -13674 4324 -13668 4340
rect -14024 4242 -13990 4288
rect -13890 4283 -13882 4288
rect -13888 4282 -13882 4283
rect -13674 4288 -13578 4324
rect -13674 4282 -13668 4288
rect -13888 4276 -13668 4282
rect -13452 4242 -13418 4370
rect -13316 4340 -13096 4346
rect -13316 4329 -13310 4340
rect -13318 4283 -13310 4329
rect -13316 4282 -13310 4283
rect -13102 4282 -13096 4340
rect -12746 4323 -12538 4376
rect -12746 4289 -12734 4323
rect -12550 4289 -12538 4323
rect -12746 4282 -12538 4289
rect -12186 4630 -11978 4636
rect -12186 4376 -12100 4630
rect -12048 4376 -11978 4630
rect -12186 4329 -11978 4376
rect -11626 4630 -11418 8038
rect -10364 6866 -10232 10106
rect -9908 7006 -9776 10690
rect -8390 10996 -6390 11410
rect -8390 10708 -8384 10996
rect -6396 10708 -6390 10996
rect -8390 9502 -6390 10708
rect -5690 10396 -3690 10408
rect -5690 10108 -5684 10396
rect -3696 10108 -3690 10396
rect -5690 9502 -3690 10108
rect -8350 9440 -8310 9502
rect -7430 9440 -7390 9502
rect -6510 9440 -6470 9502
rect -9908 6926 -9902 7006
rect -9782 6926 -9776 7006
rect -9908 6920 -9776 6926
rect -8806 9428 -8760 9440
rect -10364 6786 -10358 6866
rect -10248 6786 -10232 6866
rect -10364 6780 -10232 6786
rect -11626 4376 -11540 4630
rect -11488 4376 -11418 4630
rect -11626 4329 -11418 4376
rect -9496 4630 -9016 4636
rect -9496 4376 -9490 4630
rect -9022 4376 -9016 4630
rect -12186 4323 -11966 4329
rect -12186 4289 -12162 4323
rect -11978 4289 -11966 4323
rect -12186 4283 -11966 4289
rect -11626 4323 -11394 4329
rect -11626 4289 -11590 4323
rect -11406 4289 -11394 4323
rect -11626 4283 -11394 4289
rect -11178 4323 -10674 4330
rect -11178 4289 -11018 4323
rect -10834 4289 -10674 4323
rect -12186 4282 -11978 4283
rect -11626 4282 -11418 4283
rect -11178 4282 -10674 4289
rect -13316 4276 -13096 4282
rect -18156 1674 -18150 4230
rect -18116 1674 -18110 4230
rect -18156 1562 -18110 1674
rect -18042 4230 -17996 4242
rect -18042 1674 -18036 4230
rect -18002 1674 -17996 4230
rect -18042 1662 -17996 1674
rect -17584 4230 -17538 4242
rect -17584 1674 -17578 4230
rect -17544 1674 -17538 4230
rect -17584 1662 -17538 1674
rect -17470 4230 -17424 4242
rect -17470 1674 -17464 4230
rect -17430 1674 -17424 4230
rect -17470 1662 -17424 1674
rect -17012 4230 -16966 4242
rect -17012 1674 -17006 4230
rect -16972 4226 -16966 4230
rect -16898 4230 -16852 4242
rect -16972 1674 -16964 4226
rect -17012 1662 -16964 1674
rect -16898 1674 -16892 4230
rect -16858 1674 -16852 4230
rect -16898 1662 -16852 1674
rect -16440 4230 -16394 4242
rect -16440 1674 -16434 4230
rect -16400 4226 -16394 4230
rect -16326 4230 -16278 4242
rect -16400 1674 -16384 4226
rect -16440 1662 -16384 1674
rect -16326 1674 -16320 4230
rect -16286 4226 -16278 4230
rect -15868 4230 -15822 4242
rect -16286 1674 -16280 4226
rect -16326 1662 -16280 1674
rect -15868 1674 -15862 4230
rect -15828 4226 -15822 4230
rect -15754 4230 -15706 4242
rect -15296 4230 -15250 4242
rect -15828 1674 -15820 4226
rect -15868 1662 -15820 1674
rect -15754 1674 -15748 4230
rect -15714 1674 -15708 4230
rect -15754 1662 -15708 1674
rect -15296 1674 -15290 4230
rect -15256 4226 -15250 4230
rect -15182 4230 -15134 4242
rect -14724 4230 -14678 4242
rect -15256 1674 -15248 4226
rect -15296 1662 -15248 1674
rect -15182 1674 -15176 4230
rect -15142 1674 -15136 4230
rect -15182 1662 -15136 1674
rect -14724 1674 -14718 4230
rect -14684 1674 -14678 4230
rect -14724 1662 -14678 1674
rect -14610 4230 -14562 4242
rect -14152 4230 -14106 4242
rect -14610 1674 -14604 4230
rect -14570 1674 -14564 4230
rect -14610 1662 -14564 1674
rect -14152 1674 -14146 4230
rect -14112 1674 -14106 4230
rect -14152 1662 -14106 1674
rect -14038 4230 -13990 4242
rect -13580 4230 -13534 4242
rect -14038 1674 -14032 4230
rect -13998 1674 -13992 4230
rect -14038 1662 -13992 1674
rect -13580 1674 -13574 4230
rect -13540 1674 -13534 4230
rect -13580 1662 -13534 1674
rect -13466 4230 -13418 4242
rect -13008 4230 -12962 4242
rect -13466 1674 -13460 4230
rect -13426 1674 -13420 4230
rect -13466 1662 -13420 1674
rect -13008 1674 -13002 4230
rect -12968 1674 -12962 4230
rect -13008 1662 -12962 1674
rect -12894 4230 -12848 4242
rect -12894 1674 -12888 4230
rect -12854 1674 -12848 4230
rect -12894 1662 -12848 1674
rect -12436 4230 -12390 4242
rect -12436 1674 -12430 4230
rect -12396 1674 -12390 4230
rect -12436 1662 -12390 1674
rect -12322 4230 -12276 4242
rect -12322 1674 -12316 4230
rect -12282 1674 -12276 4230
rect -12322 1662 -12276 1674
rect -11864 4230 -11818 4242
rect -11864 1674 -11858 4230
rect -11824 1674 -11818 4230
rect -11864 1662 -11818 1674
rect -11750 4230 -11704 4242
rect -11750 1674 -11744 4230
rect -11710 1674 -11704 4230
rect -11750 1662 -11704 1674
rect -11292 4230 -11246 4242
rect -11292 1674 -11286 4230
rect -11252 1674 -11246 4230
rect -11292 1662 -11246 1674
rect -11178 4230 -11132 4282
rect -11178 1674 -11172 4230
rect -11138 1674 -11132 4230
rect -18628 1552 -18556 1562
rect -18628 1448 -18618 1552
rect -18566 1448 -18556 1552
rect -18628 1438 -18556 1448
rect -18170 1552 -18098 1562
rect -18170 1448 -18160 1552
rect -18108 1448 -18098 1552
rect -18170 1438 -18098 1448
rect -18040 1362 -17998 1662
rect -17578 1562 -17544 1662
rect -17594 1552 -17522 1562
rect -17594 1448 -17584 1552
rect -17532 1448 -17522 1552
rect -17594 1438 -17522 1448
rect -17468 1362 -17426 1662
rect -17006 1562 -16964 1662
rect -17022 1552 -16950 1562
rect -17022 1448 -17012 1552
rect -16960 1448 -16950 1552
rect -17022 1438 -16950 1448
rect -16896 1362 -16854 1662
rect -16434 1562 -16384 1662
rect -15862 1562 -15820 1662
rect -15290 1562 -15248 1662
rect -14718 1562 -14684 1662
rect -14146 1562 -14112 1662
rect -13574 1562 -13540 1662
rect -13002 1562 -12968 1662
rect -16450 1552 -16378 1562
rect -16450 1448 -16440 1552
rect -16388 1448 -16378 1552
rect -16450 1438 -16378 1448
rect -15878 1552 -15806 1562
rect -15878 1448 -15868 1552
rect -15816 1448 -15806 1552
rect -15878 1438 -15806 1448
rect -15306 1552 -15234 1562
rect -15306 1448 -15296 1552
rect -15244 1448 -15234 1552
rect -15306 1438 -15234 1448
rect -14734 1552 -14662 1562
rect -14734 1448 -14724 1552
rect -14672 1448 -14662 1552
rect -14734 1438 -14662 1448
rect -14162 1552 -14090 1562
rect -14162 1448 -14152 1552
rect -14100 1448 -14090 1552
rect -14162 1438 -14090 1448
rect -13590 1552 -13518 1562
rect -13590 1448 -13580 1552
rect -13528 1448 -13518 1552
rect -13590 1438 -13518 1448
rect -13018 1552 -12950 1562
rect -13018 1448 -13008 1552
rect -12956 1448 -12950 1552
rect -13018 1438 -12950 1448
rect -12892 1362 -12850 1662
rect -12430 1562 -12396 1662
rect -12446 1552 -12378 1562
rect -12446 1448 -12436 1552
rect -12384 1448 -12378 1552
rect -12446 1438 -12378 1448
rect -12320 1362 -12278 1662
rect -11858 1562 -11824 1662
rect -11874 1552 -11806 1562
rect -11874 1448 -11864 1552
rect -11812 1448 -11806 1552
rect -11874 1438 -11806 1448
rect -11748 1362 -11706 1662
rect -11286 1562 -11252 1662
rect -11178 1562 -11132 1674
rect -10720 4230 -10674 4282
rect -10720 1674 -10714 4230
rect -10680 1674 -10674 4230
rect -10720 1562 -10674 1674
rect -10138 4142 -10006 4154
rect -10138 1800 -10122 4142
rect -10022 1800 -10006 4142
rect -11302 1552 -11234 1562
rect -11302 1448 -11292 1552
rect -11240 1448 -11234 1552
rect -11302 1438 -11234 1448
rect -11192 1552 -11120 1562
rect -11192 1448 -11182 1552
rect -11130 1448 -11120 1552
rect -11192 1438 -11120 1448
rect -10734 1552 -10662 1562
rect -10734 1448 -10724 1552
rect -10672 1448 -10662 1552
rect -10734 1438 -10662 1448
rect -10138 1552 -10006 1800
rect -10138 1448 -10112 1552
rect -10060 1448 -10006 1552
rect -10138 1438 -10006 1448
rect -9496 1536 -9016 4376
rect -9496 1388 -9490 1536
rect -9022 1388 -9016 1536
rect -9496 1382 -9016 1388
rect -8806 1712 -8800 9428
rect -8766 1712 -8760 9428
rect -8350 9428 -8302 9440
rect -8350 9402 -8342 9428
rect -8806 1660 -8760 1712
rect -8348 1712 -8342 9402
rect -8308 1712 -8302 9428
rect -8348 1696 -8302 1712
rect -7890 9428 -7844 9440
rect -7890 1712 -7884 9428
rect -7850 1712 -7844 9428
rect -7890 1700 -7844 1712
rect -7432 9428 -7386 9440
rect -7432 1712 -7426 9428
rect -7392 1712 -7386 9428
rect -7432 1700 -7386 1712
rect -6974 9428 -6928 9440
rect -6974 1712 -6968 9428
rect -6934 1712 -6928 9428
rect -6974 1700 -6928 1712
rect -6516 9428 -6470 9440
rect -6516 1712 -6510 9428
rect -6476 1712 -6470 9428
rect -6516 1700 -6470 1712
rect -6058 9428 -6012 9440
rect -6058 1712 -6052 9428
rect -6018 1722 -6012 9428
rect -5610 9428 -5550 9502
rect -5610 9422 -5594 9428
rect -6018 1712 -6010 1722
rect -6058 1700 -6010 1712
rect -5600 1712 -5594 9422
rect -5560 9422 -5550 9428
rect -5142 9428 -5096 9440
rect -5560 1712 -5554 9422
rect -5142 1722 -5136 9428
rect -5600 1700 -5554 1712
rect -5150 1712 -5136 1722
rect -5102 1712 -5096 9428
rect -4690 9428 -4630 9502
rect -4690 9402 -4678 9428
rect -5150 1700 -5096 1712
rect -4684 1712 -4678 9402
rect -4644 9402 -4630 9428
rect -4226 9428 -4180 9440
rect -4644 1712 -4638 9402
rect -4226 1722 -4220 9428
rect -4684 1700 -4638 1712
rect -4230 1712 -4220 1722
rect -4186 1712 -4180 9428
rect -3770 9428 -3710 9502
rect -2890 9500 1810 12808
rect 9278 12640 10226 12646
rect 9278 12122 9286 12640
rect 10220 12122 10226 12640
rect 5310 11860 7310 11902
rect 5310 11410 5316 11860
rect 7304 11410 7310 11860
rect 5310 10996 7310 11410
rect 5310 10708 5316 10996
rect 7304 10708 7310 10996
rect 2610 10396 4610 10408
rect 2610 10108 2616 10396
rect 4604 10108 4610 10396
rect 2610 9502 4610 10108
rect 5310 9502 7310 10708
rect -3770 9402 -3762 9428
rect -4230 1700 -4180 1712
rect -3768 1712 -3762 9402
rect -3728 9402 -3710 9428
rect -2850 9440 -2810 9500
rect -1930 9440 -1890 9500
rect -1010 9440 -970 9500
rect -90 9440 -50 9500
rect -2850 9428 -2802 9440
rect -2850 9422 -2842 9428
rect -3728 1712 -3722 9402
rect -3768 1700 -3722 1712
rect -2848 1712 -2842 9422
rect -2808 1712 -2802 9428
rect -2848 1700 -2802 1712
rect -2390 9428 -2344 9440
rect -2390 1712 -2384 9428
rect -2350 1712 -2344 9428
rect -2390 1700 -2344 1712
rect -1932 9428 -1886 9440
rect -1932 1712 -1926 9428
rect -1892 1712 -1886 9428
rect -1932 1700 -1886 1712
rect -1474 9428 -1428 9440
rect -1474 1712 -1468 9428
rect -1434 1712 -1428 9428
rect -1474 1700 -1428 1712
rect -1016 9428 -970 9440
rect -1016 1712 -1010 9428
rect -976 1712 -970 9428
rect -1016 1700 -970 1712
rect -558 9428 -512 9440
rect -558 1712 -552 9428
rect -518 1722 -512 9428
rect -100 9428 -50 9440
rect -518 1712 -510 1722
rect -558 1700 -510 1712
rect -100 1712 -94 9428
rect -60 9402 -50 9428
rect 358 9428 404 9440
rect -60 1712 -54 9402
rect 358 1722 364 9428
rect -100 1700 -54 1712
rect 350 1712 364 1722
rect 398 1712 404 9428
rect 810 9428 870 9500
rect 810 9402 822 9428
rect 350 1700 404 1712
rect 816 1712 822 9402
rect 856 9402 870 9428
rect 1274 9428 1320 9440
rect 856 1712 862 9402
rect 1274 1722 1280 9428
rect 816 1700 862 1712
rect 1270 1712 1280 1722
rect 1314 1712 1320 9428
rect 1730 9428 1790 9500
rect 1730 9402 1738 9428
rect 1270 1700 1320 1712
rect 1732 1712 1738 9402
rect 1772 9402 1790 9428
rect 2650 9440 2690 9502
rect 3570 9440 3610 9502
rect 4490 9440 4530 9502
rect 2650 9428 2698 9440
rect 2650 9402 2658 9428
rect 1772 1712 1778 9402
rect 1732 1700 1778 1712
rect 2652 1712 2658 9402
rect 2692 1712 2698 9428
rect 2652 1700 2698 1712
rect 3110 9428 3156 9440
rect 3110 1712 3116 9428
rect 3150 1712 3156 9428
rect 3110 1700 3156 1712
rect 3568 9428 3614 9440
rect 3568 1712 3574 9428
rect 3608 1712 3614 9428
rect 3568 1700 3614 1712
rect 4026 9428 4072 9440
rect 4026 1712 4032 9428
rect 4066 1712 4072 9428
rect 4026 1700 4072 1712
rect 4484 9428 4530 9440
rect 4484 1712 4490 9428
rect 4524 1712 4530 9428
rect 4484 1700 4530 1712
rect 4942 9428 4988 9440
rect 4942 1712 4948 9428
rect 4982 1722 4988 9428
rect 5390 9428 5450 9502
rect 5390 9402 5406 9428
rect 4982 1712 4990 1722
rect 4942 1700 4990 1712
rect 5400 1712 5406 9402
rect 5440 9402 5450 9428
rect 5858 9428 5904 9440
rect 5440 1712 5446 9402
rect 5858 1722 5864 9428
rect 5400 1700 5446 1712
rect 5850 1712 5864 1722
rect 5898 1712 5904 9428
rect 6310 9428 6370 9502
rect 7230 9440 7270 9502
rect 6310 9422 6322 9428
rect 5850 1700 5904 1712
rect 6316 1712 6322 9422
rect 6356 9422 6370 9428
rect 6774 9428 6820 9440
rect 6356 1712 6362 9422
rect 6774 1722 6780 9428
rect 6316 1700 6362 1712
rect 6770 1712 6780 1722
rect 6814 1712 6820 9428
rect 7230 9428 7278 9440
rect 7230 9422 7238 9428
rect 6770 1700 6820 1712
rect 7232 1712 7238 9422
rect 7272 1712 7278 9428
rect -8806 1659 -8658 1660
rect -8466 1659 -8348 1660
rect -8190 1659 -8010 1662
rect -8806 1653 -8348 1659
rect -8806 1619 -8646 1653
rect -8462 1619 -8348 1653
rect -18930 1244 -18924 1358
rect -18730 1244 -18724 1358
rect -18930 1238 -18724 1244
rect -18054 1352 -17982 1362
rect -18054 1248 -18044 1352
rect -17992 1248 -17982 1352
rect -18054 1238 -17982 1248
rect -17482 1352 -17410 1362
rect -17482 1248 -17472 1352
rect -17420 1248 -17410 1352
rect -17482 1238 -17410 1248
rect -16910 1352 -16838 1362
rect -16910 1248 -16900 1352
rect -16848 1248 -16838 1352
rect -12906 1352 -12834 1362
rect -16910 1238 -16838 1248
rect -15680 1296 -13226 1312
rect -15680 1196 -15668 1296
rect -13326 1196 -13226 1296
rect -12906 1248 -12896 1352
rect -12844 1248 -12834 1352
rect -12906 1238 -12834 1248
rect -12334 1352 -12262 1362
rect -12334 1248 -12324 1352
rect -12272 1248 -12262 1352
rect -12334 1238 -12262 1248
rect -11762 1352 -11690 1362
rect -11762 1248 -11752 1352
rect -11700 1248 -11690 1352
rect -8806 1302 -8348 1619
rect -8200 1653 -7992 1659
rect -8200 1619 -8188 1653
rect -8004 1619 -7992 1653
rect -8200 1613 -7992 1619
rect -8190 1522 -8010 1613
rect -8190 1402 -8170 1522
rect -8030 1402 -8010 1522
rect -8190 1382 -8010 1402
rect -7890 1342 -7850 1700
rect -7730 1659 -7550 1662
rect -7270 1659 -7090 1662
rect -7742 1653 -7534 1659
rect -7742 1619 -7730 1653
rect -7546 1619 -7534 1653
rect -7742 1613 -7534 1619
rect -7284 1653 -7076 1659
rect -7284 1619 -7272 1653
rect -7088 1619 -7076 1653
rect -7284 1613 -7076 1619
rect -7730 1522 -7550 1613
rect -7730 1402 -7710 1522
rect -7570 1402 -7550 1522
rect -7730 1382 -7550 1402
rect -7270 1522 -7090 1613
rect -7270 1402 -7250 1522
rect -7110 1402 -7090 1522
rect -7270 1382 -7090 1402
rect -6970 1342 -6930 1700
rect -6810 1659 -6630 1662
rect -6350 1659 -6170 1662
rect -6826 1653 -6618 1659
rect -6826 1619 -6814 1653
rect -6630 1619 -6618 1653
rect -6826 1613 -6618 1619
rect -6368 1653 -6160 1659
rect -6368 1619 -6356 1653
rect -6172 1619 -6160 1653
rect -6368 1613 -6160 1619
rect -6810 1522 -6630 1613
rect -6810 1402 -6790 1522
rect -6650 1402 -6630 1522
rect -6810 1382 -6630 1402
rect -6350 1522 -6170 1613
rect -6350 1402 -6330 1522
rect -6190 1402 -6170 1522
rect -6350 1382 -6170 1402
rect -6050 1342 -6010 1700
rect -5890 1659 -5710 1662
rect -5430 1659 -5250 1662
rect -5910 1653 -5702 1659
rect -5910 1619 -5898 1653
rect -5714 1619 -5702 1653
rect -5910 1613 -5702 1619
rect -5452 1653 -5244 1659
rect -5452 1619 -5440 1653
rect -5256 1619 -5244 1653
rect -5452 1613 -5244 1619
rect -5890 1522 -5710 1613
rect -5890 1402 -5870 1522
rect -5730 1402 -5710 1522
rect -5890 1382 -5710 1402
rect -5430 1522 -5250 1613
rect -5430 1402 -5410 1522
rect -5270 1402 -5250 1522
rect -5430 1382 -5250 1402
rect -5150 1342 -5110 1700
rect -4970 1659 -4790 1662
rect -4510 1659 -4330 1662
rect -4994 1653 -4786 1659
rect -4994 1619 -4982 1653
rect -4798 1619 -4786 1653
rect -4994 1613 -4786 1619
rect -4536 1653 -4328 1659
rect -4536 1619 -4524 1653
rect -4340 1619 -4328 1653
rect -4536 1613 -4328 1619
rect -4970 1522 -4790 1613
rect -4970 1402 -4950 1522
rect -4810 1402 -4790 1522
rect -4970 1382 -4790 1402
rect -4510 1522 -4330 1613
rect -4510 1402 -4490 1522
rect -4350 1402 -4330 1522
rect -4510 1382 -4330 1402
rect -4230 1342 -4190 1700
rect -4050 1659 -3870 1662
rect -2690 1659 -2510 1662
rect -4078 1653 -3870 1659
rect -4078 1619 -4066 1653
rect -3882 1619 -3870 1653
rect -4078 1613 -3870 1619
rect -2700 1653 -2492 1659
rect -2700 1619 -2688 1653
rect -2504 1619 -2492 1653
rect -2700 1613 -2492 1619
rect -4050 1522 -3870 1613
rect -4050 1402 -4030 1522
rect -3890 1402 -3870 1522
rect -4050 1382 -3870 1402
rect -2690 1522 -2510 1613
rect -2690 1402 -2670 1522
rect -2530 1402 -2510 1522
rect -2690 1382 -2510 1402
rect -2390 1342 -2350 1700
rect -2230 1659 -2050 1662
rect -1770 1659 -1590 1662
rect -2242 1653 -2034 1659
rect -2242 1619 -2230 1653
rect -2046 1619 -2034 1653
rect -2242 1613 -2034 1619
rect -1784 1653 -1576 1659
rect -1784 1619 -1772 1653
rect -1588 1619 -1576 1653
rect -1784 1613 -1576 1619
rect -2230 1522 -2050 1613
rect -2230 1402 -2210 1522
rect -2070 1402 -2050 1522
rect -2230 1382 -2050 1402
rect -1770 1522 -1590 1613
rect -1770 1402 -1750 1522
rect -1610 1402 -1590 1522
rect -1770 1382 -1590 1402
rect -1470 1342 -1430 1700
rect -1310 1659 -1130 1662
rect -850 1659 -670 1662
rect -1326 1653 -1118 1659
rect -1326 1619 -1314 1653
rect -1130 1619 -1118 1653
rect -1326 1613 -1118 1619
rect -868 1653 -660 1659
rect -868 1619 -856 1653
rect -672 1619 -660 1653
rect -868 1613 -660 1619
rect -1310 1522 -1130 1613
rect -1310 1402 -1290 1522
rect -1150 1402 -1130 1522
rect -1310 1382 -1130 1402
rect -850 1522 -670 1613
rect -850 1402 -830 1522
rect -690 1402 -670 1522
rect -850 1382 -670 1402
rect -550 1342 -510 1700
rect -390 1659 -210 1662
rect 70 1659 250 1662
rect -410 1653 -202 1659
rect -410 1619 -398 1653
rect -214 1619 -202 1653
rect -410 1613 -202 1619
rect 48 1653 256 1659
rect 48 1619 60 1653
rect 244 1619 256 1653
rect 48 1613 256 1619
rect -390 1522 -210 1613
rect -390 1402 -370 1522
rect -230 1402 -210 1522
rect -390 1382 -210 1402
rect 70 1522 250 1613
rect 70 1402 90 1522
rect 230 1402 250 1522
rect 70 1382 250 1402
rect 350 1342 390 1700
rect 530 1659 710 1662
rect 990 1659 1170 1662
rect 506 1653 714 1659
rect 506 1619 518 1653
rect 702 1619 714 1653
rect 506 1613 714 1619
rect 964 1653 1172 1659
rect 964 1619 976 1653
rect 1160 1619 1172 1653
rect 964 1613 1172 1619
rect 530 1522 710 1613
rect 530 1402 550 1522
rect 690 1402 710 1522
rect 530 1382 710 1402
rect 990 1522 1170 1613
rect 990 1402 1010 1522
rect 1150 1402 1170 1522
rect 990 1382 1170 1402
rect 1270 1342 1310 1700
rect 1450 1659 1630 1662
rect 2810 1659 2990 1662
rect 1422 1653 1630 1659
rect 1422 1619 1434 1653
rect 1618 1619 1630 1653
rect 1422 1613 1630 1619
rect 2800 1653 3008 1659
rect 2800 1619 2812 1653
rect 2996 1619 3008 1653
rect 2800 1613 3008 1619
rect 1450 1522 1630 1613
rect 1450 1402 1470 1522
rect 1610 1402 1630 1522
rect 1450 1382 1630 1402
rect 2810 1522 2990 1613
rect 2810 1402 2830 1522
rect 2970 1402 2990 1522
rect 2810 1382 2990 1402
rect 3110 1342 3150 1700
rect 3270 1659 3450 1662
rect 3730 1659 3910 1662
rect 3258 1653 3466 1659
rect 3258 1619 3270 1653
rect 3454 1619 3466 1653
rect 3258 1613 3466 1619
rect 3716 1653 3924 1659
rect 3716 1619 3728 1653
rect 3912 1619 3924 1653
rect 3716 1613 3924 1619
rect 3270 1522 3450 1613
rect 3270 1402 3290 1522
rect 3430 1402 3450 1522
rect 3270 1382 3450 1402
rect 3730 1522 3910 1613
rect 3730 1402 3750 1522
rect 3890 1402 3910 1522
rect 3730 1382 3910 1402
rect 4030 1342 4070 1700
rect 4190 1659 4370 1662
rect 4650 1659 4830 1662
rect 4174 1653 4382 1659
rect 4174 1619 4186 1653
rect 4370 1619 4382 1653
rect 4174 1613 4382 1619
rect 4632 1653 4840 1659
rect 4632 1619 4644 1653
rect 4828 1619 4840 1653
rect 4632 1613 4840 1619
rect 4190 1522 4370 1613
rect 4190 1402 4210 1522
rect 4350 1402 4370 1522
rect 4190 1382 4370 1402
rect 4650 1522 4830 1613
rect 4650 1402 4670 1522
rect 4810 1402 4830 1522
rect 4650 1382 4830 1402
rect 4950 1342 4990 1700
rect 5110 1659 5290 1662
rect 5570 1659 5750 1662
rect 5090 1653 5298 1659
rect 5090 1619 5102 1653
rect 5286 1619 5298 1653
rect 5090 1613 5298 1619
rect 5548 1653 5756 1659
rect 5548 1619 5560 1653
rect 5744 1619 5756 1653
rect 5548 1613 5756 1619
rect 5110 1522 5290 1613
rect 5110 1402 5130 1522
rect 5270 1402 5290 1522
rect 5110 1382 5290 1402
rect 5570 1522 5750 1613
rect 5570 1402 5590 1522
rect 5730 1402 5750 1522
rect 5570 1382 5750 1402
rect 5850 1342 5890 1700
rect 6030 1659 6210 1662
rect 6490 1659 6670 1662
rect 6006 1653 6214 1659
rect 6006 1619 6018 1653
rect 6202 1619 6214 1653
rect 6006 1613 6214 1619
rect 6464 1653 6672 1659
rect 6464 1619 6476 1653
rect 6660 1619 6672 1653
rect 6464 1613 6672 1619
rect 6030 1522 6210 1613
rect 6030 1402 6050 1522
rect 6190 1402 6210 1522
rect 6030 1382 6210 1402
rect 6490 1522 6670 1613
rect 6490 1402 6510 1522
rect 6650 1402 6670 1522
rect 6490 1382 6670 1402
rect 6770 1342 6810 1700
rect 7232 1696 7278 1712
rect 7690 9428 7736 9440
rect 7690 1712 7696 9428
rect 7730 1712 7736 9428
rect 9278 3162 10226 12122
rect 10622 11860 11326 14498
rect 10622 11410 10628 11860
rect 11320 11410 11326 11860
rect 10622 8072 11326 11410
rect 11440 15190 12144 15196
rect 11440 14498 11446 15190
rect 12138 14498 12144 15190
rect 12340 15179 12902 15185
rect 12340 14782 12352 15179
rect 12890 14782 12902 15179
rect 12340 14776 12902 14782
rect 11440 10396 12144 14498
rect 11440 10108 11448 10396
rect 12138 10108 12144 10396
rect 11440 10102 12144 10108
rect 12740 11864 18584 11918
rect 12740 11830 12828 11864
rect 12862 11830 12928 11864
rect 12962 11830 13028 11864
rect 13062 11830 13128 11864
rect 13162 11830 13228 11864
rect 13262 11830 13328 11864
rect 13362 11830 14116 11864
rect 14150 11830 14216 11864
rect 14250 11830 14316 11864
rect 14350 11830 14416 11864
rect 14450 11830 14516 11864
rect 14550 11830 14616 11864
rect 14650 11830 15404 11864
rect 15438 11830 15504 11864
rect 15538 11830 15604 11864
rect 15638 11830 15704 11864
rect 15738 11830 15804 11864
rect 15838 11830 15904 11864
rect 15938 11830 16692 11864
rect 16726 11830 16792 11864
rect 16826 11830 16892 11864
rect 16926 11830 16992 11864
rect 17026 11830 17092 11864
rect 17126 11830 17192 11864
rect 17226 11830 17980 11864
rect 18014 11830 18080 11864
rect 18114 11830 18180 11864
rect 18214 11830 18280 11864
rect 18314 11830 18380 11864
rect 18414 11830 18480 11864
rect 18514 11830 18584 11864
rect 12740 11764 18584 11830
rect 12740 11730 12828 11764
rect 12862 11730 12928 11764
rect 12962 11730 13028 11764
rect 13062 11730 13128 11764
rect 13162 11730 13228 11764
rect 13262 11730 13328 11764
rect 13362 11730 14116 11764
rect 14150 11730 14216 11764
rect 14250 11730 14316 11764
rect 14350 11730 14416 11764
rect 14450 11730 14516 11764
rect 14550 11730 14616 11764
rect 14650 11730 15404 11764
rect 15438 11730 15504 11764
rect 15538 11730 15604 11764
rect 15638 11730 15704 11764
rect 15738 11730 15804 11764
rect 15838 11730 15904 11764
rect 15938 11730 16692 11764
rect 16726 11730 16792 11764
rect 16826 11730 16892 11764
rect 16926 11730 16992 11764
rect 17026 11730 17092 11764
rect 17126 11730 17192 11764
rect 17226 11730 17980 11764
rect 18014 11730 18080 11764
rect 18114 11730 18180 11764
rect 18214 11730 18280 11764
rect 18314 11730 18380 11764
rect 18414 11730 18480 11764
rect 18514 11730 18584 11764
rect 12740 11664 18584 11730
rect 12740 11630 12828 11664
rect 12862 11630 12928 11664
rect 12962 11630 13028 11664
rect 13062 11630 13128 11664
rect 13162 11630 13228 11664
rect 13262 11630 13328 11664
rect 13362 11630 14116 11664
rect 14150 11630 14216 11664
rect 14250 11630 14316 11664
rect 14350 11630 14416 11664
rect 14450 11630 14516 11664
rect 14550 11630 14616 11664
rect 14650 11630 15404 11664
rect 15438 11630 15504 11664
rect 15538 11630 15604 11664
rect 15638 11630 15704 11664
rect 15738 11630 15804 11664
rect 15838 11630 15904 11664
rect 15938 11630 16692 11664
rect 16726 11630 16792 11664
rect 16826 11630 16892 11664
rect 16926 11630 16992 11664
rect 17026 11630 17092 11664
rect 17126 11630 17192 11664
rect 17226 11630 17980 11664
rect 18014 11630 18080 11664
rect 18114 11630 18180 11664
rect 18214 11630 18280 11664
rect 18314 11630 18380 11664
rect 18414 11630 18480 11664
rect 18514 11630 18584 11664
rect 12740 11564 18584 11630
rect 12740 11530 12828 11564
rect 12862 11530 12928 11564
rect 12962 11530 13028 11564
rect 13062 11530 13128 11564
rect 13162 11530 13228 11564
rect 13262 11530 13328 11564
rect 13362 11530 14116 11564
rect 14150 11530 14216 11564
rect 14250 11530 14316 11564
rect 14350 11530 14416 11564
rect 14450 11530 14516 11564
rect 14550 11530 14616 11564
rect 14650 11530 15404 11564
rect 15438 11530 15504 11564
rect 15538 11530 15604 11564
rect 15638 11530 15704 11564
rect 15738 11530 15804 11564
rect 15838 11530 15904 11564
rect 15938 11530 16692 11564
rect 16726 11530 16792 11564
rect 16826 11530 16892 11564
rect 16926 11530 16992 11564
rect 17026 11530 17092 11564
rect 17126 11530 17192 11564
rect 17226 11530 17980 11564
rect 18014 11530 18080 11564
rect 18114 11530 18180 11564
rect 18214 11530 18280 11564
rect 18314 11530 18380 11564
rect 18414 11530 18480 11564
rect 18514 11530 18584 11564
rect 12740 11464 18584 11530
rect 12740 11430 12828 11464
rect 12862 11430 12928 11464
rect 12962 11430 13028 11464
rect 13062 11430 13128 11464
rect 13162 11430 13228 11464
rect 13262 11430 13328 11464
rect 13362 11430 14116 11464
rect 14150 11430 14216 11464
rect 14250 11430 14316 11464
rect 14350 11430 14416 11464
rect 14450 11430 14516 11464
rect 14550 11430 14616 11464
rect 14650 11430 15404 11464
rect 15438 11430 15504 11464
rect 15538 11430 15604 11464
rect 15638 11430 15704 11464
rect 15738 11430 15804 11464
rect 15838 11430 15904 11464
rect 15938 11430 16692 11464
rect 16726 11430 16792 11464
rect 16826 11430 16892 11464
rect 16926 11430 16992 11464
rect 17026 11430 17092 11464
rect 17126 11430 17192 11464
rect 17226 11430 17980 11464
rect 18014 11430 18080 11464
rect 18114 11430 18180 11464
rect 18214 11430 18280 11464
rect 18314 11430 18380 11464
rect 18414 11430 18480 11464
rect 18514 11430 18584 11464
rect 12740 11364 18584 11430
rect 12740 11330 12828 11364
rect 12862 11330 12928 11364
rect 12962 11330 13028 11364
rect 13062 11330 13128 11364
rect 13162 11330 13228 11364
rect 13262 11330 13328 11364
rect 13362 11330 14116 11364
rect 14150 11330 14216 11364
rect 14250 11330 14316 11364
rect 14350 11330 14416 11364
rect 14450 11330 14516 11364
rect 14550 11330 14616 11364
rect 14650 11330 15404 11364
rect 15438 11330 15504 11364
rect 15538 11330 15604 11364
rect 15638 11330 15704 11364
rect 15738 11330 15804 11364
rect 15838 11330 15904 11364
rect 15938 11330 16692 11364
rect 16726 11330 16792 11364
rect 16826 11330 16892 11364
rect 16926 11330 16992 11364
rect 17026 11330 17092 11364
rect 17126 11330 17192 11364
rect 17226 11330 17980 11364
rect 18014 11330 18080 11364
rect 18114 11330 18180 11364
rect 18214 11330 18280 11364
rect 18314 11330 18380 11364
rect 18414 11330 18480 11364
rect 18514 11330 18584 11364
rect 12740 10576 18584 11330
rect 12740 10542 12828 10576
rect 12862 10542 12928 10576
rect 12962 10542 13028 10576
rect 13062 10542 13128 10576
rect 13162 10542 13228 10576
rect 13262 10542 13328 10576
rect 13362 10542 14116 10576
rect 14150 10542 14216 10576
rect 14250 10542 14316 10576
rect 14350 10542 14416 10576
rect 14450 10542 14516 10576
rect 14550 10542 14616 10576
rect 14650 10542 15404 10576
rect 15438 10542 15504 10576
rect 15538 10542 15604 10576
rect 15638 10542 15704 10576
rect 15738 10542 15804 10576
rect 15838 10542 15904 10576
rect 15938 10542 16692 10576
rect 16726 10542 16792 10576
rect 16826 10542 16892 10576
rect 16926 10542 16992 10576
rect 17026 10542 17092 10576
rect 17126 10542 17192 10576
rect 17226 10542 17980 10576
rect 18014 10542 18080 10576
rect 18114 10542 18180 10576
rect 18214 10542 18280 10576
rect 18314 10542 18380 10576
rect 18414 10542 18480 10576
rect 18514 10542 18584 10576
rect 12740 10476 18584 10542
rect 12740 10442 12828 10476
rect 12862 10442 12928 10476
rect 12962 10442 13028 10476
rect 13062 10442 13128 10476
rect 13162 10442 13228 10476
rect 13262 10442 13328 10476
rect 13362 10442 14116 10476
rect 14150 10442 14216 10476
rect 14250 10442 14316 10476
rect 14350 10442 14416 10476
rect 14450 10442 14516 10476
rect 14550 10442 14616 10476
rect 14650 10442 15404 10476
rect 15438 10442 15504 10476
rect 15538 10442 15604 10476
rect 15638 10442 15704 10476
rect 15738 10442 15804 10476
rect 15838 10442 15904 10476
rect 15938 10442 16692 10476
rect 16726 10442 16792 10476
rect 16826 10442 16892 10476
rect 16926 10442 16992 10476
rect 17026 10442 17092 10476
rect 17126 10442 17192 10476
rect 17226 10442 17980 10476
rect 18014 10442 18080 10476
rect 18114 10442 18180 10476
rect 18214 10442 18280 10476
rect 18314 10442 18380 10476
rect 18414 10442 18480 10476
rect 18514 10442 18584 10476
rect 12740 10376 18584 10442
rect 12740 10342 12828 10376
rect 12862 10342 12928 10376
rect 12962 10342 13028 10376
rect 13062 10342 13128 10376
rect 13162 10342 13228 10376
rect 13262 10342 13328 10376
rect 13362 10342 14116 10376
rect 14150 10342 14216 10376
rect 14250 10342 14316 10376
rect 14350 10342 14416 10376
rect 14450 10342 14516 10376
rect 14550 10342 14616 10376
rect 14650 10342 15404 10376
rect 15438 10342 15504 10376
rect 15538 10342 15604 10376
rect 15638 10342 15704 10376
rect 15738 10342 15804 10376
rect 15838 10342 15904 10376
rect 15938 10342 16692 10376
rect 16726 10342 16792 10376
rect 16826 10342 16892 10376
rect 16926 10342 16992 10376
rect 17026 10342 17092 10376
rect 17126 10342 17192 10376
rect 17226 10342 17980 10376
rect 18014 10342 18080 10376
rect 18114 10342 18180 10376
rect 18214 10342 18280 10376
rect 18314 10342 18380 10376
rect 18414 10342 18480 10376
rect 18514 10342 18584 10376
rect 12740 10276 18584 10342
rect 12740 10242 12828 10276
rect 12862 10242 12928 10276
rect 12962 10242 13028 10276
rect 13062 10242 13128 10276
rect 13162 10242 13228 10276
rect 13262 10242 13328 10276
rect 13362 10242 14116 10276
rect 14150 10242 14216 10276
rect 14250 10242 14316 10276
rect 14350 10242 14416 10276
rect 14450 10242 14516 10276
rect 14550 10242 14616 10276
rect 14650 10242 15404 10276
rect 15438 10242 15504 10276
rect 15538 10242 15604 10276
rect 15638 10242 15704 10276
rect 15738 10242 15804 10276
rect 15838 10242 15904 10276
rect 15938 10242 16692 10276
rect 16726 10242 16792 10276
rect 16826 10242 16892 10276
rect 16926 10242 16992 10276
rect 17026 10242 17092 10276
rect 17126 10242 17192 10276
rect 17226 10242 17980 10276
rect 18014 10242 18080 10276
rect 18114 10242 18180 10276
rect 18214 10242 18280 10276
rect 18314 10242 18380 10276
rect 18414 10242 18480 10276
rect 18514 10242 18584 10276
rect 12740 10176 18584 10242
rect 12740 10142 12828 10176
rect 12862 10142 12928 10176
rect 12962 10142 13028 10176
rect 13062 10142 13128 10176
rect 13162 10142 13228 10176
rect 13262 10142 13328 10176
rect 13362 10142 14116 10176
rect 14150 10142 14216 10176
rect 14250 10142 14316 10176
rect 14350 10142 14416 10176
rect 14450 10142 14516 10176
rect 14550 10142 14616 10176
rect 14650 10142 15404 10176
rect 15438 10142 15504 10176
rect 15538 10142 15604 10176
rect 15638 10142 15704 10176
rect 15738 10142 15804 10176
rect 15838 10142 15904 10176
rect 15938 10142 16692 10176
rect 16726 10142 16792 10176
rect 16826 10142 16892 10176
rect 16926 10142 16992 10176
rect 17026 10142 17092 10176
rect 17126 10142 17192 10176
rect 17226 10142 17980 10176
rect 18014 10142 18080 10176
rect 18114 10142 18180 10176
rect 18214 10142 18280 10176
rect 18314 10142 18380 10176
rect 18414 10142 18480 10176
rect 18514 10142 18584 10176
rect 10622 7380 10628 8072
rect 11320 7380 11326 8072
rect 10622 7372 11326 7380
rect 12740 10076 18584 10142
rect 12740 10042 12828 10076
rect 12862 10042 12928 10076
rect 12962 10042 13028 10076
rect 13062 10042 13128 10076
rect 13162 10042 13228 10076
rect 13262 10042 13328 10076
rect 13362 10042 14116 10076
rect 14150 10042 14216 10076
rect 14250 10042 14316 10076
rect 14350 10042 14416 10076
rect 14450 10042 14516 10076
rect 14550 10042 14616 10076
rect 14650 10042 15404 10076
rect 15438 10042 15504 10076
rect 15538 10042 15604 10076
rect 15638 10042 15704 10076
rect 15738 10042 15804 10076
rect 15838 10042 15904 10076
rect 15938 10042 16692 10076
rect 16726 10042 16792 10076
rect 16826 10042 16892 10076
rect 16926 10042 16992 10076
rect 17026 10042 17092 10076
rect 17126 10042 17192 10076
rect 17226 10042 17980 10076
rect 18014 10042 18080 10076
rect 18114 10042 18180 10076
rect 18214 10042 18280 10076
rect 18314 10042 18380 10076
rect 18414 10042 18480 10076
rect 18514 10042 18584 10076
rect 12740 9288 18584 10042
rect 12740 9254 12828 9288
rect 12862 9254 12928 9288
rect 12962 9254 13028 9288
rect 13062 9254 13128 9288
rect 13162 9254 13228 9288
rect 13262 9254 13328 9288
rect 13362 9254 14116 9288
rect 14150 9254 14216 9288
rect 14250 9254 14316 9288
rect 14350 9254 14416 9288
rect 14450 9254 14516 9288
rect 14550 9254 14616 9288
rect 14650 9254 15404 9288
rect 15438 9254 15504 9288
rect 15538 9254 15604 9288
rect 15638 9254 15704 9288
rect 15738 9254 15804 9288
rect 15838 9254 15904 9288
rect 15938 9254 16692 9288
rect 16726 9254 16792 9288
rect 16826 9254 16892 9288
rect 16926 9254 16992 9288
rect 17026 9254 17092 9288
rect 17126 9254 17192 9288
rect 17226 9254 17980 9288
rect 18014 9254 18080 9288
rect 18114 9254 18180 9288
rect 18214 9254 18280 9288
rect 18314 9254 18380 9288
rect 18414 9254 18480 9288
rect 18514 9254 18584 9288
rect 12740 9188 18584 9254
rect 12740 9154 12828 9188
rect 12862 9154 12928 9188
rect 12962 9154 13028 9188
rect 13062 9154 13128 9188
rect 13162 9154 13228 9188
rect 13262 9154 13328 9188
rect 13362 9154 14116 9188
rect 14150 9154 14216 9188
rect 14250 9154 14316 9188
rect 14350 9154 14416 9188
rect 14450 9154 14516 9188
rect 14550 9154 14616 9188
rect 14650 9154 15404 9188
rect 15438 9154 15504 9188
rect 15538 9154 15604 9188
rect 15638 9154 15704 9188
rect 15738 9154 15804 9188
rect 15838 9154 15904 9188
rect 15938 9154 16692 9188
rect 16726 9154 16792 9188
rect 16826 9154 16892 9188
rect 16926 9154 16992 9188
rect 17026 9154 17092 9188
rect 17126 9154 17192 9188
rect 17226 9154 17980 9188
rect 18014 9154 18080 9188
rect 18114 9154 18180 9188
rect 18214 9154 18280 9188
rect 18314 9154 18380 9188
rect 18414 9154 18480 9188
rect 18514 9154 18584 9188
rect 12740 9088 18584 9154
rect 12740 9054 12828 9088
rect 12862 9054 12928 9088
rect 12962 9054 13028 9088
rect 13062 9054 13128 9088
rect 13162 9054 13228 9088
rect 13262 9054 13328 9088
rect 13362 9054 14116 9088
rect 14150 9054 14216 9088
rect 14250 9054 14316 9088
rect 14350 9054 14416 9088
rect 14450 9054 14516 9088
rect 14550 9054 14616 9088
rect 14650 9054 15404 9088
rect 15438 9054 15504 9088
rect 15538 9054 15604 9088
rect 15638 9054 15704 9088
rect 15738 9054 15804 9088
rect 15838 9054 15904 9088
rect 15938 9054 16692 9088
rect 16726 9054 16792 9088
rect 16826 9054 16892 9088
rect 16926 9054 16992 9088
rect 17026 9054 17092 9088
rect 17126 9054 17192 9088
rect 17226 9054 17980 9088
rect 18014 9054 18080 9088
rect 18114 9054 18180 9088
rect 18214 9054 18280 9088
rect 18314 9054 18380 9088
rect 18414 9054 18480 9088
rect 18514 9054 18584 9088
rect 12740 8988 18584 9054
rect 12740 8954 12828 8988
rect 12862 8954 12928 8988
rect 12962 8954 13028 8988
rect 13062 8954 13128 8988
rect 13162 8954 13228 8988
rect 13262 8954 13328 8988
rect 13362 8954 14116 8988
rect 14150 8954 14216 8988
rect 14250 8954 14316 8988
rect 14350 8954 14416 8988
rect 14450 8954 14516 8988
rect 14550 8954 14616 8988
rect 14650 8954 15404 8988
rect 15438 8954 15504 8988
rect 15538 8954 15604 8988
rect 15638 8954 15704 8988
rect 15738 8954 15804 8988
rect 15838 8954 15904 8988
rect 15938 8954 16692 8988
rect 16726 8954 16792 8988
rect 16826 8954 16892 8988
rect 16926 8954 16992 8988
rect 17026 8954 17092 8988
rect 17126 8954 17192 8988
rect 17226 8954 17980 8988
rect 18014 8954 18080 8988
rect 18114 8954 18180 8988
rect 18214 8954 18280 8988
rect 18314 8954 18380 8988
rect 18414 8954 18480 8988
rect 18514 8954 18584 8988
rect 12740 8888 18584 8954
rect 12740 8854 12828 8888
rect 12862 8854 12928 8888
rect 12962 8854 13028 8888
rect 13062 8854 13128 8888
rect 13162 8854 13228 8888
rect 13262 8854 13328 8888
rect 13362 8854 14116 8888
rect 14150 8854 14216 8888
rect 14250 8854 14316 8888
rect 14350 8854 14416 8888
rect 14450 8854 14516 8888
rect 14550 8854 14616 8888
rect 14650 8854 15404 8888
rect 15438 8854 15504 8888
rect 15538 8854 15604 8888
rect 15638 8854 15704 8888
rect 15738 8854 15804 8888
rect 15838 8854 15904 8888
rect 15938 8854 16692 8888
rect 16726 8854 16792 8888
rect 16826 8854 16892 8888
rect 16926 8854 16992 8888
rect 17026 8854 17092 8888
rect 17126 8854 17192 8888
rect 17226 8854 17980 8888
rect 18014 8854 18080 8888
rect 18114 8854 18180 8888
rect 18214 8854 18280 8888
rect 18314 8854 18380 8888
rect 18414 8854 18480 8888
rect 18514 8854 18584 8888
rect 12740 8788 18584 8854
rect 12740 8754 12828 8788
rect 12862 8754 12928 8788
rect 12962 8754 13028 8788
rect 13062 8754 13128 8788
rect 13162 8754 13228 8788
rect 13262 8754 13328 8788
rect 13362 8754 14116 8788
rect 14150 8754 14216 8788
rect 14250 8754 14316 8788
rect 14350 8754 14416 8788
rect 14450 8754 14516 8788
rect 14550 8754 14616 8788
rect 14650 8754 15404 8788
rect 15438 8754 15504 8788
rect 15538 8754 15604 8788
rect 15638 8754 15704 8788
rect 15738 8754 15804 8788
rect 15838 8754 15904 8788
rect 15938 8754 16692 8788
rect 16726 8754 16792 8788
rect 16826 8754 16892 8788
rect 16926 8754 16992 8788
rect 17026 8754 17092 8788
rect 17126 8754 17192 8788
rect 17226 8754 17980 8788
rect 18014 8754 18080 8788
rect 18114 8754 18180 8788
rect 18214 8754 18280 8788
rect 18314 8754 18380 8788
rect 18414 8754 18480 8788
rect 18514 8754 18584 8788
rect 12740 8136 18584 8754
rect 12740 8000 15254 8136
rect 12740 7966 12828 8000
rect 12862 7966 12928 8000
rect 12962 7966 13028 8000
rect 13062 7966 13128 8000
rect 13162 7966 13228 8000
rect 13262 7966 13328 8000
rect 13362 7966 14116 8000
rect 14150 7966 14216 8000
rect 14250 7966 14316 8000
rect 14350 7966 14416 8000
rect 14450 7966 14516 8000
rect 14550 7966 14616 8000
rect 14650 7966 15254 8000
rect 12740 7900 15254 7966
rect 12740 7866 12828 7900
rect 12862 7866 12928 7900
rect 12962 7866 13028 7900
rect 13062 7866 13128 7900
rect 13162 7866 13228 7900
rect 13262 7866 13328 7900
rect 13362 7866 14116 7900
rect 14150 7866 14216 7900
rect 14250 7866 14316 7900
rect 14350 7866 14416 7900
rect 14450 7866 14516 7900
rect 14550 7866 14616 7900
rect 14650 7866 15254 7900
rect 12740 7800 15254 7866
rect 12740 7766 12828 7800
rect 12862 7766 12928 7800
rect 12962 7766 13028 7800
rect 13062 7766 13128 7800
rect 13162 7766 13228 7800
rect 13262 7766 13328 7800
rect 13362 7766 14116 7800
rect 14150 7766 14216 7800
rect 14250 7766 14316 7800
rect 14350 7766 14416 7800
rect 14450 7766 14516 7800
rect 14550 7766 14616 7800
rect 14650 7766 15254 7800
rect 12740 7700 15254 7766
rect 12740 7666 12828 7700
rect 12862 7666 12928 7700
rect 12962 7666 13028 7700
rect 13062 7666 13128 7700
rect 13162 7666 13228 7700
rect 13262 7666 13328 7700
rect 13362 7666 14116 7700
rect 14150 7666 14216 7700
rect 14250 7666 14316 7700
rect 14350 7666 14416 7700
rect 14450 7666 14516 7700
rect 14550 7666 14616 7700
rect 14650 7666 15254 7700
rect 12740 7600 15254 7666
rect 12740 7566 12828 7600
rect 12862 7566 12928 7600
rect 12962 7566 13028 7600
rect 13062 7566 13128 7600
rect 13162 7566 13228 7600
rect 13262 7566 13328 7600
rect 13362 7566 14116 7600
rect 14150 7566 14216 7600
rect 14250 7566 14316 7600
rect 14350 7566 14416 7600
rect 14450 7566 14516 7600
rect 14550 7566 14616 7600
rect 14650 7566 15254 7600
rect 12740 7500 15254 7566
rect 12740 7466 12828 7500
rect 12862 7466 12928 7500
rect 12962 7466 13028 7500
rect 13062 7466 13128 7500
rect 13162 7466 13228 7500
rect 13262 7466 13328 7500
rect 13362 7466 14116 7500
rect 14150 7466 14216 7500
rect 14250 7466 14316 7500
rect 14350 7466 14416 7500
rect 14450 7466 14516 7500
rect 14550 7466 14616 7500
rect 14650 7466 15254 7500
rect 9278 2226 9284 3162
rect 10220 2226 10226 3162
rect 9278 2220 10226 2226
rect 12740 7318 15254 7466
rect 15312 8072 16016 8078
rect 15312 7380 15318 8072
rect 16010 7380 16016 8072
rect 15312 7374 16016 7380
rect 16074 8000 18584 8136
rect 16074 7966 16692 8000
rect 16726 7966 16792 8000
rect 16826 7966 16892 8000
rect 16926 7966 16992 8000
rect 17026 7966 17092 8000
rect 17126 7966 17192 8000
rect 17226 7966 17980 8000
rect 18014 7966 18080 8000
rect 18114 7966 18180 8000
rect 18214 7966 18280 8000
rect 18314 7966 18380 8000
rect 18414 7966 18480 8000
rect 18514 7966 18584 8000
rect 16074 7900 18584 7966
rect 16074 7866 16692 7900
rect 16726 7866 16792 7900
rect 16826 7866 16892 7900
rect 16926 7866 16992 7900
rect 17026 7866 17092 7900
rect 17126 7866 17192 7900
rect 17226 7866 17980 7900
rect 18014 7866 18080 7900
rect 18114 7866 18180 7900
rect 18214 7866 18280 7900
rect 18314 7866 18380 7900
rect 18414 7866 18480 7900
rect 18514 7866 18584 7900
rect 16074 7800 18584 7866
rect 16074 7766 16692 7800
rect 16726 7766 16792 7800
rect 16826 7766 16892 7800
rect 16926 7766 16992 7800
rect 17026 7766 17092 7800
rect 17126 7766 17192 7800
rect 17226 7766 17980 7800
rect 18014 7766 18080 7800
rect 18114 7766 18180 7800
rect 18214 7766 18280 7800
rect 18314 7766 18380 7800
rect 18414 7766 18480 7800
rect 18514 7766 18584 7800
rect 16074 7700 18584 7766
rect 16074 7666 16692 7700
rect 16726 7666 16792 7700
rect 16826 7666 16892 7700
rect 16926 7666 16992 7700
rect 17026 7666 17092 7700
rect 17126 7666 17192 7700
rect 17226 7666 17980 7700
rect 18014 7666 18080 7700
rect 18114 7666 18180 7700
rect 18214 7666 18280 7700
rect 18314 7666 18380 7700
rect 18414 7666 18480 7700
rect 18514 7666 18584 7700
rect 16074 7600 18584 7666
rect 16074 7566 16692 7600
rect 16726 7566 16792 7600
rect 16826 7566 16892 7600
rect 16926 7566 16992 7600
rect 17026 7566 17092 7600
rect 17126 7566 17192 7600
rect 17226 7566 17980 7600
rect 18014 7566 18080 7600
rect 18114 7566 18180 7600
rect 18214 7566 18280 7600
rect 18314 7566 18380 7600
rect 18414 7566 18480 7600
rect 18514 7566 18584 7600
rect 16074 7500 18584 7566
rect 16074 7466 16692 7500
rect 16726 7466 16792 7500
rect 16826 7466 16892 7500
rect 16926 7466 16992 7500
rect 17026 7466 17092 7500
rect 17126 7466 17192 7500
rect 17226 7466 17980 7500
rect 18014 7466 18080 7500
rect 18114 7466 18180 7500
rect 18214 7466 18280 7500
rect 18314 7466 18380 7500
rect 18414 7466 18480 7500
rect 18514 7466 18584 7500
rect 16074 7318 18584 7466
rect 12740 6712 18584 7318
rect 12740 6678 12828 6712
rect 12862 6678 12928 6712
rect 12962 6678 13028 6712
rect 13062 6678 13128 6712
rect 13162 6678 13228 6712
rect 13262 6678 13328 6712
rect 13362 6678 14116 6712
rect 14150 6678 14216 6712
rect 14250 6678 14316 6712
rect 14350 6678 14416 6712
rect 14450 6678 14516 6712
rect 14550 6678 14616 6712
rect 14650 6678 15404 6712
rect 15438 6678 15504 6712
rect 15538 6678 15604 6712
rect 15638 6678 15704 6712
rect 15738 6678 15804 6712
rect 15838 6678 15904 6712
rect 15938 6678 16692 6712
rect 16726 6678 16792 6712
rect 16826 6678 16892 6712
rect 16926 6678 16992 6712
rect 17026 6678 17092 6712
rect 17126 6678 17192 6712
rect 17226 6678 17980 6712
rect 18014 6678 18080 6712
rect 18114 6678 18180 6712
rect 18214 6678 18280 6712
rect 18314 6678 18380 6712
rect 18414 6678 18480 6712
rect 18514 6678 18584 6712
rect 12740 6612 18584 6678
rect 12740 6578 12828 6612
rect 12862 6578 12928 6612
rect 12962 6578 13028 6612
rect 13062 6578 13128 6612
rect 13162 6578 13228 6612
rect 13262 6578 13328 6612
rect 13362 6578 14116 6612
rect 14150 6578 14216 6612
rect 14250 6578 14316 6612
rect 14350 6578 14416 6612
rect 14450 6578 14516 6612
rect 14550 6578 14616 6612
rect 14650 6578 15404 6612
rect 15438 6578 15504 6612
rect 15538 6578 15604 6612
rect 15638 6578 15704 6612
rect 15738 6578 15804 6612
rect 15838 6578 15904 6612
rect 15938 6578 16692 6612
rect 16726 6578 16792 6612
rect 16826 6578 16892 6612
rect 16926 6578 16992 6612
rect 17026 6578 17092 6612
rect 17126 6578 17192 6612
rect 17226 6578 17980 6612
rect 18014 6578 18080 6612
rect 18114 6578 18180 6612
rect 18214 6578 18280 6612
rect 18314 6578 18380 6612
rect 18414 6578 18480 6612
rect 18514 6578 18584 6612
rect 12740 6512 18584 6578
rect 12740 6478 12828 6512
rect 12862 6478 12928 6512
rect 12962 6478 13028 6512
rect 13062 6478 13128 6512
rect 13162 6478 13228 6512
rect 13262 6478 13328 6512
rect 13362 6478 14116 6512
rect 14150 6478 14216 6512
rect 14250 6478 14316 6512
rect 14350 6478 14416 6512
rect 14450 6478 14516 6512
rect 14550 6478 14616 6512
rect 14650 6478 15404 6512
rect 15438 6478 15504 6512
rect 15538 6478 15604 6512
rect 15638 6478 15704 6512
rect 15738 6478 15804 6512
rect 15838 6478 15904 6512
rect 15938 6478 16692 6512
rect 16726 6478 16792 6512
rect 16826 6478 16892 6512
rect 16926 6478 16992 6512
rect 17026 6478 17092 6512
rect 17126 6478 17192 6512
rect 17226 6478 17980 6512
rect 18014 6478 18080 6512
rect 18114 6478 18180 6512
rect 18214 6478 18280 6512
rect 18314 6478 18380 6512
rect 18414 6478 18480 6512
rect 18514 6478 18584 6512
rect 12740 6412 18584 6478
rect 12740 6378 12828 6412
rect 12862 6378 12928 6412
rect 12962 6378 13028 6412
rect 13062 6378 13128 6412
rect 13162 6378 13228 6412
rect 13262 6378 13328 6412
rect 13362 6378 14116 6412
rect 14150 6378 14216 6412
rect 14250 6378 14316 6412
rect 14350 6378 14416 6412
rect 14450 6378 14516 6412
rect 14550 6378 14616 6412
rect 14650 6378 15404 6412
rect 15438 6378 15504 6412
rect 15538 6378 15604 6412
rect 15638 6378 15704 6412
rect 15738 6378 15804 6412
rect 15838 6378 15904 6412
rect 15938 6378 16692 6412
rect 16726 6378 16792 6412
rect 16826 6378 16892 6412
rect 16926 6378 16992 6412
rect 17026 6378 17092 6412
rect 17126 6378 17192 6412
rect 17226 6378 17980 6412
rect 18014 6378 18080 6412
rect 18114 6378 18180 6412
rect 18214 6378 18280 6412
rect 18314 6378 18380 6412
rect 18414 6378 18480 6412
rect 18514 6378 18584 6412
rect 12740 6312 18584 6378
rect 12740 6278 12828 6312
rect 12862 6278 12928 6312
rect 12962 6278 13028 6312
rect 13062 6278 13128 6312
rect 13162 6278 13228 6312
rect 13262 6278 13328 6312
rect 13362 6278 14116 6312
rect 14150 6278 14216 6312
rect 14250 6278 14316 6312
rect 14350 6278 14416 6312
rect 14450 6278 14516 6312
rect 14550 6278 14616 6312
rect 14650 6278 15404 6312
rect 15438 6278 15504 6312
rect 15538 6278 15604 6312
rect 15638 6278 15704 6312
rect 15738 6278 15804 6312
rect 15838 6278 15904 6312
rect 15938 6278 16692 6312
rect 16726 6278 16792 6312
rect 16826 6278 16892 6312
rect 16926 6278 16992 6312
rect 17026 6278 17092 6312
rect 17126 6278 17192 6312
rect 17226 6278 17980 6312
rect 18014 6278 18080 6312
rect 18114 6278 18180 6312
rect 18214 6278 18280 6312
rect 18314 6278 18380 6312
rect 18414 6278 18480 6312
rect 18514 6278 18584 6312
rect 12740 6212 18584 6278
rect 12740 6178 12828 6212
rect 12862 6178 12928 6212
rect 12962 6178 13028 6212
rect 13062 6178 13128 6212
rect 13162 6178 13228 6212
rect 13262 6178 13328 6212
rect 13362 6178 14116 6212
rect 14150 6178 14216 6212
rect 14250 6178 14316 6212
rect 14350 6178 14416 6212
rect 14450 6178 14516 6212
rect 14550 6178 14616 6212
rect 14650 6178 15404 6212
rect 15438 6178 15504 6212
rect 15538 6178 15604 6212
rect 15638 6178 15704 6212
rect 15738 6178 15804 6212
rect 15838 6178 15904 6212
rect 15938 6178 16692 6212
rect 16726 6178 16792 6212
rect 16826 6178 16892 6212
rect 16926 6178 16992 6212
rect 17026 6178 17092 6212
rect 17126 6178 17192 6212
rect 17226 6178 17980 6212
rect 18014 6178 18080 6212
rect 18114 6178 18180 6212
rect 18214 6178 18280 6212
rect 18314 6178 18380 6212
rect 18414 6178 18480 6212
rect 18514 6178 18584 6212
rect 12740 5424 18584 6178
rect 12740 5390 12828 5424
rect 12862 5390 12928 5424
rect 12962 5390 13028 5424
rect 13062 5390 13128 5424
rect 13162 5390 13228 5424
rect 13262 5390 13328 5424
rect 13362 5390 14116 5424
rect 14150 5390 14216 5424
rect 14250 5390 14316 5424
rect 14350 5390 14416 5424
rect 14450 5390 14516 5424
rect 14550 5390 14616 5424
rect 14650 5390 15404 5424
rect 15438 5390 15504 5424
rect 15538 5390 15604 5424
rect 15638 5390 15704 5424
rect 15738 5390 15804 5424
rect 15838 5390 15904 5424
rect 15938 5390 16692 5424
rect 16726 5390 16792 5424
rect 16826 5390 16892 5424
rect 16926 5390 16992 5424
rect 17026 5390 17092 5424
rect 17126 5390 17192 5424
rect 17226 5390 17980 5424
rect 18014 5390 18080 5424
rect 18114 5390 18180 5424
rect 18214 5390 18280 5424
rect 18314 5390 18380 5424
rect 18414 5390 18480 5424
rect 18514 5390 18584 5424
rect 12740 5324 18584 5390
rect 12740 5290 12828 5324
rect 12862 5290 12928 5324
rect 12962 5290 13028 5324
rect 13062 5290 13128 5324
rect 13162 5290 13228 5324
rect 13262 5290 13328 5324
rect 13362 5290 14116 5324
rect 14150 5290 14216 5324
rect 14250 5290 14316 5324
rect 14350 5290 14416 5324
rect 14450 5290 14516 5324
rect 14550 5290 14616 5324
rect 14650 5290 15404 5324
rect 15438 5290 15504 5324
rect 15538 5290 15604 5324
rect 15638 5290 15704 5324
rect 15738 5290 15804 5324
rect 15838 5290 15904 5324
rect 15938 5290 16692 5324
rect 16726 5290 16792 5324
rect 16826 5290 16892 5324
rect 16926 5290 16992 5324
rect 17026 5290 17092 5324
rect 17126 5290 17192 5324
rect 17226 5290 17980 5324
rect 18014 5290 18080 5324
rect 18114 5290 18180 5324
rect 18214 5290 18280 5324
rect 18314 5290 18380 5324
rect 18414 5290 18480 5324
rect 18514 5290 18584 5324
rect 12740 5224 18584 5290
rect 12740 5190 12828 5224
rect 12862 5190 12928 5224
rect 12962 5190 13028 5224
rect 13062 5190 13128 5224
rect 13162 5190 13228 5224
rect 13262 5190 13328 5224
rect 13362 5190 14116 5224
rect 14150 5190 14216 5224
rect 14250 5190 14316 5224
rect 14350 5190 14416 5224
rect 14450 5190 14516 5224
rect 14550 5190 14616 5224
rect 14650 5190 15404 5224
rect 15438 5190 15504 5224
rect 15538 5190 15604 5224
rect 15638 5190 15704 5224
rect 15738 5190 15804 5224
rect 15838 5190 15904 5224
rect 15938 5190 16692 5224
rect 16726 5190 16792 5224
rect 16826 5190 16892 5224
rect 16926 5190 16992 5224
rect 17026 5190 17092 5224
rect 17126 5190 17192 5224
rect 17226 5190 17980 5224
rect 18014 5190 18080 5224
rect 18114 5190 18180 5224
rect 18214 5190 18280 5224
rect 18314 5190 18380 5224
rect 18414 5190 18480 5224
rect 18514 5190 18584 5224
rect 12740 5124 18584 5190
rect 12740 5090 12828 5124
rect 12862 5090 12928 5124
rect 12962 5090 13028 5124
rect 13062 5090 13128 5124
rect 13162 5090 13228 5124
rect 13262 5090 13328 5124
rect 13362 5090 14116 5124
rect 14150 5090 14216 5124
rect 14250 5090 14316 5124
rect 14350 5090 14416 5124
rect 14450 5090 14516 5124
rect 14550 5090 14616 5124
rect 14650 5090 15404 5124
rect 15438 5090 15504 5124
rect 15538 5090 15604 5124
rect 15638 5090 15704 5124
rect 15738 5090 15804 5124
rect 15838 5090 15904 5124
rect 15938 5090 16692 5124
rect 16726 5090 16792 5124
rect 16826 5090 16892 5124
rect 16926 5090 16992 5124
rect 17026 5090 17092 5124
rect 17126 5090 17192 5124
rect 17226 5090 17980 5124
rect 18014 5090 18080 5124
rect 18114 5090 18180 5124
rect 18214 5090 18280 5124
rect 18314 5090 18380 5124
rect 18414 5090 18480 5124
rect 18514 5090 18584 5124
rect 12740 5024 18584 5090
rect 12740 4990 12828 5024
rect 12862 4990 12928 5024
rect 12962 4990 13028 5024
rect 13062 4990 13128 5024
rect 13162 4990 13228 5024
rect 13262 4990 13328 5024
rect 13362 4990 14116 5024
rect 14150 4990 14216 5024
rect 14250 4990 14316 5024
rect 14350 4990 14416 5024
rect 14450 4990 14516 5024
rect 14550 4990 14616 5024
rect 14650 4990 15404 5024
rect 15438 4990 15504 5024
rect 15538 4990 15604 5024
rect 15638 4990 15704 5024
rect 15738 4990 15804 5024
rect 15838 4990 15904 5024
rect 15938 4990 16692 5024
rect 16726 4990 16792 5024
rect 16826 4990 16892 5024
rect 16926 4990 16992 5024
rect 17026 4990 17092 5024
rect 17126 4990 17192 5024
rect 17226 4990 17980 5024
rect 18014 4990 18080 5024
rect 18114 4990 18180 5024
rect 18214 4990 18280 5024
rect 18314 4990 18380 5024
rect 18414 4990 18480 5024
rect 18514 4990 18584 5024
rect 12740 4924 18584 4990
rect 12740 4890 12828 4924
rect 12862 4890 12928 4924
rect 12962 4890 13028 4924
rect 13062 4890 13128 4924
rect 13162 4890 13228 4924
rect 13262 4890 13328 4924
rect 13362 4890 14116 4924
rect 14150 4890 14216 4924
rect 14250 4890 14316 4924
rect 14350 4890 14416 4924
rect 14450 4890 14516 4924
rect 14550 4890 14616 4924
rect 14650 4890 15404 4924
rect 15438 4890 15504 4924
rect 15538 4890 15604 4924
rect 15638 4890 15704 4924
rect 15738 4890 15804 4924
rect 15838 4890 15904 4924
rect 15938 4890 16692 4924
rect 16726 4890 16792 4924
rect 16826 4890 16892 4924
rect 16926 4890 16992 4924
rect 17026 4890 17092 4924
rect 17126 4890 17192 4924
rect 17226 4890 17980 4924
rect 18014 4890 18080 4924
rect 18114 4890 18180 4924
rect 18214 4890 18280 4924
rect 18314 4890 18380 4924
rect 18414 4890 18480 4924
rect 18514 4890 18584 4924
rect 12740 4136 18584 4890
rect 12740 4102 12828 4136
rect 12862 4102 12928 4136
rect 12962 4102 13028 4136
rect 13062 4102 13128 4136
rect 13162 4102 13228 4136
rect 13262 4102 13328 4136
rect 13362 4102 14116 4136
rect 14150 4102 14216 4136
rect 14250 4102 14316 4136
rect 14350 4102 14416 4136
rect 14450 4102 14516 4136
rect 14550 4102 14616 4136
rect 14650 4102 15404 4136
rect 15438 4102 15504 4136
rect 15538 4102 15604 4136
rect 15638 4102 15704 4136
rect 15738 4102 15804 4136
rect 15838 4102 15904 4136
rect 15938 4102 16692 4136
rect 16726 4102 16792 4136
rect 16826 4102 16892 4136
rect 16926 4102 16992 4136
rect 17026 4102 17092 4136
rect 17126 4102 17192 4136
rect 17226 4102 17980 4136
rect 18014 4102 18080 4136
rect 18114 4102 18180 4136
rect 18214 4102 18280 4136
rect 18314 4102 18380 4136
rect 18414 4102 18480 4136
rect 18514 4102 18584 4136
rect 12740 4036 18584 4102
rect 12740 4002 12828 4036
rect 12862 4002 12928 4036
rect 12962 4002 13028 4036
rect 13062 4002 13128 4036
rect 13162 4002 13228 4036
rect 13262 4002 13328 4036
rect 13362 4002 14116 4036
rect 14150 4002 14216 4036
rect 14250 4002 14316 4036
rect 14350 4002 14416 4036
rect 14450 4002 14516 4036
rect 14550 4002 14616 4036
rect 14650 4002 15404 4036
rect 15438 4002 15504 4036
rect 15538 4002 15604 4036
rect 15638 4002 15704 4036
rect 15738 4002 15804 4036
rect 15838 4002 15904 4036
rect 15938 4002 16692 4036
rect 16726 4002 16792 4036
rect 16826 4002 16892 4036
rect 16926 4002 16992 4036
rect 17026 4002 17092 4036
rect 17126 4002 17192 4036
rect 17226 4002 17980 4036
rect 18014 4002 18080 4036
rect 18114 4002 18180 4036
rect 18214 4002 18280 4036
rect 18314 4002 18380 4036
rect 18414 4002 18480 4036
rect 18514 4002 18584 4036
rect 12740 3936 18584 4002
rect 12740 3902 12828 3936
rect 12862 3902 12928 3936
rect 12962 3902 13028 3936
rect 13062 3902 13128 3936
rect 13162 3902 13228 3936
rect 13262 3902 13328 3936
rect 13362 3902 14116 3936
rect 14150 3902 14216 3936
rect 14250 3902 14316 3936
rect 14350 3902 14416 3936
rect 14450 3902 14516 3936
rect 14550 3902 14616 3936
rect 14650 3902 15404 3936
rect 15438 3902 15504 3936
rect 15538 3902 15604 3936
rect 15638 3902 15704 3936
rect 15738 3902 15804 3936
rect 15838 3902 15904 3936
rect 15938 3902 16692 3936
rect 16726 3902 16792 3936
rect 16826 3902 16892 3936
rect 16926 3902 16992 3936
rect 17026 3902 17092 3936
rect 17126 3902 17192 3936
rect 17226 3902 17980 3936
rect 18014 3902 18080 3936
rect 18114 3902 18180 3936
rect 18214 3902 18280 3936
rect 18314 3902 18380 3936
rect 18414 3902 18480 3936
rect 18514 3902 18584 3936
rect 12740 3836 18584 3902
rect 12740 3802 12828 3836
rect 12862 3802 12928 3836
rect 12962 3802 13028 3836
rect 13062 3802 13128 3836
rect 13162 3802 13228 3836
rect 13262 3802 13328 3836
rect 13362 3802 14116 3836
rect 14150 3802 14216 3836
rect 14250 3802 14316 3836
rect 14350 3802 14416 3836
rect 14450 3802 14516 3836
rect 14550 3802 14616 3836
rect 14650 3802 15404 3836
rect 15438 3802 15504 3836
rect 15538 3802 15604 3836
rect 15638 3802 15704 3836
rect 15738 3802 15804 3836
rect 15838 3802 15904 3836
rect 15938 3802 16692 3836
rect 16726 3802 16792 3836
rect 16826 3802 16892 3836
rect 16926 3802 16992 3836
rect 17026 3802 17092 3836
rect 17126 3802 17192 3836
rect 17226 3802 17980 3836
rect 18014 3802 18080 3836
rect 18114 3802 18180 3836
rect 18214 3802 18280 3836
rect 18314 3802 18380 3836
rect 18414 3802 18480 3836
rect 18514 3802 18584 3836
rect 12740 3736 18584 3802
rect 12740 3702 12828 3736
rect 12862 3702 12928 3736
rect 12962 3702 13028 3736
rect 13062 3702 13128 3736
rect 13162 3702 13228 3736
rect 13262 3702 13328 3736
rect 13362 3702 14116 3736
rect 14150 3702 14216 3736
rect 14250 3702 14316 3736
rect 14350 3702 14416 3736
rect 14450 3702 14516 3736
rect 14550 3702 14616 3736
rect 14650 3702 15404 3736
rect 15438 3702 15504 3736
rect 15538 3702 15604 3736
rect 15638 3702 15704 3736
rect 15738 3702 15804 3736
rect 15838 3702 15904 3736
rect 15938 3702 16692 3736
rect 16726 3702 16792 3736
rect 16826 3702 16892 3736
rect 16926 3702 16992 3736
rect 17026 3702 17092 3736
rect 17126 3702 17192 3736
rect 17226 3702 17980 3736
rect 18014 3702 18080 3736
rect 18114 3702 18180 3736
rect 18214 3702 18280 3736
rect 18314 3702 18380 3736
rect 18414 3702 18480 3736
rect 18514 3702 18584 3736
rect 12740 3636 18584 3702
rect 12740 3602 12828 3636
rect 12862 3602 12928 3636
rect 12962 3602 13028 3636
rect 13062 3602 13128 3636
rect 13162 3602 13228 3636
rect 13262 3602 13328 3636
rect 13362 3602 14116 3636
rect 14150 3602 14216 3636
rect 14250 3602 14316 3636
rect 14350 3602 14416 3636
rect 14450 3602 14516 3636
rect 14550 3602 14616 3636
rect 14650 3602 15404 3636
rect 15438 3602 15504 3636
rect 15538 3602 15604 3636
rect 15638 3602 15704 3636
rect 15738 3602 15804 3636
rect 15838 3602 15904 3636
rect 15938 3602 16692 3636
rect 16726 3602 16792 3636
rect 16826 3602 16892 3636
rect 16926 3602 16992 3636
rect 17026 3602 17092 3636
rect 17126 3602 17192 3636
rect 17226 3602 17980 3636
rect 18014 3602 18080 3636
rect 18114 3602 18180 3636
rect 18214 3602 18280 3636
rect 18314 3602 18380 3636
rect 18414 3602 18480 3636
rect 18514 3602 18584 3636
rect 12740 2916 18584 3602
rect 12740 2908 14036 2916
rect 12740 2232 12742 2908
rect 13424 2240 14036 2908
rect 14718 2848 18584 2916
rect 14718 2814 15404 2848
rect 15438 2814 15504 2848
rect 15538 2814 15604 2848
rect 15638 2814 15704 2848
rect 15738 2814 15804 2848
rect 15838 2814 15904 2848
rect 15938 2814 16692 2848
rect 16726 2814 16792 2848
rect 16826 2814 16892 2848
rect 16926 2814 16992 2848
rect 17026 2814 17092 2848
rect 17126 2814 17192 2848
rect 17226 2814 17980 2848
rect 18014 2814 18080 2848
rect 18114 2814 18180 2848
rect 18214 2814 18280 2848
rect 18314 2814 18380 2848
rect 18414 2814 18480 2848
rect 18514 2814 18584 2848
rect 14718 2748 18584 2814
rect 14718 2714 15404 2748
rect 15438 2714 15504 2748
rect 15538 2714 15604 2748
rect 15638 2714 15704 2748
rect 15738 2714 15804 2748
rect 15838 2714 15904 2748
rect 15938 2714 16692 2748
rect 16726 2714 16792 2748
rect 16826 2714 16892 2748
rect 16926 2714 16992 2748
rect 17026 2714 17092 2748
rect 17126 2714 17192 2748
rect 17226 2714 17980 2748
rect 18014 2714 18080 2748
rect 18114 2714 18180 2748
rect 18214 2714 18280 2748
rect 18314 2714 18380 2748
rect 18414 2714 18480 2748
rect 18514 2714 18584 2748
rect 14718 2648 18584 2714
rect 14718 2614 15404 2648
rect 15438 2614 15504 2648
rect 15538 2614 15604 2648
rect 15638 2614 15704 2648
rect 15738 2614 15804 2648
rect 15838 2614 15904 2648
rect 15938 2614 16692 2648
rect 16726 2614 16792 2648
rect 16826 2614 16892 2648
rect 16926 2614 16992 2648
rect 17026 2614 17092 2648
rect 17126 2614 17192 2648
rect 17226 2614 17980 2648
rect 18014 2614 18080 2648
rect 18114 2614 18180 2648
rect 18214 2614 18280 2648
rect 18314 2614 18380 2648
rect 18414 2614 18480 2648
rect 18514 2614 18584 2648
rect 14718 2548 18584 2614
rect 14718 2514 15404 2548
rect 15438 2514 15504 2548
rect 15538 2514 15604 2548
rect 15638 2514 15704 2548
rect 15738 2514 15804 2548
rect 15838 2514 15904 2548
rect 15938 2514 16692 2548
rect 16726 2514 16792 2548
rect 16826 2514 16892 2548
rect 16926 2514 16992 2548
rect 17026 2514 17092 2548
rect 17126 2514 17192 2548
rect 17226 2514 17980 2548
rect 18014 2514 18080 2548
rect 18114 2514 18180 2548
rect 18214 2514 18280 2548
rect 18314 2514 18380 2548
rect 18414 2514 18480 2548
rect 18514 2514 18584 2548
rect 14718 2448 18584 2514
rect 14718 2414 15404 2448
rect 15438 2414 15504 2448
rect 15538 2414 15604 2448
rect 15638 2414 15704 2448
rect 15738 2414 15804 2448
rect 15838 2414 15904 2448
rect 15938 2414 16692 2448
rect 16726 2414 16792 2448
rect 16826 2414 16892 2448
rect 16926 2414 16992 2448
rect 17026 2414 17092 2448
rect 17126 2414 17192 2448
rect 17226 2414 17980 2448
rect 18014 2414 18080 2448
rect 18114 2414 18180 2448
rect 18214 2414 18280 2448
rect 18314 2414 18380 2448
rect 18414 2414 18480 2448
rect 18514 2414 18584 2448
rect 14718 2348 18584 2414
rect 14718 2314 15404 2348
rect 15438 2314 15504 2348
rect 15538 2314 15604 2348
rect 15638 2314 15704 2348
rect 15738 2314 15804 2348
rect 15838 2314 15904 2348
rect 15938 2314 16692 2348
rect 16726 2314 16792 2348
rect 16826 2314 16892 2348
rect 16926 2314 16992 2348
rect 17026 2314 17092 2348
rect 17126 2314 17192 2348
rect 17226 2314 17980 2348
rect 18014 2314 18080 2348
rect 18114 2314 18180 2348
rect 18214 2314 18280 2348
rect 18314 2314 18380 2348
rect 18414 2314 18480 2348
rect 18514 2314 18584 2348
rect 14718 2240 18584 2314
rect 13424 2232 18584 2240
rect 12740 2218 18584 2232
rect 6950 1659 7130 1662
rect 7690 1660 7736 1712
rect 6922 1653 7130 1659
rect 6922 1619 6934 1653
rect 7118 1619 7130 1653
rect 6922 1613 7130 1619
rect 6950 1522 7130 1613
rect 6950 1402 6970 1522
rect 7110 1402 7130 1522
rect 6950 1382 7130 1402
rect 7278 1653 7736 1660
rect 7278 1619 7392 1653
rect 7576 1619 7736 1653
rect -11762 1238 -11690 1248
rect -15680 1180 -13226 1196
rect -9500 1202 -8348 1302
rect -7930 1322 -7810 1342
rect -7930 1242 -7910 1322
rect -7830 1242 -7810 1322
rect -7930 1222 -7810 1242
rect -7010 1322 -6890 1342
rect -7010 1242 -6990 1322
rect -6910 1242 -6890 1322
rect -7010 1222 -6890 1242
rect -6090 1322 -5970 1342
rect -6090 1242 -6070 1322
rect -5990 1242 -5970 1322
rect -6090 1222 -5970 1242
rect -5170 1322 -5050 1342
rect -5170 1242 -5150 1322
rect -5070 1242 -5050 1322
rect -5170 1222 -5050 1242
rect -4250 1322 -4130 1342
rect -4250 1242 -4230 1322
rect -4150 1242 -4130 1322
rect -2430 1322 -2310 1342
rect -4250 1222 -4130 1242
rect -9500 1102 -9400 1202
rect -9000 1102 -8348 1202
rect -9500 1002 -8348 1102
rect -3590 1202 -2990 1302
rect -2430 1242 -2410 1322
rect -2330 1242 -2310 1322
rect -2430 1222 -2310 1242
rect -1510 1322 -1390 1342
rect -1510 1242 -1490 1322
rect -1410 1242 -1390 1322
rect -1510 1222 -1390 1242
rect -590 1322 -470 1342
rect -590 1242 -570 1322
rect -490 1242 -470 1322
rect -590 1222 -470 1242
rect 330 1322 450 1342
rect 330 1242 350 1322
rect 430 1242 450 1322
rect 330 1222 450 1242
rect 1250 1322 1370 1342
rect 1250 1242 1270 1322
rect 1350 1242 1370 1322
rect 3070 1322 3190 1342
rect 1250 1222 1370 1242
rect -3590 1102 -3490 1202
rect -3090 1102 -2990 1202
rect -3590 1002 -2990 1102
rect 1910 1202 2510 1302
rect 3070 1242 3090 1322
rect 3170 1242 3190 1322
rect 3070 1222 3190 1242
rect 3990 1322 4110 1342
rect 3990 1242 4010 1322
rect 4090 1242 4110 1322
rect 3990 1222 4110 1242
rect 4910 1322 5030 1342
rect 4910 1242 4930 1322
rect 5010 1242 5030 1322
rect 4910 1222 5030 1242
rect 5830 1322 5950 1342
rect 5830 1242 5850 1322
rect 5930 1242 5950 1322
rect 5830 1222 5950 1242
rect 6750 1322 6870 1342
rect 6750 1242 6770 1322
rect 6850 1242 6870 1322
rect 6750 1222 6870 1242
rect 7278 1300 7736 1619
rect 1910 1102 2010 1202
rect 2410 1102 2510 1202
rect 1910 1002 2510 1102
rect 7278 1200 8466 1300
rect 7278 1100 7966 1200
rect 8366 1100 8466 1200
rect 7278 1000 8466 1100
<< via1 >>
rect -21546 25052 -10302 25066
rect -21546 24254 -21532 25052
rect -21532 24254 -10316 25052
rect -10316 24254 -10302 25052
rect -21546 24240 -10302 24254
rect 1720 22968 2278 23526
rect 3344 22968 3902 23526
rect 7434 22968 7992 23526
rect 9888 22968 10446 23526
rect 890 22168 1448 22726
rect 4162 22168 4720 22726
rect 6616 22168 7174 22726
rect 9070 22168 9628 22726
rect 11524 22168 12082 22726
rect 72 21914 630 21926
rect 72 21517 82 21914
rect 82 21517 620 21914
rect 620 21517 630 21914
rect 72 21506 630 21517
rect 890 21914 1448 21926
rect 890 21517 900 21914
rect 900 21517 1438 21914
rect 1438 21517 1448 21914
rect 890 21506 1448 21517
rect 1708 21914 2266 21926
rect 1708 21517 1718 21914
rect 1718 21517 2256 21914
rect 2256 21517 2266 21914
rect 1708 21506 2266 21517
rect 2526 21914 3084 21926
rect 2526 21517 2536 21914
rect 2536 21517 3074 21914
rect 3074 21517 3084 21914
rect 2526 21506 3084 21517
rect 3344 21914 3902 21926
rect 3344 21517 3354 21914
rect 3354 21517 3892 21914
rect 3892 21517 3902 21914
rect 3344 21506 3902 21517
rect 4162 21914 4720 21926
rect 4162 21517 4172 21914
rect 4172 21517 4710 21914
rect 4710 21517 4720 21914
rect 4162 21506 4720 21517
rect 4980 21914 5538 21926
rect 4980 21517 4990 21914
rect 4990 21517 5528 21914
rect 5528 21517 5538 21914
rect 4980 21506 5538 21517
rect 5798 21914 6356 21926
rect 5798 21517 5808 21914
rect 5808 21517 6346 21914
rect 6346 21517 6356 21914
rect 5798 21506 6356 21517
rect 6616 21914 7174 21926
rect 6616 21517 6626 21914
rect 6626 21517 7164 21914
rect 7164 21517 7174 21914
rect 6616 21506 7174 21517
rect 7434 21914 7992 21926
rect 7434 21517 7444 21914
rect 7444 21517 7982 21914
rect 7982 21517 7992 21914
rect 7434 21506 7992 21517
rect 8252 21914 8810 21926
rect 8252 21517 8262 21914
rect 8262 21517 8800 21914
rect 8800 21517 8810 21914
rect 8252 21506 8810 21517
rect 9070 21914 9628 21926
rect 9070 21517 9080 21914
rect 9080 21517 9618 21914
rect 9618 21517 9628 21914
rect 9070 21506 9628 21517
rect 9888 21914 10446 21926
rect 9888 21517 9898 21914
rect 9898 21517 10436 21914
rect 10436 21517 10446 21914
rect 9888 21506 10446 21517
rect 10706 21914 11264 21926
rect 10706 21517 10716 21914
rect 10716 21517 11254 21914
rect 11254 21517 11264 21914
rect 10706 21506 11264 21517
rect 11524 21914 12082 21926
rect 11524 21517 11534 21914
rect 11534 21517 12072 21914
rect 12072 21517 12082 21914
rect 11524 21506 12082 21517
rect 72 20706 630 21264
rect 2526 20706 3084 21264
rect 4980 20706 5538 21264
rect 8252 20706 8810 21264
rect 10706 20706 11264 21264
rect 890 16232 1448 16790
rect 4162 16232 4720 16790
rect 6616 16232 7174 16790
rect 9070 16232 9628 16790
rect 1708 15432 2266 15990
rect 3344 15432 3902 15990
rect 7434 15432 7992 15990
rect 72 15179 630 15190
rect 72 14781 82 15179
rect 82 14781 620 15179
rect 620 14781 630 15179
rect 72 14770 630 14781
rect 890 15179 1448 15190
rect 890 14782 900 15179
rect 900 14782 1438 15179
rect 1438 14782 1448 15179
rect 890 14770 1448 14782
rect 1708 15179 2266 15190
rect 1708 14782 1718 15179
rect 1718 14782 2256 15179
rect 2256 14782 2266 15179
rect 1708 14770 2266 14782
rect 2526 15179 3084 15190
rect 2526 14781 2536 15179
rect 2536 14781 3074 15179
rect 3074 14781 3084 15179
rect 2526 14770 3084 14781
rect 3344 15179 3902 15190
rect 3344 14782 3354 15179
rect 3354 14782 3892 15179
rect 3892 14782 3902 15179
rect 3344 14770 3902 14782
rect 4162 15179 4720 15190
rect 4162 14782 4172 15179
rect 4172 14782 4710 15179
rect 4710 14782 4720 15179
rect 4162 14770 4720 14782
rect 4980 15179 5538 15190
rect 4980 14781 4990 15179
rect 4990 14781 5528 15179
rect 5528 14781 5538 15179
rect 4980 14770 5538 14781
rect 5798 15179 6356 15190
rect 5798 15158 5808 15179
rect 5720 14782 5808 15158
rect 5808 14782 6346 15179
rect 6346 15158 6356 15179
rect 6346 14782 6412 15158
rect 5720 14640 6412 14782
rect 6616 15179 7174 15190
rect 6616 14782 6626 15179
rect 6626 14782 7164 15179
rect 7164 14782 7174 15179
rect 6616 14770 7174 14782
rect 7434 15179 7992 15190
rect 7434 14782 7444 15179
rect 7444 14782 7982 15179
rect 7982 14782 7992 15179
rect 7434 14770 7992 14782
rect 8252 15179 8810 15190
rect 8252 14781 8262 15179
rect 8262 14781 8800 15179
rect 8800 14781 8810 15179
rect 8252 14770 8810 14781
rect 9070 15179 9628 15190
rect 9070 14782 9080 15179
rect 9080 14782 9618 15179
rect 9618 14782 9628 15179
rect 9070 14770 9628 14782
rect 72 13970 630 14528
rect 2526 13970 3084 14528
rect 4980 13970 5538 14528
rect 8252 13970 8810 14528
rect 9810 15179 10502 15190
rect 9810 14782 9898 15179
rect 9898 14782 10436 15179
rect 10436 14782 10502 15179
rect 9810 14498 10502 14782
rect 10628 15179 11320 15190
rect 10628 14782 10716 15179
rect 10716 14782 11254 15179
rect 11254 14782 11320 15179
rect 10628 14498 11320 14782
rect -8384 11410 -6396 11860
rect -9902 10690 -9782 11104
rect -10358 10106 -10238 10398
rect -21364 4944 -21312 4996
rect -19530 4950 -19478 5002
rect -18924 4944 -18730 5002
rect -20446 4738 -20394 4790
rect -19240 1448 -19188 1552
rect -15564 6932 -15420 6986
rect -16136 6792 -15992 6846
rect -14420 6932 -14276 6986
rect -14992 6792 -14848 6846
rect -13276 6932 -13132 6986
rect -13848 6792 -13704 6846
rect -17768 4376 -17716 4630
rect -17208 4376 -17156 4630
rect -16648 4376 -16596 4630
rect -15868 4676 -15816 4780
rect -15296 4676 -15244 4780
rect -15748 4376 -15696 4630
rect -16170 4323 -15962 4340
rect -16170 4289 -16166 4323
rect -16166 4289 -15982 4323
rect -15982 4289 -15962 4323
rect -16170 4282 -15962 4289
rect -15598 4323 -15390 4336
rect -15598 4289 -15594 4323
rect -15594 4289 -15410 4323
rect -15410 4289 -15390 4323
rect -15598 4278 -15390 4289
rect -14724 4676 -14672 4780
rect -14152 4676 -14100 4780
rect -14604 4376 -14552 4630
rect -15026 4323 -14818 4340
rect -15026 4289 -15022 4323
rect -15022 4289 -14838 4323
rect -14838 4289 -14818 4323
rect -15026 4282 -14818 4289
rect -14454 4323 -14246 4340
rect -14454 4289 -14450 4323
rect -14450 4289 -14266 4323
rect -14266 4289 -14246 4323
rect -14454 4282 -14246 4289
rect -13580 4676 -13528 4780
rect -13008 4676 -12956 4780
rect -13460 4376 -13408 4630
rect -12660 4376 -12608 4630
rect -13882 4323 -13674 4340
rect -13882 4289 -13878 4323
rect -13878 4289 -13694 4323
rect -13694 4289 -13674 4323
rect -13882 4282 -13674 4289
rect -13310 4323 -13102 4340
rect -13310 4289 -13306 4323
rect -13306 4289 -13122 4323
rect -13122 4289 -13102 4323
rect -13310 4282 -13102 4289
rect -12100 4376 -12048 4630
rect -8384 10708 -6396 10996
rect -5684 10108 -3696 10396
rect -9902 6926 -9782 7006
rect -10358 6786 -10248 6866
rect -11540 4376 -11488 4630
rect -9490 4376 -9022 4630
rect -18618 1448 -18566 1552
rect -18160 1448 -18108 1552
rect -17584 1448 -17532 1552
rect -17012 1448 -16960 1552
rect -16440 1448 -16388 1552
rect -15868 1448 -15816 1552
rect -15296 1448 -15244 1552
rect -14724 1448 -14672 1552
rect -14152 1448 -14100 1552
rect -13580 1448 -13528 1552
rect -13008 1448 -12956 1552
rect -12436 1448 -12384 1552
rect -11864 1448 -11812 1552
rect -11292 1448 -11240 1552
rect -11182 1448 -11130 1552
rect -10724 1448 -10672 1552
rect -10112 1448 -10060 1552
rect -9490 1388 -9022 1536
rect 9286 12122 10220 12640
rect 5316 11410 7304 11860
rect 5316 10708 7304 10996
rect 2616 10108 4604 10396
rect -18924 1244 -18730 1358
rect -18044 1248 -17992 1352
rect -17472 1248 -17420 1352
rect -16900 1248 -16848 1352
rect -12896 1248 -12844 1352
rect -12324 1248 -12272 1352
rect -11752 1248 -11700 1352
rect -8170 1402 -8030 1522
rect -7710 1402 -7570 1522
rect -7250 1402 -7110 1522
rect -6790 1402 -6650 1522
rect -6330 1402 -6190 1522
rect -5870 1402 -5730 1522
rect -5410 1402 -5270 1522
rect -4950 1402 -4810 1522
rect -4490 1402 -4350 1522
rect -4030 1402 -3890 1522
rect -2670 1402 -2530 1522
rect -2210 1402 -2070 1522
rect -1750 1402 -1610 1522
rect -1290 1402 -1150 1522
rect -830 1402 -690 1522
rect -370 1402 -230 1522
rect 90 1402 230 1522
rect 550 1402 690 1522
rect 1010 1402 1150 1522
rect 1470 1402 1610 1522
rect 2830 1402 2970 1522
rect 3290 1402 3430 1522
rect 3750 1402 3890 1522
rect 4210 1402 4350 1522
rect 4670 1402 4810 1522
rect 5130 1402 5270 1522
rect 5590 1402 5730 1522
rect 6050 1402 6190 1522
rect 6510 1402 6650 1522
rect 10628 11410 11320 11860
rect 11446 15179 12138 15190
rect 11446 14782 11534 15179
rect 11534 14782 12072 15179
rect 12072 14782 12138 15179
rect 11446 14498 12138 14782
rect 11448 10108 12138 10396
rect 10628 7380 11320 8072
rect 9284 2226 10220 3162
rect 15318 8000 16010 8072
rect 15318 7966 15404 8000
rect 15404 7966 15438 8000
rect 15438 7966 15504 8000
rect 15504 7966 15538 8000
rect 15538 7966 15604 8000
rect 15604 7966 15638 8000
rect 15638 7966 15704 8000
rect 15704 7966 15738 8000
rect 15738 7966 15804 8000
rect 15804 7966 15838 8000
rect 15838 7966 15904 8000
rect 15904 7966 15938 8000
rect 15938 7966 16010 8000
rect 15318 7900 16010 7966
rect 15318 7866 15404 7900
rect 15404 7866 15438 7900
rect 15438 7866 15504 7900
rect 15504 7866 15538 7900
rect 15538 7866 15604 7900
rect 15604 7866 15638 7900
rect 15638 7866 15704 7900
rect 15704 7866 15738 7900
rect 15738 7866 15804 7900
rect 15804 7866 15838 7900
rect 15838 7866 15904 7900
rect 15904 7866 15938 7900
rect 15938 7866 16010 7900
rect 15318 7800 16010 7866
rect 15318 7766 15404 7800
rect 15404 7766 15438 7800
rect 15438 7766 15504 7800
rect 15504 7766 15538 7800
rect 15538 7766 15604 7800
rect 15604 7766 15638 7800
rect 15638 7766 15704 7800
rect 15704 7766 15738 7800
rect 15738 7766 15804 7800
rect 15804 7766 15838 7800
rect 15838 7766 15904 7800
rect 15904 7766 15938 7800
rect 15938 7766 16010 7800
rect 15318 7700 16010 7766
rect 15318 7666 15404 7700
rect 15404 7666 15438 7700
rect 15438 7666 15504 7700
rect 15504 7666 15538 7700
rect 15538 7666 15604 7700
rect 15604 7666 15638 7700
rect 15638 7666 15704 7700
rect 15704 7666 15738 7700
rect 15738 7666 15804 7700
rect 15804 7666 15838 7700
rect 15838 7666 15904 7700
rect 15904 7666 15938 7700
rect 15938 7666 16010 7700
rect 15318 7600 16010 7666
rect 15318 7566 15404 7600
rect 15404 7566 15438 7600
rect 15438 7566 15504 7600
rect 15504 7566 15538 7600
rect 15538 7566 15604 7600
rect 15604 7566 15638 7600
rect 15638 7566 15704 7600
rect 15704 7566 15738 7600
rect 15738 7566 15804 7600
rect 15804 7566 15838 7600
rect 15838 7566 15904 7600
rect 15904 7566 15938 7600
rect 15938 7566 16010 7600
rect 15318 7500 16010 7566
rect 15318 7466 15404 7500
rect 15404 7466 15438 7500
rect 15438 7466 15504 7500
rect 15504 7466 15538 7500
rect 15538 7466 15604 7500
rect 15604 7466 15638 7500
rect 15638 7466 15704 7500
rect 15704 7466 15738 7500
rect 15738 7466 15804 7500
rect 15804 7466 15838 7500
rect 15838 7466 15904 7500
rect 15904 7466 15938 7500
rect 15938 7466 16010 7500
rect 15318 7380 16010 7466
rect 12742 2848 13424 2908
rect 12742 2814 12828 2848
rect 12828 2814 12862 2848
rect 12862 2814 12928 2848
rect 12928 2814 12962 2848
rect 12962 2814 13028 2848
rect 13028 2814 13062 2848
rect 13062 2814 13128 2848
rect 13128 2814 13162 2848
rect 13162 2814 13228 2848
rect 13228 2814 13262 2848
rect 13262 2814 13328 2848
rect 13328 2814 13362 2848
rect 13362 2814 13424 2848
rect 12742 2748 13424 2814
rect 12742 2714 12828 2748
rect 12828 2714 12862 2748
rect 12862 2714 12928 2748
rect 12928 2714 12962 2748
rect 12962 2714 13028 2748
rect 13028 2714 13062 2748
rect 13062 2714 13128 2748
rect 13128 2714 13162 2748
rect 13162 2714 13228 2748
rect 13228 2714 13262 2748
rect 13262 2714 13328 2748
rect 13328 2714 13362 2748
rect 13362 2714 13424 2748
rect 12742 2648 13424 2714
rect 12742 2614 12828 2648
rect 12828 2614 12862 2648
rect 12862 2614 12928 2648
rect 12928 2614 12962 2648
rect 12962 2614 13028 2648
rect 13028 2614 13062 2648
rect 13062 2614 13128 2648
rect 13128 2614 13162 2648
rect 13162 2614 13228 2648
rect 13228 2614 13262 2648
rect 13262 2614 13328 2648
rect 13328 2614 13362 2648
rect 13362 2614 13424 2648
rect 12742 2548 13424 2614
rect 12742 2514 12828 2548
rect 12828 2514 12862 2548
rect 12862 2514 12928 2548
rect 12928 2514 12962 2548
rect 12962 2514 13028 2548
rect 13028 2514 13062 2548
rect 13062 2514 13128 2548
rect 13128 2514 13162 2548
rect 13162 2514 13228 2548
rect 13228 2514 13262 2548
rect 13262 2514 13328 2548
rect 13328 2514 13362 2548
rect 13362 2514 13424 2548
rect 12742 2448 13424 2514
rect 12742 2414 12828 2448
rect 12828 2414 12862 2448
rect 12862 2414 12928 2448
rect 12928 2414 12962 2448
rect 12962 2414 13028 2448
rect 13028 2414 13062 2448
rect 13062 2414 13128 2448
rect 13128 2414 13162 2448
rect 13162 2414 13228 2448
rect 13228 2414 13262 2448
rect 13262 2414 13328 2448
rect 13328 2414 13362 2448
rect 13362 2414 13424 2448
rect 12742 2348 13424 2414
rect 12742 2314 12828 2348
rect 12828 2314 12862 2348
rect 12862 2314 12928 2348
rect 12928 2314 12962 2348
rect 12962 2314 13028 2348
rect 13028 2314 13062 2348
rect 13062 2314 13128 2348
rect 13128 2314 13162 2348
rect 13162 2314 13228 2348
rect 13228 2314 13262 2348
rect 13262 2314 13328 2348
rect 13328 2314 13362 2348
rect 13362 2314 13424 2348
rect 12742 2232 13424 2314
rect 14036 2848 14718 2916
rect 14036 2814 14116 2848
rect 14116 2814 14150 2848
rect 14150 2814 14216 2848
rect 14216 2814 14250 2848
rect 14250 2814 14316 2848
rect 14316 2814 14350 2848
rect 14350 2814 14416 2848
rect 14416 2814 14450 2848
rect 14450 2814 14516 2848
rect 14516 2814 14550 2848
rect 14550 2814 14616 2848
rect 14616 2814 14650 2848
rect 14650 2814 14718 2848
rect 14036 2748 14718 2814
rect 14036 2714 14116 2748
rect 14116 2714 14150 2748
rect 14150 2714 14216 2748
rect 14216 2714 14250 2748
rect 14250 2714 14316 2748
rect 14316 2714 14350 2748
rect 14350 2714 14416 2748
rect 14416 2714 14450 2748
rect 14450 2714 14516 2748
rect 14516 2714 14550 2748
rect 14550 2714 14616 2748
rect 14616 2714 14650 2748
rect 14650 2714 14718 2748
rect 14036 2648 14718 2714
rect 14036 2614 14116 2648
rect 14116 2614 14150 2648
rect 14150 2614 14216 2648
rect 14216 2614 14250 2648
rect 14250 2614 14316 2648
rect 14316 2614 14350 2648
rect 14350 2614 14416 2648
rect 14416 2614 14450 2648
rect 14450 2614 14516 2648
rect 14516 2614 14550 2648
rect 14550 2614 14616 2648
rect 14616 2614 14650 2648
rect 14650 2614 14718 2648
rect 14036 2548 14718 2614
rect 14036 2514 14116 2548
rect 14116 2514 14150 2548
rect 14150 2514 14216 2548
rect 14216 2514 14250 2548
rect 14250 2514 14316 2548
rect 14316 2514 14350 2548
rect 14350 2514 14416 2548
rect 14416 2514 14450 2548
rect 14450 2514 14516 2548
rect 14516 2514 14550 2548
rect 14550 2514 14616 2548
rect 14616 2514 14650 2548
rect 14650 2514 14718 2548
rect 14036 2448 14718 2514
rect 14036 2414 14116 2448
rect 14116 2414 14150 2448
rect 14150 2414 14216 2448
rect 14216 2414 14250 2448
rect 14250 2414 14316 2448
rect 14316 2414 14350 2448
rect 14350 2414 14416 2448
rect 14416 2414 14450 2448
rect 14450 2414 14516 2448
rect 14516 2414 14550 2448
rect 14550 2414 14616 2448
rect 14616 2414 14650 2448
rect 14650 2414 14718 2448
rect 14036 2348 14718 2414
rect 14036 2314 14116 2348
rect 14116 2314 14150 2348
rect 14150 2314 14216 2348
rect 14216 2314 14250 2348
rect 14250 2314 14316 2348
rect 14316 2314 14350 2348
rect 14350 2314 14416 2348
rect 14416 2314 14450 2348
rect 14450 2314 14516 2348
rect 14516 2314 14550 2348
rect 14550 2314 14616 2348
rect 14616 2314 14650 2348
rect 14650 2314 14718 2348
rect 14036 2240 14718 2314
rect 6970 1402 7110 1522
rect -7910 1242 -7830 1322
rect -6990 1242 -6910 1322
rect -6070 1242 -5990 1322
rect -5150 1242 -5070 1322
rect -4230 1242 -4150 1322
rect -9400 1102 -9000 1202
rect -2410 1242 -2330 1322
rect -1490 1242 -1410 1322
rect -570 1242 -490 1322
rect 350 1242 430 1322
rect 1270 1242 1350 1322
rect -3490 1102 -3090 1202
rect 3090 1242 3170 1322
rect 4010 1242 4090 1322
rect 4930 1242 5010 1322
rect 5850 1242 5930 1322
rect 6770 1242 6850 1322
rect 2010 1102 2410 1202
rect 7966 1100 8366 1200
<< metal2 >>
rect -21561 25072 -10287 25081
rect -21561 24234 -21552 25072
rect -10296 24234 -10287 25072
rect -21561 24225 -10287 24234
rect 1714 23526 2284 23532
rect 1714 22968 1720 23526
rect 2278 22968 2284 23526
rect 884 22726 1454 22732
rect 884 22168 890 22726
rect 1448 22168 1454 22726
rect 66 21926 636 21932
rect 66 21506 72 21926
rect 630 21506 636 21926
rect 66 21264 636 21506
rect 884 21926 1454 22168
rect 1714 21932 2284 22968
rect 3338 23526 3908 23532
rect 3338 22968 3344 23526
rect 3902 22968 3908 23526
rect 884 21506 890 21926
rect 1448 21506 1454 21926
rect 884 21500 1454 21506
rect 1702 21926 2284 21932
rect 1702 21506 1708 21926
rect 2266 21518 2284 21926
rect 2520 21926 3090 21932
rect 2266 21506 2272 21518
rect 1702 21500 2272 21506
rect 2520 21506 2526 21926
rect 3084 21506 3090 21926
rect 66 20706 72 21264
rect 630 20706 636 21264
rect 66 20700 636 20706
rect 2520 21264 3090 21506
rect 3338 21926 3908 22968
rect 7428 23526 7998 23532
rect 7428 22968 7434 23526
rect 7992 22968 7998 23526
rect 3338 21506 3344 21926
rect 3902 21506 3908 21926
rect 3338 21500 3908 21506
rect 4156 22726 4726 22732
rect 4156 22168 4162 22726
rect 4720 22168 4726 22726
rect 4156 21926 4726 22168
rect 6610 22726 7180 22732
rect 6610 22168 6616 22726
rect 7174 22168 7180 22726
rect 4156 21506 4162 21926
rect 4720 21506 4726 21926
rect 4156 21500 4726 21506
rect 4974 21926 5544 21932
rect 4974 21506 4980 21926
rect 5538 21506 5544 21926
rect 2520 20706 2526 21264
rect 3084 20706 3090 21264
rect 2520 20700 3090 20706
rect 4974 21264 5544 21506
rect 4974 20706 4980 21264
rect 5538 20706 5544 21264
rect 4974 20700 5544 20706
rect 5792 21926 6362 21932
rect 5792 21506 5798 21926
rect 6356 21506 6362 21926
rect 5792 19070 6362 21506
rect 6610 21926 7180 22168
rect 6610 21506 6616 21926
rect 7174 21506 7180 21926
rect 6610 21500 7180 21506
rect 7428 21926 7998 22968
rect 9888 23526 10452 23532
rect 10446 22968 10452 23526
rect 9888 22962 10452 22968
rect 9064 22726 9634 22732
rect 9064 22168 9070 22726
rect 9628 22168 9634 22726
rect 7428 21506 7434 21926
rect 7992 21506 7998 21926
rect 7428 21500 7998 21506
rect 8246 21926 8816 21932
rect 8246 21506 8252 21926
rect 8810 21506 8816 21926
rect 8246 21264 8816 21506
rect 9064 21926 9634 22168
rect 9064 21506 9070 21926
rect 9628 21506 9634 21926
rect 9064 21500 9634 21506
rect 9882 21926 10452 22962
rect 11518 22726 12088 22732
rect 11518 22168 11524 22726
rect 12082 22168 12088 22726
rect 9882 21506 9888 21926
rect 10446 21506 10452 21926
rect 9882 21500 10452 21506
rect 10700 21926 11270 21932
rect 10700 21506 10706 21926
rect 11264 21506 11270 21926
rect 8246 20706 8252 21264
rect 8810 20706 8816 21264
rect 8246 20700 8816 20706
rect 10700 21264 11270 21506
rect 11518 21926 12088 22168
rect 11518 21506 11524 21926
rect 12082 21506 12088 21926
rect 11518 21500 12088 21506
rect 10700 20706 10706 21264
rect 11264 20706 11270 21264
rect 10700 20700 11270 20706
rect 5792 18500 12076 19070
rect 884 16790 1454 16796
rect 884 16232 890 16790
rect 1448 16232 1454 16790
rect 66 15190 636 15196
rect 66 14770 72 15190
rect 630 14770 636 15190
rect 66 14528 636 14770
rect 884 15190 1454 16232
rect 4156 16790 4726 16796
rect 4156 16232 4162 16790
rect 4720 16232 4726 16790
rect 884 14770 890 15190
rect 1448 14770 1454 15190
rect 884 14764 1454 14770
rect 1702 15990 2272 15996
rect 1702 15432 1708 15990
rect 2266 15432 2272 15990
rect 1702 15190 2272 15432
rect 3338 15990 3908 15996
rect 3338 15432 3344 15990
rect 3902 15432 3908 15990
rect 1702 14770 1708 15190
rect 2266 14770 2272 15190
rect 1702 14764 2272 14770
rect 2520 15190 3090 15196
rect 2520 14770 2526 15190
rect 3084 14770 3090 15190
rect 66 13970 72 14528
rect 630 13970 636 14528
rect 2520 14528 3090 14770
rect 3338 15190 3908 15432
rect 3338 14770 3344 15190
rect 3902 14770 3908 15190
rect 3338 14764 3908 14770
rect 4156 15190 4726 16232
rect 6610 16790 7180 16796
rect 6610 16232 6616 16790
rect 7174 16232 7180 16790
rect 4156 14770 4162 15190
rect 4720 14770 4726 15190
rect 4156 14764 4726 14770
rect 4974 15190 5544 15196
rect 4974 14770 4980 15190
rect 5538 14770 5544 15190
rect 5792 15190 6362 15196
rect 5792 15158 5798 15190
rect 6356 15158 6362 15190
rect 6610 15190 7180 16232
rect 9064 16790 9634 16796
rect 9064 16232 9070 16790
rect 9628 16232 9634 16790
rect 2520 13970 2526 14528
rect 3084 13970 3090 14528
rect 4974 14528 5544 14770
rect 4974 13970 4980 14528
rect 5538 13970 5544 14528
rect 5714 14640 5720 15158
rect 6412 14640 6418 15158
rect 6610 14770 6616 15190
rect 7174 14770 7180 15190
rect 6610 14764 7180 14770
rect 7428 15990 7998 15996
rect 7428 15432 7434 15990
rect 7992 15432 7998 15990
rect 7428 15190 7998 15432
rect 7428 14770 7434 15190
rect 7992 14770 7998 15190
rect 7428 14764 7998 14770
rect 8246 15190 8816 15196
rect 8246 14770 8252 15190
rect 8810 14770 8816 15190
rect 66 13964 630 13970
rect 2520 13964 3084 13970
rect 4974 13964 5538 13970
rect 5714 13892 6418 14640
rect 8246 14528 8816 14770
rect 9064 15190 9634 16232
rect 11506 15196 12076 18500
rect 9064 14770 9070 15190
rect 9628 14770 9634 15190
rect 9064 14764 9634 14770
rect 9804 15190 10508 15196
rect 8246 13970 8252 14528
rect 8810 13970 8816 14528
rect 9804 14498 9810 15190
rect 10502 14498 10508 15190
rect 10622 15190 11326 15196
rect 10622 14498 10628 15190
rect 11320 14498 11326 15190
rect 11440 15190 12144 15196
rect 11440 14498 11446 15190
rect 12138 14498 12144 15190
rect 9804 14492 10508 14498
rect 11440 14492 12144 14498
rect 8246 13964 8816 13970
rect 5714 12646 6416 13892
rect 5714 12640 10226 12646
rect 5714 12122 9286 12640
rect 10220 12122 10226 12640
rect 5714 12116 10226 12122
rect -9906 11860 11340 11868
rect -9906 11786 -8384 11860
rect -6396 11786 5316 11860
rect 7304 11786 10628 11860
rect -9906 11110 -9252 11786
rect 11320 11410 11340 11860
rect -9908 11104 -9252 11110
rect -9908 10690 -9902 11104
rect -9782 10802 -9252 11104
rect 11070 10802 11340 11410
rect -9782 10708 -8384 10802
rect -6396 10708 5316 10802
rect 7304 10708 11340 10802
rect -9782 10690 11340 10708
rect -9908 10686 11340 10690
rect -9908 10684 -9776 10686
rect -10364 10398 12144 10402
rect -10364 10106 -10358 10398
rect -10238 10396 12144 10398
rect -10238 10108 -5684 10396
rect -3696 10108 2616 10396
rect 4604 10108 11448 10396
rect 12138 10108 12144 10396
rect -10238 10106 12144 10108
rect -10364 9802 12144 10106
rect 10622 8072 16016 8078
rect 10622 7380 10628 8072
rect 11320 7380 15318 8072
rect 16010 7380 16016 8072
rect 10622 7374 16016 7380
rect -15584 6986 -9902 7006
rect -15584 6932 -15564 6986
rect -15420 6932 -14420 6986
rect -14276 6932 -13276 6986
rect -13132 6932 -9902 6986
rect -15584 6926 -9902 6932
rect -9782 6926 -9776 7006
rect -16156 6846 -10358 6866
rect -16156 6792 -16136 6846
rect -15992 6792 -14992 6846
rect -14848 6792 -13848 6846
rect -13704 6792 -10358 6846
rect -16156 6786 -10358 6792
rect -10248 6786 -10242 6866
rect -21370 5002 -18724 5008
rect -21370 4996 -19530 5002
rect -21370 4944 -21364 4996
rect -21312 4950 -19530 4996
rect -19478 4950 -18924 5002
rect -21312 4944 -18924 4950
rect -18730 4944 -18724 5002
rect -21370 4938 -18724 4944
rect -21317 4790 -12946 4798
rect -21317 4738 -20446 4790
rect -20394 4780 -12946 4790
rect -20394 4738 -15868 4780
rect -21317 4676 -15868 4738
rect -15816 4676 -15296 4780
rect -15244 4676 -14724 4780
rect -14672 4676 -14152 4780
rect -14100 4676 -13580 4780
rect -13528 4676 -13008 4780
rect -12956 4676 -12946 4780
rect -21317 4664 -12946 4676
rect -18620 4630 -9016 4636
rect -18620 4629 -17768 4630
rect -18620 4377 -18600 4629
rect -18000 4377 -17768 4629
rect -18620 4376 -17768 4377
rect -17716 4376 -17208 4630
rect -17156 4376 -16648 4630
rect -16596 4376 -15748 4630
rect -15696 4376 -14604 4630
rect -14552 4376 -13460 4630
rect -13408 4376 -12660 4630
rect -12608 4376 -12100 4630
rect -12048 4376 -11540 4630
rect -11488 4629 -9490 4630
rect -11488 4377 -10109 4629
rect -9509 4377 -9490 4629
rect -11488 4376 -9490 4377
rect -9022 4376 -9016 4630
rect -18620 4370 -9016 4376
rect -16176 4340 -13096 4342
rect -16176 4282 -16170 4340
rect -15962 4336 -15026 4340
rect -15962 4282 -15598 4336
rect -16176 4278 -15598 4282
rect -15390 4282 -15026 4336
rect -14818 4282 -14454 4340
rect -14246 4282 -13882 4340
rect -13674 4282 -13310 4340
rect -13102 4282 -13096 4340
rect -15390 4278 -13096 4282
rect -16176 4276 -13096 4278
rect -16176 4272 -15130 4276
rect 9278 3162 14768 3168
rect 9278 2226 9284 3162
rect 10220 2916 14768 3162
rect 10220 2908 14036 2916
rect 10220 2232 12742 2908
rect 13424 2240 14036 2908
rect 14718 2240 14768 2916
rect 13424 2232 14768 2240
rect 10220 2226 14768 2232
rect 9278 2220 14768 2226
rect -19268 1556 -10002 1562
rect -19268 1442 -19258 1556
rect -10012 1442 -10002 1556
rect -19268 1438 -10002 1442
rect -9496 1536 7130 1542
rect -9496 1388 -9490 1536
rect -9022 1522 7130 1536
rect -9022 1402 -8170 1522
rect -8030 1402 -7710 1522
rect -7570 1402 -7250 1522
rect -7110 1402 -6790 1522
rect -6650 1402 -6330 1522
rect -6190 1402 -5870 1522
rect -5730 1402 -5410 1522
rect -5270 1402 -4950 1522
rect -4810 1402 -4490 1522
rect -4350 1402 -4030 1522
rect -3890 1402 -2670 1522
rect -2530 1402 -2210 1522
rect -2070 1402 -1750 1522
rect -1610 1402 -1290 1522
rect -1150 1402 -830 1522
rect -690 1402 -370 1522
rect -230 1402 90 1522
rect 230 1402 550 1522
rect 690 1402 1010 1522
rect 1150 1402 1470 1522
rect 1610 1402 2830 1522
rect 2970 1402 3290 1522
rect 3430 1402 3750 1522
rect 3890 1402 4210 1522
rect 4350 1402 4670 1522
rect 4810 1402 5130 1522
rect 5270 1402 5590 1522
rect 5730 1402 6050 1522
rect 6190 1402 6510 1522
rect 6650 1402 6970 1522
rect 7110 1402 7130 1522
rect -9022 1388 7130 1402
rect -9496 1382 7130 1388
rect -18930 1362 -18724 1364
rect -18930 1358 -11690 1362
rect -18930 1244 -18924 1358
rect -18730 1352 -11690 1358
rect -18730 1248 -18044 1352
rect -17992 1248 -17472 1352
rect -17420 1248 -16900 1352
rect -16848 1248 -12896 1352
rect -12844 1248 -12324 1352
rect -12272 1248 -11752 1352
rect -11700 1248 -11690 1352
rect -7930 1334 -7810 1342
rect -7010 1334 -6890 1342
rect -6090 1334 -5970 1342
rect -5170 1334 -5050 1342
rect -4250 1334 -4130 1342
rect -2430 1334 -2310 1342
rect -1510 1334 -1390 1342
rect -590 1334 -470 1342
rect 330 1334 450 1342
rect 1250 1334 1370 1342
rect 3070 1334 3190 1342
rect 3990 1334 4110 1342
rect 4910 1334 5030 1342
rect 5830 1334 5950 1342
rect 6750 1334 6870 1342
rect -18730 1244 -11690 1248
rect -18930 1238 -11690 1244
rect -9504 1324 8454 1334
rect -9504 1006 -9494 1324
rect 8444 1300 8454 1324
rect 8444 1006 8466 1300
rect -9504 1000 8466 1006
rect -9504 998 8454 1000
<< via2 >>
rect -21552 25066 -10296 25072
rect -21552 24240 -21546 25066
rect -21546 24240 -10302 25066
rect -10302 24240 -10296 25066
rect -21552 24234 -10296 24240
rect -9252 11410 -8384 11786
rect -8384 11410 -6396 11786
rect -6396 11410 5316 11786
rect 5316 11410 7304 11786
rect 7304 11410 10628 11786
rect 10628 11410 11070 11786
rect -9252 10996 11070 11410
rect -9252 10802 -8384 10996
rect -8384 10802 -6396 10996
rect -6396 10802 5316 10996
rect 5316 10802 7304 10996
rect 7304 10802 11070 10996
rect -18600 4377 -18000 4629
rect -10109 4377 -9509 4629
rect -19258 1552 -10012 1556
rect -19258 1448 -19240 1552
rect -19240 1448 -19188 1552
rect -19188 1448 -18618 1552
rect -18618 1448 -18566 1552
rect -18566 1448 -18160 1552
rect -18160 1448 -18108 1552
rect -18108 1448 -17584 1552
rect -17584 1448 -17532 1552
rect -17532 1448 -17012 1552
rect -17012 1448 -16960 1552
rect -16960 1448 -16440 1552
rect -16440 1448 -16388 1552
rect -16388 1448 -15868 1552
rect -15868 1448 -15816 1552
rect -15816 1448 -15296 1552
rect -15296 1448 -15244 1552
rect -15244 1448 -14724 1552
rect -14724 1448 -14672 1552
rect -14672 1448 -14152 1552
rect -14152 1448 -14100 1552
rect -14100 1448 -13580 1552
rect -13580 1448 -13528 1552
rect -13528 1448 -13008 1552
rect -13008 1448 -12956 1552
rect -12956 1448 -12436 1552
rect -12436 1448 -12384 1552
rect -12384 1448 -11864 1552
rect -11864 1448 -11812 1552
rect -11812 1448 -11292 1552
rect -11292 1448 -11240 1552
rect -11240 1448 -11182 1552
rect -11182 1448 -11130 1552
rect -11130 1448 -10724 1552
rect -10724 1448 -10672 1552
rect -10672 1448 -10112 1552
rect -10112 1448 -10060 1552
rect -10060 1448 -10012 1552
rect -19258 1442 -10012 1448
rect -9494 1322 8444 1324
rect -9494 1242 -7910 1322
rect -7910 1242 -7830 1322
rect -7830 1242 -6990 1322
rect -6990 1242 -6910 1322
rect -6910 1242 -6070 1322
rect -6070 1242 -5990 1322
rect -5990 1242 -5150 1322
rect -5150 1242 -5070 1322
rect -5070 1242 -4230 1322
rect -4230 1242 -4150 1322
rect -4150 1242 -2410 1322
rect -2410 1242 -2330 1322
rect -2330 1242 -1490 1322
rect -1490 1242 -1410 1322
rect -1410 1242 -570 1322
rect -570 1242 -490 1322
rect -490 1242 350 1322
rect 350 1242 430 1322
rect 430 1242 1270 1322
rect 1270 1242 1350 1322
rect 1350 1242 3090 1322
rect 3090 1242 3170 1322
rect 3170 1242 4010 1322
rect 4010 1242 4090 1322
rect 4090 1242 4930 1322
rect 4930 1242 5010 1322
rect 5010 1242 5850 1322
rect 5850 1242 5930 1322
rect 5930 1242 6770 1322
rect 6770 1242 6850 1322
rect 6850 1242 8444 1322
rect -9494 1202 8444 1242
rect -9494 1102 -9400 1202
rect -9400 1102 -9000 1202
rect -9000 1102 -3490 1202
rect -3490 1102 -3090 1202
rect -3090 1102 2010 1202
rect 2010 1102 2410 1202
rect 2410 1200 8444 1202
rect 2410 1102 7966 1200
rect -9494 1100 7966 1102
rect 7966 1100 8366 1200
rect 8366 1100 8444 1200
rect -9494 1006 8444 1100
<< metal3 >>
rect -21567 25081 -10281 25087
rect -21567 24225 -21561 25081
rect -10287 24225 -10281 25081
rect -21567 24219 -10281 24225
rect -17888 16638 -10718 16666
rect -17888 16094 -17273 16638
rect -17209 16094 -16554 16638
rect -16490 16094 -15835 16638
rect -15771 16094 -15116 16638
rect -15052 16094 -14397 16638
rect -14333 16094 -13678 16638
rect -13614 16094 -12959 16638
rect -12895 16094 -12240 16638
rect -12176 16094 -11521 16638
rect -11457 16094 -10802 16638
rect -10738 16094 -10718 16638
rect -17888 15938 -10718 16094
rect -17888 15394 -17273 15938
rect -17209 15394 -16554 15938
rect -16490 15394 -15835 15938
rect -15771 15394 -15116 15938
rect -15052 15394 -14397 15938
rect -14333 15394 -13678 15938
rect -13614 15394 -12959 15938
rect -12895 15394 -12240 15938
rect -12176 15394 -11521 15938
rect -11457 15394 -10802 15938
rect -10738 15394 -10718 15938
rect -17888 15238 -10718 15394
rect -17888 14694 -17273 15238
rect -17209 14694 -16554 15238
rect -16490 14694 -15835 15238
rect -15771 14694 -15116 15238
rect -15052 14694 -14397 15238
rect -14333 14694 -13678 15238
rect -13614 14694 -12959 15238
rect -12895 14694 -12240 15238
rect -12176 14694 -11521 15238
rect -11457 14694 -10802 15238
rect -10738 14694 -10718 15238
rect -17888 14538 -10718 14694
rect -17888 13994 -17273 14538
rect -17209 13994 -16554 14538
rect -16490 13994 -15835 14538
rect -15771 13994 -15116 14538
rect -15052 13994 -14397 14538
rect -14333 13994 -13678 14538
rect -13614 13994 -12959 14538
rect -12895 13994 -12240 14538
rect -12176 13994 -11521 14538
rect -11457 13994 -10802 14538
rect -10738 13994 -10718 14538
rect -17888 13838 -10718 13994
rect -17888 13294 -17273 13838
rect -17209 13294 -16554 13838
rect -16490 13294 -15835 13838
rect -15771 13294 -15116 13838
rect -15052 13294 -14397 13838
rect -14333 13294 -13678 13838
rect -13614 13294 -12959 13838
rect -12895 13294 -12240 13838
rect -12176 13294 -11521 13838
rect -11457 13294 -10802 13838
rect -10738 13294 -10718 13838
rect -17888 13138 -10718 13294
rect -17888 12594 -17273 13138
rect -17209 12594 -16554 13138
rect -16490 12594 -15835 13138
rect -15771 12594 -15116 13138
rect -15052 12594 -14397 13138
rect -14333 12594 -13678 13138
rect -13614 12594 -12959 13138
rect -12895 12594 -12240 13138
rect -12176 12594 -11521 13138
rect -11457 12594 -10802 13138
rect -10738 12594 -10718 13138
rect -17888 12438 -10718 12594
rect -17888 11894 -17273 12438
rect -17209 11894 -16554 12438
rect -16490 11894 -15835 12438
rect -15771 11894 -15116 12438
rect -15052 11894 -14397 12438
rect -14333 11894 -13678 12438
rect -13614 11894 -12959 12438
rect -12895 11894 -12240 12438
rect -12176 11894 -11521 12438
rect -11457 11894 -10802 12438
rect -10738 11894 -10718 12438
rect -17888 11738 -10718 11894
rect -17888 11194 -17273 11738
rect -17209 11194 -16554 11738
rect -16490 11194 -15835 11738
rect -15771 11194 -15116 11738
rect -15052 11194 -14397 11738
rect -14333 11194 -13678 11738
rect -13614 11194 -12959 11738
rect -12895 11194 -12240 11738
rect -12176 11194 -11521 11738
rect -11457 11194 -10802 11738
rect -10738 11194 -10718 11738
rect -17888 11038 -10718 11194
rect -17888 10494 -17273 11038
rect -17209 10494 -16554 11038
rect -16490 10494 -15835 11038
rect -15771 10494 -15116 11038
rect -15052 10494 -14397 11038
rect -14333 10494 -13678 11038
rect -13614 10494 -12959 11038
rect -12895 10494 -12240 11038
rect -12176 10494 -11521 11038
rect -11457 10494 -10802 11038
rect -10738 10494 -10718 11038
rect -9257 11786 11075 11791
rect -9257 10802 -9252 11786
rect 11070 10802 11075 11786
rect -9257 10797 11075 10802
rect -17888 10338 -10718 10494
rect -17888 9794 -17273 10338
rect -17209 9794 -16554 10338
rect -16490 9794 -15835 10338
rect -15771 9794 -15116 10338
rect -15052 9794 -14397 10338
rect -14333 9794 -13678 10338
rect -13614 9794 -12959 10338
rect -12895 9794 -12240 10338
rect -12176 9794 -11521 10338
rect -11457 9794 -10802 10338
rect -10738 9794 -10718 10338
rect -18620 4643 -17980 4649
rect -18620 4363 -18614 4643
rect -17986 4363 -17980 4643
rect -18620 4357 -17980 4363
rect -17888 1562 -10718 9794
rect -10129 4643 -9489 4649
rect -10129 4363 -10123 4643
rect -9495 4363 -9489 4643
rect -10129 4357 -9489 4363
rect -19266 1556 8465 1562
rect -19266 1442 -19258 1556
rect -10012 1442 8465 1556
rect -20266 1340 8465 1442
rect -20266 1324 8466 1340
rect -20266 1006 -9494 1324
rect 8444 1006 8466 1324
rect -20266 1000 8466 1006
rect -17888 966 -10718 1000
<< via3 >>
rect -21561 25072 -10287 25081
rect -21561 24234 -21552 25072
rect -21552 24234 -10296 25072
rect -10296 24234 -10287 25072
rect -21561 24225 -10287 24234
rect -17273 16094 -17209 16638
rect -16554 16094 -16490 16638
rect -15835 16094 -15771 16638
rect -15116 16094 -15052 16638
rect -14397 16094 -14333 16638
rect -13678 16094 -13614 16638
rect -12959 16094 -12895 16638
rect -12240 16094 -12176 16638
rect -11521 16094 -11457 16638
rect -10802 16094 -10738 16638
rect -17273 15394 -17209 15938
rect -16554 15394 -16490 15938
rect -15835 15394 -15771 15938
rect -15116 15394 -15052 15938
rect -14397 15394 -14333 15938
rect -13678 15394 -13614 15938
rect -12959 15394 -12895 15938
rect -12240 15394 -12176 15938
rect -11521 15394 -11457 15938
rect -10802 15394 -10738 15938
rect -17273 14694 -17209 15238
rect -16554 14694 -16490 15238
rect -15835 14694 -15771 15238
rect -15116 14694 -15052 15238
rect -14397 14694 -14333 15238
rect -13678 14694 -13614 15238
rect -12959 14694 -12895 15238
rect -12240 14694 -12176 15238
rect -11521 14694 -11457 15238
rect -10802 14694 -10738 15238
rect -17273 13994 -17209 14538
rect -16554 13994 -16490 14538
rect -15835 13994 -15771 14538
rect -15116 13994 -15052 14538
rect -14397 13994 -14333 14538
rect -13678 13994 -13614 14538
rect -12959 13994 -12895 14538
rect -12240 13994 -12176 14538
rect -11521 13994 -11457 14538
rect -10802 13994 -10738 14538
rect -17273 13294 -17209 13838
rect -16554 13294 -16490 13838
rect -15835 13294 -15771 13838
rect -15116 13294 -15052 13838
rect -14397 13294 -14333 13838
rect -13678 13294 -13614 13838
rect -12959 13294 -12895 13838
rect -12240 13294 -12176 13838
rect -11521 13294 -11457 13838
rect -10802 13294 -10738 13838
rect -17273 12594 -17209 13138
rect -16554 12594 -16490 13138
rect -15835 12594 -15771 13138
rect -15116 12594 -15052 13138
rect -14397 12594 -14333 13138
rect -13678 12594 -13614 13138
rect -12959 12594 -12895 13138
rect -12240 12594 -12176 13138
rect -11521 12594 -11457 13138
rect -10802 12594 -10738 13138
rect -17273 11894 -17209 12438
rect -16554 11894 -16490 12438
rect -15835 11894 -15771 12438
rect -15116 11894 -15052 12438
rect -14397 11894 -14333 12438
rect -13678 11894 -13614 12438
rect -12959 11894 -12895 12438
rect -12240 11894 -12176 12438
rect -11521 11894 -11457 12438
rect -10802 11894 -10738 12438
rect -17273 11194 -17209 11738
rect -16554 11194 -16490 11738
rect -15835 11194 -15771 11738
rect -15116 11194 -15052 11738
rect -14397 11194 -14333 11738
rect -13678 11194 -13614 11738
rect -12959 11194 -12895 11738
rect -12240 11194 -12176 11738
rect -11521 11194 -11457 11738
rect -10802 11194 -10738 11738
rect -17273 10494 -17209 11038
rect -16554 10494 -16490 11038
rect -15835 10494 -15771 11038
rect -15116 10494 -15052 11038
rect -14397 10494 -14333 11038
rect -13678 10494 -13614 11038
rect -12959 10494 -12895 11038
rect -12240 10494 -12176 11038
rect -11521 10494 -11457 11038
rect -10802 10494 -10738 11038
rect -9246 10808 11064 11780
rect -17273 9794 -17209 10338
rect -16554 9794 -16490 10338
rect -15835 9794 -15771 10338
rect -15116 9794 -15052 10338
rect -14397 9794 -14333 10338
rect -13678 9794 -13614 10338
rect -12959 9794 -12895 10338
rect -12240 9794 -12176 10338
rect -11521 9794 -11457 10338
rect -10802 9794 -10738 10338
rect -18614 4629 -17986 4643
rect -18614 4377 -18600 4629
rect -18600 4377 -18000 4629
rect -18000 4377 -17986 4629
rect -18614 4363 -17986 4377
rect -10123 4629 -9495 4643
rect -10123 4377 -10109 4629
rect -10109 4377 -9509 4629
rect -9509 4377 -9495 4629
rect -10123 4363 -9495 4377
<< mimcap >>
rect -17788 16526 -17388 16566
rect -17788 16206 -17748 16526
rect -17428 16206 -17388 16526
rect -17788 16166 -17388 16206
rect -17069 16526 -16669 16566
rect -17069 16206 -17029 16526
rect -16709 16206 -16669 16526
rect -17069 16166 -16669 16206
rect -16350 16526 -15950 16566
rect -16350 16206 -16310 16526
rect -15990 16206 -15950 16526
rect -16350 16166 -15950 16206
rect -15631 16526 -15231 16566
rect -15631 16206 -15591 16526
rect -15271 16206 -15231 16526
rect -15631 16166 -15231 16206
rect -14912 16526 -14512 16566
rect -14912 16206 -14872 16526
rect -14552 16206 -14512 16526
rect -14912 16166 -14512 16206
rect -14193 16526 -13793 16566
rect -14193 16206 -14153 16526
rect -13833 16206 -13793 16526
rect -14193 16166 -13793 16206
rect -13474 16526 -13074 16566
rect -13474 16206 -13434 16526
rect -13114 16206 -13074 16526
rect -13474 16166 -13074 16206
rect -12755 16526 -12355 16566
rect -12755 16206 -12715 16526
rect -12395 16206 -12355 16526
rect -12755 16166 -12355 16206
rect -12036 16526 -11636 16566
rect -12036 16206 -11996 16526
rect -11676 16206 -11636 16526
rect -12036 16166 -11636 16206
rect -11317 16526 -10917 16566
rect -11317 16206 -11277 16526
rect -10957 16206 -10917 16526
rect -11317 16166 -10917 16206
rect -17788 15826 -17388 15866
rect -17788 15506 -17748 15826
rect -17428 15506 -17388 15826
rect -17788 15466 -17388 15506
rect -17069 15826 -16669 15866
rect -17069 15506 -17029 15826
rect -16709 15506 -16669 15826
rect -17069 15466 -16669 15506
rect -16350 15826 -15950 15866
rect -16350 15506 -16310 15826
rect -15990 15506 -15950 15826
rect -16350 15466 -15950 15506
rect -15631 15826 -15231 15866
rect -15631 15506 -15591 15826
rect -15271 15506 -15231 15826
rect -15631 15466 -15231 15506
rect -14912 15826 -14512 15866
rect -14912 15506 -14872 15826
rect -14552 15506 -14512 15826
rect -14912 15466 -14512 15506
rect -14193 15826 -13793 15866
rect -14193 15506 -14153 15826
rect -13833 15506 -13793 15826
rect -14193 15466 -13793 15506
rect -13474 15826 -13074 15866
rect -13474 15506 -13434 15826
rect -13114 15506 -13074 15826
rect -13474 15466 -13074 15506
rect -12755 15826 -12355 15866
rect -12755 15506 -12715 15826
rect -12395 15506 -12355 15826
rect -12755 15466 -12355 15506
rect -12036 15826 -11636 15866
rect -12036 15506 -11996 15826
rect -11676 15506 -11636 15826
rect -12036 15466 -11636 15506
rect -11317 15826 -10917 15866
rect -11317 15506 -11277 15826
rect -10957 15506 -10917 15826
rect -11317 15466 -10917 15506
rect -17788 15126 -17388 15166
rect -17788 14806 -17748 15126
rect -17428 14806 -17388 15126
rect -17788 14766 -17388 14806
rect -17069 15126 -16669 15166
rect -17069 14806 -17029 15126
rect -16709 14806 -16669 15126
rect -17069 14766 -16669 14806
rect -16350 15126 -15950 15166
rect -16350 14806 -16310 15126
rect -15990 14806 -15950 15126
rect -16350 14766 -15950 14806
rect -15631 15126 -15231 15166
rect -15631 14806 -15591 15126
rect -15271 14806 -15231 15126
rect -15631 14766 -15231 14806
rect -14912 15126 -14512 15166
rect -14912 14806 -14872 15126
rect -14552 14806 -14512 15126
rect -14912 14766 -14512 14806
rect -14193 15126 -13793 15166
rect -14193 14806 -14153 15126
rect -13833 14806 -13793 15126
rect -14193 14766 -13793 14806
rect -13474 15126 -13074 15166
rect -13474 14806 -13434 15126
rect -13114 14806 -13074 15126
rect -13474 14766 -13074 14806
rect -12755 15126 -12355 15166
rect -12755 14806 -12715 15126
rect -12395 14806 -12355 15126
rect -12755 14766 -12355 14806
rect -12036 15126 -11636 15166
rect -12036 14806 -11996 15126
rect -11676 14806 -11636 15126
rect -12036 14766 -11636 14806
rect -11317 15126 -10917 15166
rect -11317 14806 -11277 15126
rect -10957 14806 -10917 15126
rect -11317 14766 -10917 14806
rect -17788 14426 -17388 14466
rect -17788 14106 -17748 14426
rect -17428 14106 -17388 14426
rect -17788 14066 -17388 14106
rect -17069 14426 -16669 14466
rect -17069 14106 -17029 14426
rect -16709 14106 -16669 14426
rect -17069 14066 -16669 14106
rect -16350 14426 -15950 14466
rect -16350 14106 -16310 14426
rect -15990 14106 -15950 14426
rect -16350 14066 -15950 14106
rect -15631 14426 -15231 14466
rect -15631 14106 -15591 14426
rect -15271 14106 -15231 14426
rect -15631 14066 -15231 14106
rect -14912 14426 -14512 14466
rect -14912 14106 -14872 14426
rect -14552 14106 -14512 14426
rect -14912 14066 -14512 14106
rect -14193 14426 -13793 14466
rect -14193 14106 -14153 14426
rect -13833 14106 -13793 14426
rect -14193 14066 -13793 14106
rect -13474 14426 -13074 14466
rect -13474 14106 -13434 14426
rect -13114 14106 -13074 14426
rect -13474 14066 -13074 14106
rect -12755 14426 -12355 14466
rect -12755 14106 -12715 14426
rect -12395 14106 -12355 14426
rect -12755 14066 -12355 14106
rect -12036 14426 -11636 14466
rect -12036 14106 -11996 14426
rect -11676 14106 -11636 14426
rect -12036 14066 -11636 14106
rect -11317 14426 -10917 14466
rect -11317 14106 -11277 14426
rect -10957 14106 -10917 14426
rect -11317 14066 -10917 14106
rect -17788 13726 -17388 13766
rect -17788 13406 -17748 13726
rect -17428 13406 -17388 13726
rect -17788 13366 -17388 13406
rect -17069 13726 -16669 13766
rect -17069 13406 -17029 13726
rect -16709 13406 -16669 13726
rect -17069 13366 -16669 13406
rect -16350 13726 -15950 13766
rect -16350 13406 -16310 13726
rect -15990 13406 -15950 13726
rect -16350 13366 -15950 13406
rect -15631 13726 -15231 13766
rect -15631 13406 -15591 13726
rect -15271 13406 -15231 13726
rect -15631 13366 -15231 13406
rect -14912 13726 -14512 13766
rect -14912 13406 -14872 13726
rect -14552 13406 -14512 13726
rect -14912 13366 -14512 13406
rect -14193 13726 -13793 13766
rect -14193 13406 -14153 13726
rect -13833 13406 -13793 13726
rect -14193 13366 -13793 13406
rect -13474 13726 -13074 13766
rect -13474 13406 -13434 13726
rect -13114 13406 -13074 13726
rect -13474 13366 -13074 13406
rect -12755 13726 -12355 13766
rect -12755 13406 -12715 13726
rect -12395 13406 -12355 13726
rect -12755 13366 -12355 13406
rect -12036 13726 -11636 13766
rect -12036 13406 -11996 13726
rect -11676 13406 -11636 13726
rect -12036 13366 -11636 13406
rect -11317 13726 -10917 13766
rect -11317 13406 -11277 13726
rect -10957 13406 -10917 13726
rect -11317 13366 -10917 13406
rect -17788 13026 -17388 13066
rect -17788 12706 -17748 13026
rect -17428 12706 -17388 13026
rect -17788 12666 -17388 12706
rect -17069 13026 -16669 13066
rect -17069 12706 -17029 13026
rect -16709 12706 -16669 13026
rect -17069 12666 -16669 12706
rect -16350 13026 -15950 13066
rect -16350 12706 -16310 13026
rect -15990 12706 -15950 13026
rect -16350 12666 -15950 12706
rect -15631 13026 -15231 13066
rect -15631 12706 -15591 13026
rect -15271 12706 -15231 13026
rect -15631 12666 -15231 12706
rect -14912 13026 -14512 13066
rect -14912 12706 -14872 13026
rect -14552 12706 -14512 13026
rect -14912 12666 -14512 12706
rect -14193 13026 -13793 13066
rect -14193 12706 -14153 13026
rect -13833 12706 -13793 13026
rect -14193 12666 -13793 12706
rect -13474 13026 -13074 13066
rect -13474 12706 -13434 13026
rect -13114 12706 -13074 13026
rect -13474 12666 -13074 12706
rect -12755 13026 -12355 13066
rect -12755 12706 -12715 13026
rect -12395 12706 -12355 13026
rect -12755 12666 -12355 12706
rect -12036 13026 -11636 13066
rect -12036 12706 -11996 13026
rect -11676 12706 -11636 13026
rect -12036 12666 -11636 12706
rect -11317 13026 -10917 13066
rect -11317 12706 -11277 13026
rect -10957 12706 -10917 13026
rect -11317 12666 -10917 12706
rect -17788 12326 -17388 12366
rect -17788 12006 -17748 12326
rect -17428 12006 -17388 12326
rect -17788 11966 -17388 12006
rect -17069 12326 -16669 12366
rect -17069 12006 -17029 12326
rect -16709 12006 -16669 12326
rect -17069 11966 -16669 12006
rect -16350 12326 -15950 12366
rect -16350 12006 -16310 12326
rect -15990 12006 -15950 12326
rect -16350 11966 -15950 12006
rect -15631 12326 -15231 12366
rect -15631 12006 -15591 12326
rect -15271 12006 -15231 12326
rect -15631 11966 -15231 12006
rect -14912 12326 -14512 12366
rect -14912 12006 -14872 12326
rect -14552 12006 -14512 12326
rect -14912 11966 -14512 12006
rect -14193 12326 -13793 12366
rect -14193 12006 -14153 12326
rect -13833 12006 -13793 12326
rect -14193 11966 -13793 12006
rect -13474 12326 -13074 12366
rect -13474 12006 -13434 12326
rect -13114 12006 -13074 12326
rect -13474 11966 -13074 12006
rect -12755 12326 -12355 12366
rect -12755 12006 -12715 12326
rect -12395 12006 -12355 12326
rect -12755 11966 -12355 12006
rect -12036 12326 -11636 12366
rect -12036 12006 -11996 12326
rect -11676 12006 -11636 12326
rect -12036 11966 -11636 12006
rect -11317 12326 -10917 12366
rect -11317 12006 -11277 12326
rect -10957 12006 -10917 12326
rect -11317 11966 -10917 12006
rect -17788 11626 -17388 11666
rect -17788 11306 -17748 11626
rect -17428 11306 -17388 11626
rect -17788 11266 -17388 11306
rect -17069 11626 -16669 11666
rect -17069 11306 -17029 11626
rect -16709 11306 -16669 11626
rect -17069 11266 -16669 11306
rect -16350 11626 -15950 11666
rect -16350 11306 -16310 11626
rect -15990 11306 -15950 11626
rect -16350 11266 -15950 11306
rect -15631 11626 -15231 11666
rect -15631 11306 -15591 11626
rect -15271 11306 -15231 11626
rect -15631 11266 -15231 11306
rect -14912 11626 -14512 11666
rect -14912 11306 -14872 11626
rect -14552 11306 -14512 11626
rect -14912 11266 -14512 11306
rect -14193 11626 -13793 11666
rect -14193 11306 -14153 11626
rect -13833 11306 -13793 11626
rect -14193 11266 -13793 11306
rect -13474 11626 -13074 11666
rect -13474 11306 -13434 11626
rect -13114 11306 -13074 11626
rect -13474 11266 -13074 11306
rect -12755 11626 -12355 11666
rect -12755 11306 -12715 11626
rect -12395 11306 -12355 11626
rect -12755 11266 -12355 11306
rect -12036 11626 -11636 11666
rect -12036 11306 -11996 11626
rect -11676 11306 -11636 11626
rect -12036 11266 -11636 11306
rect -11317 11626 -10917 11666
rect -11317 11306 -11277 11626
rect -10957 11306 -10917 11626
rect -11317 11266 -10917 11306
rect -17788 10926 -17388 10966
rect -17788 10606 -17748 10926
rect -17428 10606 -17388 10926
rect -17788 10566 -17388 10606
rect -17069 10926 -16669 10966
rect -17069 10606 -17029 10926
rect -16709 10606 -16669 10926
rect -17069 10566 -16669 10606
rect -16350 10926 -15950 10966
rect -16350 10606 -16310 10926
rect -15990 10606 -15950 10926
rect -16350 10566 -15950 10606
rect -15631 10926 -15231 10966
rect -15631 10606 -15591 10926
rect -15271 10606 -15231 10926
rect -15631 10566 -15231 10606
rect -14912 10926 -14512 10966
rect -14912 10606 -14872 10926
rect -14552 10606 -14512 10926
rect -14912 10566 -14512 10606
rect -14193 10926 -13793 10966
rect -14193 10606 -14153 10926
rect -13833 10606 -13793 10926
rect -14193 10566 -13793 10606
rect -13474 10926 -13074 10966
rect -13474 10606 -13434 10926
rect -13114 10606 -13074 10926
rect -13474 10566 -13074 10606
rect -12755 10926 -12355 10966
rect -12755 10606 -12715 10926
rect -12395 10606 -12355 10926
rect -12755 10566 -12355 10606
rect -12036 10926 -11636 10966
rect -12036 10606 -11996 10926
rect -11676 10606 -11636 10926
rect -12036 10566 -11636 10606
rect -11317 10926 -10917 10966
rect -11317 10606 -11277 10926
rect -10957 10606 -10917 10926
rect -11317 10566 -10917 10606
rect -17788 10226 -17388 10266
rect -17788 9906 -17748 10226
rect -17428 9906 -17388 10226
rect -17788 9866 -17388 9906
rect -17069 10226 -16669 10266
rect -17069 9906 -17029 10226
rect -16709 9906 -16669 10226
rect -17069 9866 -16669 9906
rect -16350 10226 -15950 10266
rect -16350 9906 -16310 10226
rect -15990 9906 -15950 10226
rect -16350 9866 -15950 9906
rect -15631 10226 -15231 10266
rect -15631 9906 -15591 10226
rect -15271 9906 -15231 10226
rect -15631 9866 -15231 9906
rect -14912 10226 -14512 10266
rect -14912 9906 -14872 10226
rect -14552 9906 -14512 10226
rect -14912 9866 -14512 9906
rect -14193 10226 -13793 10266
rect -14193 9906 -14153 10226
rect -13833 9906 -13793 10226
rect -14193 9866 -13793 9906
rect -13474 10226 -13074 10266
rect -13474 9906 -13434 10226
rect -13114 9906 -13074 10226
rect -13474 9866 -13074 9906
rect -12755 10226 -12355 10266
rect -12755 9906 -12715 10226
rect -12395 9906 -12355 10226
rect -12755 9866 -12355 9906
rect -12036 10226 -11636 10266
rect -12036 9906 -11996 10226
rect -11676 9906 -11636 10226
rect -12036 9866 -11636 9906
rect -11317 10226 -10917 10266
rect -11317 9906 -11277 10226
rect -10957 9906 -10917 10226
rect -11317 9866 -10917 9906
<< mimcapcontact >>
rect -17748 16206 -17428 16526
rect -17029 16206 -16709 16526
rect -16310 16206 -15990 16526
rect -15591 16206 -15271 16526
rect -14872 16206 -14552 16526
rect -14153 16206 -13833 16526
rect -13434 16206 -13114 16526
rect -12715 16206 -12395 16526
rect -11996 16206 -11676 16526
rect -11277 16206 -10957 16526
rect -17748 15506 -17428 15826
rect -17029 15506 -16709 15826
rect -16310 15506 -15990 15826
rect -15591 15506 -15271 15826
rect -14872 15506 -14552 15826
rect -14153 15506 -13833 15826
rect -13434 15506 -13114 15826
rect -12715 15506 -12395 15826
rect -11996 15506 -11676 15826
rect -11277 15506 -10957 15826
rect -17748 14806 -17428 15126
rect -17029 14806 -16709 15126
rect -16310 14806 -15990 15126
rect -15591 14806 -15271 15126
rect -14872 14806 -14552 15126
rect -14153 14806 -13833 15126
rect -13434 14806 -13114 15126
rect -12715 14806 -12395 15126
rect -11996 14806 -11676 15126
rect -11277 14806 -10957 15126
rect -17748 14106 -17428 14426
rect -17029 14106 -16709 14426
rect -16310 14106 -15990 14426
rect -15591 14106 -15271 14426
rect -14872 14106 -14552 14426
rect -14153 14106 -13833 14426
rect -13434 14106 -13114 14426
rect -12715 14106 -12395 14426
rect -11996 14106 -11676 14426
rect -11277 14106 -10957 14426
rect -17748 13406 -17428 13726
rect -17029 13406 -16709 13726
rect -16310 13406 -15990 13726
rect -15591 13406 -15271 13726
rect -14872 13406 -14552 13726
rect -14153 13406 -13833 13726
rect -13434 13406 -13114 13726
rect -12715 13406 -12395 13726
rect -11996 13406 -11676 13726
rect -11277 13406 -10957 13726
rect -17748 12706 -17428 13026
rect -17029 12706 -16709 13026
rect -16310 12706 -15990 13026
rect -15591 12706 -15271 13026
rect -14872 12706 -14552 13026
rect -14153 12706 -13833 13026
rect -13434 12706 -13114 13026
rect -12715 12706 -12395 13026
rect -11996 12706 -11676 13026
rect -11277 12706 -10957 13026
rect -17748 12006 -17428 12326
rect -17029 12006 -16709 12326
rect -16310 12006 -15990 12326
rect -15591 12006 -15271 12326
rect -14872 12006 -14552 12326
rect -14153 12006 -13833 12326
rect -13434 12006 -13114 12326
rect -12715 12006 -12395 12326
rect -11996 12006 -11676 12326
rect -11277 12006 -10957 12326
rect -17748 11306 -17428 11626
rect -17029 11306 -16709 11626
rect -16310 11306 -15990 11626
rect -15591 11306 -15271 11626
rect -14872 11306 -14552 11626
rect -14153 11306 -13833 11626
rect -13434 11306 -13114 11626
rect -12715 11306 -12395 11626
rect -11996 11306 -11676 11626
rect -11277 11306 -10957 11626
rect -17748 10606 -17428 10926
rect -17029 10606 -16709 10926
rect -16310 10606 -15990 10926
rect -15591 10606 -15271 10926
rect -14872 10606 -14552 10926
rect -14153 10606 -13833 10926
rect -13434 10606 -13114 10926
rect -12715 10606 -12395 10926
rect -11996 10606 -11676 10926
rect -11277 10606 -10957 10926
rect -17748 9906 -17428 10226
rect -17029 9906 -16709 10226
rect -16310 9906 -15990 10226
rect -15591 9906 -15271 10226
rect -14872 9906 -14552 10226
rect -14153 9906 -13833 10226
rect -13434 9906 -13114 10226
rect -12715 9906 -12395 10226
rect -11996 9906 -11676 10226
rect -11277 9906 -10957 10226
<< metal4 >>
rect -21578 25081 -10252 25118
rect -21578 24225 -21561 25081
rect -10287 24225 -10252 25081
rect -21578 16956 -10252 24225
rect -21532 16950 -10252 16956
rect -17289 16638 -17193 16654
rect -17788 16526 -17388 16566
rect -17788 16206 -17748 16526
rect -17428 16206 -17388 16526
rect -17788 15826 -17388 16206
rect -17289 16094 -17273 16638
rect -17209 16094 -17193 16638
rect -16570 16638 -16474 16654
rect -17289 16078 -17193 16094
rect -17068 16526 -16668 16566
rect -17068 16206 -17029 16526
rect -16709 16206 -16668 16526
rect -17788 15506 -17748 15826
rect -17428 15506 -17388 15826
rect -17788 15126 -17388 15506
rect -17289 15938 -17193 15954
rect -17289 15394 -17273 15938
rect -17209 15394 -17193 15938
rect -17289 15378 -17193 15394
rect -17068 15826 -16668 16206
rect -16570 16094 -16554 16638
rect -16490 16094 -16474 16638
rect -15851 16638 -15755 16654
rect -16570 16078 -16474 16094
rect -16348 16526 -15948 16566
rect -16348 16206 -16310 16526
rect -15990 16206 -15948 16526
rect -17068 15506 -17029 15826
rect -16709 15506 -16668 15826
rect -17788 14806 -17748 15126
rect -17428 14806 -17388 15126
rect -17788 14426 -17388 14806
rect -17289 15238 -17193 15254
rect -17289 14694 -17273 15238
rect -17209 14694 -17193 15238
rect -17289 14678 -17193 14694
rect -17068 15126 -16668 15506
rect -16570 15938 -16474 15954
rect -16570 15394 -16554 15938
rect -16490 15394 -16474 15938
rect -16570 15378 -16474 15394
rect -16348 15826 -15948 16206
rect -15851 16094 -15835 16638
rect -15771 16094 -15755 16638
rect -15132 16638 -15036 16654
rect -15851 16078 -15755 16094
rect -15628 16526 -15228 16566
rect -15628 16206 -15591 16526
rect -15271 16206 -15228 16526
rect -16348 15506 -16310 15826
rect -15990 15506 -15948 15826
rect -17068 14806 -17029 15126
rect -16709 14806 -16668 15126
rect -17788 14106 -17748 14426
rect -17428 14106 -17388 14426
rect -17788 13726 -17388 14106
rect -17289 14538 -17193 14554
rect -17289 13994 -17273 14538
rect -17209 13994 -17193 14538
rect -17289 13978 -17193 13994
rect -17068 14426 -16668 14806
rect -16570 15238 -16474 15254
rect -16570 14694 -16554 15238
rect -16490 14694 -16474 15238
rect -16570 14678 -16474 14694
rect -16348 15126 -15948 15506
rect -15851 15938 -15755 15954
rect -15851 15394 -15835 15938
rect -15771 15394 -15755 15938
rect -15851 15378 -15755 15394
rect -15628 15826 -15228 16206
rect -15132 16094 -15116 16638
rect -15052 16094 -15036 16638
rect -14413 16638 -14317 16654
rect -15132 16078 -15036 16094
rect -14908 16526 -14508 16566
rect -14908 16206 -14872 16526
rect -14552 16206 -14508 16526
rect -15628 15506 -15591 15826
rect -15271 15506 -15228 15826
rect -16348 14806 -16310 15126
rect -15990 14806 -15948 15126
rect -17068 14106 -17029 14426
rect -16709 14106 -16668 14426
rect -17788 13406 -17748 13726
rect -17428 13406 -17388 13726
rect -17788 13026 -17388 13406
rect -17289 13838 -17193 13854
rect -17289 13294 -17273 13838
rect -17209 13294 -17193 13838
rect -17289 13278 -17193 13294
rect -17068 13726 -16668 14106
rect -16570 14538 -16474 14554
rect -16570 13994 -16554 14538
rect -16490 13994 -16474 14538
rect -16570 13978 -16474 13994
rect -16348 14426 -15948 14806
rect -15851 15238 -15755 15254
rect -15851 14694 -15835 15238
rect -15771 14694 -15755 15238
rect -15851 14678 -15755 14694
rect -15628 15126 -15228 15506
rect -15132 15938 -15036 15954
rect -15132 15394 -15116 15938
rect -15052 15394 -15036 15938
rect -15132 15378 -15036 15394
rect -14908 15826 -14508 16206
rect -14413 16094 -14397 16638
rect -14333 16094 -14317 16638
rect -13694 16638 -13598 16654
rect -14413 16078 -14317 16094
rect -14188 16526 -13788 16566
rect -14188 16206 -14153 16526
rect -13833 16206 -13788 16526
rect -14908 15506 -14872 15826
rect -14552 15506 -14508 15826
rect -15628 14806 -15591 15126
rect -15271 14806 -15228 15126
rect -16348 14106 -16310 14426
rect -15990 14106 -15948 14426
rect -17068 13406 -17029 13726
rect -16709 13406 -16668 13726
rect -17788 12706 -17748 13026
rect -17428 12706 -17388 13026
rect -17788 12326 -17388 12706
rect -17289 13138 -17193 13154
rect -17289 12594 -17273 13138
rect -17209 12594 -17193 13138
rect -17289 12578 -17193 12594
rect -17068 13026 -16668 13406
rect -16570 13838 -16474 13854
rect -16570 13294 -16554 13838
rect -16490 13294 -16474 13838
rect -16570 13278 -16474 13294
rect -16348 13726 -15948 14106
rect -15851 14538 -15755 14554
rect -15851 13994 -15835 14538
rect -15771 13994 -15755 14538
rect -15851 13978 -15755 13994
rect -15628 14426 -15228 14806
rect -15132 15238 -15036 15254
rect -15132 14694 -15116 15238
rect -15052 14694 -15036 15238
rect -15132 14678 -15036 14694
rect -14908 15126 -14508 15506
rect -14413 15938 -14317 15954
rect -14413 15394 -14397 15938
rect -14333 15394 -14317 15938
rect -14413 15378 -14317 15394
rect -14188 15826 -13788 16206
rect -13694 16094 -13678 16638
rect -13614 16094 -13598 16638
rect -12975 16638 -12879 16654
rect -13694 16078 -13598 16094
rect -13468 16526 -13068 16566
rect -13468 16206 -13434 16526
rect -13114 16206 -13068 16526
rect -14188 15506 -14153 15826
rect -13833 15506 -13788 15826
rect -14908 14806 -14872 15126
rect -14552 14806 -14508 15126
rect -15628 14106 -15591 14426
rect -15271 14106 -15228 14426
rect -16348 13406 -16310 13726
rect -15990 13406 -15948 13726
rect -17068 12706 -17029 13026
rect -16709 12706 -16668 13026
rect -17788 12006 -17748 12326
rect -17428 12006 -17388 12326
rect -17788 11626 -17388 12006
rect -17289 12438 -17193 12454
rect -17289 11894 -17273 12438
rect -17209 11894 -17193 12438
rect -17289 11878 -17193 11894
rect -17068 12326 -16668 12706
rect -16570 13138 -16474 13154
rect -16570 12594 -16554 13138
rect -16490 12594 -16474 13138
rect -16570 12578 -16474 12594
rect -16348 13026 -15948 13406
rect -15851 13838 -15755 13854
rect -15851 13294 -15835 13838
rect -15771 13294 -15755 13838
rect -15851 13278 -15755 13294
rect -15628 13726 -15228 14106
rect -15132 14538 -15036 14554
rect -15132 13994 -15116 14538
rect -15052 13994 -15036 14538
rect -15132 13978 -15036 13994
rect -14908 14426 -14508 14806
rect -14413 15238 -14317 15254
rect -14413 14694 -14397 15238
rect -14333 14694 -14317 15238
rect -14413 14678 -14317 14694
rect -14188 15126 -13788 15506
rect -13694 15938 -13598 15954
rect -13694 15394 -13678 15938
rect -13614 15394 -13598 15938
rect -13694 15378 -13598 15394
rect -13468 15826 -13068 16206
rect -12975 16094 -12959 16638
rect -12895 16094 -12879 16638
rect -12256 16638 -12160 16654
rect -12975 16078 -12879 16094
rect -12748 16526 -12348 16566
rect -12748 16206 -12715 16526
rect -12395 16206 -12348 16526
rect -13468 15506 -13434 15826
rect -13114 15506 -13068 15826
rect -14188 14806 -14153 15126
rect -13833 14806 -13788 15126
rect -14908 14106 -14872 14426
rect -14552 14106 -14508 14426
rect -15628 13406 -15591 13726
rect -15271 13406 -15228 13726
rect -16348 12706 -16310 13026
rect -15990 12706 -15948 13026
rect -17068 12006 -17029 12326
rect -16709 12006 -16668 12326
rect -17788 11306 -17748 11626
rect -17428 11306 -17388 11626
rect -17788 10926 -17388 11306
rect -17289 11738 -17193 11754
rect -17289 11194 -17273 11738
rect -17209 11194 -17193 11738
rect -17289 11178 -17193 11194
rect -17068 11626 -16668 12006
rect -16570 12438 -16474 12454
rect -16570 11894 -16554 12438
rect -16490 11894 -16474 12438
rect -16570 11878 -16474 11894
rect -16348 12326 -15948 12706
rect -15851 13138 -15755 13154
rect -15851 12594 -15835 13138
rect -15771 12594 -15755 13138
rect -15851 12578 -15755 12594
rect -15628 13026 -15228 13406
rect -15132 13838 -15036 13854
rect -15132 13294 -15116 13838
rect -15052 13294 -15036 13838
rect -15132 13278 -15036 13294
rect -14908 13726 -14508 14106
rect -14413 14538 -14317 14554
rect -14413 13994 -14397 14538
rect -14333 13994 -14317 14538
rect -14413 13978 -14317 13994
rect -14188 14426 -13788 14806
rect -13694 15238 -13598 15254
rect -13694 14694 -13678 15238
rect -13614 14694 -13598 15238
rect -13694 14678 -13598 14694
rect -13468 15126 -13068 15506
rect -12975 15938 -12879 15954
rect -12975 15394 -12959 15938
rect -12895 15394 -12879 15938
rect -12975 15378 -12879 15394
rect -12748 15826 -12348 16206
rect -12256 16094 -12240 16638
rect -12176 16094 -12160 16638
rect -11537 16638 -11441 16654
rect -12256 16078 -12160 16094
rect -12028 16526 -11628 16566
rect -12028 16206 -11996 16526
rect -11676 16206 -11628 16526
rect -12748 15506 -12715 15826
rect -12395 15506 -12348 15826
rect -13468 14806 -13434 15126
rect -13114 14806 -13068 15126
rect -14188 14106 -14153 14426
rect -13833 14106 -13788 14426
rect -14908 13406 -14872 13726
rect -14552 13406 -14508 13726
rect -15628 12706 -15591 13026
rect -15271 12706 -15228 13026
rect -16348 12006 -16310 12326
rect -15990 12006 -15948 12326
rect -17068 11306 -17029 11626
rect -16709 11306 -16668 11626
rect -17788 10606 -17748 10926
rect -17428 10606 -17388 10926
rect -17788 10226 -17388 10606
rect -17289 11038 -17193 11054
rect -17289 10494 -17273 11038
rect -17209 10494 -17193 11038
rect -17289 10478 -17193 10494
rect -17068 10926 -16668 11306
rect -16570 11738 -16474 11754
rect -16570 11194 -16554 11738
rect -16490 11194 -16474 11738
rect -16570 11178 -16474 11194
rect -16348 11626 -15948 12006
rect -15851 12438 -15755 12454
rect -15851 11894 -15835 12438
rect -15771 11894 -15755 12438
rect -15851 11878 -15755 11894
rect -15628 12326 -15228 12706
rect -15132 13138 -15036 13154
rect -15132 12594 -15116 13138
rect -15052 12594 -15036 13138
rect -15132 12578 -15036 12594
rect -14908 13026 -14508 13406
rect -14413 13838 -14317 13854
rect -14413 13294 -14397 13838
rect -14333 13294 -14317 13838
rect -14413 13278 -14317 13294
rect -14188 13726 -13788 14106
rect -13694 14538 -13598 14554
rect -13694 13994 -13678 14538
rect -13614 13994 -13598 14538
rect -13694 13978 -13598 13994
rect -13468 14426 -13068 14806
rect -12975 15238 -12879 15254
rect -12975 14694 -12959 15238
rect -12895 14694 -12879 15238
rect -12975 14678 -12879 14694
rect -12748 15126 -12348 15506
rect -12256 15938 -12160 15954
rect -12256 15394 -12240 15938
rect -12176 15394 -12160 15938
rect -12256 15378 -12160 15394
rect -12028 15826 -11628 16206
rect -11537 16094 -11521 16638
rect -11457 16094 -11441 16638
rect -10818 16638 -10722 16654
rect -11317 16526 -10908 16566
rect -11317 16206 -11277 16526
rect -10957 16206 -10908 16526
rect -11317 16166 -10908 16206
rect -11537 16078 -11441 16094
rect -12028 15506 -11996 15826
rect -11676 15506 -11628 15826
rect -12748 14806 -12715 15126
rect -12395 14806 -12348 15126
rect -13468 14106 -13434 14426
rect -13114 14106 -13068 14426
rect -14188 13406 -14153 13726
rect -13833 13406 -13788 13726
rect -14908 12706 -14872 13026
rect -14552 12706 -14508 13026
rect -15628 12006 -15591 12326
rect -15271 12006 -15228 12326
rect -16348 11306 -16310 11626
rect -15990 11306 -15948 11626
rect -17068 10606 -17029 10926
rect -16709 10606 -16668 10926
rect -17788 9906 -17748 10226
rect -17428 9906 -17388 10226
rect -17788 9698 -17388 9906
rect -17289 10338 -17193 10354
rect -17289 9794 -17273 10338
rect -17209 9794 -17193 10338
rect -17289 9778 -17193 9794
rect -17068 10226 -16668 10606
rect -16570 11038 -16474 11054
rect -16570 10494 -16554 11038
rect -16490 10494 -16474 11038
rect -16570 10478 -16474 10494
rect -16348 10926 -15948 11306
rect -15851 11738 -15755 11754
rect -15851 11194 -15835 11738
rect -15771 11194 -15755 11738
rect -15851 11178 -15755 11194
rect -15628 11626 -15228 12006
rect -15132 12438 -15036 12454
rect -15132 11894 -15116 12438
rect -15052 11894 -15036 12438
rect -15132 11878 -15036 11894
rect -14908 12326 -14508 12706
rect -14413 13138 -14317 13154
rect -14413 12594 -14397 13138
rect -14333 12594 -14317 13138
rect -14413 12578 -14317 12594
rect -14188 13026 -13788 13406
rect -13694 13838 -13598 13854
rect -13694 13294 -13678 13838
rect -13614 13294 -13598 13838
rect -13694 13278 -13598 13294
rect -13468 13726 -13068 14106
rect -12975 14538 -12879 14554
rect -12975 13994 -12959 14538
rect -12895 13994 -12879 14538
rect -12975 13978 -12879 13994
rect -12748 14426 -12348 14806
rect -12256 15238 -12160 15254
rect -12256 14694 -12240 15238
rect -12176 14694 -12160 15238
rect -12256 14678 -12160 14694
rect -12028 15126 -11628 15506
rect -11537 15938 -11441 15954
rect -11537 15394 -11521 15938
rect -11457 15394 -11441 15938
rect -11537 15378 -11441 15394
rect -11308 15826 -10908 16166
rect -10818 16094 -10802 16638
rect -10738 16094 -10722 16638
rect -10818 16078 -10722 16094
rect -11308 15506 -11277 15826
rect -10957 15506 -10908 15826
rect -12028 14806 -11996 15126
rect -11676 14806 -11628 15126
rect -12748 14106 -12715 14426
rect -12395 14106 -12348 14426
rect -13468 13406 -13434 13726
rect -13114 13406 -13068 13726
rect -14188 12706 -14153 13026
rect -13833 12706 -13788 13026
rect -14908 12006 -14872 12326
rect -14552 12006 -14508 12326
rect -15628 11306 -15591 11626
rect -15271 11306 -15228 11626
rect -16348 10606 -16310 10926
rect -15990 10606 -15948 10926
rect -17068 9906 -17029 10226
rect -16709 9906 -16668 10226
rect -17068 9698 -16668 9906
rect -16570 10338 -16474 10354
rect -16570 9794 -16554 10338
rect -16490 9794 -16474 10338
rect -16570 9778 -16474 9794
rect -16348 10226 -15948 10606
rect -15851 11038 -15755 11054
rect -15851 10494 -15835 11038
rect -15771 10494 -15755 11038
rect -15851 10478 -15755 10494
rect -15628 10926 -15228 11306
rect -15132 11738 -15036 11754
rect -15132 11194 -15116 11738
rect -15052 11194 -15036 11738
rect -15132 11178 -15036 11194
rect -14908 11626 -14508 12006
rect -14413 12438 -14317 12454
rect -14413 11894 -14397 12438
rect -14333 11894 -14317 12438
rect -14413 11878 -14317 11894
rect -14188 12326 -13788 12706
rect -13694 13138 -13598 13154
rect -13694 12594 -13678 13138
rect -13614 12594 -13598 13138
rect -13694 12578 -13598 12594
rect -13468 13026 -13068 13406
rect -12975 13838 -12879 13854
rect -12975 13294 -12959 13838
rect -12895 13294 -12879 13838
rect -12975 13278 -12879 13294
rect -12748 13726 -12348 14106
rect -12256 14538 -12160 14554
rect -12256 13994 -12240 14538
rect -12176 13994 -12160 14538
rect -12256 13978 -12160 13994
rect -12028 14426 -11628 14806
rect -11537 15238 -11441 15254
rect -11537 14694 -11521 15238
rect -11457 14694 -11441 15238
rect -11537 14678 -11441 14694
rect -11308 15126 -10908 15506
rect -10818 15938 -10722 15954
rect -10818 15394 -10802 15938
rect -10738 15394 -10722 15938
rect -10818 15378 -10722 15394
rect -11308 14806 -11277 15126
rect -10957 14806 -10908 15126
rect -12028 14106 -11996 14426
rect -11676 14106 -11628 14426
rect -12748 13406 -12715 13726
rect -12395 13406 -12348 13726
rect -13468 12706 -13434 13026
rect -13114 12706 -13068 13026
rect -14188 12006 -14153 12326
rect -13833 12006 -13788 12326
rect -14908 11306 -14872 11626
rect -14552 11306 -14508 11626
rect -15628 10606 -15591 10926
rect -15271 10606 -15228 10926
rect -16348 9906 -16310 10226
rect -15990 9906 -15948 10226
rect -16348 9698 -15948 9906
rect -15851 10338 -15755 10354
rect -15851 9794 -15835 10338
rect -15771 9794 -15755 10338
rect -15851 9778 -15755 9794
rect -15628 10226 -15228 10606
rect -15132 11038 -15036 11054
rect -15132 10494 -15116 11038
rect -15052 10494 -15036 11038
rect -15132 10478 -15036 10494
rect -14908 10926 -14508 11306
rect -14413 11738 -14317 11754
rect -14413 11194 -14397 11738
rect -14333 11194 -14317 11738
rect -14413 11178 -14317 11194
rect -14188 11626 -13788 12006
rect -13694 12438 -13598 12454
rect -13694 11894 -13678 12438
rect -13614 11894 -13598 12438
rect -13694 11878 -13598 11894
rect -13468 12326 -13068 12706
rect -12975 13138 -12879 13154
rect -12975 12594 -12959 13138
rect -12895 12594 -12879 13138
rect -12975 12578 -12879 12594
rect -12748 13026 -12348 13406
rect -12256 13838 -12160 13854
rect -12256 13294 -12240 13838
rect -12176 13294 -12160 13838
rect -12256 13278 -12160 13294
rect -12028 13726 -11628 14106
rect -11537 14538 -11441 14554
rect -11537 13994 -11521 14538
rect -11457 13994 -11441 14538
rect -11537 13978 -11441 13994
rect -11308 14426 -10908 14806
rect -10818 15238 -10722 15254
rect -10818 14694 -10802 15238
rect -10738 14694 -10722 15238
rect -10818 14678 -10722 14694
rect -11308 14106 -11277 14426
rect -10957 14106 -10908 14426
rect -12028 13406 -11996 13726
rect -11676 13406 -11628 13726
rect -12748 12706 -12715 13026
rect -12395 12706 -12348 13026
rect -13468 12006 -13434 12326
rect -13114 12006 -13068 12326
rect -14188 11306 -14153 11626
rect -13833 11306 -13788 11626
rect -14908 10606 -14872 10926
rect -14552 10606 -14508 10926
rect -15628 9906 -15591 10226
rect -15271 9906 -15228 10226
rect -15628 9698 -15228 9906
rect -15132 10338 -15036 10354
rect -15132 9794 -15116 10338
rect -15052 9794 -15036 10338
rect -15132 9778 -15036 9794
rect -14908 10226 -14508 10606
rect -14413 11038 -14317 11054
rect -14413 10494 -14397 11038
rect -14333 10494 -14317 11038
rect -14413 10478 -14317 10494
rect -14188 10926 -13788 11306
rect -13694 11738 -13598 11754
rect -13694 11194 -13678 11738
rect -13614 11194 -13598 11738
rect -13694 11178 -13598 11194
rect -13468 11626 -13068 12006
rect -12975 12438 -12879 12454
rect -12975 11894 -12959 12438
rect -12895 11894 -12879 12438
rect -12975 11878 -12879 11894
rect -12748 12326 -12348 12706
rect -12256 13138 -12160 13154
rect -12256 12594 -12240 13138
rect -12176 12594 -12160 13138
rect -12256 12578 -12160 12594
rect -12028 13026 -11628 13406
rect -11537 13838 -11441 13854
rect -11537 13294 -11521 13838
rect -11457 13294 -11441 13838
rect -11537 13278 -11441 13294
rect -11308 13726 -10908 14106
rect -10818 14538 -10722 14554
rect -10818 13994 -10802 14538
rect -10738 13994 -10722 14538
rect -10818 13978 -10722 13994
rect -11308 13406 -11277 13726
rect -10957 13406 -10908 13726
rect -12028 12706 -11996 13026
rect -11676 12706 -11628 13026
rect -12748 12006 -12715 12326
rect -12395 12006 -12348 12326
rect -13468 11306 -13434 11626
rect -13114 11306 -13068 11626
rect -14188 10606 -14153 10926
rect -13833 10606 -13788 10926
rect -14908 9906 -14872 10226
rect -14552 9906 -14508 10226
rect -14908 9698 -14508 9906
rect -14413 10338 -14317 10354
rect -14413 9794 -14397 10338
rect -14333 9794 -14317 10338
rect -14413 9778 -14317 9794
rect -14188 10226 -13788 10606
rect -13694 11038 -13598 11054
rect -13694 10494 -13678 11038
rect -13614 10494 -13598 11038
rect -13694 10478 -13598 10494
rect -13468 10926 -13068 11306
rect -12975 11738 -12879 11754
rect -12975 11194 -12959 11738
rect -12895 11194 -12879 11738
rect -12975 11178 -12879 11194
rect -12748 11626 -12348 12006
rect -12256 12438 -12160 12454
rect -12256 11894 -12240 12438
rect -12176 11894 -12160 12438
rect -12256 11878 -12160 11894
rect -12028 12326 -11628 12706
rect -11537 13138 -11441 13154
rect -11537 12594 -11521 13138
rect -11457 12594 -11441 13138
rect -11537 12578 -11441 12594
rect -11308 13026 -10908 13406
rect -10818 13838 -10722 13854
rect -10818 13294 -10802 13838
rect -10738 13294 -10722 13838
rect -10818 13278 -10722 13294
rect -11308 12706 -11277 13026
rect -10957 12706 -10908 13026
rect -12028 12006 -11996 12326
rect -11676 12006 -11628 12326
rect -12748 11306 -12715 11626
rect -12395 11306 -12348 11626
rect -13468 10606 -13434 10926
rect -13114 10606 -13068 10926
rect -14188 9906 -14153 10226
rect -13833 9906 -13788 10226
rect -14188 9698 -13788 9906
rect -13694 10338 -13598 10354
rect -13694 9794 -13678 10338
rect -13614 9794 -13598 10338
rect -13694 9778 -13598 9794
rect -13468 10226 -13068 10606
rect -12975 11038 -12879 11054
rect -12975 10494 -12959 11038
rect -12895 10494 -12879 11038
rect -12975 10478 -12879 10494
rect -12748 10926 -12348 11306
rect -12256 11738 -12160 11754
rect -12256 11194 -12240 11738
rect -12176 11194 -12160 11738
rect -12256 11178 -12160 11194
rect -12028 11626 -11628 12006
rect -11537 12438 -11441 12454
rect -11537 11894 -11521 12438
rect -11457 11894 -11441 12438
rect -11537 11878 -11441 11894
rect -11308 12326 -10908 12706
rect -10818 13138 -10722 13154
rect -10818 12594 -10802 13138
rect -10738 12594 -10722 13138
rect -10818 12578 -10722 12594
rect -11308 12006 -11277 12326
rect -10957 12006 -10908 12326
rect -12028 11306 -11996 11626
rect -11676 11306 -11628 11626
rect -12748 10606 -12715 10926
rect -12395 10606 -12348 10926
rect -13468 9906 -13434 10226
rect -13114 9906 -13068 10226
rect -13468 9698 -13068 9906
rect -12975 10338 -12879 10354
rect -12975 9794 -12959 10338
rect -12895 9794 -12879 10338
rect -12975 9778 -12879 9794
rect -12748 10226 -12348 10606
rect -12256 11038 -12160 11054
rect -12256 10494 -12240 11038
rect -12176 10494 -12160 11038
rect -12256 10478 -12160 10494
rect -12028 10926 -11628 11306
rect -11537 11738 -11441 11754
rect -11537 11194 -11521 11738
rect -11457 11194 -11441 11738
rect -11537 11178 -11441 11194
rect -11308 11626 -10908 12006
rect -10818 12438 -10722 12454
rect -10818 11894 -10802 12438
rect -10738 11894 -10722 12438
rect -10818 11878 -10722 11894
rect -9247 11780 11065 11781
rect -11308 11306 -11277 11626
rect -10957 11306 -10908 11626
rect -12028 10606 -11996 10926
rect -11676 10606 -11628 10926
rect -12748 9906 -12715 10226
rect -12395 9906 -12348 10226
rect -12748 9698 -12348 9906
rect -12256 10338 -12160 10354
rect -12256 9794 -12240 10338
rect -12176 9794 -12160 10338
rect -12256 9778 -12160 9794
rect -12028 10226 -11628 10606
rect -11537 11038 -11441 11054
rect -11537 10494 -11521 11038
rect -11457 10494 -11441 11038
rect -11537 10478 -11441 10494
rect -11308 10926 -10908 11306
rect -10818 11738 -10722 11754
rect -10818 11194 -10802 11738
rect -10738 11194 -10722 11738
rect -10818 11178 -10722 11194
rect -11308 10606 -11277 10926
rect -10957 10606 -10908 10926
rect -12028 9906 -11996 10226
rect -11676 9906 -11628 10226
rect -12028 9698 -11628 9906
rect -11537 10338 -11441 10354
rect -11537 9794 -11521 10338
rect -11457 9794 -11441 10338
rect -11537 9778 -11441 9794
rect -11308 10226 -10908 10606
rect -10818 11038 -10722 11054
rect -10818 10494 -10802 11038
rect -10738 10494 -10722 11038
rect -9247 10808 -9246 11780
rect 11064 10808 11065 11780
rect -9247 10807 11065 10808
rect -10818 10478 -10722 10494
rect -11308 9906 -11277 10226
rect -10957 9906 -10908 10226
rect -11308 9706 -10908 9906
rect -10818 10338 -10722 10354
rect -10818 9794 -10802 10338
rect -10738 9794 -10722 10338
rect -10818 9778 -10722 9794
rect -11308 9698 -10888 9706
rect -17788 9691 -10888 9698
rect -18614 4645 -9482 9691
rect -18616 4643 -9482 4645
rect -18616 4363 -18614 4643
rect -17986 4363 -10123 4643
rect -9495 4363 -9482 4643
rect -18616 4361 -9482 4363
rect -18614 4360 -9482 4361
<< via4 >>
rect -9246 10808 11064 11780
<< mimcap2 >>
rect -21478 23766 -21078 23806
rect -21478 23446 -21438 23766
rect -21118 23446 -21078 23766
rect -21478 23406 -21078 23446
rect -20356 23766 -19956 23806
rect -20356 23446 -20316 23766
rect -19996 23446 -19956 23766
rect -20356 23406 -19956 23446
rect -19234 23766 -18834 23806
rect -19234 23446 -19194 23766
rect -18874 23446 -18834 23766
rect -19234 23406 -18834 23446
rect -18112 23766 -17712 23806
rect -18112 23446 -18072 23766
rect -17752 23446 -17712 23766
rect -18112 23406 -17712 23446
rect -16990 23766 -16590 23806
rect -16990 23446 -16950 23766
rect -16630 23446 -16590 23766
rect -16990 23406 -16590 23446
rect -15868 23766 -15468 23806
rect -15868 23446 -15828 23766
rect -15508 23446 -15468 23766
rect -15868 23406 -15468 23446
rect -14746 23766 -14346 23806
rect -14746 23446 -14706 23766
rect -14386 23446 -14346 23766
rect -14746 23406 -14346 23446
rect -13624 23766 -13224 23806
rect -13624 23446 -13584 23766
rect -13264 23446 -13224 23766
rect -13624 23406 -13224 23446
rect -12502 23766 -12102 23806
rect -12502 23446 -12462 23766
rect -12142 23446 -12102 23766
rect -12502 23406 -12102 23446
rect -11380 23766 -10980 23806
rect -11380 23446 -11340 23766
rect -11020 23446 -10980 23766
rect -11380 23406 -10980 23446
rect -21478 23066 -21078 23106
rect -21478 22746 -21438 23066
rect -21118 22746 -21078 23066
rect -21478 22706 -21078 22746
rect -20356 23066 -19956 23106
rect -20356 22746 -20316 23066
rect -19996 22746 -19956 23066
rect -20356 22706 -19956 22746
rect -19234 23066 -18834 23106
rect -19234 22746 -19194 23066
rect -18874 22746 -18834 23066
rect -19234 22706 -18834 22746
rect -18112 23066 -17712 23106
rect -18112 22746 -18072 23066
rect -17752 22746 -17712 23066
rect -18112 22706 -17712 22746
rect -16990 23066 -16590 23106
rect -16990 22746 -16950 23066
rect -16630 22746 -16590 23066
rect -16990 22706 -16590 22746
rect -15868 23066 -15468 23106
rect -15868 22746 -15828 23066
rect -15508 22746 -15468 23066
rect -15868 22706 -15468 22746
rect -14746 23066 -14346 23106
rect -14746 22746 -14706 23066
rect -14386 22746 -14346 23066
rect -14746 22706 -14346 22746
rect -13624 23066 -13224 23106
rect -13624 22746 -13584 23066
rect -13264 22746 -13224 23066
rect -13624 22706 -13224 22746
rect -12502 23066 -12102 23106
rect -12502 22746 -12462 23066
rect -12142 22746 -12102 23066
rect -12502 22706 -12102 22746
rect -11380 23066 -10980 23106
rect -11380 22746 -11340 23066
rect -11020 22746 -10980 23066
rect -11380 22706 -10980 22746
rect -21478 22366 -21078 22406
rect -21478 22046 -21438 22366
rect -21118 22046 -21078 22366
rect -21478 22006 -21078 22046
rect -20356 22366 -19956 22406
rect -20356 22046 -20316 22366
rect -19996 22046 -19956 22366
rect -20356 22006 -19956 22046
rect -19234 22366 -18834 22406
rect -19234 22046 -19194 22366
rect -18874 22046 -18834 22366
rect -19234 22006 -18834 22046
rect -18112 22366 -17712 22406
rect -18112 22046 -18072 22366
rect -17752 22046 -17712 22366
rect -18112 22006 -17712 22046
rect -16990 22366 -16590 22406
rect -16990 22046 -16950 22366
rect -16630 22046 -16590 22366
rect -16990 22006 -16590 22046
rect -15868 22366 -15468 22406
rect -15868 22046 -15828 22366
rect -15508 22046 -15468 22366
rect -15868 22006 -15468 22046
rect -14746 22366 -14346 22406
rect -14746 22046 -14706 22366
rect -14386 22046 -14346 22366
rect -14746 22006 -14346 22046
rect -13624 22366 -13224 22406
rect -13624 22046 -13584 22366
rect -13264 22046 -13224 22366
rect -13624 22006 -13224 22046
rect -12502 22366 -12102 22406
rect -12502 22046 -12462 22366
rect -12142 22046 -12102 22366
rect -12502 22006 -12102 22046
rect -11380 22366 -10980 22406
rect -11380 22046 -11340 22366
rect -11020 22046 -10980 22366
rect -11380 22006 -10980 22046
rect -21478 21666 -21078 21706
rect -21478 21346 -21438 21666
rect -21118 21346 -21078 21666
rect -21478 21306 -21078 21346
rect -20356 21666 -19956 21706
rect -20356 21346 -20316 21666
rect -19996 21346 -19956 21666
rect -20356 21306 -19956 21346
rect -19234 21666 -18834 21706
rect -19234 21346 -19194 21666
rect -18874 21346 -18834 21666
rect -19234 21306 -18834 21346
rect -18112 21666 -17712 21706
rect -18112 21346 -18072 21666
rect -17752 21346 -17712 21666
rect -18112 21306 -17712 21346
rect -16990 21666 -16590 21706
rect -16990 21346 -16950 21666
rect -16630 21346 -16590 21666
rect -16990 21306 -16590 21346
rect -15868 21666 -15468 21706
rect -15868 21346 -15828 21666
rect -15508 21346 -15468 21666
rect -15868 21306 -15468 21346
rect -14746 21666 -14346 21706
rect -14746 21346 -14706 21666
rect -14386 21346 -14346 21666
rect -14746 21306 -14346 21346
rect -13624 21666 -13224 21706
rect -13624 21346 -13584 21666
rect -13264 21346 -13224 21666
rect -13624 21306 -13224 21346
rect -12502 21666 -12102 21706
rect -12502 21346 -12462 21666
rect -12142 21346 -12102 21666
rect -12502 21306 -12102 21346
rect -11380 21666 -10980 21706
rect -11380 21346 -11340 21666
rect -11020 21346 -10980 21666
rect -11380 21306 -10980 21346
rect -21478 20966 -21078 21006
rect -21478 20646 -21438 20966
rect -21118 20646 -21078 20966
rect -21478 20606 -21078 20646
rect -20356 20966 -19956 21006
rect -20356 20646 -20316 20966
rect -19996 20646 -19956 20966
rect -20356 20606 -19956 20646
rect -19234 20966 -18834 21006
rect -19234 20646 -19194 20966
rect -18874 20646 -18834 20966
rect -19234 20606 -18834 20646
rect -18112 20966 -17712 21006
rect -18112 20646 -18072 20966
rect -17752 20646 -17712 20966
rect -18112 20606 -17712 20646
rect -16990 20966 -16590 21006
rect -16990 20646 -16950 20966
rect -16630 20646 -16590 20966
rect -16990 20606 -16590 20646
rect -15868 20966 -15468 21006
rect -15868 20646 -15828 20966
rect -15508 20646 -15468 20966
rect -15868 20606 -15468 20646
rect -14746 20966 -14346 21006
rect -14746 20646 -14706 20966
rect -14386 20646 -14346 20966
rect -14746 20606 -14346 20646
rect -13624 20966 -13224 21006
rect -13624 20646 -13584 20966
rect -13264 20646 -13224 20966
rect -13624 20606 -13224 20646
rect -12502 20966 -12102 21006
rect -12502 20646 -12462 20966
rect -12142 20646 -12102 20966
rect -12502 20606 -12102 20646
rect -11380 20966 -10980 21006
rect -11380 20646 -11340 20966
rect -11020 20646 -10980 20966
rect -11380 20606 -10980 20646
rect -21478 20266 -21078 20306
rect -21478 19946 -21438 20266
rect -21118 19946 -21078 20266
rect -21478 19906 -21078 19946
rect -20356 20266 -19956 20306
rect -20356 19946 -20316 20266
rect -19996 19946 -19956 20266
rect -20356 19906 -19956 19946
rect -19234 20266 -18834 20306
rect -19234 19946 -19194 20266
rect -18874 19946 -18834 20266
rect -19234 19906 -18834 19946
rect -18112 20266 -17712 20306
rect -18112 19946 -18072 20266
rect -17752 19946 -17712 20266
rect -18112 19906 -17712 19946
rect -16990 20266 -16590 20306
rect -16990 19946 -16950 20266
rect -16630 19946 -16590 20266
rect -16990 19906 -16590 19946
rect -15868 20266 -15468 20306
rect -15868 19946 -15828 20266
rect -15508 19946 -15468 20266
rect -15868 19906 -15468 19946
rect -14746 20266 -14346 20306
rect -14746 19946 -14706 20266
rect -14386 19946 -14346 20266
rect -14746 19906 -14346 19946
rect -13624 20266 -13224 20306
rect -13624 19946 -13584 20266
rect -13264 19946 -13224 20266
rect -13624 19906 -13224 19946
rect -12502 20266 -12102 20306
rect -12502 19946 -12462 20266
rect -12142 19946 -12102 20266
rect -12502 19906 -12102 19946
rect -11380 20266 -10980 20306
rect -11380 19946 -11340 20266
rect -11020 19946 -10980 20266
rect -11380 19906 -10980 19946
rect -21478 19566 -21078 19606
rect -21478 19246 -21438 19566
rect -21118 19246 -21078 19566
rect -21478 19206 -21078 19246
rect -20356 19566 -19956 19606
rect -20356 19246 -20316 19566
rect -19996 19246 -19956 19566
rect -20356 19206 -19956 19246
rect -19234 19566 -18834 19606
rect -19234 19246 -19194 19566
rect -18874 19246 -18834 19566
rect -19234 19206 -18834 19246
rect -18112 19566 -17712 19606
rect -18112 19246 -18072 19566
rect -17752 19246 -17712 19566
rect -18112 19206 -17712 19246
rect -16990 19566 -16590 19606
rect -16990 19246 -16950 19566
rect -16630 19246 -16590 19566
rect -16990 19206 -16590 19246
rect -15868 19566 -15468 19606
rect -15868 19246 -15828 19566
rect -15508 19246 -15468 19566
rect -15868 19206 -15468 19246
rect -14746 19566 -14346 19606
rect -14746 19246 -14706 19566
rect -14386 19246 -14346 19566
rect -14746 19206 -14346 19246
rect -13624 19566 -13224 19606
rect -13624 19246 -13584 19566
rect -13264 19246 -13224 19566
rect -13624 19206 -13224 19246
rect -12502 19566 -12102 19606
rect -12502 19246 -12462 19566
rect -12142 19246 -12102 19566
rect -12502 19206 -12102 19246
rect -11380 19566 -10980 19606
rect -11380 19246 -11340 19566
rect -11020 19246 -10980 19566
rect -11380 19206 -10980 19246
rect -21478 18866 -21078 18906
rect -21478 18546 -21438 18866
rect -21118 18546 -21078 18866
rect -21478 18506 -21078 18546
rect -20356 18866 -19956 18906
rect -20356 18546 -20316 18866
rect -19996 18546 -19956 18866
rect -20356 18506 -19956 18546
rect -19234 18866 -18834 18906
rect -19234 18546 -19194 18866
rect -18874 18546 -18834 18866
rect -19234 18506 -18834 18546
rect -18112 18866 -17712 18906
rect -18112 18546 -18072 18866
rect -17752 18546 -17712 18866
rect -18112 18506 -17712 18546
rect -16990 18866 -16590 18906
rect -16990 18546 -16950 18866
rect -16630 18546 -16590 18866
rect -16990 18506 -16590 18546
rect -15868 18866 -15468 18906
rect -15868 18546 -15828 18866
rect -15508 18546 -15468 18866
rect -15868 18506 -15468 18546
rect -14746 18866 -14346 18906
rect -14746 18546 -14706 18866
rect -14386 18546 -14346 18866
rect -14746 18506 -14346 18546
rect -13624 18866 -13224 18906
rect -13624 18546 -13584 18866
rect -13264 18546 -13224 18866
rect -13624 18506 -13224 18546
rect -12502 18866 -12102 18906
rect -12502 18546 -12462 18866
rect -12142 18546 -12102 18866
rect -12502 18506 -12102 18546
rect -11380 18866 -10980 18906
rect -11380 18546 -11340 18866
rect -11020 18546 -10980 18866
rect -11380 18506 -10980 18546
rect -21478 18166 -21078 18206
rect -21478 17846 -21438 18166
rect -21118 17846 -21078 18166
rect -21478 17806 -21078 17846
rect -20356 18166 -19956 18206
rect -20356 17846 -20316 18166
rect -19996 17846 -19956 18166
rect -20356 17806 -19956 17846
rect -19234 18166 -18834 18206
rect -19234 17846 -19194 18166
rect -18874 17846 -18834 18166
rect -19234 17806 -18834 17846
rect -18112 18166 -17712 18206
rect -18112 17846 -18072 18166
rect -17752 17846 -17712 18166
rect -18112 17806 -17712 17846
rect -16990 18166 -16590 18206
rect -16990 17846 -16950 18166
rect -16630 17846 -16590 18166
rect -16990 17806 -16590 17846
rect -15868 18166 -15468 18206
rect -15868 17846 -15828 18166
rect -15508 17846 -15468 18166
rect -15868 17806 -15468 17846
rect -14746 18166 -14346 18206
rect -14746 17846 -14706 18166
rect -14386 17846 -14346 18166
rect -14746 17806 -14346 17846
rect -13624 18166 -13224 18206
rect -13624 17846 -13584 18166
rect -13264 17846 -13224 18166
rect -13624 17806 -13224 17846
rect -12502 18166 -12102 18206
rect -12502 17846 -12462 18166
rect -12142 17846 -12102 18166
rect -12502 17806 -12102 17846
rect -11380 18166 -10980 18206
rect -11380 17846 -11340 18166
rect -11020 17846 -10980 18166
rect -11380 17806 -10980 17846
rect -21478 17466 -21078 17506
rect -21478 17146 -21438 17466
rect -21118 17146 -21078 17466
rect -21478 17106 -21078 17146
rect -20356 17466 -19956 17506
rect -20356 17146 -20316 17466
rect -19996 17146 -19956 17466
rect -20356 17106 -19956 17146
rect -19234 17466 -18834 17506
rect -19234 17146 -19194 17466
rect -18874 17146 -18834 17466
rect -19234 17106 -18834 17146
rect -18112 17466 -17712 17506
rect -18112 17146 -18072 17466
rect -17752 17146 -17712 17466
rect -18112 17106 -17712 17146
rect -16990 17466 -16590 17506
rect -16990 17146 -16950 17466
rect -16630 17146 -16590 17466
rect -16990 17106 -16590 17146
rect -15868 17466 -15468 17506
rect -15868 17146 -15828 17466
rect -15508 17146 -15468 17466
rect -15868 17106 -15468 17146
rect -14746 17466 -14346 17506
rect -14746 17146 -14706 17466
rect -14386 17146 -14346 17466
rect -14746 17106 -14346 17146
rect -13624 17466 -13224 17506
rect -13624 17146 -13584 17466
rect -13264 17146 -13224 17466
rect -13624 17106 -13224 17146
rect -12502 17466 -12102 17506
rect -12502 17146 -12462 17466
rect -12142 17146 -12102 17466
rect -12502 17106 -12102 17146
rect -11380 17466 -10980 17506
rect -11380 17146 -11340 17466
rect -11020 17146 -10980 17466
rect -11380 17106 -10980 17146
<< mimcap2contact >>
rect -21438 23446 -21118 23766
rect -20316 23446 -19996 23766
rect -19194 23446 -18874 23766
rect -18072 23446 -17752 23766
rect -16950 23446 -16630 23766
rect -15828 23446 -15508 23766
rect -14706 23446 -14386 23766
rect -13584 23446 -13264 23766
rect -12462 23446 -12142 23766
rect -11340 23446 -11020 23766
rect -21438 22746 -21118 23066
rect -20316 22746 -19996 23066
rect -19194 22746 -18874 23066
rect -18072 22746 -17752 23066
rect -16950 22746 -16630 23066
rect -15828 22746 -15508 23066
rect -14706 22746 -14386 23066
rect -13584 22746 -13264 23066
rect -12462 22746 -12142 23066
rect -11340 22746 -11020 23066
rect -21438 22046 -21118 22366
rect -20316 22046 -19996 22366
rect -19194 22046 -18874 22366
rect -18072 22046 -17752 22366
rect -16950 22046 -16630 22366
rect -15828 22046 -15508 22366
rect -14706 22046 -14386 22366
rect -13584 22046 -13264 22366
rect -12462 22046 -12142 22366
rect -11340 22046 -11020 22366
rect -21438 21346 -21118 21666
rect -20316 21346 -19996 21666
rect -19194 21346 -18874 21666
rect -18072 21346 -17752 21666
rect -16950 21346 -16630 21666
rect -15828 21346 -15508 21666
rect -14706 21346 -14386 21666
rect -13584 21346 -13264 21666
rect -12462 21346 -12142 21666
rect -11340 21346 -11020 21666
rect -21438 20646 -21118 20966
rect -20316 20646 -19996 20966
rect -19194 20646 -18874 20966
rect -18072 20646 -17752 20966
rect -16950 20646 -16630 20966
rect -15828 20646 -15508 20966
rect -14706 20646 -14386 20966
rect -13584 20646 -13264 20966
rect -12462 20646 -12142 20966
rect -11340 20646 -11020 20966
rect -21438 19946 -21118 20266
rect -20316 19946 -19996 20266
rect -19194 19946 -18874 20266
rect -18072 19946 -17752 20266
rect -16950 19946 -16630 20266
rect -15828 19946 -15508 20266
rect -14706 19946 -14386 20266
rect -13584 19946 -13264 20266
rect -12462 19946 -12142 20266
rect -11340 19946 -11020 20266
rect -21438 19246 -21118 19566
rect -20316 19246 -19996 19566
rect -19194 19246 -18874 19566
rect -18072 19246 -17752 19566
rect -16950 19246 -16630 19566
rect -15828 19246 -15508 19566
rect -14706 19246 -14386 19566
rect -13584 19246 -13264 19566
rect -12462 19246 -12142 19566
rect -11340 19246 -11020 19566
rect -21438 18546 -21118 18866
rect -20316 18546 -19996 18866
rect -19194 18546 -18874 18866
rect -18072 18546 -17752 18866
rect -16950 18546 -16630 18866
rect -15828 18546 -15508 18866
rect -14706 18546 -14386 18866
rect -13584 18546 -13264 18866
rect -12462 18546 -12142 18866
rect -11340 18546 -11020 18866
rect -21438 17846 -21118 18166
rect -20316 17846 -19996 18166
rect -19194 17846 -18874 18166
rect -18072 17846 -17752 18166
rect -16950 17846 -16630 18166
rect -15828 17846 -15508 18166
rect -14706 17846 -14386 18166
rect -13584 17846 -13264 18166
rect -12462 17846 -12142 18166
rect -11340 17846 -11020 18166
rect -21438 17146 -21118 17466
rect -20316 17146 -19996 17466
rect -19194 17146 -18874 17466
rect -18072 17146 -17752 17466
rect -16950 17146 -16630 17466
rect -15828 17146 -15508 17466
rect -14706 17146 -14386 17466
rect -13584 17146 -13264 17466
rect -12462 17146 -12142 17466
rect -11340 17146 -11020 17466
<< metal5 >>
rect -21532 23950 11082 24225
rect -21532 23766 11238 23950
rect -21532 23446 -21438 23766
rect -21118 23446 -20316 23766
rect -19996 23446 -19194 23766
rect -18874 23446 -18072 23766
rect -17752 23446 -16950 23766
rect -16630 23446 -15828 23766
rect -15508 23446 -14706 23766
rect -14386 23446 -13584 23766
rect -13264 23446 -12462 23766
rect -12142 23446 -11340 23766
rect -11020 23446 11238 23766
rect -21532 23066 11238 23446
rect -21532 22746 -21438 23066
rect -21118 22746 -20316 23066
rect -19996 22746 -19194 23066
rect -18874 22746 -18072 23066
rect -17752 22746 -16950 23066
rect -16630 22746 -15828 23066
rect -15508 22746 -14706 23066
rect -14386 22746 -13584 23066
rect -13264 22746 -12462 23066
rect -12142 22746 -11340 23066
rect -11020 22746 11238 23066
rect -21532 22366 11238 22746
rect -21532 22046 -21438 22366
rect -21118 22046 -20316 22366
rect -19996 22046 -19194 22366
rect -18874 22046 -18072 22366
rect -17752 22046 -16950 22366
rect -16630 22046 -15828 22366
rect -15508 22046 -14706 22366
rect -14386 22046 -13584 22366
rect -13264 22046 -12462 22366
rect -12142 22046 -11340 22366
rect -11020 22046 11238 22366
rect -21532 21666 11238 22046
rect -21532 21346 -21438 21666
rect -21118 21346 -20316 21666
rect -19996 21346 -19194 21666
rect -18874 21346 -18072 21666
rect -17752 21346 -16950 21666
rect -16630 21346 -15828 21666
rect -15508 21346 -14706 21666
rect -14386 21346 -13584 21666
rect -13264 21346 -12462 21666
rect -12142 21346 -11340 21666
rect -11020 21346 11238 21666
rect -21532 20966 11238 21346
rect -21532 20646 -21438 20966
rect -21118 20646 -20316 20966
rect -19996 20646 -19194 20966
rect -18874 20646 -18072 20966
rect -17752 20646 -16950 20966
rect -16630 20646 -15828 20966
rect -15508 20646 -14706 20966
rect -14386 20646 -13584 20966
rect -13264 20646 -12462 20966
rect -12142 20646 -11340 20966
rect -11020 20646 11238 20966
rect -21532 20266 11238 20646
rect -21532 19946 -21438 20266
rect -21118 19946 -20316 20266
rect -19996 19946 -19194 20266
rect -18874 19946 -18072 20266
rect -17752 19946 -16950 20266
rect -16630 19946 -15828 20266
rect -15508 19946 -14706 20266
rect -14386 19946 -13584 20266
rect -13264 19946 -12462 20266
rect -12142 19946 -11340 20266
rect -11020 19946 11238 20266
rect -21532 19566 11238 19946
rect -21532 19246 -21438 19566
rect -21118 19246 -20316 19566
rect -19996 19246 -19194 19566
rect -18874 19246 -18072 19566
rect -17752 19246 -16950 19566
rect -16630 19246 -15828 19566
rect -15508 19246 -14706 19566
rect -14386 19246 -13584 19566
rect -13264 19246 -12462 19566
rect -12142 19246 -11340 19566
rect -11020 19246 11238 19566
rect -21532 18866 11238 19246
rect -21532 18546 -21438 18866
rect -21118 18546 -20316 18866
rect -19996 18546 -19194 18866
rect -18874 18546 -18072 18866
rect -17752 18546 -16950 18866
rect -16630 18546 -15828 18866
rect -15508 18546 -14706 18866
rect -14386 18546 -13584 18866
rect -13264 18546 -12462 18866
rect -12142 18546 -11340 18866
rect -11020 18546 11238 18866
rect -21532 18166 11238 18546
rect -21532 17846 -21438 18166
rect -21118 17846 -20316 18166
rect -19996 17846 -19194 18166
rect -18874 17846 -18072 18166
rect -17752 17846 -16950 18166
rect -16630 17846 -15828 18166
rect -15508 17846 -14706 18166
rect -14386 17846 -13584 18166
rect -13264 17846 -12462 18166
rect -12142 17846 -11340 18166
rect -11020 17846 11238 18166
rect -21532 17466 11238 17846
rect -21532 17146 -21438 17466
rect -21118 17146 -20316 17466
rect -19996 17146 -19194 17466
rect -18874 17146 -18072 17466
rect -17752 17146 -16950 17466
rect -16630 17146 -15828 17466
rect -15508 17146 -14706 17466
rect -14386 17146 -13584 17466
rect -13264 17146 -12462 17466
rect -12142 17146 -11340 17466
rect -11020 17146 11238 17466
rect -21532 11780 11238 17146
rect -21532 10808 -9246 11780
rect 11064 10808 11238 11780
rect -21532 10748 11238 10808
rect -9246 10710 11238 10748
<< res2p85 >>
rect -8934 16850 -8360 20178
rect -8116 16850 -7542 20178
rect -7298 16850 -6724 20178
rect -5662 17260 -5088 21564
rect -4844 17260 -4270 21564
rect -4026 17260 -3452 21564
rect -3208 17260 -2634 21564
rect -754 15194 -180 21502
rect 64 15194 638 21502
rect 882 15194 1456 21502
rect 1700 15194 2274 21502
rect 2518 15194 3092 21502
rect 3336 15194 3910 21502
rect 4154 15194 4728 21502
rect 4972 15194 5546 21502
rect 5790 15194 6364 21502
rect 6608 15194 7182 21502
rect 7426 15194 8000 21502
rect 8244 15194 8818 21502
rect 9062 15194 9636 21502
rect 9880 15194 10454 21502
rect 10698 15194 11272 21502
rect 11516 15194 12090 21502
rect 12334 15194 12908 21502
<< labels >>
flabel metal1 -19254 8502 -18792 8700 1 FreeSans 1600 0 0 0 porst
port 0 n
flabel metal1 -2858 12824 1810 13500 1 FreeSans 1600 0 0 0 Vbg
port 1 n
flabel metal3 -20266 1000 -19556 1422 1 FreeSans 1600 0 0 0 VDD!
flabel metal2 -21312 4728 -19530 4798 1 FreeSans 800 0 0 0 ampcurrentsource_0/Vq
flabel metal2 -21312 4938 -19530 5008 1 FreeSans 800 0 0 0 ampcurrentsource_0/Vx
flabel locali -20452 5698 -20370 5726 1 FreeSans 800 0 0 0 ampcurrentsource_0/GND!
rlabel via1 -8118 1418 -8072 1462 5 currentmirror_0/Vgate
rlabel metal3 -7396 1062 -7262 1180 5 currentmirror_0/VDD!
flabel metal1 -590 9602 -290 9702 5 FreeSans 1600 0 0 0 currentmirror_0/Vbg
flabel metal2 -590 10202 -390 10302 5 FreeSans 1600 0 0 0 currentmirror_0/Vb
flabel metal2 -590 10802 -390 10902 5 FreeSans 1600 0 0 0 currentmirror_0/Va
flabel metal2 11606 2220 12742 3168 7 FreeSans 1600 0 0 0 bandgapcorev3_0/Vbneg
flabel locali -4664 16814 -3560 17104 1 FreeSans 800 90 0 0 bandgapcorev3_0/GND!
flabel metal2 884 21500 1454 21932 1 FreeSans 800 90 0 0 bandgapcorev3_0/VbEnd
flabel metal2 1702 14764 2272 15196 1 FreeSans 800 90 0 0 bandgapcorev3_0/VbgEnd
flabel metal2 66 20700 636 21932 1 FreeSans 800 90 0 0 bandgapcorev3_0/VaEnd
flabel metal2 9810 14498 10502 15190 1 FreeSans 1600 90 0 0 bandgapcorev3_0/Vbg
flabel metal2 11440 14492 12144 15196 1 FreeSans 1600 90 0 0 bandgapcorev3_0/Vb
flabel metal1 10622 13926 11326 14498 3 FreeSans 1600 0 0 0 bandgapcorev3_0/Va
flabel locali 18108 11530 18356 11634 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,0]/Emitter
flabel locali 18196 10959 18297 11008 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,0]/Collector
flabel locali 18202 11118 18320 11158 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,0]/Base
flabel locali 16820 11530 17068 11634 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,1]/Emitter
flabel locali 16908 10959 17009 11008 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,1]/Collector
flabel locali 16914 11118 17032 11158 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,1]/Base
flabel locali 15532 11530 15780 11634 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,2]/Emitter
flabel locali 15620 10959 15721 11008 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,2]/Collector
flabel locali 15626 11118 15744 11158 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,2]/Base
flabel locali 14244 11530 14492 11634 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,3]/Emitter
flabel locali 14332 10959 14433 11008 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,3]/Collector
flabel locali 14338 11118 14456 11158 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,3]/Base
flabel locali 12956 11530 13204 11634 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,4]/Emitter
flabel locali 13044 10959 13145 11008 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,4]/Collector
flabel locali 13050 11118 13168 11158 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,4]/Base
flabel locali 18108 10242 18356 10346 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,0]/Emitter
flabel locali 18196 9671 18297 9720 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,0]/Collector
flabel locali 18202 9830 18320 9870 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,0]/Base
flabel locali 16820 10242 17068 10346 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,1]/Emitter
flabel locali 16908 9671 17009 9720 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,1]/Collector
flabel locali 16914 9830 17032 9870 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,1]/Base
flabel locali 15532 10242 15780 10346 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,2]/Emitter
flabel locali 15620 9671 15721 9720 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,2]/Collector
flabel locali 15626 9830 15744 9870 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,2]/Base
flabel locali 14244 10242 14492 10346 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,3]/Emitter
flabel locali 14332 9671 14433 9720 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,3]/Collector
flabel locali 14338 9830 14456 9870 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,3]/Base
flabel locali 12956 10242 13204 10346 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,4]/Emitter
flabel locali 13044 9671 13145 9720 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,4]/Collector
flabel locali 13050 9830 13168 9870 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,4]/Base
flabel locali 18108 8954 18356 9058 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,0]/Emitter
flabel locali 18196 8383 18297 8432 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,0]/Collector
flabel locali 18202 8542 18320 8582 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,0]/Base
flabel locali 16820 8954 17068 9058 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,1]/Emitter
flabel locali 16908 8383 17009 8432 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,1]/Collector
flabel locali 16914 8542 17032 8582 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,1]/Base
flabel locali 15532 8954 15780 9058 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,2]/Emitter
flabel locali 15620 8383 15721 8432 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,2]/Collector
flabel locali 15626 8542 15744 8582 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,2]/Base
flabel locali 14244 8954 14492 9058 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,3]/Emitter
flabel locali 14332 8383 14433 8432 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,3]/Collector
flabel locali 14338 8542 14456 8582 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,3]/Base
flabel locali 12956 8954 13204 9058 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,4]/Emitter
flabel locali 13044 8383 13145 8432 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,4]/Collector
flabel locali 13050 8542 13168 8582 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,4]/Base
flabel locali 18108 7666 18356 7770 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,0]/Emitter
flabel locali 18196 7095 18297 7144 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,0]/Collector
flabel locali 18202 7254 18320 7294 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,0]/Base
flabel locali 16820 7666 17068 7770 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,1]/Emitter
flabel locali 16908 7095 17009 7144 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,1]/Collector
flabel locali 16914 7254 17032 7294 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,1]/Base
flabel locali 15532 7666 15780 7770 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,2]/Emitter
flabel locali 15620 7095 15721 7144 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,2]/Collector
flabel locali 15626 7254 15744 7294 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,2]/Base
flabel locali 14244 7666 14492 7770 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,3]/Emitter
flabel locali 14332 7095 14433 7144 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,3]/Collector
flabel locali 14338 7254 14456 7294 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,3]/Base
flabel locali 12956 7666 13204 7770 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,4]/Emitter
flabel locali 13044 7095 13145 7144 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,4]/Collector
flabel locali 13050 7254 13168 7294 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,4]/Base
flabel locali 18108 6378 18356 6482 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,0]/Emitter
flabel locali 18196 5807 18297 5856 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,0]/Collector
flabel locali 18202 5966 18320 6006 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,0]/Base
flabel locali 16820 6378 17068 6482 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,1]/Emitter
flabel locali 16908 5807 17009 5856 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,1]/Collector
flabel locali 16914 5966 17032 6006 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,1]/Base
flabel locali 15532 6378 15780 6482 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,2]/Emitter
flabel locali 15620 5807 15721 5856 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,2]/Collector
flabel locali 15626 5966 15744 6006 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,2]/Base
flabel locali 14244 6378 14492 6482 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,3]/Emitter
flabel locali 14332 5807 14433 5856 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,3]/Collector
flabel locali 14338 5966 14456 6006 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,3]/Base
flabel locali 12956 6378 13204 6482 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,4]/Emitter
flabel locali 13044 5807 13145 5856 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,4]/Collector
flabel locali 13050 5966 13168 6006 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,4]/Base
flabel locali 18108 5090 18356 5194 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,0]/Emitter
flabel locali 18196 4519 18297 4568 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,0]/Collector
flabel locali 18202 4678 18320 4718 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,0]/Base
flabel locali 16820 5090 17068 5194 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,1]/Emitter
flabel locali 16908 4519 17009 4568 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,1]/Collector
flabel locali 16914 4678 17032 4718 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,1]/Base
flabel locali 15532 5090 15780 5194 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,2]/Emitter
flabel locali 15620 4519 15721 4568 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,2]/Collector
flabel locali 15626 4678 15744 4718 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,2]/Base
flabel locali 14244 5090 14492 5194 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,3]/Emitter
flabel locali 14332 4519 14433 4568 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,3]/Collector
flabel locali 14338 4678 14456 4718 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,3]/Base
flabel locali 12956 5090 13204 5194 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,4]/Emitter
flabel locali 13044 4519 13145 4568 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,4]/Collector
flabel locali 13050 4678 13168 4718 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,4]/Base
flabel locali 18108 3802 18356 3906 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,0]/Emitter
flabel locali 18196 3231 18297 3280 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,0]/Collector
flabel locali 18202 3390 18320 3430 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,0]/Base
flabel locali 16820 3802 17068 3906 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,1]/Emitter
flabel locali 16908 3231 17009 3280 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,1]/Collector
flabel locali 16914 3390 17032 3430 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,1]/Base
flabel locali 15532 3802 15780 3906 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,2]/Emitter
flabel locali 15620 3231 15721 3280 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,2]/Collector
flabel locali 15626 3390 15744 3430 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,2]/Base
flabel locali 14244 3802 14492 3906 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,3]/Emitter
flabel locali 14332 3231 14433 3280 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,3]/Collector
flabel locali 14338 3390 14456 3430 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,3]/Base
flabel locali 12956 3802 13204 3906 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,4]/Emitter
flabel locali 13044 3231 13145 3280 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,4]/Collector
flabel locali 13050 3390 13168 3430 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,4]/Base
flabel locali 18108 2514 18356 2618 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,0]/Emitter
flabel locali 18196 1943 18297 1992 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,0]/Collector
flabel locali 18202 2102 18320 2142 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,0]/Base
flabel locali 16820 2514 17068 2618 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,1]/Emitter
flabel locali 16908 1943 17009 1992 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,1]/Collector
flabel locali 16914 2102 17032 2142 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,1]/Base
flabel locali 15532 2514 15780 2618 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,2]/Emitter
flabel locali 15620 1943 15721 1992 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,2]/Collector
flabel locali 15626 2102 15744 2142 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,2]/Base
flabel locali 14244 2514 14492 2618 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,3]/Emitter
flabel locali 14332 1943 14433 1992 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,3]/Collector
flabel locali 14338 2102 14456 2142 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,3]/Base
flabel locali 12956 2514 13204 2618 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,4]/Emitter
flabel locali 13044 1943 13145 1992 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,4]/Collector
flabel locali 13050 2102 13168 2142 0 FreeSans 400 0 0 0 bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,4]/Base
flabel metal2 -14560 1438 -14544 1562 5 FreeSans 800 0 0 0 amplifier_0/VDD!
flabel metal2 -13906 4666 -13890 4790 5 FreeSans 800 0 0 0 amplifier_0/Vq
flabel metal2 -13964 6926 -13948 7006 5 FreeSans 800 0 0 0 amplifier_0/Va
flabel metal2 -14736 6786 -14720 6866 5 FreeSans 800 0 0 0 amplifier_0/Vb
flabel metal2 -13230 4370 -13136 4636 5 FreeSans 800 0 0 0 amplifier_0/Vgate
flabel metal2 -14954 4370 -14860 4636 5 FreeSans 800 0 0 0 amplifier_0/Vgate
flabel metal1 -16312 4384 -16278 4476 5 FreeSans 800 0 0 0 amplifier_0/vg
flabel metal2 -12212 1238 -12190 1362 5 FreeSans 800 0 0 0 amplifier_0/Vx
flabel psubdiffcont -17434 5042 -17334 6642 5 FreeSans 800 0 0 0 amplifier_0/GND!
flabel psubdiff -11984 6642 -11784 6742 5 FreeSans 800 180 0 0 amplifier_0/GND!
<< end >>
