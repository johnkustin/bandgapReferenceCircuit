magic
tech sky130A
magscale 1 2
timestamp 1620776712
<< locali >>
rect 8400 -5000 8600 5300
rect 9500 -5000 9900 5200
rect 10800 -5000 11200 5200
rect 12100 -5000 12500 5200
rect 13300 -5000 13800 5300
rect 14600 5100 14800 5300
rect 14600 4300 14700 5100
rect 14600 -5000 14800 4300
<< viali >>
rect 14700 4300 14800 5100
<< metal1 >>
rect 8102 11700 8572 11826
rect 8102 11500 8200 11700
rect 8500 11500 8572 11700
rect 8102 11394 8572 11500
rect 9800 8100 11400 8200
rect 8102 5900 8172 6600
rect 8502 6492 8572 6600
rect 8444 6486 8630 6492
rect 8444 6300 8450 6486
rect 8624 6400 8630 6486
rect 9800 6400 9900 8100
rect 11302 6500 11372 6600
rect 14102 6568 14172 6600
rect 14088 6548 14188 6568
rect 8624 6300 9900 6400
rect 8444 6294 8630 6300
rect 8102 5686 9400 5900
rect 8102 5500 8450 5686
rect 8624 5500 9400 5686
rect 8102 4300 9400 5500
rect 11000 5000 11700 6500
rect 14088 6488 14108 6548
rect 14168 6488 14188 6548
rect 14088 6468 14188 6488
rect 14800 5200 15400 5300
rect 14600 5100 15400 5200
rect 10000 3900 14500 5000
rect 14600 4300 14700 5100
rect 14800 4300 15000 5100
rect 14600 4100 15000 4300
rect 15300 4100 15400 5100
rect 14800 3900 15400 4100
rect 10000 3700 14600 3900
rect 8700 -4700 14600 3700
<< via1 >>
rect 8200 11500 8500 11700
rect 8450 6300 8624 6486
rect 8450 5500 8624 5686
rect 14108 6488 14168 6548
rect 15000 4100 15300 5100
<< metal2 >>
rect 8100 11700 15500 11800
rect 8100 11500 8200 11700
rect 8500 11500 15500 11700
rect 8100 11400 15500 11500
rect 14900 8348 15500 11400
rect 14758 8248 15500 8348
rect 14900 7884 15500 8248
rect 14758 7784 15500 7884
rect 14900 6568 15500 7784
rect 14088 6548 15500 6568
rect 8444 6486 8630 6492
rect 8444 6300 8450 6486
rect 8624 6300 8630 6486
rect 14088 6488 14108 6548
rect 14168 6488 15500 6548
rect 14088 6468 15500 6488
rect 8444 6294 8630 6300
rect 8444 5686 8630 5692
rect 8444 5500 8450 5686
rect 8624 5500 8630 5686
rect 8444 5494 8630 5500
rect 14900 5100 15500 6468
rect 14900 4100 15000 5100
rect 15300 4100 15500 5100
rect 14900 3900 15500 4100
use sky130_fd_pr__res_xhigh_po_0p35_3LWQVB  sky130_fd_pr__res_xhigh_po_0p35_3LWQVB_0
timestamp 1620775510
transform 1 0 11335 0 1 7402
box -37 -808 37 808
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 7 1288
timestamp 1620596431
transform 1 0 8374 0 1 -5042
box 26 26 1314 1314
use sky130_fd_pr__res_xhigh_po_0p35_ZG99VC  sky130_fd_pr__res_xhigh_po_0p35_ZG99VC_1
timestamp 1620775510
transform 1 0 8137 0 1 9210
box -37 -2616 37 2616
use sky130_fd_pr__res_xhigh_po_0p35_ZG99VC  sky130_fd_pr__res_xhigh_po_0p35_ZG99VC_0
timestamp 1620775510
transform 1 0 8537 0 1 9210
box -37 -2616 37 2616
<< labels >>
flabel metal2 14900 6100 15400 6400 1 FreeSans 1600 0 0 0 GND!
port 2 n
flabel metal1 11240 5360 11440 5580 1 FreeSans 800 0 0 0 Vbneg
flabel metal1 8700 5500 9000 5800 1 FreeSans 1600 0 0 0 Va
port 1 n
flabel via1 8458 6304 8606 6468 1 FreeSans 1600 0 0 0 Vb
port 0 n
<< end >>
