magic
tech sky130A
magscale 1 2
timestamp 1621270741
<< error_p >>
rect -4538 3331 -4498 3450
rect -4478 3331 -4438 3450
rect -4338 3334 -4156 3500
rect -4796 3289 -4438 3331
rect -4796 3011 -4754 3289
rect -4682 3011 -4438 3289
rect -4796 2969 -4438 3011
rect -4538 2850 -4498 2969
rect -4478 2850 -4438 2969
rect -4362 2966 -4156 3334
rect -3416 3331 -3376 3450
rect -3356 3331 -3316 3450
rect -3216 3334 -3034 3500
rect -3674 3289 -3316 3331
rect -3674 3011 -3632 3289
rect -3560 3011 -3316 3289
rect -3674 2969 -3316 3011
rect -4538 2631 -4498 2750
rect -4478 2631 -4438 2750
rect -4338 2634 -4156 2966
rect -3416 2850 -3376 2969
rect -3356 2850 -3316 2969
rect -3240 2966 -3034 3334
rect -2294 3331 -2254 3450
rect -2234 3331 -2194 3450
rect -2094 3334 -1912 3500
rect -2552 3289 -2194 3331
rect -2552 3011 -2510 3289
rect -2438 3011 -2194 3289
rect -2552 2969 -2194 3011
rect -4796 2589 -4438 2631
rect -4796 2311 -4754 2589
rect -4682 2311 -4438 2589
rect -4796 2269 -4438 2311
rect -4538 2150 -4498 2269
rect -4478 2150 -4438 2269
rect -4362 2266 -4156 2634
rect -3416 2631 -3376 2750
rect -3356 2631 -3316 2750
rect -3216 2634 -3034 2966
rect -2294 2850 -2254 2969
rect -2234 2850 -2194 2969
rect -2118 2966 -1912 3334
rect -1172 3331 -1132 3450
rect -1112 3331 -1072 3450
rect -972 3334 -790 3500
rect -1430 3289 -1072 3331
rect -1430 3011 -1388 3289
rect -1316 3011 -1072 3289
rect -1430 2969 -1072 3011
rect -3674 2589 -3316 2631
rect -3674 2311 -3632 2589
rect -3560 2311 -3316 2589
rect -3674 2269 -3316 2311
rect -4538 1931 -4498 2050
rect -4478 1931 -4438 2050
rect -4338 1934 -4156 2266
rect -3416 2150 -3376 2269
rect -3356 2150 -3316 2269
rect -3240 2266 -3034 2634
rect -2294 2631 -2254 2750
rect -2234 2631 -2194 2750
rect -2094 2634 -1912 2966
rect -1172 2850 -1132 2969
rect -1112 2850 -1072 2969
rect -996 2966 -790 3334
rect -50 3331 -10 3450
rect 10 3331 50 3450
rect 150 3334 332 3500
rect -308 3289 50 3331
rect -308 3011 -266 3289
rect -194 3011 50 3289
rect -308 2969 50 3011
rect -2552 2589 -2194 2631
rect -2552 2311 -2510 2589
rect -2438 2311 -2194 2589
rect -2552 2269 -2194 2311
rect -4796 1889 -4438 1931
rect -4796 1611 -4754 1889
rect -4682 1611 -4438 1889
rect -4796 1569 -4438 1611
rect -4538 1450 -4498 1569
rect -4478 1450 -4438 1569
rect -4362 1566 -4156 1934
rect -3416 1931 -3376 2050
rect -3356 1931 -3316 2050
rect -3216 1934 -3034 2266
rect -2294 2150 -2254 2269
rect -2234 2150 -2194 2269
rect -2118 2266 -1912 2634
rect -1172 2631 -1132 2750
rect -1112 2631 -1072 2750
rect -972 2634 -790 2966
rect -50 2850 -10 2969
rect 10 2850 50 2969
rect 126 2966 332 3334
rect 1072 3331 1112 3450
rect 1132 3331 1172 3450
rect 1272 3334 1454 3500
rect 814 3289 1172 3331
rect 814 3011 856 3289
rect 928 3011 1172 3289
rect 814 2969 1172 3011
rect -1430 2589 -1072 2631
rect -1430 2311 -1388 2589
rect -1316 2311 -1072 2589
rect -1430 2269 -1072 2311
rect -3674 1889 -3316 1931
rect -3674 1611 -3632 1889
rect -3560 1611 -3316 1889
rect -3674 1569 -3316 1611
rect -4538 1231 -4498 1350
rect -4478 1231 -4438 1350
rect -4338 1234 -4156 1566
rect -3416 1450 -3376 1569
rect -3356 1450 -3316 1569
rect -3240 1566 -3034 1934
rect -2294 1931 -2254 2050
rect -2234 1931 -2194 2050
rect -2094 1934 -1912 2266
rect -1172 2150 -1132 2269
rect -1112 2150 -1072 2269
rect -996 2266 -790 2634
rect -50 2631 -10 2750
rect 10 2631 50 2750
rect 150 2634 332 2966
rect 1072 2850 1112 2969
rect 1132 2850 1172 2969
rect 1248 2966 1454 3334
rect 2194 3331 2234 3450
rect 2254 3331 2294 3450
rect 2394 3334 2576 3500
rect 1936 3289 2294 3331
rect 1936 3011 1978 3289
rect 2050 3011 2294 3289
rect 1936 2969 2294 3011
rect -308 2589 50 2631
rect -308 2311 -266 2589
rect -194 2311 50 2589
rect -308 2269 50 2311
rect -2552 1889 -2194 1931
rect -2552 1611 -2510 1889
rect -2438 1611 -2194 1889
rect -2552 1569 -2194 1611
rect -4796 1189 -4438 1231
rect -4796 911 -4754 1189
rect -4682 911 -4438 1189
rect -4796 869 -4438 911
rect -4538 750 -4498 869
rect -4478 750 -4438 869
rect -4362 866 -4156 1234
rect -3416 1231 -3376 1350
rect -3356 1231 -3316 1350
rect -3216 1234 -3034 1566
rect -2294 1450 -2254 1569
rect -2234 1450 -2194 1569
rect -2118 1566 -1912 1934
rect -1172 1931 -1132 2050
rect -1112 1931 -1072 2050
rect -972 1934 -790 2266
rect -50 2150 -10 2269
rect 10 2150 50 2269
rect 126 2266 332 2634
rect 1072 2631 1112 2750
rect 1132 2631 1172 2750
rect 1272 2634 1454 2966
rect 2194 2850 2234 2969
rect 2254 2850 2294 2969
rect 2370 2966 2576 3334
rect 3316 3331 3356 3450
rect 3376 3331 3416 3450
rect 3516 3334 3698 3500
rect 3058 3289 3416 3331
rect 3058 3011 3100 3289
rect 3172 3011 3416 3289
rect 3058 2969 3416 3011
rect 814 2589 1172 2631
rect 814 2311 856 2589
rect 928 2311 1172 2589
rect 814 2269 1172 2311
rect -1430 1889 -1072 1931
rect -1430 1611 -1388 1889
rect -1316 1611 -1072 1889
rect -1430 1569 -1072 1611
rect -3674 1189 -3316 1231
rect -3674 911 -3632 1189
rect -3560 911 -3316 1189
rect -3674 869 -3316 911
rect -4538 531 -4498 650
rect -4478 531 -4438 650
rect -4338 534 -4156 866
rect -3416 750 -3376 869
rect -3356 750 -3316 869
rect -3240 866 -3034 1234
rect -2294 1231 -2254 1350
rect -2234 1231 -2194 1350
rect -2094 1234 -1912 1566
rect -1172 1450 -1132 1569
rect -1112 1450 -1072 1569
rect -996 1566 -790 1934
rect -50 1931 -10 2050
rect 10 1931 50 2050
rect 150 1934 332 2266
rect 1072 2150 1112 2269
rect 1132 2150 1172 2269
rect 1248 2266 1454 2634
rect 2194 2631 2234 2750
rect 2254 2631 2294 2750
rect 2394 2634 2576 2966
rect 3316 2850 3356 2969
rect 3376 2850 3416 2969
rect 3492 2966 3698 3334
rect 4438 3331 4478 3450
rect 4498 3331 4538 3450
rect 4638 3334 4820 3500
rect 4180 3289 4538 3331
rect 4180 3011 4222 3289
rect 4294 3011 4538 3289
rect 4180 2969 4538 3011
rect 1936 2589 2294 2631
rect 1936 2311 1978 2589
rect 2050 2311 2294 2589
rect 1936 2269 2294 2311
rect -308 1889 50 1931
rect -308 1611 -266 1889
rect -194 1611 50 1889
rect -308 1569 50 1611
rect -2552 1189 -2194 1231
rect -2552 911 -2510 1189
rect -2438 911 -2194 1189
rect -2552 869 -2194 911
rect -4796 489 -4438 531
rect -4796 211 -4754 489
rect -4682 211 -4438 489
rect -4796 169 -4438 211
rect -4538 50 -4498 169
rect -4478 50 -4438 169
rect -4362 166 -4156 534
rect -3416 531 -3376 650
rect -3356 531 -3316 650
rect -3216 534 -3034 866
rect -2294 750 -2254 869
rect -2234 750 -2194 869
rect -2118 866 -1912 1234
rect -1172 1231 -1132 1350
rect -1112 1231 -1072 1350
rect -972 1234 -790 1566
rect -50 1450 -10 1569
rect 10 1450 50 1569
rect 126 1566 332 1934
rect 1072 1931 1112 2050
rect 1132 1931 1172 2050
rect 1272 1934 1454 2266
rect 2194 2150 2234 2269
rect 2254 2150 2294 2269
rect 2370 2266 2576 2634
rect 3316 2631 3356 2750
rect 3376 2631 3416 2750
rect 3516 2634 3698 2966
rect 4438 2850 4478 2969
rect 4498 2850 4538 2969
rect 4614 2966 4820 3334
rect 5302 3289 5622 3331
rect 5302 3011 5344 3289
rect 5302 2969 5622 3011
rect 3058 2589 3416 2631
rect 3058 2311 3100 2589
rect 3172 2311 3416 2589
rect 3058 2269 3416 2311
rect 814 1889 1172 1931
rect 814 1611 856 1889
rect 928 1611 1172 1889
rect 814 1569 1172 1611
rect -1430 1189 -1072 1231
rect -1430 911 -1388 1189
rect -1316 911 -1072 1189
rect -1430 869 -1072 911
rect -3674 489 -3316 531
rect -3674 211 -3632 489
rect -3560 211 -3316 489
rect -3674 169 -3316 211
rect -4538 -169 -4498 -50
rect -4478 -169 -4438 -50
rect -4338 -166 -4156 166
rect -3416 50 -3376 169
rect -3356 50 -3316 169
rect -3240 166 -3034 534
rect -2294 531 -2254 650
rect -2234 531 -2194 650
rect -2094 534 -1912 866
rect -1172 750 -1132 869
rect -1112 750 -1072 869
rect -996 866 -790 1234
rect -50 1231 -10 1350
rect 10 1231 50 1350
rect 150 1234 332 1566
rect 1072 1450 1112 1569
rect 1132 1450 1172 1569
rect 1248 1566 1454 1934
rect 2194 1931 2234 2050
rect 2254 1931 2294 2050
rect 2394 1934 2576 2266
rect 3316 2150 3356 2269
rect 3376 2150 3416 2269
rect 3492 2266 3698 2634
rect 4438 2631 4478 2750
rect 4498 2631 4538 2750
rect 4638 2634 4820 2966
rect 4180 2589 4538 2631
rect 4180 2311 4222 2589
rect 4294 2311 4538 2589
rect 4180 2269 4538 2311
rect 1936 1889 2294 1931
rect 1936 1611 1978 1889
rect 2050 1611 2294 1889
rect 1936 1569 2294 1611
rect -308 1189 50 1231
rect -308 911 -266 1189
rect -194 911 50 1189
rect -308 869 50 911
rect -2552 489 -2194 531
rect -2552 211 -2510 489
rect -2438 211 -2194 489
rect -2552 169 -2194 211
rect -4796 -211 -4438 -169
rect -4796 -489 -4754 -211
rect -4682 -489 -4438 -211
rect -4796 -531 -4438 -489
rect -4538 -650 -4498 -531
rect -4478 -650 -4438 -531
rect -4362 -534 -4156 -166
rect -3416 -169 -3376 -50
rect -3356 -169 -3316 -50
rect -3216 -166 -3034 166
rect -2294 50 -2254 169
rect -2234 50 -2194 169
rect -2118 166 -1912 534
rect -1172 531 -1132 650
rect -1112 531 -1072 650
rect -972 534 -790 866
rect -50 750 -10 869
rect 10 750 50 869
rect 126 866 332 1234
rect 1072 1231 1112 1350
rect 1132 1231 1172 1350
rect 1272 1234 1454 1566
rect 2194 1450 2234 1569
rect 2254 1450 2294 1569
rect 2370 1566 2576 1934
rect 3316 1931 3356 2050
rect 3376 1931 3416 2050
rect 3516 1934 3698 2266
rect 4438 2150 4478 2269
rect 4498 2150 4538 2269
rect 4614 2266 4820 2634
rect 5302 2589 5622 2631
rect 5302 2311 5344 2589
rect 5302 2269 5622 2311
rect 3058 1889 3416 1931
rect 3058 1611 3100 1889
rect 3172 1611 3416 1889
rect 3058 1569 3416 1611
rect 814 1189 1172 1231
rect 814 911 856 1189
rect 928 911 1172 1189
rect 814 869 1172 911
rect -1430 489 -1072 531
rect -1430 211 -1388 489
rect -1316 211 -1072 489
rect -1430 169 -1072 211
rect -3674 -211 -3316 -169
rect -3674 -489 -3632 -211
rect -3560 -489 -3316 -211
rect -3674 -531 -3316 -489
rect -4538 -869 -4498 -750
rect -4478 -869 -4438 -750
rect -4338 -866 -4156 -534
rect -3416 -650 -3376 -531
rect -3356 -650 -3316 -531
rect -3240 -534 -3034 -166
rect -2294 -169 -2254 -50
rect -2234 -169 -2194 -50
rect -2094 -166 -1912 166
rect -1172 50 -1132 169
rect -1112 50 -1072 169
rect -996 166 -790 534
rect -50 531 -10 650
rect 10 531 50 650
rect 150 534 332 866
rect 1072 750 1112 869
rect 1132 750 1172 869
rect 1248 866 1454 1234
rect 2194 1231 2234 1350
rect 2254 1231 2294 1350
rect 2394 1234 2576 1566
rect 3316 1450 3356 1569
rect 3376 1450 3416 1569
rect 3492 1566 3698 1934
rect 4438 1931 4478 2050
rect 4498 1931 4538 2050
rect 4638 1934 4820 2266
rect 4180 1889 4538 1931
rect 4180 1611 4222 1889
rect 4294 1611 4538 1889
rect 4180 1569 4538 1611
rect 1936 1189 2294 1231
rect 1936 911 1978 1189
rect 2050 911 2294 1189
rect 1936 869 2294 911
rect -308 489 50 531
rect -308 211 -266 489
rect -194 211 50 489
rect -308 169 50 211
rect -2552 -211 -2194 -169
rect -2552 -489 -2510 -211
rect -2438 -489 -2194 -211
rect -2552 -531 -2194 -489
rect -4796 -911 -4438 -869
rect -4796 -1189 -4754 -911
rect -4682 -1189 -4438 -911
rect -4796 -1231 -4438 -1189
rect -4538 -1350 -4498 -1231
rect -4478 -1350 -4438 -1231
rect -4362 -1234 -4156 -866
rect -3416 -869 -3376 -750
rect -3356 -869 -3316 -750
rect -3216 -866 -3034 -534
rect -2294 -650 -2254 -531
rect -2234 -650 -2194 -531
rect -2118 -534 -1912 -166
rect -1172 -169 -1132 -50
rect -1112 -169 -1072 -50
rect -972 -166 -790 166
rect -50 50 -10 169
rect 10 50 50 169
rect 126 166 332 534
rect 1072 531 1112 650
rect 1132 531 1172 650
rect 1272 534 1454 866
rect 2194 750 2234 869
rect 2254 750 2294 869
rect 2370 866 2576 1234
rect 3316 1231 3356 1350
rect 3376 1231 3416 1350
rect 3516 1234 3698 1566
rect 4438 1450 4478 1569
rect 4498 1450 4538 1569
rect 4614 1566 4820 1934
rect 5302 1889 5622 1931
rect 5302 1611 5344 1889
rect 5302 1569 5622 1611
rect 3058 1189 3416 1231
rect 3058 911 3100 1189
rect 3172 911 3416 1189
rect 3058 869 3416 911
rect 814 489 1172 531
rect 814 211 856 489
rect 928 211 1172 489
rect 814 169 1172 211
rect -1430 -211 -1072 -169
rect -1430 -489 -1388 -211
rect -1316 -489 -1072 -211
rect -1430 -531 -1072 -489
rect -3674 -911 -3316 -869
rect -3674 -1189 -3632 -911
rect -3560 -1189 -3316 -911
rect -3674 -1231 -3316 -1189
rect -4538 -1569 -4498 -1450
rect -4478 -1569 -4438 -1450
rect -4338 -1566 -4156 -1234
rect -3416 -1350 -3376 -1231
rect -3356 -1350 -3316 -1231
rect -3240 -1234 -3034 -866
rect -2294 -869 -2254 -750
rect -2234 -869 -2194 -750
rect -2094 -866 -1912 -534
rect -1172 -650 -1132 -531
rect -1112 -650 -1072 -531
rect -996 -534 -790 -166
rect -50 -169 -10 -50
rect 10 -169 50 -50
rect 150 -166 332 166
rect 1072 50 1112 169
rect 1132 50 1172 169
rect 1248 166 1454 534
rect 2194 531 2234 650
rect 2254 531 2294 650
rect 2394 534 2576 866
rect 3316 750 3356 869
rect 3376 750 3416 869
rect 3492 866 3698 1234
rect 4438 1231 4478 1350
rect 4498 1231 4538 1350
rect 4638 1234 4820 1566
rect 4180 1189 4538 1231
rect 4180 911 4222 1189
rect 4294 911 4538 1189
rect 4180 869 4538 911
rect 1936 489 2294 531
rect 1936 211 1978 489
rect 2050 211 2294 489
rect 1936 169 2294 211
rect -308 -211 50 -169
rect -308 -489 -266 -211
rect -194 -489 50 -211
rect -308 -531 50 -489
rect -2552 -911 -2194 -869
rect -2552 -1189 -2510 -911
rect -2438 -1189 -2194 -911
rect -2552 -1231 -2194 -1189
rect -4796 -1611 -4438 -1569
rect -4796 -1889 -4754 -1611
rect -4682 -1889 -4438 -1611
rect -4796 -1931 -4438 -1889
rect -4538 -2050 -4498 -1931
rect -4478 -2050 -4438 -1931
rect -4362 -1934 -4156 -1566
rect -3416 -1569 -3376 -1450
rect -3356 -1569 -3316 -1450
rect -3216 -1566 -3034 -1234
rect -2294 -1350 -2254 -1231
rect -2234 -1350 -2194 -1231
rect -2118 -1234 -1912 -866
rect -1172 -869 -1132 -750
rect -1112 -869 -1072 -750
rect -972 -866 -790 -534
rect -50 -650 -10 -531
rect 10 -650 50 -531
rect 126 -534 332 -166
rect 1072 -169 1112 -50
rect 1132 -169 1172 -50
rect 1272 -166 1454 166
rect 2194 50 2234 169
rect 2254 50 2294 169
rect 2370 166 2576 534
rect 3316 531 3356 650
rect 3376 531 3416 650
rect 3516 534 3698 866
rect 4438 750 4478 869
rect 4498 750 4538 869
rect 4614 866 4820 1234
rect 5302 1189 5622 1231
rect 5302 911 5344 1189
rect 5302 869 5622 911
rect 3058 489 3416 531
rect 3058 211 3100 489
rect 3172 211 3416 489
rect 3058 169 3416 211
rect 814 -211 1172 -169
rect 814 -489 856 -211
rect 928 -489 1172 -211
rect 814 -531 1172 -489
rect -1430 -911 -1072 -869
rect -1430 -1189 -1388 -911
rect -1316 -1189 -1072 -911
rect -1430 -1231 -1072 -1189
rect -3674 -1611 -3316 -1569
rect -3674 -1889 -3632 -1611
rect -3560 -1889 -3316 -1611
rect -3674 -1931 -3316 -1889
rect -4538 -2269 -4498 -2150
rect -4478 -2269 -4438 -2150
rect -4338 -2266 -4156 -1934
rect -3416 -2050 -3376 -1931
rect -3356 -2050 -3316 -1931
rect -3240 -1934 -3034 -1566
rect -2294 -1569 -2254 -1450
rect -2234 -1569 -2194 -1450
rect -2094 -1566 -1912 -1234
rect -1172 -1350 -1132 -1231
rect -1112 -1350 -1072 -1231
rect -996 -1234 -790 -866
rect -50 -869 -10 -750
rect 10 -869 50 -750
rect 150 -866 332 -534
rect 1072 -650 1112 -531
rect 1132 -650 1172 -531
rect 1248 -534 1454 -166
rect 2194 -169 2234 -50
rect 2254 -169 2294 -50
rect 2394 -166 2576 166
rect 3316 50 3356 169
rect 3376 50 3416 169
rect 3492 166 3698 534
rect 4438 531 4478 650
rect 4498 531 4538 650
rect 4638 534 4820 866
rect 4180 489 4538 531
rect 4180 211 4222 489
rect 4294 211 4538 489
rect 4180 169 4538 211
rect 1936 -211 2294 -169
rect 1936 -489 1978 -211
rect 2050 -489 2294 -211
rect 1936 -531 2294 -489
rect -308 -911 50 -869
rect -308 -1189 -266 -911
rect -194 -1189 50 -911
rect -308 -1231 50 -1189
rect -2552 -1611 -2194 -1569
rect -2552 -1889 -2510 -1611
rect -2438 -1889 -2194 -1611
rect -2552 -1931 -2194 -1889
rect -4796 -2311 -4438 -2269
rect -4796 -2589 -4754 -2311
rect -4682 -2589 -4438 -2311
rect -4796 -2631 -4438 -2589
rect -4538 -2750 -4498 -2631
rect -4478 -2750 -4438 -2631
rect -4362 -2634 -4156 -2266
rect -3416 -2269 -3376 -2150
rect -3356 -2269 -3316 -2150
rect -3216 -2266 -3034 -1934
rect -2294 -2050 -2254 -1931
rect -2234 -2050 -2194 -1931
rect -2118 -1934 -1912 -1566
rect -1172 -1569 -1132 -1450
rect -1112 -1569 -1072 -1450
rect -972 -1566 -790 -1234
rect -50 -1350 -10 -1231
rect 10 -1350 50 -1231
rect 126 -1234 332 -866
rect 1072 -869 1112 -750
rect 1132 -869 1172 -750
rect 1272 -866 1454 -534
rect 2194 -650 2234 -531
rect 2254 -650 2294 -531
rect 2370 -534 2576 -166
rect 3316 -169 3356 -50
rect 3376 -169 3416 -50
rect 3516 -166 3698 166
rect 4438 50 4478 169
rect 4498 50 4538 169
rect 4614 166 4820 534
rect 5302 489 5622 531
rect 5302 211 5344 489
rect 5302 169 5622 211
rect 3058 -211 3416 -169
rect 3058 -489 3100 -211
rect 3172 -489 3416 -211
rect 3058 -531 3416 -489
rect 814 -911 1172 -869
rect 814 -1189 856 -911
rect 928 -1189 1172 -911
rect 814 -1231 1172 -1189
rect -1430 -1611 -1072 -1569
rect -1430 -1889 -1388 -1611
rect -1316 -1889 -1072 -1611
rect -1430 -1931 -1072 -1889
rect -3674 -2311 -3316 -2269
rect -3674 -2589 -3632 -2311
rect -3560 -2589 -3316 -2311
rect -3674 -2631 -3316 -2589
rect -4538 -2969 -4498 -2850
rect -4478 -2969 -4438 -2850
rect -4338 -2966 -4156 -2634
rect -3416 -2750 -3376 -2631
rect -3356 -2750 -3316 -2631
rect -3240 -2634 -3034 -2266
rect -2294 -2269 -2254 -2150
rect -2234 -2269 -2194 -2150
rect -2094 -2266 -1912 -1934
rect -1172 -2050 -1132 -1931
rect -1112 -2050 -1072 -1931
rect -996 -1934 -790 -1566
rect -50 -1569 -10 -1450
rect 10 -1569 50 -1450
rect 150 -1566 332 -1234
rect 1072 -1350 1112 -1231
rect 1132 -1350 1172 -1231
rect 1248 -1234 1454 -866
rect 2194 -869 2234 -750
rect 2254 -869 2294 -750
rect 2394 -866 2576 -534
rect 3316 -650 3356 -531
rect 3376 -650 3416 -531
rect 3492 -534 3698 -166
rect 4438 -169 4478 -50
rect 4498 -169 4538 -50
rect 4638 -166 4820 166
rect 4180 -211 4538 -169
rect 4180 -489 4222 -211
rect 4294 -489 4538 -211
rect 4180 -531 4538 -489
rect 1936 -911 2294 -869
rect 1936 -1189 1978 -911
rect 2050 -1189 2294 -911
rect 1936 -1231 2294 -1189
rect -308 -1611 50 -1569
rect -308 -1889 -266 -1611
rect -194 -1889 50 -1611
rect -308 -1931 50 -1889
rect -2552 -2311 -2194 -2269
rect -2552 -2589 -2510 -2311
rect -2438 -2589 -2194 -2311
rect -2552 -2631 -2194 -2589
rect -4796 -3011 -4438 -2969
rect -4796 -3289 -4754 -3011
rect -4682 -3289 -4438 -3011
rect -4796 -3331 -4438 -3289
rect -4538 -3450 -4498 -3331
rect -4478 -3450 -4438 -3331
rect -4362 -3334 -4156 -2966
rect -3416 -2969 -3376 -2850
rect -3356 -2969 -3316 -2850
rect -3216 -2966 -3034 -2634
rect -2294 -2750 -2254 -2631
rect -2234 -2750 -2194 -2631
rect -2118 -2634 -1912 -2266
rect -1172 -2269 -1132 -2150
rect -1112 -2269 -1072 -2150
rect -972 -2266 -790 -1934
rect -50 -2050 -10 -1931
rect 10 -2050 50 -1931
rect 126 -1934 332 -1566
rect 1072 -1569 1112 -1450
rect 1132 -1569 1172 -1450
rect 1272 -1566 1454 -1234
rect 2194 -1350 2234 -1231
rect 2254 -1350 2294 -1231
rect 2370 -1234 2576 -866
rect 3316 -869 3356 -750
rect 3376 -869 3416 -750
rect 3516 -866 3698 -534
rect 4438 -650 4478 -531
rect 4498 -650 4538 -531
rect 4614 -534 4820 -166
rect 5302 -211 5622 -169
rect 5302 -489 5344 -211
rect 5302 -531 5622 -489
rect 3058 -911 3416 -869
rect 3058 -1189 3100 -911
rect 3172 -1189 3416 -911
rect 3058 -1231 3416 -1189
rect 814 -1611 1172 -1569
rect 814 -1889 856 -1611
rect 928 -1889 1172 -1611
rect 814 -1931 1172 -1889
rect -1430 -2311 -1072 -2269
rect -1430 -2589 -1388 -2311
rect -1316 -2589 -1072 -2311
rect -1430 -2631 -1072 -2589
rect -3674 -3011 -3316 -2969
rect -3674 -3289 -3632 -3011
rect -3560 -3289 -3316 -3011
rect -3674 -3331 -3316 -3289
rect -4338 -3500 -4156 -3334
rect -3416 -3450 -3376 -3331
rect -3356 -3450 -3316 -3331
rect -3240 -3334 -3034 -2966
rect -2294 -2969 -2254 -2850
rect -2234 -2969 -2194 -2850
rect -2094 -2966 -1912 -2634
rect -1172 -2750 -1132 -2631
rect -1112 -2750 -1072 -2631
rect -996 -2634 -790 -2266
rect -50 -2269 -10 -2150
rect 10 -2269 50 -2150
rect 150 -2266 332 -1934
rect 1072 -2050 1112 -1931
rect 1132 -2050 1172 -1931
rect 1248 -1934 1454 -1566
rect 2194 -1569 2234 -1450
rect 2254 -1569 2294 -1450
rect 2394 -1566 2576 -1234
rect 3316 -1350 3356 -1231
rect 3376 -1350 3416 -1231
rect 3492 -1234 3698 -866
rect 4438 -869 4478 -750
rect 4498 -869 4538 -750
rect 4638 -866 4820 -534
rect 4180 -911 4538 -869
rect 4180 -1189 4222 -911
rect 4294 -1189 4538 -911
rect 4180 -1231 4538 -1189
rect 1936 -1611 2294 -1569
rect 1936 -1889 1978 -1611
rect 2050 -1889 2294 -1611
rect 1936 -1931 2294 -1889
rect -308 -2311 50 -2269
rect -308 -2589 -266 -2311
rect -194 -2589 50 -2311
rect -308 -2631 50 -2589
rect -2552 -3011 -2194 -2969
rect -2552 -3289 -2510 -3011
rect -2438 -3289 -2194 -3011
rect -2552 -3331 -2194 -3289
rect -3216 -3500 -3034 -3334
rect -2294 -3450 -2254 -3331
rect -2234 -3450 -2194 -3331
rect -2118 -3334 -1912 -2966
rect -1172 -2969 -1132 -2850
rect -1112 -2969 -1072 -2850
rect -972 -2966 -790 -2634
rect -50 -2750 -10 -2631
rect 10 -2750 50 -2631
rect 126 -2634 332 -2266
rect 1072 -2269 1112 -2150
rect 1132 -2269 1172 -2150
rect 1272 -2266 1454 -1934
rect 2194 -2050 2234 -1931
rect 2254 -2050 2294 -1931
rect 2370 -1934 2576 -1566
rect 3316 -1569 3356 -1450
rect 3376 -1569 3416 -1450
rect 3516 -1566 3698 -1234
rect 4438 -1350 4478 -1231
rect 4498 -1350 4538 -1231
rect 4614 -1234 4820 -866
rect 5302 -911 5622 -869
rect 5302 -1189 5344 -911
rect 5302 -1231 5622 -1189
rect 3058 -1611 3416 -1569
rect 3058 -1889 3100 -1611
rect 3172 -1889 3416 -1611
rect 3058 -1931 3416 -1889
rect 814 -2311 1172 -2269
rect 814 -2589 856 -2311
rect 928 -2589 1172 -2311
rect 814 -2631 1172 -2589
rect -1430 -3011 -1072 -2969
rect -1430 -3289 -1388 -3011
rect -1316 -3289 -1072 -3011
rect -1430 -3331 -1072 -3289
rect -2094 -3500 -1912 -3334
rect -1172 -3450 -1132 -3331
rect -1112 -3450 -1072 -3331
rect -996 -3334 -790 -2966
rect -50 -2969 -10 -2850
rect 10 -2969 50 -2850
rect 150 -2966 332 -2634
rect 1072 -2750 1112 -2631
rect 1132 -2750 1172 -2631
rect 1248 -2634 1454 -2266
rect 2194 -2269 2234 -2150
rect 2254 -2269 2294 -2150
rect 2394 -2266 2576 -1934
rect 3316 -2050 3356 -1931
rect 3376 -2050 3416 -1931
rect 3492 -1934 3698 -1566
rect 4438 -1569 4478 -1450
rect 4498 -1569 4538 -1450
rect 4638 -1566 4820 -1234
rect 4180 -1611 4538 -1569
rect 4180 -1889 4222 -1611
rect 4294 -1889 4538 -1611
rect 4180 -1931 4538 -1889
rect 1936 -2311 2294 -2269
rect 1936 -2589 1978 -2311
rect 2050 -2589 2294 -2311
rect 1936 -2631 2294 -2589
rect -308 -3011 50 -2969
rect -308 -3289 -266 -3011
rect -194 -3289 50 -3011
rect -308 -3331 50 -3289
rect -972 -3500 -790 -3334
rect -50 -3450 -10 -3331
rect 10 -3450 50 -3331
rect 126 -3334 332 -2966
rect 1072 -2969 1112 -2850
rect 1132 -2969 1172 -2850
rect 1272 -2966 1454 -2634
rect 2194 -2750 2234 -2631
rect 2254 -2750 2294 -2631
rect 2370 -2634 2576 -2266
rect 3316 -2269 3356 -2150
rect 3376 -2269 3416 -2150
rect 3516 -2266 3698 -1934
rect 4438 -2050 4478 -1931
rect 4498 -2050 4538 -1931
rect 4614 -1934 4820 -1566
rect 5302 -1611 5622 -1569
rect 5302 -1889 5344 -1611
rect 5302 -1931 5622 -1889
rect 3058 -2311 3416 -2269
rect 3058 -2589 3100 -2311
rect 3172 -2589 3416 -2311
rect 3058 -2631 3416 -2589
rect 814 -3011 1172 -2969
rect 814 -3289 856 -3011
rect 928 -3289 1172 -3011
rect 814 -3331 1172 -3289
rect 150 -3500 332 -3334
rect 1072 -3450 1112 -3331
rect 1132 -3450 1172 -3331
rect 1248 -3334 1454 -2966
rect 2194 -2969 2234 -2850
rect 2254 -2969 2294 -2850
rect 2394 -2966 2576 -2634
rect 3316 -2750 3356 -2631
rect 3376 -2750 3416 -2631
rect 3492 -2634 3698 -2266
rect 4438 -2269 4478 -2150
rect 4498 -2269 4538 -2150
rect 4638 -2266 4820 -1934
rect 4180 -2311 4538 -2269
rect 4180 -2589 4222 -2311
rect 4294 -2589 4538 -2311
rect 4180 -2631 4538 -2589
rect 1936 -3011 2294 -2969
rect 1936 -3289 1978 -3011
rect 2050 -3289 2294 -3011
rect 1936 -3331 2294 -3289
rect 1272 -3500 1454 -3334
rect 2194 -3450 2234 -3331
rect 2254 -3450 2294 -3331
rect 2370 -3334 2576 -2966
rect 3316 -2969 3356 -2850
rect 3376 -2969 3416 -2850
rect 3516 -2966 3698 -2634
rect 4438 -2750 4478 -2631
rect 4498 -2750 4538 -2631
rect 4614 -2634 4820 -2266
rect 5302 -2311 5622 -2269
rect 5302 -2589 5344 -2311
rect 5302 -2631 5622 -2589
rect 3058 -3011 3416 -2969
rect 3058 -3289 3100 -3011
rect 3172 -3289 3416 -3011
rect 3058 -3331 3416 -3289
rect 2394 -3500 2576 -3334
rect 3316 -3450 3356 -3331
rect 3376 -3450 3416 -3331
rect 3492 -3334 3698 -2966
rect 4438 -2969 4478 -2850
rect 4498 -2969 4538 -2850
rect 4638 -2966 4820 -2634
rect 4180 -3011 4538 -2969
rect 4180 -3289 4222 -3011
rect 4294 -3289 4538 -3011
rect 4180 -3331 4538 -3289
rect 3516 -3500 3698 -3334
rect 4438 -3450 4478 -3331
rect 4498 -3450 4538 -3331
rect 4614 -3334 4820 -2966
rect 5302 -3011 5622 -2969
rect 5302 -3289 5344 -3011
rect 5302 -3331 5622 -3289
rect 4638 -3500 4820 -3334
<< metal4 >>
rect -5600 3289 -4498 3450
rect -5600 3011 -4754 3289
rect -4518 3011 -4498 3289
rect -5600 2850 -4498 3011
rect -4478 3289 -3376 3450
rect -4478 3011 -3632 3289
rect -3396 3011 -3376 3289
rect -4478 2850 -3376 3011
rect -3356 3289 -2254 3450
rect -3356 3011 -2510 3289
rect -2274 3011 -2254 3289
rect -3356 2850 -2254 3011
rect -2234 3289 -1132 3450
rect -2234 3011 -1388 3289
rect -1152 3011 -1132 3289
rect -2234 2850 -1132 3011
rect -1112 3289 -10 3450
rect -1112 3011 -266 3289
rect -30 3011 -10 3289
rect -1112 2850 -10 3011
rect 10 3289 1112 3450
rect 10 3011 856 3289
rect 1092 3011 1112 3289
rect 10 2850 1112 3011
rect 1132 3289 2234 3450
rect 1132 3011 1978 3289
rect 2214 3011 2234 3289
rect 1132 2850 2234 3011
rect 2254 3289 3356 3450
rect 2254 3011 3100 3289
rect 3336 3011 3356 3289
rect 2254 2850 3356 3011
rect 3376 3289 4478 3450
rect 3376 3011 4222 3289
rect 4458 3011 4478 3289
rect 3376 2850 4478 3011
rect 4498 3289 5600 3450
rect 4498 3011 5344 3289
rect 5580 3011 5600 3289
rect 4498 2850 5600 3011
rect -5600 2589 -4498 2750
rect -5600 2311 -4754 2589
rect -4518 2311 -4498 2589
rect -5600 2150 -4498 2311
rect -4478 2589 -3376 2750
rect -4478 2311 -3632 2589
rect -3396 2311 -3376 2589
rect -4478 2150 -3376 2311
rect -3356 2589 -2254 2750
rect -3356 2311 -2510 2589
rect -2274 2311 -2254 2589
rect -3356 2150 -2254 2311
rect -2234 2589 -1132 2750
rect -2234 2311 -1388 2589
rect -1152 2311 -1132 2589
rect -2234 2150 -1132 2311
rect -1112 2589 -10 2750
rect -1112 2311 -266 2589
rect -30 2311 -10 2589
rect -1112 2150 -10 2311
rect 10 2589 1112 2750
rect 10 2311 856 2589
rect 1092 2311 1112 2589
rect 10 2150 1112 2311
rect 1132 2589 2234 2750
rect 1132 2311 1978 2589
rect 2214 2311 2234 2589
rect 1132 2150 2234 2311
rect 2254 2589 3356 2750
rect 2254 2311 3100 2589
rect 3336 2311 3356 2589
rect 2254 2150 3356 2311
rect 3376 2589 4478 2750
rect 3376 2311 4222 2589
rect 4458 2311 4478 2589
rect 3376 2150 4478 2311
rect 4498 2589 5600 2750
rect 4498 2311 5344 2589
rect 5580 2311 5600 2589
rect 4498 2150 5600 2311
rect -5600 1889 -4498 2050
rect -5600 1611 -4754 1889
rect -4518 1611 -4498 1889
rect -5600 1450 -4498 1611
rect -4478 1889 -3376 2050
rect -4478 1611 -3632 1889
rect -3396 1611 -3376 1889
rect -4478 1450 -3376 1611
rect -3356 1889 -2254 2050
rect -3356 1611 -2510 1889
rect -2274 1611 -2254 1889
rect -3356 1450 -2254 1611
rect -2234 1889 -1132 2050
rect -2234 1611 -1388 1889
rect -1152 1611 -1132 1889
rect -2234 1450 -1132 1611
rect -1112 1889 -10 2050
rect -1112 1611 -266 1889
rect -30 1611 -10 1889
rect -1112 1450 -10 1611
rect 10 1889 1112 2050
rect 10 1611 856 1889
rect 1092 1611 1112 1889
rect 10 1450 1112 1611
rect 1132 1889 2234 2050
rect 1132 1611 1978 1889
rect 2214 1611 2234 1889
rect 1132 1450 2234 1611
rect 2254 1889 3356 2050
rect 2254 1611 3100 1889
rect 3336 1611 3356 1889
rect 2254 1450 3356 1611
rect 3376 1889 4478 2050
rect 3376 1611 4222 1889
rect 4458 1611 4478 1889
rect 3376 1450 4478 1611
rect 4498 1889 5600 2050
rect 4498 1611 5344 1889
rect 5580 1611 5600 1889
rect 4498 1450 5600 1611
rect -5600 1189 -4498 1350
rect -5600 911 -4754 1189
rect -4518 911 -4498 1189
rect -5600 750 -4498 911
rect -4478 1189 -3376 1350
rect -4478 911 -3632 1189
rect -3396 911 -3376 1189
rect -4478 750 -3376 911
rect -3356 1189 -2254 1350
rect -3356 911 -2510 1189
rect -2274 911 -2254 1189
rect -3356 750 -2254 911
rect -2234 1189 -1132 1350
rect -2234 911 -1388 1189
rect -1152 911 -1132 1189
rect -2234 750 -1132 911
rect -1112 1189 -10 1350
rect -1112 911 -266 1189
rect -30 911 -10 1189
rect -1112 750 -10 911
rect 10 1189 1112 1350
rect 10 911 856 1189
rect 1092 911 1112 1189
rect 10 750 1112 911
rect 1132 1189 2234 1350
rect 1132 911 1978 1189
rect 2214 911 2234 1189
rect 1132 750 2234 911
rect 2254 1189 3356 1350
rect 2254 911 3100 1189
rect 3336 911 3356 1189
rect 2254 750 3356 911
rect 3376 1189 4478 1350
rect 3376 911 4222 1189
rect 4458 911 4478 1189
rect 3376 750 4478 911
rect 4498 1189 5600 1350
rect 4498 911 5344 1189
rect 5580 911 5600 1189
rect 4498 750 5600 911
rect -5600 489 -4498 650
rect -5600 211 -4754 489
rect -4518 211 -4498 489
rect -5600 50 -4498 211
rect -4478 489 -3376 650
rect -4478 211 -3632 489
rect -3396 211 -3376 489
rect -4478 50 -3376 211
rect -3356 489 -2254 650
rect -3356 211 -2510 489
rect -2274 211 -2254 489
rect -3356 50 -2254 211
rect -2234 489 -1132 650
rect -2234 211 -1388 489
rect -1152 211 -1132 489
rect -2234 50 -1132 211
rect -1112 489 -10 650
rect -1112 211 -266 489
rect -30 211 -10 489
rect -1112 50 -10 211
rect 10 489 1112 650
rect 10 211 856 489
rect 1092 211 1112 489
rect 10 50 1112 211
rect 1132 489 2234 650
rect 1132 211 1978 489
rect 2214 211 2234 489
rect 1132 50 2234 211
rect 2254 489 3356 650
rect 2254 211 3100 489
rect 3336 211 3356 489
rect 2254 50 3356 211
rect 3376 489 4478 650
rect 3376 211 4222 489
rect 4458 211 4478 489
rect 3376 50 4478 211
rect 4498 489 5600 650
rect 4498 211 5344 489
rect 5580 211 5600 489
rect 4498 50 5600 211
rect -5600 -211 -4498 -50
rect -5600 -489 -4754 -211
rect -4518 -489 -4498 -211
rect -5600 -650 -4498 -489
rect -4478 -211 -3376 -50
rect -4478 -489 -3632 -211
rect -3396 -489 -3376 -211
rect -4478 -650 -3376 -489
rect -3356 -211 -2254 -50
rect -3356 -489 -2510 -211
rect -2274 -489 -2254 -211
rect -3356 -650 -2254 -489
rect -2234 -211 -1132 -50
rect -2234 -489 -1388 -211
rect -1152 -489 -1132 -211
rect -2234 -650 -1132 -489
rect -1112 -211 -10 -50
rect -1112 -489 -266 -211
rect -30 -489 -10 -211
rect -1112 -650 -10 -489
rect 10 -211 1112 -50
rect 10 -489 856 -211
rect 1092 -489 1112 -211
rect 10 -650 1112 -489
rect 1132 -211 2234 -50
rect 1132 -489 1978 -211
rect 2214 -489 2234 -211
rect 1132 -650 2234 -489
rect 2254 -211 3356 -50
rect 2254 -489 3100 -211
rect 3336 -489 3356 -211
rect 2254 -650 3356 -489
rect 3376 -211 4478 -50
rect 3376 -489 4222 -211
rect 4458 -489 4478 -211
rect 3376 -650 4478 -489
rect 4498 -211 5600 -50
rect 4498 -489 5344 -211
rect 5580 -489 5600 -211
rect 4498 -650 5600 -489
rect -5600 -911 -4498 -750
rect -5600 -1189 -4754 -911
rect -4518 -1189 -4498 -911
rect -5600 -1350 -4498 -1189
rect -4478 -911 -3376 -750
rect -4478 -1189 -3632 -911
rect -3396 -1189 -3376 -911
rect -4478 -1350 -3376 -1189
rect -3356 -911 -2254 -750
rect -3356 -1189 -2510 -911
rect -2274 -1189 -2254 -911
rect -3356 -1350 -2254 -1189
rect -2234 -911 -1132 -750
rect -2234 -1189 -1388 -911
rect -1152 -1189 -1132 -911
rect -2234 -1350 -1132 -1189
rect -1112 -911 -10 -750
rect -1112 -1189 -266 -911
rect -30 -1189 -10 -911
rect -1112 -1350 -10 -1189
rect 10 -911 1112 -750
rect 10 -1189 856 -911
rect 1092 -1189 1112 -911
rect 10 -1350 1112 -1189
rect 1132 -911 2234 -750
rect 1132 -1189 1978 -911
rect 2214 -1189 2234 -911
rect 1132 -1350 2234 -1189
rect 2254 -911 3356 -750
rect 2254 -1189 3100 -911
rect 3336 -1189 3356 -911
rect 2254 -1350 3356 -1189
rect 3376 -911 4478 -750
rect 3376 -1189 4222 -911
rect 4458 -1189 4478 -911
rect 3376 -1350 4478 -1189
rect 4498 -911 5600 -750
rect 4498 -1189 5344 -911
rect 5580 -1189 5600 -911
rect 4498 -1350 5600 -1189
rect -5600 -1611 -4498 -1450
rect -5600 -1889 -4754 -1611
rect -4518 -1889 -4498 -1611
rect -5600 -2050 -4498 -1889
rect -4478 -1611 -3376 -1450
rect -4478 -1889 -3632 -1611
rect -3396 -1889 -3376 -1611
rect -4478 -2050 -3376 -1889
rect -3356 -1611 -2254 -1450
rect -3356 -1889 -2510 -1611
rect -2274 -1889 -2254 -1611
rect -3356 -2050 -2254 -1889
rect -2234 -1611 -1132 -1450
rect -2234 -1889 -1388 -1611
rect -1152 -1889 -1132 -1611
rect -2234 -2050 -1132 -1889
rect -1112 -1611 -10 -1450
rect -1112 -1889 -266 -1611
rect -30 -1889 -10 -1611
rect -1112 -2050 -10 -1889
rect 10 -1611 1112 -1450
rect 10 -1889 856 -1611
rect 1092 -1889 1112 -1611
rect 10 -2050 1112 -1889
rect 1132 -1611 2234 -1450
rect 1132 -1889 1978 -1611
rect 2214 -1889 2234 -1611
rect 1132 -2050 2234 -1889
rect 2254 -1611 3356 -1450
rect 2254 -1889 3100 -1611
rect 3336 -1889 3356 -1611
rect 2254 -2050 3356 -1889
rect 3376 -1611 4478 -1450
rect 3376 -1889 4222 -1611
rect 4458 -1889 4478 -1611
rect 3376 -2050 4478 -1889
rect 4498 -1611 5600 -1450
rect 4498 -1889 5344 -1611
rect 5580 -1889 5600 -1611
rect 4498 -2050 5600 -1889
rect -5600 -2311 -4498 -2150
rect -5600 -2589 -4754 -2311
rect -4518 -2589 -4498 -2311
rect -5600 -2750 -4498 -2589
rect -4478 -2311 -3376 -2150
rect -4478 -2589 -3632 -2311
rect -3396 -2589 -3376 -2311
rect -4478 -2750 -3376 -2589
rect -3356 -2311 -2254 -2150
rect -3356 -2589 -2510 -2311
rect -2274 -2589 -2254 -2311
rect -3356 -2750 -2254 -2589
rect -2234 -2311 -1132 -2150
rect -2234 -2589 -1388 -2311
rect -1152 -2589 -1132 -2311
rect -2234 -2750 -1132 -2589
rect -1112 -2311 -10 -2150
rect -1112 -2589 -266 -2311
rect -30 -2589 -10 -2311
rect -1112 -2750 -10 -2589
rect 10 -2311 1112 -2150
rect 10 -2589 856 -2311
rect 1092 -2589 1112 -2311
rect 10 -2750 1112 -2589
rect 1132 -2311 2234 -2150
rect 1132 -2589 1978 -2311
rect 2214 -2589 2234 -2311
rect 1132 -2750 2234 -2589
rect 2254 -2311 3356 -2150
rect 2254 -2589 3100 -2311
rect 3336 -2589 3356 -2311
rect 2254 -2750 3356 -2589
rect 3376 -2311 4478 -2150
rect 3376 -2589 4222 -2311
rect 4458 -2589 4478 -2311
rect 3376 -2750 4478 -2589
rect 4498 -2311 5600 -2150
rect 4498 -2589 5344 -2311
rect 5580 -2589 5600 -2311
rect 4498 -2750 5600 -2589
rect -5600 -3011 -4498 -2850
rect -5600 -3289 -4754 -3011
rect -4518 -3289 -4498 -3011
rect -5600 -3450 -4498 -3289
rect -4478 -3011 -3376 -2850
rect -4478 -3289 -3632 -3011
rect -3396 -3289 -3376 -3011
rect -4478 -3450 -3376 -3289
rect -3356 -3011 -2254 -2850
rect -3356 -3289 -2510 -3011
rect -2274 -3289 -2254 -3011
rect -3356 -3450 -2254 -3289
rect -2234 -3011 -1132 -2850
rect -2234 -3289 -1388 -3011
rect -1152 -3289 -1132 -3011
rect -2234 -3450 -1132 -3289
rect -1112 -3011 -10 -2850
rect -1112 -3289 -266 -3011
rect -30 -3289 -10 -3011
rect -1112 -3450 -10 -3289
rect 10 -3011 1112 -2850
rect 10 -3289 856 -3011
rect 1092 -3289 1112 -3011
rect 10 -3450 1112 -3289
rect 1132 -3011 2234 -2850
rect 1132 -3289 1978 -3011
rect 2214 -3289 2234 -3011
rect 1132 -3450 2234 -3289
rect 2254 -3011 3356 -2850
rect 2254 -3289 3100 -3011
rect 3336 -3289 3356 -3011
rect 2254 -3450 3356 -3289
rect 3376 -3011 4478 -2850
rect 3376 -3289 4222 -3011
rect 4458 -3289 4478 -3011
rect 3376 -3450 4478 -3289
rect 4498 -3011 5600 -2850
rect 4498 -3289 5344 -3011
rect 5580 -3289 5600 -3011
rect 4498 -3450 5600 -3289
<< via4 >>
rect -4754 3011 -4518 3289
rect -3632 3011 -3396 3289
rect -2510 3011 -2274 3289
rect -1388 3011 -1152 3289
rect -266 3011 -30 3289
rect 856 3011 1092 3289
rect 1978 3011 2214 3289
rect 3100 3011 3336 3289
rect 4222 3011 4458 3289
rect 5344 3011 5580 3289
rect -4754 2311 -4518 2589
rect -3632 2311 -3396 2589
rect -2510 2311 -2274 2589
rect -1388 2311 -1152 2589
rect -266 2311 -30 2589
rect 856 2311 1092 2589
rect 1978 2311 2214 2589
rect 3100 2311 3336 2589
rect 4222 2311 4458 2589
rect 5344 2311 5580 2589
rect -4754 1611 -4518 1889
rect -3632 1611 -3396 1889
rect -2510 1611 -2274 1889
rect -1388 1611 -1152 1889
rect -266 1611 -30 1889
rect 856 1611 1092 1889
rect 1978 1611 2214 1889
rect 3100 1611 3336 1889
rect 4222 1611 4458 1889
rect 5344 1611 5580 1889
rect -4754 911 -4518 1189
rect -3632 911 -3396 1189
rect -2510 911 -2274 1189
rect -1388 911 -1152 1189
rect -266 911 -30 1189
rect 856 911 1092 1189
rect 1978 911 2214 1189
rect 3100 911 3336 1189
rect 4222 911 4458 1189
rect 5344 911 5580 1189
rect -4754 211 -4518 489
rect -3632 211 -3396 489
rect -2510 211 -2274 489
rect -1388 211 -1152 489
rect -266 211 -30 489
rect 856 211 1092 489
rect 1978 211 2214 489
rect 3100 211 3336 489
rect 4222 211 4458 489
rect 5344 211 5580 489
rect -4754 -489 -4518 -211
rect -3632 -489 -3396 -211
rect -2510 -489 -2274 -211
rect -1388 -489 -1152 -211
rect -266 -489 -30 -211
rect 856 -489 1092 -211
rect 1978 -489 2214 -211
rect 3100 -489 3336 -211
rect 4222 -489 4458 -211
rect 5344 -489 5580 -211
rect -4754 -1189 -4518 -911
rect -3632 -1189 -3396 -911
rect -2510 -1189 -2274 -911
rect -1388 -1189 -1152 -911
rect -266 -1189 -30 -911
rect 856 -1189 1092 -911
rect 1978 -1189 2214 -911
rect 3100 -1189 3336 -911
rect 4222 -1189 4458 -911
rect 5344 -1189 5580 -911
rect -4754 -1889 -4518 -1611
rect -3632 -1889 -3396 -1611
rect -2510 -1889 -2274 -1611
rect -1388 -1889 -1152 -1611
rect -266 -1889 -30 -1611
rect 856 -1889 1092 -1611
rect 1978 -1889 2214 -1611
rect 3100 -1889 3336 -1611
rect 4222 -1889 4458 -1611
rect 5344 -1889 5580 -1611
rect -4754 -2589 -4518 -2311
rect -3632 -2589 -3396 -2311
rect -2510 -2589 -2274 -2311
rect -1388 -2589 -1152 -2311
rect -266 -2589 -30 -2311
rect 856 -2589 1092 -2311
rect 1978 -2589 2214 -2311
rect 3100 -2589 3336 -2311
rect 4222 -2589 4458 -2311
rect 5344 -2589 5580 -2311
rect -4754 -3289 -4518 -3011
rect -3632 -3289 -3396 -3011
rect -2510 -3289 -2274 -3011
rect -1388 -3289 -1152 -3011
rect -266 -3289 -30 -3011
rect 856 -3289 1092 -3011
rect 1978 -3289 2214 -3011
rect 3100 -3289 3336 -3011
rect 4222 -3289 4458 -3011
rect 5344 -3289 5580 -3011
<< mimcap2 >>
rect -5500 3310 -5100 3350
rect -5500 2990 -5460 3310
rect -5140 2990 -5100 3310
rect -5500 2950 -5100 2990
rect -4378 3310 -3978 3350
rect -4378 2990 -4338 3310
rect -4018 2990 -3978 3310
rect -4378 2950 -3978 2990
rect -3256 3310 -2856 3350
rect -3256 2990 -3216 3310
rect -2896 2990 -2856 3310
rect -3256 2950 -2856 2990
rect -2134 3310 -1734 3350
rect -2134 2990 -2094 3310
rect -1774 2990 -1734 3310
rect -2134 2950 -1734 2990
rect -1012 3310 -612 3350
rect -1012 2990 -972 3310
rect -652 2990 -612 3310
rect -1012 2950 -612 2990
rect 110 3310 510 3350
rect 110 2990 150 3310
rect 470 2990 510 3310
rect 110 2950 510 2990
rect 1232 3310 1632 3350
rect 1232 2990 1272 3310
rect 1592 2990 1632 3310
rect 1232 2950 1632 2990
rect 2354 3310 2754 3350
rect 2354 2990 2394 3310
rect 2714 2990 2754 3310
rect 2354 2950 2754 2990
rect 3476 3310 3876 3350
rect 3476 2990 3516 3310
rect 3836 2990 3876 3310
rect 3476 2950 3876 2990
rect 4598 3310 4998 3350
rect 4598 2990 4638 3310
rect 4958 2990 4998 3310
rect 4598 2950 4998 2990
rect -5500 2610 -5100 2650
rect -5500 2290 -5460 2610
rect -5140 2290 -5100 2610
rect -5500 2250 -5100 2290
rect -4378 2610 -3978 2650
rect -4378 2290 -4338 2610
rect -4018 2290 -3978 2610
rect -4378 2250 -3978 2290
rect -3256 2610 -2856 2650
rect -3256 2290 -3216 2610
rect -2896 2290 -2856 2610
rect -3256 2250 -2856 2290
rect -2134 2610 -1734 2650
rect -2134 2290 -2094 2610
rect -1774 2290 -1734 2610
rect -2134 2250 -1734 2290
rect -1012 2610 -612 2650
rect -1012 2290 -972 2610
rect -652 2290 -612 2610
rect -1012 2250 -612 2290
rect 110 2610 510 2650
rect 110 2290 150 2610
rect 470 2290 510 2610
rect 110 2250 510 2290
rect 1232 2610 1632 2650
rect 1232 2290 1272 2610
rect 1592 2290 1632 2610
rect 1232 2250 1632 2290
rect 2354 2610 2754 2650
rect 2354 2290 2394 2610
rect 2714 2290 2754 2610
rect 2354 2250 2754 2290
rect 3476 2610 3876 2650
rect 3476 2290 3516 2610
rect 3836 2290 3876 2610
rect 3476 2250 3876 2290
rect 4598 2610 4998 2650
rect 4598 2290 4638 2610
rect 4958 2290 4998 2610
rect 4598 2250 4998 2290
rect -5500 1910 -5100 1950
rect -5500 1590 -5460 1910
rect -5140 1590 -5100 1910
rect -5500 1550 -5100 1590
rect -4378 1910 -3978 1950
rect -4378 1590 -4338 1910
rect -4018 1590 -3978 1910
rect -4378 1550 -3978 1590
rect -3256 1910 -2856 1950
rect -3256 1590 -3216 1910
rect -2896 1590 -2856 1910
rect -3256 1550 -2856 1590
rect -2134 1910 -1734 1950
rect -2134 1590 -2094 1910
rect -1774 1590 -1734 1910
rect -2134 1550 -1734 1590
rect -1012 1910 -612 1950
rect -1012 1590 -972 1910
rect -652 1590 -612 1910
rect -1012 1550 -612 1590
rect 110 1910 510 1950
rect 110 1590 150 1910
rect 470 1590 510 1910
rect 110 1550 510 1590
rect 1232 1910 1632 1950
rect 1232 1590 1272 1910
rect 1592 1590 1632 1910
rect 1232 1550 1632 1590
rect 2354 1910 2754 1950
rect 2354 1590 2394 1910
rect 2714 1590 2754 1910
rect 2354 1550 2754 1590
rect 3476 1910 3876 1950
rect 3476 1590 3516 1910
rect 3836 1590 3876 1910
rect 3476 1550 3876 1590
rect 4598 1910 4998 1950
rect 4598 1590 4638 1910
rect 4958 1590 4998 1910
rect 4598 1550 4998 1590
rect -5500 1210 -5100 1250
rect -5500 890 -5460 1210
rect -5140 890 -5100 1210
rect -5500 850 -5100 890
rect -4378 1210 -3978 1250
rect -4378 890 -4338 1210
rect -4018 890 -3978 1210
rect -4378 850 -3978 890
rect -3256 1210 -2856 1250
rect -3256 890 -3216 1210
rect -2896 890 -2856 1210
rect -3256 850 -2856 890
rect -2134 1210 -1734 1250
rect -2134 890 -2094 1210
rect -1774 890 -1734 1210
rect -2134 850 -1734 890
rect -1012 1210 -612 1250
rect -1012 890 -972 1210
rect -652 890 -612 1210
rect -1012 850 -612 890
rect 110 1210 510 1250
rect 110 890 150 1210
rect 470 890 510 1210
rect 110 850 510 890
rect 1232 1210 1632 1250
rect 1232 890 1272 1210
rect 1592 890 1632 1210
rect 1232 850 1632 890
rect 2354 1210 2754 1250
rect 2354 890 2394 1210
rect 2714 890 2754 1210
rect 2354 850 2754 890
rect 3476 1210 3876 1250
rect 3476 890 3516 1210
rect 3836 890 3876 1210
rect 3476 850 3876 890
rect 4598 1210 4998 1250
rect 4598 890 4638 1210
rect 4958 890 4998 1210
rect 4598 850 4998 890
rect -5500 510 -5100 550
rect -5500 190 -5460 510
rect -5140 190 -5100 510
rect -5500 150 -5100 190
rect -4378 510 -3978 550
rect -4378 190 -4338 510
rect -4018 190 -3978 510
rect -4378 150 -3978 190
rect -3256 510 -2856 550
rect -3256 190 -3216 510
rect -2896 190 -2856 510
rect -3256 150 -2856 190
rect -2134 510 -1734 550
rect -2134 190 -2094 510
rect -1774 190 -1734 510
rect -2134 150 -1734 190
rect -1012 510 -612 550
rect -1012 190 -972 510
rect -652 190 -612 510
rect -1012 150 -612 190
rect 110 510 510 550
rect 110 190 150 510
rect 470 190 510 510
rect 110 150 510 190
rect 1232 510 1632 550
rect 1232 190 1272 510
rect 1592 190 1632 510
rect 1232 150 1632 190
rect 2354 510 2754 550
rect 2354 190 2394 510
rect 2714 190 2754 510
rect 2354 150 2754 190
rect 3476 510 3876 550
rect 3476 190 3516 510
rect 3836 190 3876 510
rect 3476 150 3876 190
rect 4598 510 4998 550
rect 4598 190 4638 510
rect 4958 190 4998 510
rect 4598 150 4998 190
rect -5500 -190 -5100 -150
rect -5500 -510 -5460 -190
rect -5140 -510 -5100 -190
rect -5500 -550 -5100 -510
rect -4378 -190 -3978 -150
rect -4378 -510 -4338 -190
rect -4018 -510 -3978 -190
rect -4378 -550 -3978 -510
rect -3256 -190 -2856 -150
rect -3256 -510 -3216 -190
rect -2896 -510 -2856 -190
rect -3256 -550 -2856 -510
rect -2134 -190 -1734 -150
rect -2134 -510 -2094 -190
rect -1774 -510 -1734 -190
rect -2134 -550 -1734 -510
rect -1012 -190 -612 -150
rect -1012 -510 -972 -190
rect -652 -510 -612 -190
rect -1012 -550 -612 -510
rect 110 -190 510 -150
rect 110 -510 150 -190
rect 470 -510 510 -190
rect 110 -550 510 -510
rect 1232 -190 1632 -150
rect 1232 -510 1272 -190
rect 1592 -510 1632 -190
rect 1232 -550 1632 -510
rect 2354 -190 2754 -150
rect 2354 -510 2394 -190
rect 2714 -510 2754 -190
rect 2354 -550 2754 -510
rect 3476 -190 3876 -150
rect 3476 -510 3516 -190
rect 3836 -510 3876 -190
rect 3476 -550 3876 -510
rect 4598 -190 4998 -150
rect 4598 -510 4638 -190
rect 4958 -510 4998 -190
rect 4598 -550 4998 -510
rect -5500 -890 -5100 -850
rect -5500 -1210 -5460 -890
rect -5140 -1210 -5100 -890
rect -5500 -1250 -5100 -1210
rect -4378 -890 -3978 -850
rect -4378 -1210 -4338 -890
rect -4018 -1210 -3978 -890
rect -4378 -1250 -3978 -1210
rect -3256 -890 -2856 -850
rect -3256 -1210 -3216 -890
rect -2896 -1210 -2856 -890
rect -3256 -1250 -2856 -1210
rect -2134 -890 -1734 -850
rect -2134 -1210 -2094 -890
rect -1774 -1210 -1734 -890
rect -2134 -1250 -1734 -1210
rect -1012 -890 -612 -850
rect -1012 -1210 -972 -890
rect -652 -1210 -612 -890
rect -1012 -1250 -612 -1210
rect 110 -890 510 -850
rect 110 -1210 150 -890
rect 470 -1210 510 -890
rect 110 -1250 510 -1210
rect 1232 -890 1632 -850
rect 1232 -1210 1272 -890
rect 1592 -1210 1632 -890
rect 1232 -1250 1632 -1210
rect 2354 -890 2754 -850
rect 2354 -1210 2394 -890
rect 2714 -1210 2754 -890
rect 2354 -1250 2754 -1210
rect 3476 -890 3876 -850
rect 3476 -1210 3516 -890
rect 3836 -1210 3876 -890
rect 3476 -1250 3876 -1210
rect 4598 -890 4998 -850
rect 4598 -1210 4638 -890
rect 4958 -1210 4998 -890
rect 4598 -1250 4998 -1210
rect -5500 -1590 -5100 -1550
rect -5500 -1910 -5460 -1590
rect -5140 -1910 -5100 -1590
rect -5500 -1950 -5100 -1910
rect -4378 -1590 -3978 -1550
rect -4378 -1910 -4338 -1590
rect -4018 -1910 -3978 -1590
rect -4378 -1950 -3978 -1910
rect -3256 -1590 -2856 -1550
rect -3256 -1910 -3216 -1590
rect -2896 -1910 -2856 -1590
rect -3256 -1950 -2856 -1910
rect -2134 -1590 -1734 -1550
rect -2134 -1910 -2094 -1590
rect -1774 -1910 -1734 -1590
rect -2134 -1950 -1734 -1910
rect -1012 -1590 -612 -1550
rect -1012 -1910 -972 -1590
rect -652 -1910 -612 -1590
rect -1012 -1950 -612 -1910
rect 110 -1590 510 -1550
rect 110 -1910 150 -1590
rect 470 -1910 510 -1590
rect 110 -1950 510 -1910
rect 1232 -1590 1632 -1550
rect 1232 -1910 1272 -1590
rect 1592 -1910 1632 -1590
rect 1232 -1950 1632 -1910
rect 2354 -1590 2754 -1550
rect 2354 -1910 2394 -1590
rect 2714 -1910 2754 -1590
rect 2354 -1950 2754 -1910
rect 3476 -1590 3876 -1550
rect 3476 -1910 3516 -1590
rect 3836 -1910 3876 -1590
rect 3476 -1950 3876 -1910
rect 4598 -1590 4998 -1550
rect 4598 -1910 4638 -1590
rect 4958 -1910 4998 -1590
rect 4598 -1950 4998 -1910
rect -5500 -2290 -5100 -2250
rect -5500 -2610 -5460 -2290
rect -5140 -2610 -5100 -2290
rect -5500 -2650 -5100 -2610
rect -4378 -2290 -3978 -2250
rect -4378 -2610 -4338 -2290
rect -4018 -2610 -3978 -2290
rect -4378 -2650 -3978 -2610
rect -3256 -2290 -2856 -2250
rect -3256 -2610 -3216 -2290
rect -2896 -2610 -2856 -2290
rect -3256 -2650 -2856 -2610
rect -2134 -2290 -1734 -2250
rect -2134 -2610 -2094 -2290
rect -1774 -2610 -1734 -2290
rect -2134 -2650 -1734 -2610
rect -1012 -2290 -612 -2250
rect -1012 -2610 -972 -2290
rect -652 -2610 -612 -2290
rect -1012 -2650 -612 -2610
rect 110 -2290 510 -2250
rect 110 -2610 150 -2290
rect 470 -2610 510 -2290
rect 110 -2650 510 -2610
rect 1232 -2290 1632 -2250
rect 1232 -2610 1272 -2290
rect 1592 -2610 1632 -2290
rect 1232 -2650 1632 -2610
rect 2354 -2290 2754 -2250
rect 2354 -2610 2394 -2290
rect 2714 -2610 2754 -2290
rect 2354 -2650 2754 -2610
rect 3476 -2290 3876 -2250
rect 3476 -2610 3516 -2290
rect 3836 -2610 3876 -2290
rect 3476 -2650 3876 -2610
rect 4598 -2290 4998 -2250
rect 4598 -2610 4638 -2290
rect 4958 -2610 4998 -2290
rect 4598 -2650 4998 -2610
rect -5500 -2990 -5100 -2950
rect -5500 -3310 -5460 -2990
rect -5140 -3310 -5100 -2990
rect -5500 -3350 -5100 -3310
rect -4378 -2990 -3978 -2950
rect -4378 -3310 -4338 -2990
rect -4018 -3310 -3978 -2990
rect -4378 -3350 -3978 -3310
rect -3256 -2990 -2856 -2950
rect -3256 -3310 -3216 -2990
rect -2896 -3310 -2856 -2990
rect -3256 -3350 -2856 -3310
rect -2134 -2990 -1734 -2950
rect -2134 -3310 -2094 -2990
rect -1774 -3310 -1734 -2990
rect -2134 -3350 -1734 -3310
rect -1012 -2990 -612 -2950
rect -1012 -3310 -972 -2990
rect -652 -3310 -612 -2990
rect -1012 -3350 -612 -3310
rect 110 -2990 510 -2950
rect 110 -3310 150 -2990
rect 470 -3310 510 -2990
rect 110 -3350 510 -3310
rect 1232 -2990 1632 -2950
rect 1232 -3310 1272 -2990
rect 1592 -3310 1632 -2990
rect 1232 -3350 1632 -3310
rect 2354 -2990 2754 -2950
rect 2354 -3310 2394 -2990
rect 2714 -3310 2754 -2990
rect 2354 -3350 2754 -3310
rect 3476 -2990 3876 -2950
rect 3476 -3310 3516 -2990
rect 3836 -3310 3876 -2990
rect 3476 -3350 3876 -3310
rect 4598 -2990 4998 -2950
rect 4598 -3310 4638 -2990
rect 4958 -3310 4998 -2990
rect 4598 -3350 4998 -3310
<< mimcap2contact >>
rect -5460 2990 -5140 3310
rect -4338 2990 -4018 3310
rect -3216 2990 -2896 3310
rect -2094 2990 -1774 3310
rect -972 2990 -652 3310
rect 150 2990 470 3310
rect 1272 2990 1592 3310
rect 2394 2990 2714 3310
rect 3516 2990 3836 3310
rect 4638 2990 4958 3310
rect -5460 2290 -5140 2610
rect -4338 2290 -4018 2610
rect -3216 2290 -2896 2610
rect -2094 2290 -1774 2610
rect -972 2290 -652 2610
rect 150 2290 470 2610
rect 1272 2290 1592 2610
rect 2394 2290 2714 2610
rect 3516 2290 3836 2610
rect 4638 2290 4958 2610
rect -5460 1590 -5140 1910
rect -4338 1590 -4018 1910
rect -3216 1590 -2896 1910
rect -2094 1590 -1774 1910
rect -972 1590 -652 1910
rect 150 1590 470 1910
rect 1272 1590 1592 1910
rect 2394 1590 2714 1910
rect 3516 1590 3836 1910
rect 4638 1590 4958 1910
rect -5460 890 -5140 1210
rect -4338 890 -4018 1210
rect -3216 890 -2896 1210
rect -2094 890 -1774 1210
rect -972 890 -652 1210
rect 150 890 470 1210
rect 1272 890 1592 1210
rect 2394 890 2714 1210
rect 3516 890 3836 1210
rect 4638 890 4958 1210
rect -5460 190 -5140 510
rect -4338 190 -4018 510
rect -3216 190 -2896 510
rect -2094 190 -1774 510
rect -972 190 -652 510
rect 150 190 470 510
rect 1272 190 1592 510
rect 2394 190 2714 510
rect 3516 190 3836 510
rect 4638 190 4958 510
rect -5460 -510 -5140 -190
rect -4338 -510 -4018 -190
rect -3216 -510 -2896 -190
rect -2094 -510 -1774 -190
rect -972 -510 -652 -190
rect 150 -510 470 -190
rect 1272 -510 1592 -190
rect 2394 -510 2714 -190
rect 3516 -510 3836 -190
rect 4638 -510 4958 -190
rect -5460 -1210 -5140 -890
rect -4338 -1210 -4018 -890
rect -3216 -1210 -2896 -890
rect -2094 -1210 -1774 -890
rect -972 -1210 -652 -890
rect 150 -1210 470 -890
rect 1272 -1210 1592 -890
rect 2394 -1210 2714 -890
rect 3516 -1210 3836 -890
rect 4638 -1210 4958 -890
rect -5460 -1910 -5140 -1590
rect -4338 -1910 -4018 -1590
rect -3216 -1910 -2896 -1590
rect -2094 -1910 -1774 -1590
rect -972 -1910 -652 -1590
rect 150 -1910 470 -1590
rect 1272 -1910 1592 -1590
rect 2394 -1910 2714 -1590
rect 3516 -1910 3836 -1590
rect 4638 -1910 4958 -1590
rect -5460 -2610 -5140 -2290
rect -4338 -2610 -4018 -2290
rect -3216 -2610 -2896 -2290
rect -2094 -2610 -1774 -2290
rect -972 -2610 -652 -2290
rect 150 -2610 470 -2290
rect 1272 -2610 1592 -2290
rect 2394 -2610 2714 -2290
rect 3516 -2610 3836 -2290
rect 4638 -2610 4958 -2290
rect -5460 -3310 -5140 -2990
rect -4338 -3310 -4018 -2990
rect -3216 -3310 -2896 -2990
rect -2094 -3310 -1774 -2990
rect -972 -3310 -652 -2990
rect 150 -3310 470 -2990
rect 1272 -3310 1592 -2990
rect 2394 -3310 2714 -2990
rect 3516 -3310 3836 -2990
rect 4638 -3310 4958 -2990
<< metal5 >>
rect -5460 3334 -5140 3500
rect -4338 3334 -4018 3500
rect -3216 3334 -2896 3500
rect -2094 3334 -1774 3500
rect -972 3334 -652 3500
rect 150 3334 470 3500
rect 1272 3334 1592 3500
rect 2394 3334 2714 3500
rect 3516 3334 3836 3500
rect 4638 3334 4958 3500
rect -5484 3310 -5116 3334
rect -5484 2990 -5460 3310
rect -5140 2990 -5116 3310
rect -5484 2966 -5116 2990
rect -4796 3289 -4476 3331
rect -4796 3011 -4754 3289
rect -4518 3011 -4476 3289
rect -4796 2969 -4476 3011
rect -4362 3310 -3994 3334
rect -4362 2990 -4338 3310
rect -4018 2990 -3994 3310
rect -4362 2966 -3994 2990
rect -3674 3289 -3354 3331
rect -3674 3011 -3632 3289
rect -3396 3011 -3354 3289
rect -3674 2969 -3354 3011
rect -3240 3310 -2872 3334
rect -3240 2990 -3216 3310
rect -2896 2990 -2872 3310
rect -3240 2966 -2872 2990
rect -2552 3289 -2232 3331
rect -2552 3011 -2510 3289
rect -2274 3011 -2232 3289
rect -2552 2969 -2232 3011
rect -2118 3310 -1750 3334
rect -2118 2990 -2094 3310
rect -1774 2990 -1750 3310
rect -2118 2966 -1750 2990
rect -1430 3289 -1110 3331
rect -1430 3011 -1388 3289
rect -1152 3011 -1110 3289
rect -1430 2969 -1110 3011
rect -996 3310 -628 3334
rect -996 2990 -972 3310
rect -652 2990 -628 3310
rect -996 2966 -628 2990
rect -308 3289 12 3331
rect -308 3011 -266 3289
rect -30 3011 12 3289
rect -308 2969 12 3011
rect 126 3310 494 3334
rect 126 2990 150 3310
rect 470 2990 494 3310
rect 126 2966 494 2990
rect 814 3289 1134 3331
rect 814 3011 856 3289
rect 1092 3011 1134 3289
rect 814 2969 1134 3011
rect 1248 3310 1616 3334
rect 1248 2990 1272 3310
rect 1592 2990 1616 3310
rect 1248 2966 1616 2990
rect 1936 3289 2256 3331
rect 1936 3011 1978 3289
rect 2214 3011 2256 3289
rect 1936 2969 2256 3011
rect 2370 3310 2738 3334
rect 2370 2990 2394 3310
rect 2714 2990 2738 3310
rect 2370 2966 2738 2990
rect 3058 3289 3378 3331
rect 3058 3011 3100 3289
rect 3336 3011 3378 3289
rect 3058 2969 3378 3011
rect 3492 3310 3860 3334
rect 3492 2990 3516 3310
rect 3836 2990 3860 3310
rect 3492 2966 3860 2990
rect 4180 3289 4500 3331
rect 4180 3011 4222 3289
rect 4458 3011 4500 3289
rect 4180 2969 4500 3011
rect 4614 3310 4982 3334
rect 4614 2990 4638 3310
rect 4958 2990 4982 3310
rect 4614 2966 4982 2990
rect 5302 3289 5622 3331
rect 5302 3011 5344 3289
rect 5580 3011 5622 3289
rect 5302 2969 5622 3011
rect -5460 2634 -5140 2966
rect -4338 2634 -4018 2966
rect -3216 2634 -2896 2966
rect -2094 2634 -1774 2966
rect -972 2634 -652 2966
rect 150 2634 470 2966
rect 1272 2634 1592 2966
rect 2394 2634 2714 2966
rect 3516 2634 3836 2966
rect 4638 2634 4958 2966
rect -5484 2610 -5116 2634
rect -5484 2290 -5460 2610
rect -5140 2290 -5116 2610
rect -5484 2266 -5116 2290
rect -4796 2589 -4476 2631
rect -4796 2311 -4754 2589
rect -4518 2311 -4476 2589
rect -4796 2269 -4476 2311
rect -4362 2610 -3994 2634
rect -4362 2290 -4338 2610
rect -4018 2290 -3994 2610
rect -4362 2266 -3994 2290
rect -3674 2589 -3354 2631
rect -3674 2311 -3632 2589
rect -3396 2311 -3354 2589
rect -3674 2269 -3354 2311
rect -3240 2610 -2872 2634
rect -3240 2290 -3216 2610
rect -2896 2290 -2872 2610
rect -3240 2266 -2872 2290
rect -2552 2589 -2232 2631
rect -2552 2311 -2510 2589
rect -2274 2311 -2232 2589
rect -2552 2269 -2232 2311
rect -2118 2610 -1750 2634
rect -2118 2290 -2094 2610
rect -1774 2290 -1750 2610
rect -2118 2266 -1750 2290
rect -1430 2589 -1110 2631
rect -1430 2311 -1388 2589
rect -1152 2311 -1110 2589
rect -1430 2269 -1110 2311
rect -996 2610 -628 2634
rect -996 2290 -972 2610
rect -652 2290 -628 2610
rect -996 2266 -628 2290
rect -308 2589 12 2631
rect -308 2311 -266 2589
rect -30 2311 12 2589
rect -308 2269 12 2311
rect 126 2610 494 2634
rect 126 2290 150 2610
rect 470 2290 494 2610
rect 126 2266 494 2290
rect 814 2589 1134 2631
rect 814 2311 856 2589
rect 1092 2311 1134 2589
rect 814 2269 1134 2311
rect 1248 2610 1616 2634
rect 1248 2290 1272 2610
rect 1592 2290 1616 2610
rect 1248 2266 1616 2290
rect 1936 2589 2256 2631
rect 1936 2311 1978 2589
rect 2214 2311 2256 2589
rect 1936 2269 2256 2311
rect 2370 2610 2738 2634
rect 2370 2290 2394 2610
rect 2714 2290 2738 2610
rect 2370 2266 2738 2290
rect 3058 2589 3378 2631
rect 3058 2311 3100 2589
rect 3336 2311 3378 2589
rect 3058 2269 3378 2311
rect 3492 2610 3860 2634
rect 3492 2290 3516 2610
rect 3836 2290 3860 2610
rect 3492 2266 3860 2290
rect 4180 2589 4500 2631
rect 4180 2311 4222 2589
rect 4458 2311 4500 2589
rect 4180 2269 4500 2311
rect 4614 2610 4982 2634
rect 4614 2290 4638 2610
rect 4958 2290 4982 2610
rect 4614 2266 4982 2290
rect 5302 2589 5622 2631
rect 5302 2311 5344 2589
rect 5580 2311 5622 2589
rect 5302 2269 5622 2311
rect -5460 1934 -5140 2266
rect -4338 1934 -4018 2266
rect -3216 1934 -2896 2266
rect -2094 1934 -1774 2266
rect -972 1934 -652 2266
rect 150 1934 470 2266
rect 1272 1934 1592 2266
rect 2394 1934 2714 2266
rect 3516 1934 3836 2266
rect 4638 1934 4958 2266
rect -5484 1910 -5116 1934
rect -5484 1590 -5460 1910
rect -5140 1590 -5116 1910
rect -5484 1566 -5116 1590
rect -4796 1889 -4476 1931
rect -4796 1611 -4754 1889
rect -4518 1611 -4476 1889
rect -4796 1569 -4476 1611
rect -4362 1910 -3994 1934
rect -4362 1590 -4338 1910
rect -4018 1590 -3994 1910
rect -4362 1566 -3994 1590
rect -3674 1889 -3354 1931
rect -3674 1611 -3632 1889
rect -3396 1611 -3354 1889
rect -3674 1569 -3354 1611
rect -3240 1910 -2872 1934
rect -3240 1590 -3216 1910
rect -2896 1590 -2872 1910
rect -3240 1566 -2872 1590
rect -2552 1889 -2232 1931
rect -2552 1611 -2510 1889
rect -2274 1611 -2232 1889
rect -2552 1569 -2232 1611
rect -2118 1910 -1750 1934
rect -2118 1590 -2094 1910
rect -1774 1590 -1750 1910
rect -2118 1566 -1750 1590
rect -1430 1889 -1110 1931
rect -1430 1611 -1388 1889
rect -1152 1611 -1110 1889
rect -1430 1569 -1110 1611
rect -996 1910 -628 1934
rect -996 1590 -972 1910
rect -652 1590 -628 1910
rect -996 1566 -628 1590
rect -308 1889 12 1931
rect -308 1611 -266 1889
rect -30 1611 12 1889
rect -308 1569 12 1611
rect 126 1910 494 1934
rect 126 1590 150 1910
rect 470 1590 494 1910
rect 126 1566 494 1590
rect 814 1889 1134 1931
rect 814 1611 856 1889
rect 1092 1611 1134 1889
rect 814 1569 1134 1611
rect 1248 1910 1616 1934
rect 1248 1590 1272 1910
rect 1592 1590 1616 1910
rect 1248 1566 1616 1590
rect 1936 1889 2256 1931
rect 1936 1611 1978 1889
rect 2214 1611 2256 1889
rect 1936 1569 2256 1611
rect 2370 1910 2738 1934
rect 2370 1590 2394 1910
rect 2714 1590 2738 1910
rect 2370 1566 2738 1590
rect 3058 1889 3378 1931
rect 3058 1611 3100 1889
rect 3336 1611 3378 1889
rect 3058 1569 3378 1611
rect 3492 1910 3860 1934
rect 3492 1590 3516 1910
rect 3836 1590 3860 1910
rect 3492 1566 3860 1590
rect 4180 1889 4500 1931
rect 4180 1611 4222 1889
rect 4458 1611 4500 1889
rect 4180 1569 4500 1611
rect 4614 1910 4982 1934
rect 4614 1590 4638 1910
rect 4958 1590 4982 1910
rect 4614 1566 4982 1590
rect 5302 1889 5622 1931
rect 5302 1611 5344 1889
rect 5580 1611 5622 1889
rect 5302 1569 5622 1611
rect -5460 1234 -5140 1566
rect -4338 1234 -4018 1566
rect -3216 1234 -2896 1566
rect -2094 1234 -1774 1566
rect -972 1234 -652 1566
rect 150 1234 470 1566
rect 1272 1234 1592 1566
rect 2394 1234 2714 1566
rect 3516 1234 3836 1566
rect 4638 1234 4958 1566
rect -5484 1210 -5116 1234
rect -5484 890 -5460 1210
rect -5140 890 -5116 1210
rect -5484 866 -5116 890
rect -4796 1189 -4476 1231
rect -4796 911 -4754 1189
rect -4518 911 -4476 1189
rect -4796 869 -4476 911
rect -4362 1210 -3994 1234
rect -4362 890 -4338 1210
rect -4018 890 -3994 1210
rect -4362 866 -3994 890
rect -3674 1189 -3354 1231
rect -3674 911 -3632 1189
rect -3396 911 -3354 1189
rect -3674 869 -3354 911
rect -3240 1210 -2872 1234
rect -3240 890 -3216 1210
rect -2896 890 -2872 1210
rect -3240 866 -2872 890
rect -2552 1189 -2232 1231
rect -2552 911 -2510 1189
rect -2274 911 -2232 1189
rect -2552 869 -2232 911
rect -2118 1210 -1750 1234
rect -2118 890 -2094 1210
rect -1774 890 -1750 1210
rect -2118 866 -1750 890
rect -1430 1189 -1110 1231
rect -1430 911 -1388 1189
rect -1152 911 -1110 1189
rect -1430 869 -1110 911
rect -996 1210 -628 1234
rect -996 890 -972 1210
rect -652 890 -628 1210
rect -996 866 -628 890
rect -308 1189 12 1231
rect -308 911 -266 1189
rect -30 911 12 1189
rect -308 869 12 911
rect 126 1210 494 1234
rect 126 890 150 1210
rect 470 890 494 1210
rect 126 866 494 890
rect 814 1189 1134 1231
rect 814 911 856 1189
rect 1092 911 1134 1189
rect 814 869 1134 911
rect 1248 1210 1616 1234
rect 1248 890 1272 1210
rect 1592 890 1616 1210
rect 1248 866 1616 890
rect 1936 1189 2256 1231
rect 1936 911 1978 1189
rect 2214 911 2256 1189
rect 1936 869 2256 911
rect 2370 1210 2738 1234
rect 2370 890 2394 1210
rect 2714 890 2738 1210
rect 2370 866 2738 890
rect 3058 1189 3378 1231
rect 3058 911 3100 1189
rect 3336 911 3378 1189
rect 3058 869 3378 911
rect 3492 1210 3860 1234
rect 3492 890 3516 1210
rect 3836 890 3860 1210
rect 3492 866 3860 890
rect 4180 1189 4500 1231
rect 4180 911 4222 1189
rect 4458 911 4500 1189
rect 4180 869 4500 911
rect 4614 1210 4982 1234
rect 4614 890 4638 1210
rect 4958 890 4982 1210
rect 4614 866 4982 890
rect 5302 1189 5622 1231
rect 5302 911 5344 1189
rect 5580 911 5622 1189
rect 5302 869 5622 911
rect -5460 534 -5140 866
rect -4338 534 -4018 866
rect -3216 534 -2896 866
rect -2094 534 -1774 866
rect -972 534 -652 866
rect 150 534 470 866
rect 1272 534 1592 866
rect 2394 534 2714 866
rect 3516 534 3836 866
rect 4638 534 4958 866
rect -5484 510 -5116 534
rect -5484 190 -5460 510
rect -5140 190 -5116 510
rect -5484 166 -5116 190
rect -4796 489 -4476 531
rect -4796 211 -4754 489
rect -4518 211 -4476 489
rect -4796 169 -4476 211
rect -4362 510 -3994 534
rect -4362 190 -4338 510
rect -4018 190 -3994 510
rect -4362 166 -3994 190
rect -3674 489 -3354 531
rect -3674 211 -3632 489
rect -3396 211 -3354 489
rect -3674 169 -3354 211
rect -3240 510 -2872 534
rect -3240 190 -3216 510
rect -2896 190 -2872 510
rect -3240 166 -2872 190
rect -2552 489 -2232 531
rect -2552 211 -2510 489
rect -2274 211 -2232 489
rect -2552 169 -2232 211
rect -2118 510 -1750 534
rect -2118 190 -2094 510
rect -1774 190 -1750 510
rect -2118 166 -1750 190
rect -1430 489 -1110 531
rect -1430 211 -1388 489
rect -1152 211 -1110 489
rect -1430 169 -1110 211
rect -996 510 -628 534
rect -996 190 -972 510
rect -652 190 -628 510
rect -996 166 -628 190
rect -308 489 12 531
rect -308 211 -266 489
rect -30 211 12 489
rect -308 169 12 211
rect 126 510 494 534
rect 126 190 150 510
rect 470 190 494 510
rect 126 166 494 190
rect 814 489 1134 531
rect 814 211 856 489
rect 1092 211 1134 489
rect 814 169 1134 211
rect 1248 510 1616 534
rect 1248 190 1272 510
rect 1592 190 1616 510
rect 1248 166 1616 190
rect 1936 489 2256 531
rect 1936 211 1978 489
rect 2214 211 2256 489
rect 1936 169 2256 211
rect 2370 510 2738 534
rect 2370 190 2394 510
rect 2714 190 2738 510
rect 2370 166 2738 190
rect 3058 489 3378 531
rect 3058 211 3100 489
rect 3336 211 3378 489
rect 3058 169 3378 211
rect 3492 510 3860 534
rect 3492 190 3516 510
rect 3836 190 3860 510
rect 3492 166 3860 190
rect 4180 489 4500 531
rect 4180 211 4222 489
rect 4458 211 4500 489
rect 4180 169 4500 211
rect 4614 510 4982 534
rect 4614 190 4638 510
rect 4958 190 4982 510
rect 4614 166 4982 190
rect 5302 489 5622 531
rect 5302 211 5344 489
rect 5580 211 5622 489
rect 5302 169 5622 211
rect -5460 -166 -5140 166
rect -4338 -166 -4018 166
rect -3216 -166 -2896 166
rect -2094 -166 -1774 166
rect -972 -166 -652 166
rect 150 -166 470 166
rect 1272 -166 1592 166
rect 2394 -166 2714 166
rect 3516 -166 3836 166
rect 4638 -166 4958 166
rect -5484 -190 -5116 -166
rect -5484 -510 -5460 -190
rect -5140 -510 -5116 -190
rect -5484 -534 -5116 -510
rect -4796 -211 -4476 -169
rect -4796 -489 -4754 -211
rect -4518 -489 -4476 -211
rect -4796 -531 -4476 -489
rect -4362 -190 -3994 -166
rect -4362 -510 -4338 -190
rect -4018 -510 -3994 -190
rect -4362 -534 -3994 -510
rect -3674 -211 -3354 -169
rect -3674 -489 -3632 -211
rect -3396 -489 -3354 -211
rect -3674 -531 -3354 -489
rect -3240 -190 -2872 -166
rect -3240 -510 -3216 -190
rect -2896 -510 -2872 -190
rect -3240 -534 -2872 -510
rect -2552 -211 -2232 -169
rect -2552 -489 -2510 -211
rect -2274 -489 -2232 -211
rect -2552 -531 -2232 -489
rect -2118 -190 -1750 -166
rect -2118 -510 -2094 -190
rect -1774 -510 -1750 -190
rect -2118 -534 -1750 -510
rect -1430 -211 -1110 -169
rect -1430 -489 -1388 -211
rect -1152 -489 -1110 -211
rect -1430 -531 -1110 -489
rect -996 -190 -628 -166
rect -996 -510 -972 -190
rect -652 -510 -628 -190
rect -996 -534 -628 -510
rect -308 -211 12 -169
rect -308 -489 -266 -211
rect -30 -489 12 -211
rect -308 -531 12 -489
rect 126 -190 494 -166
rect 126 -510 150 -190
rect 470 -510 494 -190
rect 126 -534 494 -510
rect 814 -211 1134 -169
rect 814 -489 856 -211
rect 1092 -489 1134 -211
rect 814 -531 1134 -489
rect 1248 -190 1616 -166
rect 1248 -510 1272 -190
rect 1592 -510 1616 -190
rect 1248 -534 1616 -510
rect 1936 -211 2256 -169
rect 1936 -489 1978 -211
rect 2214 -489 2256 -211
rect 1936 -531 2256 -489
rect 2370 -190 2738 -166
rect 2370 -510 2394 -190
rect 2714 -510 2738 -190
rect 2370 -534 2738 -510
rect 3058 -211 3378 -169
rect 3058 -489 3100 -211
rect 3336 -489 3378 -211
rect 3058 -531 3378 -489
rect 3492 -190 3860 -166
rect 3492 -510 3516 -190
rect 3836 -510 3860 -190
rect 3492 -534 3860 -510
rect 4180 -211 4500 -169
rect 4180 -489 4222 -211
rect 4458 -489 4500 -211
rect 4180 -531 4500 -489
rect 4614 -190 4982 -166
rect 4614 -510 4638 -190
rect 4958 -510 4982 -190
rect 4614 -534 4982 -510
rect 5302 -211 5622 -169
rect 5302 -489 5344 -211
rect 5580 -489 5622 -211
rect 5302 -531 5622 -489
rect -5460 -866 -5140 -534
rect -4338 -866 -4018 -534
rect -3216 -866 -2896 -534
rect -2094 -866 -1774 -534
rect -972 -866 -652 -534
rect 150 -866 470 -534
rect 1272 -866 1592 -534
rect 2394 -866 2714 -534
rect 3516 -866 3836 -534
rect 4638 -866 4958 -534
rect -5484 -890 -5116 -866
rect -5484 -1210 -5460 -890
rect -5140 -1210 -5116 -890
rect -5484 -1234 -5116 -1210
rect -4796 -911 -4476 -869
rect -4796 -1189 -4754 -911
rect -4518 -1189 -4476 -911
rect -4796 -1231 -4476 -1189
rect -4362 -890 -3994 -866
rect -4362 -1210 -4338 -890
rect -4018 -1210 -3994 -890
rect -4362 -1234 -3994 -1210
rect -3674 -911 -3354 -869
rect -3674 -1189 -3632 -911
rect -3396 -1189 -3354 -911
rect -3674 -1231 -3354 -1189
rect -3240 -890 -2872 -866
rect -3240 -1210 -3216 -890
rect -2896 -1210 -2872 -890
rect -3240 -1234 -2872 -1210
rect -2552 -911 -2232 -869
rect -2552 -1189 -2510 -911
rect -2274 -1189 -2232 -911
rect -2552 -1231 -2232 -1189
rect -2118 -890 -1750 -866
rect -2118 -1210 -2094 -890
rect -1774 -1210 -1750 -890
rect -2118 -1234 -1750 -1210
rect -1430 -911 -1110 -869
rect -1430 -1189 -1388 -911
rect -1152 -1189 -1110 -911
rect -1430 -1231 -1110 -1189
rect -996 -890 -628 -866
rect -996 -1210 -972 -890
rect -652 -1210 -628 -890
rect -996 -1234 -628 -1210
rect -308 -911 12 -869
rect -308 -1189 -266 -911
rect -30 -1189 12 -911
rect -308 -1231 12 -1189
rect 126 -890 494 -866
rect 126 -1210 150 -890
rect 470 -1210 494 -890
rect 126 -1234 494 -1210
rect 814 -911 1134 -869
rect 814 -1189 856 -911
rect 1092 -1189 1134 -911
rect 814 -1231 1134 -1189
rect 1248 -890 1616 -866
rect 1248 -1210 1272 -890
rect 1592 -1210 1616 -890
rect 1248 -1234 1616 -1210
rect 1936 -911 2256 -869
rect 1936 -1189 1978 -911
rect 2214 -1189 2256 -911
rect 1936 -1231 2256 -1189
rect 2370 -890 2738 -866
rect 2370 -1210 2394 -890
rect 2714 -1210 2738 -890
rect 2370 -1234 2738 -1210
rect 3058 -911 3378 -869
rect 3058 -1189 3100 -911
rect 3336 -1189 3378 -911
rect 3058 -1231 3378 -1189
rect 3492 -890 3860 -866
rect 3492 -1210 3516 -890
rect 3836 -1210 3860 -890
rect 3492 -1234 3860 -1210
rect 4180 -911 4500 -869
rect 4180 -1189 4222 -911
rect 4458 -1189 4500 -911
rect 4180 -1231 4500 -1189
rect 4614 -890 4982 -866
rect 4614 -1210 4638 -890
rect 4958 -1210 4982 -890
rect 4614 -1234 4982 -1210
rect 5302 -911 5622 -869
rect 5302 -1189 5344 -911
rect 5580 -1189 5622 -911
rect 5302 -1231 5622 -1189
rect -5460 -1566 -5140 -1234
rect -4338 -1566 -4018 -1234
rect -3216 -1566 -2896 -1234
rect -2094 -1566 -1774 -1234
rect -972 -1566 -652 -1234
rect 150 -1566 470 -1234
rect 1272 -1566 1592 -1234
rect 2394 -1566 2714 -1234
rect 3516 -1566 3836 -1234
rect 4638 -1566 4958 -1234
rect -5484 -1590 -5116 -1566
rect -5484 -1910 -5460 -1590
rect -5140 -1910 -5116 -1590
rect -5484 -1934 -5116 -1910
rect -4796 -1611 -4476 -1569
rect -4796 -1889 -4754 -1611
rect -4518 -1889 -4476 -1611
rect -4796 -1931 -4476 -1889
rect -4362 -1590 -3994 -1566
rect -4362 -1910 -4338 -1590
rect -4018 -1910 -3994 -1590
rect -4362 -1934 -3994 -1910
rect -3674 -1611 -3354 -1569
rect -3674 -1889 -3632 -1611
rect -3396 -1889 -3354 -1611
rect -3674 -1931 -3354 -1889
rect -3240 -1590 -2872 -1566
rect -3240 -1910 -3216 -1590
rect -2896 -1910 -2872 -1590
rect -3240 -1934 -2872 -1910
rect -2552 -1611 -2232 -1569
rect -2552 -1889 -2510 -1611
rect -2274 -1889 -2232 -1611
rect -2552 -1931 -2232 -1889
rect -2118 -1590 -1750 -1566
rect -2118 -1910 -2094 -1590
rect -1774 -1910 -1750 -1590
rect -2118 -1934 -1750 -1910
rect -1430 -1611 -1110 -1569
rect -1430 -1889 -1388 -1611
rect -1152 -1889 -1110 -1611
rect -1430 -1931 -1110 -1889
rect -996 -1590 -628 -1566
rect -996 -1910 -972 -1590
rect -652 -1910 -628 -1590
rect -996 -1934 -628 -1910
rect -308 -1611 12 -1569
rect -308 -1889 -266 -1611
rect -30 -1889 12 -1611
rect -308 -1931 12 -1889
rect 126 -1590 494 -1566
rect 126 -1910 150 -1590
rect 470 -1910 494 -1590
rect 126 -1934 494 -1910
rect 814 -1611 1134 -1569
rect 814 -1889 856 -1611
rect 1092 -1889 1134 -1611
rect 814 -1931 1134 -1889
rect 1248 -1590 1616 -1566
rect 1248 -1910 1272 -1590
rect 1592 -1910 1616 -1590
rect 1248 -1934 1616 -1910
rect 1936 -1611 2256 -1569
rect 1936 -1889 1978 -1611
rect 2214 -1889 2256 -1611
rect 1936 -1931 2256 -1889
rect 2370 -1590 2738 -1566
rect 2370 -1910 2394 -1590
rect 2714 -1910 2738 -1590
rect 2370 -1934 2738 -1910
rect 3058 -1611 3378 -1569
rect 3058 -1889 3100 -1611
rect 3336 -1889 3378 -1611
rect 3058 -1931 3378 -1889
rect 3492 -1590 3860 -1566
rect 3492 -1910 3516 -1590
rect 3836 -1910 3860 -1590
rect 3492 -1934 3860 -1910
rect 4180 -1611 4500 -1569
rect 4180 -1889 4222 -1611
rect 4458 -1889 4500 -1611
rect 4180 -1931 4500 -1889
rect 4614 -1590 4982 -1566
rect 4614 -1910 4638 -1590
rect 4958 -1910 4982 -1590
rect 4614 -1934 4982 -1910
rect 5302 -1611 5622 -1569
rect 5302 -1889 5344 -1611
rect 5580 -1889 5622 -1611
rect 5302 -1931 5622 -1889
rect -5460 -2266 -5140 -1934
rect -4338 -2266 -4018 -1934
rect -3216 -2266 -2896 -1934
rect -2094 -2266 -1774 -1934
rect -972 -2266 -652 -1934
rect 150 -2266 470 -1934
rect 1272 -2266 1592 -1934
rect 2394 -2266 2714 -1934
rect 3516 -2266 3836 -1934
rect 4638 -2266 4958 -1934
rect -5484 -2290 -5116 -2266
rect -5484 -2610 -5460 -2290
rect -5140 -2610 -5116 -2290
rect -5484 -2634 -5116 -2610
rect -4796 -2311 -4476 -2269
rect -4796 -2589 -4754 -2311
rect -4518 -2589 -4476 -2311
rect -4796 -2631 -4476 -2589
rect -4362 -2290 -3994 -2266
rect -4362 -2610 -4338 -2290
rect -4018 -2610 -3994 -2290
rect -4362 -2634 -3994 -2610
rect -3674 -2311 -3354 -2269
rect -3674 -2589 -3632 -2311
rect -3396 -2589 -3354 -2311
rect -3674 -2631 -3354 -2589
rect -3240 -2290 -2872 -2266
rect -3240 -2610 -3216 -2290
rect -2896 -2610 -2872 -2290
rect -3240 -2634 -2872 -2610
rect -2552 -2311 -2232 -2269
rect -2552 -2589 -2510 -2311
rect -2274 -2589 -2232 -2311
rect -2552 -2631 -2232 -2589
rect -2118 -2290 -1750 -2266
rect -2118 -2610 -2094 -2290
rect -1774 -2610 -1750 -2290
rect -2118 -2634 -1750 -2610
rect -1430 -2311 -1110 -2269
rect -1430 -2589 -1388 -2311
rect -1152 -2589 -1110 -2311
rect -1430 -2631 -1110 -2589
rect -996 -2290 -628 -2266
rect -996 -2610 -972 -2290
rect -652 -2610 -628 -2290
rect -996 -2634 -628 -2610
rect -308 -2311 12 -2269
rect -308 -2589 -266 -2311
rect -30 -2589 12 -2311
rect -308 -2631 12 -2589
rect 126 -2290 494 -2266
rect 126 -2610 150 -2290
rect 470 -2610 494 -2290
rect 126 -2634 494 -2610
rect 814 -2311 1134 -2269
rect 814 -2589 856 -2311
rect 1092 -2589 1134 -2311
rect 814 -2631 1134 -2589
rect 1248 -2290 1616 -2266
rect 1248 -2610 1272 -2290
rect 1592 -2610 1616 -2290
rect 1248 -2634 1616 -2610
rect 1936 -2311 2256 -2269
rect 1936 -2589 1978 -2311
rect 2214 -2589 2256 -2311
rect 1936 -2631 2256 -2589
rect 2370 -2290 2738 -2266
rect 2370 -2610 2394 -2290
rect 2714 -2610 2738 -2290
rect 2370 -2634 2738 -2610
rect 3058 -2311 3378 -2269
rect 3058 -2589 3100 -2311
rect 3336 -2589 3378 -2311
rect 3058 -2631 3378 -2589
rect 3492 -2290 3860 -2266
rect 3492 -2610 3516 -2290
rect 3836 -2610 3860 -2290
rect 3492 -2634 3860 -2610
rect 4180 -2311 4500 -2269
rect 4180 -2589 4222 -2311
rect 4458 -2589 4500 -2311
rect 4180 -2631 4500 -2589
rect 4614 -2290 4982 -2266
rect 4614 -2610 4638 -2290
rect 4958 -2610 4982 -2290
rect 4614 -2634 4982 -2610
rect 5302 -2311 5622 -2269
rect 5302 -2589 5344 -2311
rect 5580 -2589 5622 -2311
rect 5302 -2631 5622 -2589
rect -5460 -2966 -5140 -2634
rect -4338 -2966 -4018 -2634
rect -3216 -2966 -2896 -2634
rect -2094 -2966 -1774 -2634
rect -972 -2966 -652 -2634
rect 150 -2966 470 -2634
rect 1272 -2966 1592 -2634
rect 2394 -2966 2714 -2634
rect 3516 -2966 3836 -2634
rect 4638 -2966 4958 -2634
rect -5484 -2990 -5116 -2966
rect -5484 -3310 -5460 -2990
rect -5140 -3310 -5116 -2990
rect -5484 -3334 -5116 -3310
rect -4796 -3011 -4476 -2969
rect -4796 -3289 -4754 -3011
rect -4518 -3289 -4476 -3011
rect -4796 -3331 -4476 -3289
rect -4362 -2990 -3994 -2966
rect -4362 -3310 -4338 -2990
rect -4018 -3310 -3994 -2990
rect -4362 -3334 -3994 -3310
rect -3674 -3011 -3354 -2969
rect -3674 -3289 -3632 -3011
rect -3396 -3289 -3354 -3011
rect -3674 -3331 -3354 -3289
rect -3240 -2990 -2872 -2966
rect -3240 -3310 -3216 -2990
rect -2896 -3310 -2872 -2990
rect -3240 -3334 -2872 -3310
rect -2552 -3011 -2232 -2969
rect -2552 -3289 -2510 -3011
rect -2274 -3289 -2232 -3011
rect -2552 -3331 -2232 -3289
rect -2118 -2990 -1750 -2966
rect -2118 -3310 -2094 -2990
rect -1774 -3310 -1750 -2990
rect -2118 -3334 -1750 -3310
rect -1430 -3011 -1110 -2969
rect -1430 -3289 -1388 -3011
rect -1152 -3289 -1110 -3011
rect -1430 -3331 -1110 -3289
rect -996 -2990 -628 -2966
rect -996 -3310 -972 -2990
rect -652 -3310 -628 -2990
rect -996 -3334 -628 -3310
rect -308 -3011 12 -2969
rect -308 -3289 -266 -3011
rect -30 -3289 12 -3011
rect -308 -3331 12 -3289
rect 126 -2990 494 -2966
rect 126 -3310 150 -2990
rect 470 -3310 494 -2990
rect 126 -3334 494 -3310
rect 814 -3011 1134 -2969
rect 814 -3289 856 -3011
rect 1092 -3289 1134 -3011
rect 814 -3331 1134 -3289
rect 1248 -2990 1616 -2966
rect 1248 -3310 1272 -2990
rect 1592 -3310 1616 -2990
rect 1248 -3334 1616 -3310
rect 1936 -3011 2256 -2969
rect 1936 -3289 1978 -3011
rect 2214 -3289 2256 -3011
rect 1936 -3331 2256 -3289
rect 2370 -2990 2738 -2966
rect 2370 -3310 2394 -2990
rect 2714 -3310 2738 -2990
rect 2370 -3334 2738 -3310
rect 3058 -3011 3378 -2969
rect 3058 -3289 3100 -3011
rect 3336 -3289 3378 -3011
rect 3058 -3331 3378 -3289
rect 3492 -2990 3860 -2966
rect 3492 -3310 3516 -2990
rect 3836 -3310 3860 -2990
rect 3492 -3334 3860 -3310
rect 4180 -3011 4500 -2969
rect 4180 -3289 4222 -3011
rect 4458 -3289 4500 -3011
rect 4180 -3331 4500 -3289
rect 4614 -2990 4982 -2966
rect 4614 -3310 4638 -2990
rect 4958 -3310 4982 -2990
rect 4614 -3334 4982 -3310
rect 5302 -3011 5622 -2969
rect 5302 -3289 5344 -3011
rect 5580 -3289 5622 -3011
rect 5302 -3331 5622 -3289
rect -5460 -3500 -5140 -3334
rect -4338 -3500 -4018 -3334
rect -3216 -3500 -2896 -3334
rect -2094 -3500 -1774 -3334
rect -972 -3500 -652 -3334
rect 150 -3500 470 -3334
rect 1272 -3500 1592 -3334
rect 2394 -3500 2714 -3334
rect 3516 -3500 3836 -3334
rect 4638 -3500 4958 -3334
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX 4498 2850 5098 3450
string parameters w 2.00 l 2.00 val 5.36 carea 1.00 cperi 0.17 nx 10 ny 10 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 1 ccov 100
string library sky130
<< end >>
