magic
tech sky130A
magscale 1 2
timestamp 1620885654
<< xpolycontact >>
rect -35 304 35 736
rect -35 -736 35 -304
<< xpolyres >>
rect -35 -304 35 304
<< viali >>
rect -19 321 19 718
rect -19 -718 19 -321
<< metal1 >>
rect -25 718 25 730
rect -25 321 -19 718
rect 19 321 25 718
rect -25 309 25 321
rect -25 -321 25 -309
rect -25 -718 -19 -321
rect 19 -718 25 -321
rect -25 -730 25 -718
<< res0p35 >>
rect -37 -306 37 306
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 3.042 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 17.492k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
