magic
tech sky130A
magscale 1 2
timestamp 1621270775
<< error_p >>
rect -2584 -3968 2584 3934
<< nwell >>
rect -2584 -3968 2584 3934
<< pmoslvt >>
rect -2490 -3906 -2090 3834
rect -2032 -3906 -1632 3834
rect -1574 -3906 -1174 3834
rect -1116 -3906 -716 3834
rect -658 -3906 -258 3834
rect -200 -3906 200 3834
rect 258 -3906 658 3834
rect 716 -3906 1116 3834
rect 1174 -3906 1574 3834
rect 1632 -3906 2032 3834
rect 2090 -3906 2490 3834
<< pdiff >>
rect -2548 3822 -2490 3834
rect -2548 -3894 -2536 3822
rect -2502 -3894 -2490 3822
rect -2548 -3906 -2490 -3894
rect -2090 3822 -2032 3834
rect -2090 -3894 -2078 3822
rect -2044 -3894 -2032 3822
rect -2090 -3906 -2032 -3894
rect -1632 3822 -1574 3834
rect -1632 -3894 -1620 3822
rect -1586 -3894 -1574 3822
rect -1632 -3906 -1574 -3894
rect -1174 3822 -1116 3834
rect -1174 -3894 -1162 3822
rect -1128 -3894 -1116 3822
rect -1174 -3906 -1116 -3894
rect -716 3822 -658 3834
rect -716 -3894 -704 3822
rect -670 -3894 -658 3822
rect -716 -3906 -658 -3894
rect -258 3822 -200 3834
rect -258 -3894 -246 3822
rect -212 -3894 -200 3822
rect -258 -3906 -200 -3894
rect 200 3822 258 3834
rect 200 -3894 212 3822
rect 246 -3894 258 3822
rect 200 -3906 258 -3894
rect 658 3822 716 3834
rect 658 -3894 670 3822
rect 704 -3894 716 3822
rect 658 -3906 716 -3894
rect 1116 3822 1174 3834
rect 1116 -3894 1128 3822
rect 1162 -3894 1174 3822
rect 1116 -3906 1174 -3894
rect 1574 3822 1632 3834
rect 1574 -3894 1586 3822
rect 1620 -3894 1632 3822
rect 1574 -3906 1632 -3894
rect 2032 3822 2090 3834
rect 2032 -3894 2044 3822
rect 2078 -3894 2090 3822
rect 2032 -3906 2090 -3894
rect 2490 3822 2548 3834
rect 2490 -3894 2502 3822
rect 2536 -3894 2548 3822
rect 2490 -3906 2548 -3894
<< pdiffc >>
rect -2536 -3894 -2502 3822
rect -2078 -3894 -2044 3822
rect -1620 -3894 -1586 3822
rect -1162 -3894 -1128 3822
rect -704 -3894 -670 3822
rect -246 -3894 -212 3822
rect 212 -3894 246 3822
rect 670 -3894 704 3822
rect 1128 -3894 1162 3822
rect 1586 -3894 1620 3822
rect 2044 -3894 2078 3822
rect 2502 -3894 2536 3822
<< poly >>
rect -2490 3915 -2090 3931
rect -2490 3881 -2474 3915
rect -2106 3881 -2090 3915
rect -2490 3834 -2090 3881
rect -2032 3915 -1632 3931
rect -2032 3881 -2016 3915
rect -1648 3881 -1632 3915
rect -2032 3834 -1632 3881
rect -1574 3915 -1174 3931
rect -1574 3881 -1558 3915
rect -1190 3881 -1174 3915
rect -1574 3834 -1174 3881
rect -1116 3915 -716 3931
rect -1116 3881 -1100 3915
rect -732 3881 -716 3915
rect -1116 3834 -716 3881
rect -658 3915 -258 3931
rect -658 3881 -642 3915
rect -274 3881 -258 3915
rect -658 3834 -258 3881
rect -200 3915 200 3931
rect -200 3881 -184 3915
rect 184 3881 200 3915
rect -200 3834 200 3881
rect 258 3915 658 3931
rect 258 3881 274 3915
rect 642 3881 658 3915
rect 258 3834 658 3881
rect 716 3915 1116 3931
rect 716 3881 732 3915
rect 1100 3881 1116 3915
rect 716 3834 1116 3881
rect 1174 3915 1574 3931
rect 1174 3881 1190 3915
rect 1558 3881 1574 3915
rect 1174 3834 1574 3881
rect 1632 3915 2032 3931
rect 1632 3881 1648 3915
rect 2016 3881 2032 3915
rect 1632 3834 2032 3881
rect 2090 3915 2490 3931
rect 2090 3881 2106 3915
rect 2474 3881 2490 3915
rect 2090 3834 2490 3881
rect -2490 -3932 -2090 -3906
rect -2032 -3932 -1632 -3906
rect -1574 -3932 -1174 -3906
rect -1116 -3932 -716 -3906
rect -658 -3932 -258 -3906
rect -200 -3932 200 -3906
rect 258 -3932 658 -3906
rect 716 -3932 1116 -3906
rect 1174 -3932 1574 -3906
rect 1632 -3932 2032 -3906
rect 2090 -3932 2490 -3906
<< polycont >>
rect -2474 3881 -2106 3915
rect -2016 3881 -1648 3915
rect -1558 3881 -1190 3915
rect -1100 3881 -732 3915
rect -642 3881 -274 3915
rect -184 3881 184 3915
rect 274 3881 642 3915
rect 732 3881 1100 3915
rect 1190 3881 1558 3915
rect 1648 3881 2016 3915
rect 2106 3881 2474 3915
<< locali >>
rect -2490 3881 -2474 3915
rect -2106 3881 -2090 3915
rect -2032 3881 -2016 3915
rect -1648 3881 -1632 3915
rect -1574 3881 -1558 3915
rect -1190 3881 -1174 3915
rect -1116 3881 -1100 3915
rect -732 3881 -716 3915
rect -658 3881 -642 3915
rect -274 3881 -258 3915
rect -200 3881 -184 3915
rect 184 3881 200 3915
rect 258 3881 274 3915
rect 642 3881 658 3915
rect 716 3881 732 3915
rect 1100 3881 1116 3915
rect 1174 3881 1190 3915
rect 1558 3881 1574 3915
rect 1632 3881 1648 3915
rect 2016 3881 2032 3915
rect 2090 3881 2106 3915
rect 2474 3881 2490 3915
rect -2536 3822 -2502 3838
rect -2536 -3910 -2502 -3894
rect -2078 3822 -2044 3838
rect -2078 -3910 -2044 -3894
rect -1620 3822 -1586 3838
rect -1620 -3910 -1586 -3894
rect -1162 3822 -1128 3838
rect -1162 -3910 -1128 -3894
rect -704 3822 -670 3838
rect -704 -3910 -670 -3894
rect -246 3822 -212 3838
rect -246 -3910 -212 -3894
rect 212 3822 246 3838
rect 212 -3910 246 -3894
rect 670 3822 704 3838
rect 670 -3910 704 -3894
rect 1128 3822 1162 3838
rect 1128 -3910 1162 -3894
rect 1586 3822 1620 3838
rect 1586 -3910 1620 -3894
rect 2044 3822 2078 3838
rect 2044 -3910 2078 -3894
rect 2502 3822 2536 3838
rect 2502 -3910 2536 -3894
<< viali >>
rect -2382 3881 -2198 3915
rect -1924 3881 -1740 3915
rect -1466 3881 -1282 3915
rect -1008 3881 -824 3915
rect -550 3881 -366 3915
rect -92 3881 92 3915
rect 366 3881 550 3915
rect 824 3881 1008 3915
rect 1282 3881 1466 3915
rect 1740 3881 1924 3915
rect 2198 3881 2382 3915
rect -2536 -3894 -2502 3822
rect -2078 -3894 -2044 3822
rect -1620 -3894 -1586 3822
rect -1162 -3894 -1128 3822
rect -704 -3894 -670 3822
rect -246 -3894 -212 3822
rect 212 -3894 246 3822
rect 670 -3894 704 3822
rect 1128 -3894 1162 3822
rect 1586 -3894 1620 3822
rect 2044 -3894 2078 3822
rect 2502 -3894 2536 3822
<< metal1 >>
rect -2394 3915 -2186 3921
rect -2394 3881 -2382 3915
rect -2198 3881 -2186 3915
rect -2394 3875 -2186 3881
rect -1936 3915 -1728 3921
rect -1936 3881 -1924 3915
rect -1740 3881 -1728 3915
rect -1936 3875 -1728 3881
rect -1478 3915 -1270 3921
rect -1478 3881 -1466 3915
rect -1282 3881 -1270 3915
rect -1478 3875 -1270 3881
rect -1020 3915 -812 3921
rect -1020 3881 -1008 3915
rect -824 3881 -812 3915
rect -1020 3875 -812 3881
rect -562 3915 -354 3921
rect -562 3881 -550 3915
rect -366 3881 -354 3915
rect -562 3875 -354 3881
rect -104 3915 104 3921
rect -104 3881 -92 3915
rect 92 3881 104 3915
rect -104 3875 104 3881
rect 354 3915 562 3921
rect 354 3881 366 3915
rect 550 3881 562 3915
rect 354 3875 562 3881
rect 812 3915 1020 3921
rect 812 3881 824 3915
rect 1008 3881 1020 3915
rect 812 3875 1020 3881
rect 1270 3915 1478 3921
rect 1270 3881 1282 3915
rect 1466 3881 1478 3915
rect 1270 3875 1478 3881
rect 1728 3915 1936 3921
rect 1728 3881 1740 3915
rect 1924 3881 1936 3915
rect 1728 3875 1936 3881
rect 2186 3915 2394 3921
rect 2186 3881 2198 3915
rect 2382 3881 2394 3915
rect 2186 3875 2394 3881
rect -2542 3822 -2496 3834
rect -2542 -3894 -2536 3822
rect -2502 -3894 -2496 3822
rect -2542 -3906 -2496 -3894
rect -2084 3822 -2038 3834
rect -2084 -3894 -2078 3822
rect -2044 -3894 -2038 3822
rect -2084 -3906 -2038 -3894
rect -1626 3822 -1580 3834
rect -1626 -3894 -1620 3822
rect -1586 -3894 -1580 3822
rect -1626 -3906 -1580 -3894
rect -1168 3822 -1122 3834
rect -1168 -3894 -1162 3822
rect -1128 -3894 -1122 3822
rect -1168 -3906 -1122 -3894
rect -710 3822 -664 3834
rect -710 -3894 -704 3822
rect -670 -3894 -664 3822
rect -710 -3906 -664 -3894
rect -252 3822 -206 3834
rect -252 -3894 -246 3822
rect -212 -3894 -206 3822
rect -252 -3906 -206 -3894
rect 206 3822 252 3834
rect 206 -3894 212 3822
rect 246 -3894 252 3822
rect 206 -3906 252 -3894
rect 664 3822 710 3834
rect 664 -3894 670 3822
rect 704 -3894 710 3822
rect 664 -3906 710 -3894
rect 1122 3822 1168 3834
rect 1122 -3894 1128 3822
rect 1162 -3894 1168 3822
rect 1122 -3906 1168 -3894
rect 1580 3822 1626 3834
rect 1580 -3894 1586 3822
rect 1620 -3894 1626 3822
rect 1580 -3906 1626 -3894
rect 2038 3822 2084 3834
rect 2038 -3894 2044 3822
rect 2078 -3894 2084 3822
rect 2038 -3906 2084 -3894
rect 2496 3822 2542 3834
rect 2496 -3894 2502 3822
rect 2536 -3894 2542 3822
rect 2496 -3906 2542 -3894
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 38.7 l 2 m 1 nf 11 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
