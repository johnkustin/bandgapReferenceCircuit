magic
tech sky130A
magscale 1 2
timestamp 1621317379
<< nwell >>
rect -9600 9500 7778 9502
rect -19400 1000 -9872 4342
rect -9600 1602 8666 9500
rect -9600 1600 -3680 1602
rect -2890 1600 1820 1602
rect 2610 1600 8666 1602
<< pmoslvt >>
rect -18562 1662 -18162 4242
rect -17990 1662 -17590 4242
rect -17418 1662 -17018 4242
rect -16846 1662 -16446 4242
rect -16274 1662 -15874 4242
rect -15702 1662 -15302 4242
rect -15130 1662 -14730 4242
rect -14558 1662 -14158 4242
rect -13986 1662 -13586 4242
rect -13414 1662 -13014 4242
rect -12842 1662 -12442 4242
rect -12270 1662 -11870 4242
rect -11698 1662 -11298 4242
rect -11126 1662 -10726 4242
rect -8754 1700 -8354 9440
rect -8296 1700 -7896 9440
rect -7838 1700 -7438 9440
rect -7380 1700 -6980 9440
rect -6922 1700 -6522 9440
rect -6464 1700 -6064 9440
rect -6006 1700 -5606 9440
rect -5548 1700 -5148 9440
rect -5090 1700 -4690 9440
rect -4632 1700 -4232 9440
rect -4174 1700 -3774 9440
rect -2796 1700 -2396 9440
rect -2338 1700 -1938 9440
rect -1880 1700 -1480 9440
rect -1422 1700 -1022 9440
rect -964 1700 -564 9440
rect -506 1700 -106 9440
rect -48 1700 352 9440
rect 410 1700 810 9440
rect 868 1700 1268 9440
rect 1326 1700 1726 9440
rect 2704 1700 3104 9440
rect 3162 1700 3562 9440
rect 3620 1700 4020 9440
rect 4078 1700 4478 9440
rect 4536 1700 4936 9440
rect 4994 1700 5394 9440
rect 5452 1700 5852 9440
rect 5910 1700 6310 9440
rect 6368 1700 6768 9440
rect 6826 1700 7226 9440
rect 7284 1700 7684 9440
<< nmoslvt >>
rect -17176 8406 -11776 8806
rect -21766 5132 -21366 5532
rect -21308 5132 -20908 5532
rect -20850 5132 -20450 5532
rect -20392 5132 -19992 5532
rect -19934 5132 -19534 5532
rect -19476 5132 -19076 5532
rect -16836 4854 -16436 6654
rect -16264 4854 -15864 6654
rect -15692 4854 -15292 6654
rect -15120 4854 -14720 6654
rect -14548 4854 -14148 6654
rect -13976 4854 -13576 6654
rect -13404 4854 -13004 6654
rect -12832 4854 -12432 6654
<< ndiff >>
rect -17176 8852 -11776 8864
rect -17176 8818 -17164 8852
rect -11788 8818 -11776 8852
rect -17176 8806 -11776 8818
rect -17176 8394 -11776 8406
rect -17176 8360 -17164 8394
rect -11788 8360 -11776 8394
rect -17176 8348 -11776 8360
rect -21824 5520 -21766 5532
rect -21824 5144 -21812 5520
rect -21778 5144 -21766 5520
rect -21824 5132 -21766 5144
rect -21366 5520 -21308 5532
rect -21366 5144 -21354 5520
rect -21320 5144 -21308 5520
rect -21366 5132 -21308 5144
rect -20908 5520 -20850 5532
rect -20908 5144 -20896 5520
rect -20862 5144 -20850 5520
rect -20908 5132 -20850 5144
rect -20450 5520 -20392 5532
rect -20450 5144 -20438 5520
rect -20404 5144 -20392 5520
rect -20450 5132 -20392 5144
rect -19992 5520 -19934 5532
rect -19992 5144 -19980 5520
rect -19946 5144 -19934 5520
rect -19992 5132 -19934 5144
rect -19534 5520 -19476 5532
rect -19534 5144 -19522 5520
rect -19488 5144 -19476 5520
rect -19534 5132 -19476 5144
rect -19076 5520 -19018 5532
rect -19076 5144 -19064 5520
rect -19030 5144 -19018 5520
rect -19076 5132 -19018 5144
rect -16894 6642 -16836 6654
rect -16894 4866 -16882 6642
rect -16848 4866 -16836 6642
rect -16894 4854 -16836 4866
rect -16436 6642 -16378 6654
rect -16436 4866 -16424 6642
rect -16390 4866 -16378 6642
rect -16436 4854 -16378 4866
rect -16322 6642 -16264 6654
rect -16322 4866 -16310 6642
rect -16276 4866 -16264 6642
rect -16322 4854 -16264 4866
rect -15864 6642 -15806 6654
rect -15864 4866 -15852 6642
rect -15818 4866 -15806 6642
rect -15864 4854 -15806 4866
rect -15750 6642 -15692 6654
rect -15750 4866 -15738 6642
rect -15704 4866 -15692 6642
rect -15750 4854 -15692 4866
rect -15292 6642 -15234 6654
rect -15292 4866 -15280 6642
rect -15246 4866 -15234 6642
rect -15292 4854 -15234 4866
rect -15178 6642 -15120 6654
rect -15178 4866 -15166 6642
rect -15132 4866 -15120 6642
rect -15178 4854 -15120 4866
rect -14720 6642 -14662 6654
rect -14720 4866 -14708 6642
rect -14674 4866 -14662 6642
rect -14720 4854 -14662 4866
rect -14606 6642 -14548 6654
rect -14606 4866 -14594 6642
rect -14560 4866 -14548 6642
rect -14606 4854 -14548 4866
rect -14148 6642 -14090 6654
rect -14148 4866 -14136 6642
rect -14102 4866 -14090 6642
rect -14148 4854 -14090 4866
rect -14034 6642 -13976 6654
rect -14034 4866 -14022 6642
rect -13988 4866 -13976 6642
rect -14034 4854 -13976 4866
rect -13576 6642 -13518 6654
rect -13576 4866 -13564 6642
rect -13530 4866 -13518 6642
rect -13576 4854 -13518 4866
rect -13462 6642 -13404 6654
rect -13462 4866 -13450 6642
rect -13416 4866 -13404 6642
rect -13462 4854 -13404 4866
rect -13004 6642 -12946 6654
rect -13004 4866 -12992 6642
rect -12958 4866 -12946 6642
rect -13004 4854 -12946 4866
rect -12890 6642 -12832 6654
rect -12890 4866 -12878 6642
rect -12844 4866 -12832 6642
rect -12890 4854 -12832 4866
rect -12432 6642 -12374 6654
rect -12432 4866 -12420 6642
rect -12386 4866 -12374 6642
rect -12432 4854 -12374 4866
<< pdiff >>
rect -8812 9428 -8754 9440
rect -18620 4230 -18562 4242
rect -18620 1674 -18608 4230
rect -18574 1674 -18562 4230
rect -18620 1662 -18562 1674
rect -18162 4230 -18104 4242
rect -18162 1674 -18150 4230
rect -18116 1674 -18104 4230
rect -18162 1662 -18104 1674
rect -18048 4230 -17990 4242
rect -18048 1674 -18036 4230
rect -18002 1674 -17990 4230
rect -18048 1662 -17990 1674
rect -17590 4230 -17532 4242
rect -17590 1674 -17578 4230
rect -17544 1674 -17532 4230
rect -17590 1662 -17532 1674
rect -17476 4230 -17418 4242
rect -17476 1674 -17464 4230
rect -17430 1674 -17418 4230
rect -17476 1662 -17418 1674
rect -17018 4230 -16960 4242
rect -17018 1674 -17006 4230
rect -16972 1674 -16960 4230
rect -17018 1662 -16960 1674
rect -16904 4230 -16846 4242
rect -16904 1674 -16892 4230
rect -16858 1674 -16846 4230
rect -16904 1662 -16846 1674
rect -16446 4230 -16388 4242
rect -16446 1674 -16434 4230
rect -16400 1674 -16388 4230
rect -16446 1662 -16388 1674
rect -16332 4230 -16274 4242
rect -16332 1674 -16320 4230
rect -16286 1674 -16274 4230
rect -16332 1662 -16274 1674
rect -15874 4230 -15816 4242
rect -15874 1674 -15862 4230
rect -15828 1674 -15816 4230
rect -15874 1662 -15816 1674
rect -15760 4230 -15702 4242
rect -15760 1674 -15748 4230
rect -15714 1674 -15702 4230
rect -15760 1662 -15702 1674
rect -15302 4230 -15244 4242
rect -15302 1674 -15290 4230
rect -15256 1674 -15244 4230
rect -15302 1662 -15244 1674
rect -15188 4230 -15130 4242
rect -15188 1674 -15176 4230
rect -15142 1674 -15130 4230
rect -15188 1662 -15130 1674
rect -14730 4230 -14672 4242
rect -14730 1674 -14718 4230
rect -14684 1674 -14672 4230
rect -14730 1662 -14672 1674
rect -14616 4230 -14558 4242
rect -14616 1674 -14604 4230
rect -14570 1674 -14558 4230
rect -14616 1662 -14558 1674
rect -14158 4230 -14100 4242
rect -14158 1674 -14146 4230
rect -14112 1674 -14100 4230
rect -14158 1662 -14100 1674
rect -14044 4230 -13986 4242
rect -14044 1674 -14032 4230
rect -13998 1674 -13986 4230
rect -14044 1662 -13986 1674
rect -13586 4230 -13528 4242
rect -13586 1674 -13574 4230
rect -13540 1674 -13528 4230
rect -13586 1662 -13528 1674
rect -13472 4230 -13414 4242
rect -13472 1674 -13460 4230
rect -13426 1674 -13414 4230
rect -13472 1662 -13414 1674
rect -13014 4230 -12956 4242
rect -13014 1674 -13002 4230
rect -12968 1674 -12956 4230
rect -13014 1662 -12956 1674
rect -12900 4230 -12842 4242
rect -12900 1674 -12888 4230
rect -12854 1674 -12842 4230
rect -12900 1662 -12842 1674
rect -12442 4230 -12384 4242
rect -12442 1674 -12430 4230
rect -12396 1674 -12384 4230
rect -12442 1662 -12384 1674
rect -12328 4230 -12270 4242
rect -12328 1674 -12316 4230
rect -12282 1674 -12270 4230
rect -12328 1662 -12270 1674
rect -11870 4230 -11812 4242
rect -11870 1674 -11858 4230
rect -11824 1674 -11812 4230
rect -11870 1662 -11812 1674
rect -11756 4230 -11698 4242
rect -11756 1674 -11744 4230
rect -11710 1674 -11698 4230
rect -11756 1662 -11698 1674
rect -11298 4230 -11240 4242
rect -11298 1674 -11286 4230
rect -11252 1674 -11240 4230
rect -11298 1662 -11240 1674
rect -11184 4230 -11126 4242
rect -11184 1674 -11172 4230
rect -11138 1674 -11126 4230
rect -11184 1662 -11126 1674
rect -10726 4230 -10668 4242
rect -10726 1674 -10714 4230
rect -10680 1674 -10668 4230
rect -8812 1712 -8800 9428
rect -8766 1712 -8754 9428
rect -8812 1700 -8754 1712
rect -8354 9428 -8296 9440
rect -8354 1712 -8342 9428
rect -8308 1712 -8296 9428
rect -8354 1700 -8296 1712
rect -7896 9428 -7838 9440
rect -7896 1712 -7884 9428
rect -7850 1712 -7838 9428
rect -7896 1700 -7838 1712
rect -7438 9428 -7380 9440
rect -7438 1712 -7426 9428
rect -7392 1712 -7380 9428
rect -7438 1700 -7380 1712
rect -6980 9428 -6922 9440
rect -6980 1712 -6968 9428
rect -6934 1712 -6922 9428
rect -6980 1700 -6922 1712
rect -6522 9428 -6464 9440
rect -6522 1712 -6510 9428
rect -6476 1712 -6464 9428
rect -6522 1700 -6464 1712
rect -6064 9428 -6006 9440
rect -6064 1712 -6052 9428
rect -6018 1712 -6006 9428
rect -6064 1700 -6006 1712
rect -5606 9428 -5548 9440
rect -5606 1712 -5594 9428
rect -5560 1712 -5548 9428
rect -5606 1700 -5548 1712
rect -5148 9428 -5090 9440
rect -5148 1712 -5136 9428
rect -5102 1712 -5090 9428
rect -5148 1700 -5090 1712
rect -4690 9428 -4632 9440
rect -4690 1712 -4678 9428
rect -4644 1712 -4632 9428
rect -4690 1700 -4632 1712
rect -4232 9428 -4174 9440
rect -4232 1712 -4220 9428
rect -4186 1712 -4174 9428
rect -4232 1700 -4174 1712
rect -3774 9428 -3716 9440
rect -3774 1712 -3762 9428
rect -3728 1712 -3716 9428
rect -2854 9428 -2796 9440
rect -3774 1700 -3716 1712
rect -2854 1712 -2842 9428
rect -2808 1712 -2796 9428
rect -2854 1700 -2796 1712
rect -2396 9428 -2338 9440
rect -2396 1712 -2384 9428
rect -2350 1712 -2338 9428
rect -2396 1700 -2338 1712
rect -1938 9428 -1880 9440
rect -1938 1712 -1926 9428
rect -1892 1712 -1880 9428
rect -1938 1700 -1880 1712
rect -1480 9428 -1422 9440
rect -1480 1712 -1468 9428
rect -1434 1712 -1422 9428
rect -1480 1700 -1422 1712
rect -1022 9428 -964 9440
rect -1022 1712 -1010 9428
rect -976 1712 -964 9428
rect -1022 1700 -964 1712
rect -564 9428 -506 9440
rect -564 1712 -552 9428
rect -518 1712 -506 9428
rect -564 1700 -506 1712
rect -106 9428 -48 9440
rect -106 1712 -94 9428
rect -60 1712 -48 9428
rect -106 1700 -48 1712
rect 352 9428 410 9440
rect 352 1712 364 9428
rect 398 1712 410 9428
rect 352 1700 410 1712
rect 810 9428 868 9440
rect 810 1712 822 9428
rect 856 1712 868 9428
rect 810 1700 868 1712
rect 1268 9428 1326 9440
rect 1268 1712 1280 9428
rect 1314 1712 1326 9428
rect 1268 1700 1326 1712
rect 1726 9428 1784 9440
rect 1726 1712 1738 9428
rect 1772 1712 1784 9428
rect 2646 9428 2704 9440
rect 1726 1700 1784 1712
rect 2646 1712 2658 9428
rect 2692 1712 2704 9428
rect 2646 1700 2704 1712
rect 3104 9428 3162 9440
rect 3104 1712 3116 9428
rect 3150 1712 3162 9428
rect 3104 1700 3162 1712
rect 3562 9428 3620 9440
rect 3562 1712 3574 9428
rect 3608 1712 3620 9428
rect 3562 1700 3620 1712
rect 4020 9428 4078 9440
rect 4020 1712 4032 9428
rect 4066 1712 4078 9428
rect 4020 1700 4078 1712
rect 4478 9428 4536 9440
rect 4478 1712 4490 9428
rect 4524 1712 4536 9428
rect 4478 1700 4536 1712
rect 4936 9428 4994 9440
rect 4936 1712 4948 9428
rect 4982 1712 4994 9428
rect 4936 1700 4994 1712
rect 5394 9428 5452 9440
rect 5394 1712 5406 9428
rect 5440 1712 5452 9428
rect 5394 1700 5452 1712
rect 5852 9428 5910 9440
rect 5852 1712 5864 9428
rect 5898 1712 5910 9428
rect 5852 1700 5910 1712
rect 6310 9428 6368 9440
rect 6310 1712 6322 9428
rect 6356 1712 6368 9428
rect 6310 1700 6368 1712
rect 6768 9428 6826 9440
rect 6768 1712 6780 9428
rect 6814 1712 6826 9428
rect 6768 1700 6826 1712
rect 7226 9428 7284 9440
rect 7226 1712 7238 9428
rect 7272 1712 7284 9428
rect 7226 1700 7284 1712
rect 7684 9428 7742 9440
rect 7684 1712 7696 9428
rect 7730 1712 7742 9428
rect 7684 1700 7742 1712
rect -10726 1662 -10668 1674
<< ndiffc >>
rect -17164 8818 -11788 8852
rect -17164 8360 -11788 8394
rect -21812 5144 -21778 5520
rect -21354 5144 -21320 5520
rect -20896 5144 -20862 5520
rect -20438 5144 -20404 5520
rect -19980 5144 -19946 5520
rect -19522 5144 -19488 5520
rect -19064 5144 -19030 5520
rect -16882 4866 -16848 6642
rect -16424 4866 -16390 6642
rect -16310 4866 -16276 6642
rect -15852 4866 -15818 6642
rect -15738 4866 -15704 6642
rect -15280 4866 -15246 6642
rect -15166 4866 -15132 6642
rect -14708 4866 -14674 6642
rect -14594 4866 -14560 6642
rect -14136 4866 -14102 6642
rect -14022 4866 -13988 6642
rect -13564 4866 -13530 6642
rect -13450 4866 -13416 6642
rect -12992 4866 -12958 6642
rect -12878 4866 -12844 6642
rect -12420 4866 -12386 6642
<< pdiffc >>
rect -18608 1674 -18574 4230
rect -18150 1674 -18116 4230
rect -18036 1674 -18002 4230
rect -17578 1674 -17544 4230
rect -17464 1674 -17430 4230
rect -17006 1674 -16972 4230
rect -16892 1674 -16858 4230
rect -16434 1674 -16400 4230
rect -16320 1674 -16286 4230
rect -15862 1674 -15828 4230
rect -15748 1674 -15714 4230
rect -15290 1674 -15256 4230
rect -15176 1674 -15142 4230
rect -14718 1674 -14684 4230
rect -14604 1674 -14570 4230
rect -14146 1674 -14112 4230
rect -14032 1674 -13998 4230
rect -13574 1674 -13540 4230
rect -13460 1674 -13426 4230
rect -13002 1674 -12968 4230
rect -12888 1674 -12854 4230
rect -12430 1674 -12396 4230
rect -12316 1674 -12282 4230
rect -11858 1674 -11824 4230
rect -11744 1674 -11710 4230
rect -11286 1674 -11252 4230
rect -11172 1674 -11138 4230
rect -10714 1674 -10680 4230
rect -8800 1712 -8766 9428
rect -8342 1712 -8308 9428
rect -7884 1712 -7850 9428
rect -7426 1712 -7392 9428
rect -6968 1712 -6934 9428
rect -6510 1712 -6476 9428
rect -6052 1712 -6018 9428
rect -5594 1712 -5560 9428
rect -5136 1712 -5102 9428
rect -4678 1712 -4644 9428
rect -4220 1712 -4186 9428
rect -3762 1712 -3728 9428
rect -2842 1712 -2808 9428
rect -2384 1712 -2350 9428
rect -1926 1712 -1892 9428
rect -1468 1712 -1434 9428
rect -1010 1712 -976 9428
rect -552 1712 -518 9428
rect -94 1712 -60 9428
rect 364 1712 398 9428
rect 822 1712 856 9428
rect 1280 1712 1314 9428
rect 1738 1712 1772 9428
rect 2658 1712 2692 9428
rect 3116 1712 3150 9428
rect 3574 1712 3608 9428
rect 4032 1712 4066 9428
rect 4490 1712 4524 9428
rect 4948 1712 4982 9428
rect 5406 1712 5440 9428
rect 5864 1712 5898 9428
rect 6322 1712 6356 9428
rect 6780 1712 6814 9428
rect 7238 1712 7272 9428
rect 7696 1712 7730 9428
<< psubdiff >>
rect -21540 25036 -10308 25060
rect -21540 24270 -21516 25036
rect -10332 24270 -10308 25036
rect -21540 24246 -10308 24270
rect -9780 21500 -9162 21524
rect -9780 15196 -9756 21500
rect -9186 15196 -9162 21500
rect -6536 21500 -5918 21524
rect -9780 15172 -9162 15196
rect -6536 15196 -6512 21500
rect -5942 15196 -5918 21500
rect -1576 21500 -958 21524
rect -6536 15172 -5918 15196
rect -1576 15196 -1552 21500
rect -982 15196 -958 21500
rect -1576 15172 -958 15196
rect 13112 21500 13730 21524
rect 13112 15196 13136 21500
rect 13706 15196 13730 21500
rect 13112 15172 13730 15196
rect -17906 9382 -11406 9406
rect -17906 9050 -17882 9382
rect -11430 9050 -11406 9382
rect -17906 9026 -11406 9050
rect -17484 6642 -17284 6742
rect -22332 5836 -18512 5860
rect -22332 5760 -20918 5836
rect -19926 5760 -18512 5836
rect -22332 5736 -18512 5760
rect -22328 5682 -21880 5736
rect -22328 5106 -22304 5682
rect -21904 5106 -21880 5682
rect -18962 5682 -18514 5736
rect -18962 5106 -18938 5682
rect -18538 5106 -18514 5682
rect -22328 5082 -21880 5106
rect -18962 5082 -18514 5106
rect -17484 5042 -17434 6642
rect -17334 5042 -17284 6642
rect -17484 4942 -17284 5042
rect -11984 6642 -11784 6742
rect -11984 5042 -11934 6642
rect -11834 5042 -11784 6642
rect -11984 4942 -11784 5042
<< nsubdiff >>
rect -9500 9102 -8900 9302
rect -19300 4142 -19100 4242
rect -19300 1800 -19250 4142
rect -19150 1800 -19100 4142
rect -19300 1700 -19100 1800
rect -10172 4142 -9972 4242
rect -10172 1800 -10122 4142
rect -10022 1800 -9972 4142
rect -9500 2102 -9300 9102
rect -9100 2102 -8900 9102
rect -9500 1902 -8900 2102
rect -10172 1700 -9972 1800
rect -3590 9102 -2990 9302
rect -3590 2102 -3390 9102
rect -3190 2102 -2990 9102
rect -3590 1902 -2990 2102
rect 1910 9102 2510 9302
rect 1910 2102 2110 9102
rect 2310 2102 2510 9102
rect 1910 1902 2510 2102
rect 7866 9100 8466 9300
rect 7866 2100 8066 9100
rect 8266 2100 8466 9100
rect 7866 1900 8466 2100
rect -15768 1296 -13226 1346
rect -15768 1196 -15668 1296
rect -13326 1196 -13226 1296
rect -15768 1146 -13226 1196
<< psubdiffcont >>
rect -21516 24270 -10332 25036
rect -9756 15196 -9186 21500
rect -6512 15196 -5942 21500
rect -1552 15196 -982 21500
rect 13136 15196 13706 21500
rect -17882 9050 -11430 9382
rect -20918 5760 -19926 5836
rect -22304 5106 -21904 5682
rect -18938 5106 -18538 5682
rect -17434 5042 -17334 6642
rect -11934 5042 -11834 6642
<< nsubdiffcont >>
rect -19250 1800 -19150 4142
rect -10122 1800 -10022 4142
rect -9300 2102 -9100 9102
rect -3390 2102 -3190 9102
rect 2110 2102 2310 9102
rect 8066 2100 8266 9100
rect -15668 1196 -13326 1296
<< poly >>
rect -8754 9440 -8354 9466
rect -8296 9440 -7896 9466
rect -7838 9440 -7438 9466
rect -7380 9440 -6980 9466
rect -6922 9440 -6522 9466
rect -6464 9440 -6064 9466
rect -6006 9440 -5606 9466
rect -5548 9440 -5148 9466
rect -5090 9440 -4690 9466
rect -4632 9440 -4232 9466
rect -4174 9440 -3774 9466
rect -2796 9440 -2396 9466
rect -2338 9440 -1938 9466
rect -1880 9440 -1480 9466
rect -1422 9440 -1022 9466
rect -964 9440 -564 9466
rect -506 9440 -106 9466
rect -48 9440 352 9466
rect 410 9440 810 9466
rect 868 9440 1268 9466
rect 1326 9440 1726 9466
rect 2704 9440 3104 9466
rect 3162 9440 3562 9466
rect 3620 9440 4020 9466
rect 4078 9440 4478 9466
rect 4536 9440 4936 9466
rect 4994 9440 5394 9466
rect 5452 9440 5852 9466
rect 5910 9440 6310 9466
rect 6368 9440 6768 9466
rect 6826 9440 7226 9466
rect 7284 9440 7684 9466
rect -17264 8790 -17176 8806
rect -17264 8422 -17248 8790
rect -17214 8422 -17176 8790
rect -17264 8406 -17176 8422
rect -11776 8406 -11750 8806
rect -16836 6726 -16436 6742
rect -16836 6692 -16820 6726
rect -16452 6692 -16436 6726
rect -16836 6654 -16436 6692
rect -16264 6726 -15864 6742
rect -16264 6692 -16248 6726
rect -15880 6692 -15864 6726
rect -16264 6654 -15864 6692
rect -15692 6726 -15292 6742
rect -15692 6692 -15676 6726
rect -15308 6692 -15292 6726
rect -15692 6654 -15292 6692
rect -15120 6726 -14720 6742
rect -15120 6692 -15104 6726
rect -14736 6692 -14720 6726
rect -15120 6654 -14720 6692
rect -14548 6726 -14148 6742
rect -14548 6692 -14532 6726
rect -14164 6692 -14148 6726
rect -14548 6654 -14148 6692
rect -13976 6726 -13576 6742
rect -13976 6692 -13960 6726
rect -13592 6692 -13576 6726
rect -13976 6654 -13576 6692
rect -13404 6726 -13004 6742
rect -13404 6692 -13388 6726
rect -13020 6692 -13004 6726
rect -13404 6654 -13004 6692
rect -12832 6726 -12432 6742
rect -12832 6692 -12816 6726
rect -12448 6692 -12432 6726
rect -12832 6654 -12432 6692
rect -21766 5604 -21366 5620
rect -21766 5570 -21750 5604
rect -21382 5570 -21366 5604
rect -21766 5532 -21366 5570
rect -21308 5604 -20908 5620
rect -21308 5570 -21292 5604
rect -20924 5570 -20908 5604
rect -21308 5532 -20908 5570
rect -20850 5604 -20450 5620
rect -20850 5570 -20834 5604
rect -20466 5570 -20450 5604
rect -20850 5532 -20450 5570
rect -20392 5604 -19992 5620
rect -20392 5570 -20376 5604
rect -20008 5570 -19992 5604
rect -20392 5532 -19992 5570
rect -19934 5604 -19534 5620
rect -19934 5570 -19918 5604
rect -19550 5570 -19534 5604
rect -19934 5532 -19534 5570
rect -19476 5604 -19076 5620
rect -19476 5570 -19460 5604
rect -19092 5570 -19076 5604
rect -19476 5532 -19076 5570
rect -21766 5106 -21366 5132
rect -21308 5106 -20908 5132
rect -20850 5106 -20450 5132
rect -20392 5106 -19992 5132
rect -19934 5106 -19534 5132
rect -19476 5106 -19076 5132
rect -16836 4828 -16436 4854
rect -16264 4828 -15864 4854
rect -15692 4828 -15292 4854
rect -15120 4828 -14720 4854
rect -14548 4828 -14148 4854
rect -13976 4828 -13576 4854
rect -13404 4828 -13004 4854
rect -12832 4828 -12432 4854
rect -18562 4323 -18162 4339
rect -18562 4289 -18546 4323
rect -18178 4289 -18162 4323
rect -18562 4242 -18162 4289
rect -17990 4323 -17590 4339
rect -17990 4289 -17974 4323
rect -17606 4289 -17590 4323
rect -17990 4242 -17590 4289
rect -17418 4323 -17018 4339
rect -17418 4289 -17402 4323
rect -17034 4289 -17018 4323
rect -17418 4242 -17018 4289
rect -16846 4323 -16446 4339
rect -16846 4289 -16830 4323
rect -16462 4289 -16446 4323
rect -16846 4242 -16446 4289
rect -16274 4323 -15874 4339
rect -16274 4289 -16258 4323
rect -15890 4289 -15874 4323
rect -16274 4242 -15874 4289
rect -15702 4323 -15302 4339
rect -15702 4289 -15686 4323
rect -15318 4289 -15302 4323
rect -15702 4242 -15302 4289
rect -15130 4323 -14730 4339
rect -15130 4289 -15114 4323
rect -14746 4289 -14730 4323
rect -15130 4242 -14730 4289
rect -14558 4323 -14158 4339
rect -14558 4289 -14542 4323
rect -14174 4289 -14158 4323
rect -14558 4242 -14158 4289
rect -13986 4323 -13586 4339
rect -13986 4289 -13970 4323
rect -13602 4289 -13586 4323
rect -13986 4242 -13586 4289
rect -13414 4323 -13014 4339
rect -13414 4289 -13398 4323
rect -13030 4289 -13014 4323
rect -13414 4242 -13014 4289
rect -12842 4323 -12442 4339
rect -12842 4289 -12826 4323
rect -12458 4289 -12442 4323
rect -12842 4242 -12442 4289
rect -12270 4323 -11870 4339
rect -12270 4289 -12254 4323
rect -11886 4289 -11870 4323
rect -12270 4242 -11870 4289
rect -11698 4323 -11298 4339
rect -11698 4289 -11682 4323
rect -11314 4289 -11298 4323
rect -11698 4242 -11298 4289
rect -11126 4323 -10726 4339
rect -11126 4289 -11110 4323
rect -10742 4289 -10726 4323
rect -11126 4242 -10726 4289
rect -18562 1636 -18162 1662
rect -17990 1636 -17590 1662
rect -17418 1636 -17018 1662
rect -16846 1636 -16446 1662
rect -16274 1636 -15874 1662
rect -15702 1636 -15302 1662
rect -15130 1636 -14730 1662
rect -14558 1636 -14158 1662
rect -13986 1636 -13586 1662
rect -13414 1636 -13014 1662
rect -12842 1636 -12442 1662
rect -12270 1636 -11870 1662
rect -11698 1636 -11298 1662
rect -11126 1636 -10726 1662
rect -8754 1653 -8354 1700
rect -8754 1619 -8738 1653
rect -8370 1619 -8354 1653
rect -8754 1603 -8354 1619
rect -8296 1653 -7896 1700
rect -8296 1619 -8280 1653
rect -7912 1619 -7896 1653
rect -8296 1603 -7896 1619
rect -7838 1653 -7438 1700
rect -7838 1619 -7822 1653
rect -7454 1619 -7438 1653
rect -7838 1603 -7438 1619
rect -7380 1653 -6980 1700
rect -7380 1619 -7364 1653
rect -6996 1619 -6980 1653
rect -7380 1603 -6980 1619
rect -6922 1653 -6522 1700
rect -6922 1619 -6906 1653
rect -6538 1619 -6522 1653
rect -6922 1603 -6522 1619
rect -6464 1653 -6064 1700
rect -6464 1619 -6448 1653
rect -6080 1619 -6064 1653
rect -6464 1603 -6064 1619
rect -6006 1653 -5606 1700
rect -6006 1619 -5990 1653
rect -5622 1619 -5606 1653
rect -6006 1603 -5606 1619
rect -5548 1653 -5148 1700
rect -5548 1619 -5532 1653
rect -5164 1619 -5148 1653
rect -5548 1603 -5148 1619
rect -5090 1653 -4690 1700
rect -5090 1619 -5074 1653
rect -4706 1619 -4690 1653
rect -5090 1603 -4690 1619
rect -4632 1653 -4232 1700
rect -4632 1619 -4616 1653
rect -4248 1619 -4232 1653
rect -4632 1603 -4232 1619
rect -4174 1653 -3774 1700
rect -4174 1619 -4158 1653
rect -3790 1619 -3774 1653
rect -4174 1603 -3774 1619
rect -2796 1653 -2396 1700
rect -2796 1619 -2780 1653
rect -2412 1619 -2396 1653
rect -2796 1603 -2396 1619
rect -2338 1653 -1938 1700
rect -2338 1619 -2322 1653
rect -1954 1619 -1938 1653
rect -2338 1603 -1938 1619
rect -1880 1653 -1480 1700
rect -1880 1619 -1864 1653
rect -1496 1619 -1480 1653
rect -1880 1603 -1480 1619
rect -1422 1653 -1022 1700
rect -1422 1619 -1406 1653
rect -1038 1619 -1022 1653
rect -1422 1603 -1022 1619
rect -964 1653 -564 1700
rect -964 1619 -948 1653
rect -580 1619 -564 1653
rect -964 1603 -564 1619
rect -506 1653 -106 1700
rect -506 1619 -490 1653
rect -122 1619 -106 1653
rect -506 1603 -106 1619
rect -48 1653 352 1700
rect -48 1619 -32 1653
rect 336 1619 352 1653
rect -48 1603 352 1619
rect 410 1653 810 1700
rect 410 1619 426 1653
rect 794 1619 810 1653
rect 410 1603 810 1619
rect 868 1653 1268 1700
rect 868 1619 884 1653
rect 1252 1619 1268 1653
rect 868 1603 1268 1619
rect 1326 1653 1726 1700
rect 1326 1619 1342 1653
rect 1710 1619 1726 1653
rect 1326 1603 1726 1619
rect 2704 1653 3104 1700
rect 2704 1619 2720 1653
rect 3088 1619 3104 1653
rect 2704 1603 3104 1619
rect 3162 1653 3562 1700
rect 3162 1619 3178 1653
rect 3546 1619 3562 1653
rect 3162 1603 3562 1619
rect 3620 1653 4020 1700
rect 3620 1619 3636 1653
rect 4004 1619 4020 1653
rect 3620 1603 4020 1619
rect 4078 1653 4478 1700
rect 4078 1619 4094 1653
rect 4462 1619 4478 1653
rect 4078 1603 4478 1619
rect 4536 1653 4936 1700
rect 4536 1619 4552 1653
rect 4920 1619 4936 1653
rect 4536 1603 4936 1619
rect 4994 1653 5394 1700
rect 4994 1619 5010 1653
rect 5378 1619 5394 1653
rect 4994 1603 5394 1619
rect 5452 1653 5852 1700
rect 5452 1619 5468 1653
rect 5836 1619 5852 1653
rect 5452 1603 5852 1619
rect 5910 1653 6310 1700
rect 5910 1619 5926 1653
rect 6294 1619 6310 1653
rect 5910 1603 6310 1619
rect 6368 1653 6768 1700
rect 6368 1619 6384 1653
rect 6752 1619 6768 1653
rect 6368 1603 6768 1619
rect 6826 1653 7226 1700
rect 6826 1619 6842 1653
rect 7210 1619 7226 1653
rect 6826 1603 7226 1619
rect 7284 1653 7684 1700
rect 7284 1619 7300 1653
rect 7668 1619 7684 1653
rect 7284 1603 7684 1619
<< polycont >>
rect -17248 8422 -17214 8790
rect -16820 6692 -16452 6726
rect -16248 6692 -15880 6726
rect -15676 6692 -15308 6726
rect -15104 6692 -14736 6726
rect -14532 6692 -14164 6726
rect -13960 6692 -13592 6726
rect -13388 6692 -13020 6726
rect -12816 6692 -12448 6726
rect -21750 5570 -21382 5604
rect -21292 5570 -20924 5604
rect -20834 5570 -20466 5604
rect -20376 5570 -20008 5604
rect -19918 5570 -19550 5604
rect -19460 5570 -19092 5604
rect -18546 4289 -18178 4323
rect -17974 4289 -17606 4323
rect -17402 4289 -17034 4323
rect -16830 4289 -16462 4323
rect -16258 4289 -15890 4323
rect -15686 4289 -15318 4323
rect -15114 4289 -14746 4323
rect -14542 4289 -14174 4323
rect -13970 4289 -13602 4323
rect -13398 4289 -13030 4323
rect -12826 4289 -12458 4323
rect -12254 4289 -11886 4323
rect -11682 4289 -11314 4323
rect -11110 4289 -10742 4323
rect -8738 1619 -8370 1653
rect -8280 1619 -7912 1653
rect -7822 1619 -7454 1653
rect -7364 1619 -6996 1653
rect -6906 1619 -6538 1653
rect -6448 1619 -6080 1653
rect -5990 1619 -5622 1653
rect -5532 1619 -5164 1653
rect -5074 1619 -4706 1653
rect -4616 1619 -4248 1653
rect -4158 1619 -3790 1653
rect -2780 1619 -2412 1653
rect -2322 1619 -1954 1653
rect -1864 1619 -1496 1653
rect -1406 1619 -1038 1653
rect -948 1619 -580 1653
rect -490 1619 -122 1653
rect -32 1619 336 1653
rect 426 1619 794 1653
rect 884 1619 1252 1653
rect 1342 1619 1710 1653
rect 2720 1619 3088 1653
rect 3178 1619 3546 1653
rect 3636 1619 4004 1653
rect 4094 1619 4462 1653
rect 4552 1619 4920 1653
rect 5010 1619 5378 1653
rect 5468 1619 5836 1653
rect 5926 1619 6294 1653
rect 6384 1619 6752 1653
rect 6842 1619 7210 1653
rect 7300 1619 7668 1653
<< xpolycontact >>
rect -5660 21562 -5090 21994
rect -8932 20176 -8362 20608
rect -8932 16420 -8362 16852
rect -8114 20176 -7544 20608
rect -8114 16420 -7544 16852
rect -7296 20176 -6726 20608
rect -7296 16420 -6726 16852
rect -5660 16830 -5090 17262
rect -4842 21562 -4272 21994
rect -4842 16830 -4272 17262
rect -4024 21562 -3454 21994
rect -4024 16830 -3454 17262
rect -3206 21562 -2636 21994
rect -3206 16830 -2636 17262
rect -752 21500 -182 21932
rect -752 14764 -182 15196
rect 66 21500 636 21932
rect 66 14764 636 15196
rect 884 21500 1454 21932
rect 884 14764 1454 15196
rect 1702 21500 2272 21932
rect 1702 14764 2272 15196
rect 2520 21500 3090 21932
rect 2520 14764 3090 15196
rect 3338 21500 3908 21932
rect 3338 14764 3908 15196
rect 4156 21500 4726 21932
rect 4156 14764 4726 15196
rect 4974 21500 5544 21932
rect 4974 14764 5544 15196
rect 5792 21500 6362 21932
rect 5792 14764 6362 15196
rect 6610 21500 7180 21932
rect 6610 14764 7180 15196
rect 7428 21500 7998 21932
rect 7428 14764 7998 15196
rect 8246 21500 8816 21932
rect 8246 14764 8816 15196
rect 9064 21500 9634 21932
rect 9064 14764 9634 15196
rect 9882 21500 10452 21932
rect 9882 14764 10452 15196
rect 10700 21500 11270 21932
rect 10700 14764 11270 15196
rect 11518 21500 12088 21932
rect 11518 14764 12088 15196
rect 12336 21500 12906 21932
rect 12336 14764 12906 15196
<< xpolyres >>
rect -8932 16852 -8362 20176
rect -8114 16852 -7544 20176
rect -7296 16852 -6726 20176
rect -5660 17262 -5090 21562
rect -4842 17262 -4272 21562
rect -4024 17262 -3454 21562
rect -3206 17262 -2636 21562
rect -752 15196 -182 21500
rect 66 15196 636 21500
rect 884 15196 1454 21500
rect 1702 15196 2272 21500
rect 2520 15196 3090 21500
rect 3338 15196 3908 21500
rect 4156 15196 4726 21500
rect 4974 15196 5544 21500
rect 5792 15196 6362 21500
rect 6610 15196 7180 21500
rect 7428 15196 7998 21500
rect 8246 15196 8816 21500
rect 9064 15196 9634 21500
rect 9882 15196 10452 21500
rect 10700 15196 11270 21500
rect 11518 15196 12088 21500
rect 12336 15196 12906 21500
<< locali >>
rect -6534 21562 -5660 21994
rect -2636 21932 -182 21994
rect -2636 21562 -752 21932
rect -6534 21516 -5930 21562
rect -9772 21500 -9170 21516
rect -9772 20608 -9756 21500
rect -9782 20166 -9756 20608
rect -9772 16106 -9756 20166
rect -9776 15602 -9756 16106
rect -9772 15196 -9756 15602
rect -9186 20608 -9170 21500
rect -6534 21500 -5926 21516
rect -3206 21500 -752 21562
rect 12906 21500 13730 21932
rect -6534 21004 -6512 21500
rect -6528 20608 -6512 21004
rect -9186 20176 -8932 20608
rect -8362 20176 -8114 20608
rect -7544 20176 -7296 20608
rect -6726 20176 -6512 20608
rect -9186 20166 -6512 20176
rect -9186 16106 -9170 20166
rect -6528 16852 -6512 20166
rect -5942 17258 -5926 21500
rect -1568 17262 -1552 21500
rect -6726 16420 -6512 16852
rect -8932 16110 -8362 16420
rect -6528 16110 -6512 16420
rect -5942 16830 -5660 17258
rect -5090 16830 -4984 17262
rect -3322 16830 -3206 17262
rect -2636 16830 -1552 17262
rect -5942 16732 -4984 16830
rect -3322 16732 -1552 16830
rect -8932 16106 -6512 16110
rect -9186 15602 -6512 16106
rect -9186 15196 -9170 15602
rect -9772 15180 -9170 15196
rect -6528 15196 -6512 15602
rect -5942 16110 -5926 16732
rect -5942 15602 -5916 16110
rect -5942 15196 -5926 15602
rect -1568 15196 -1552 16732
rect -982 15196 -966 21500
rect 13120 15196 13136 21500
rect 13706 15196 13722 21500
rect -6528 15180 -5926 15196
rect -1576 14764 -752 15196
rect 12906 14764 13730 15196
rect -8800 9428 -8766 9444
rect -17898 9388 -11414 9398
rect -17898 9044 -17888 9388
rect -11424 9044 -11414 9388
rect -17898 9034 -11414 9044
rect -9500 9102 -8900 9302
rect -17180 8818 -17164 8852
rect -11788 8818 -11772 8852
rect -17248 8790 -17214 8806
rect -17248 8406 -17214 8422
rect -17180 8360 -17164 8394
rect -11788 8360 -11772 8394
rect -16836 6692 -16820 6726
rect -16452 6692 -16436 6726
rect -16264 6692 -16248 6726
rect -15880 6692 -15864 6726
rect -15692 6692 -15676 6726
rect -15308 6692 -15292 6726
rect -15120 6692 -15104 6726
rect -14736 6692 -14720 6726
rect -14548 6692 -14532 6726
rect -14164 6692 -14148 6726
rect -13976 6692 -13960 6726
rect -13592 6692 -13576 6726
rect -13404 6692 -13388 6726
rect -13020 6692 -13004 6726
rect -12832 6692 -12816 6726
rect -12448 6692 -12432 6726
rect -17450 6642 -17318 6658
rect -20934 5836 -19910 5852
rect -20934 5760 -20918 5836
rect -19926 5760 -19910 5836
rect -20934 5720 -19910 5760
rect -22320 5682 -21888 5698
rect -22320 5106 -22304 5682
rect -21904 5604 -21888 5682
rect -20934 5668 -20906 5720
rect -20854 5668 -19990 5720
rect -19938 5668 -19910 5720
rect -20934 5656 -19910 5668
rect -18954 5682 -18522 5698
rect -18954 5604 -18938 5682
rect -21904 5570 -21750 5604
rect -21382 5570 -21366 5604
rect -21308 5570 -21292 5604
rect -20924 5570 -20834 5604
rect -20466 5570 -20376 5604
rect -20008 5570 -19918 5604
rect -19550 5570 -19534 5604
rect -19476 5570 -19460 5604
rect -19092 5570 -18938 5604
rect -21904 5520 -21778 5570
rect -21904 5144 -21812 5520
rect -21904 5128 -21778 5144
rect -21354 5520 -21320 5536
rect -21354 5128 -21320 5144
rect -20896 5520 -20862 5536
rect -20896 5128 -20862 5144
rect -20438 5520 -20404 5536
rect -20438 5128 -20404 5144
rect -19980 5520 -19946 5536
rect -19980 5128 -19946 5144
rect -19522 5520 -19488 5536
rect -19522 5128 -19488 5144
rect -19064 5520 -18938 5570
rect -19030 5144 -18938 5520
rect -19064 5128 -18938 5144
rect -21904 5106 -21888 5128
rect -22320 5090 -21888 5106
rect -18954 5106 -18938 5128
rect -18538 5106 -18522 5682
rect -18954 5090 -18522 5106
rect -17450 5042 -17434 6642
rect -17334 5042 -17318 6642
rect -17450 5026 -17318 5042
rect -16882 6642 -16848 6658
rect -16882 4850 -16848 4866
rect -16424 6642 -16390 6658
rect -16424 4850 -16390 4866
rect -16310 6642 -16276 6658
rect -16310 4850 -16276 4866
rect -15852 6642 -15818 6658
rect -15852 4850 -15818 4866
rect -15738 6642 -15704 6658
rect -15738 4850 -15704 4866
rect -15280 6642 -15246 6658
rect -15280 4850 -15246 4866
rect -15166 6642 -15132 6658
rect -15166 4850 -15132 4866
rect -14708 6642 -14674 6658
rect -14708 4850 -14674 4866
rect -14594 6642 -14560 6658
rect -14594 4850 -14560 4866
rect -14136 6642 -14102 6658
rect -14136 4850 -14102 4866
rect -14022 6642 -13988 6658
rect -14022 4850 -13988 4866
rect -13564 6642 -13530 6658
rect -13564 4850 -13530 4866
rect -13450 6642 -13416 6658
rect -13450 4850 -13416 4866
rect -12992 6642 -12958 6658
rect -12992 4850 -12958 4866
rect -12878 6642 -12844 6658
rect -12878 4850 -12844 4866
rect -12420 6642 -12386 6658
rect -11950 6642 -11818 6658
rect -11950 5042 -11934 6642
rect -11834 5042 -11818 6642
rect -11950 5026 -11818 5042
rect -12420 4850 -12386 4866
rect -18562 4289 -18546 4323
rect -18178 4289 -18162 4323
rect -17990 4289 -17974 4323
rect -17606 4289 -17590 4323
rect -17418 4289 -17402 4323
rect -17034 4289 -17018 4323
rect -16846 4289 -16830 4323
rect -16462 4289 -16446 4323
rect -16274 4289 -16258 4323
rect -15890 4289 -15874 4323
rect -15702 4289 -15686 4323
rect -15318 4289 -15302 4323
rect -15130 4289 -15114 4323
rect -14746 4289 -14730 4323
rect -14558 4289 -14542 4323
rect -14174 4289 -14158 4323
rect -13986 4289 -13970 4323
rect -13602 4289 -13586 4323
rect -13414 4289 -13398 4323
rect -13030 4289 -13014 4323
rect -12842 4289 -12826 4323
rect -12458 4289 -12442 4323
rect -12270 4289 -12254 4323
rect -11886 4289 -11870 4323
rect -11698 4289 -11682 4323
rect -11314 4289 -11298 4323
rect -11126 4289 -11110 4323
rect -10742 4289 -10726 4323
rect -18608 4230 -18574 4246
rect -19266 4142 -19134 4154
rect -19266 1800 -19250 4142
rect -19150 1800 -19134 4142
rect -19266 1784 -19134 1800
rect -18608 1658 -18574 1674
rect -18150 4230 -18116 4246
rect -18150 1658 -18116 1674
rect -18036 4230 -18002 4246
rect -18036 1658 -18002 1674
rect -17578 4230 -17544 4246
rect -17578 1658 -17544 1674
rect -17464 4230 -17430 4246
rect -17464 1658 -17430 1674
rect -17006 4230 -16972 4246
rect -17006 1658 -16972 1674
rect -16892 4230 -16858 4246
rect -16892 1658 -16858 1674
rect -16434 4230 -16400 4246
rect -16434 1658 -16400 1674
rect -16320 4230 -16286 4246
rect -16320 1658 -16286 1674
rect -15862 4230 -15828 4246
rect -15862 1658 -15828 1674
rect -15748 4230 -15714 4246
rect -15748 1658 -15714 1674
rect -15290 4230 -15256 4246
rect -15290 1658 -15256 1674
rect -15176 4230 -15142 4246
rect -15176 1658 -15142 1674
rect -14718 4230 -14684 4246
rect -14718 1658 -14684 1674
rect -14604 4230 -14570 4246
rect -14604 1658 -14570 1674
rect -14146 4230 -14112 4246
rect -14146 1658 -14112 1674
rect -14032 4230 -13998 4246
rect -14032 1658 -13998 1674
rect -13574 4230 -13540 4246
rect -13574 1658 -13540 1674
rect -13460 4230 -13426 4246
rect -13460 1658 -13426 1674
rect -13002 4230 -12968 4246
rect -13002 1658 -12968 1674
rect -12888 4230 -12854 4246
rect -12888 1658 -12854 1674
rect -12430 4230 -12396 4246
rect -12430 1658 -12396 1674
rect -12316 4230 -12282 4246
rect -12316 1658 -12282 1674
rect -11858 4230 -11824 4246
rect -11858 1658 -11824 1674
rect -11744 4230 -11710 4246
rect -11744 1658 -11710 1674
rect -11286 4230 -11252 4246
rect -11286 1658 -11252 1674
rect -11172 4230 -11138 4246
rect -11172 1658 -11138 1674
rect -10714 4230 -10680 4246
rect -10138 4142 -10006 4154
rect -10138 1800 -10122 4142
rect -10022 1800 -10006 4142
rect -10138 1784 -10006 1800
rect -9500 2102 -9300 9102
rect -9100 2102 -8900 9102
rect -10714 1658 -10680 1674
rect -15680 1296 -13310 1312
rect -15680 1196 -15668 1296
rect -13326 1196 -13310 1296
rect -15680 1180 -13310 1196
rect -9500 1202 -8900 2102
rect -8800 1696 -8766 1712
rect -8342 9428 -8308 9444
rect -8342 1696 -8308 1712
rect -7884 9428 -7850 9444
rect -7884 1696 -7850 1712
rect -7426 9428 -7392 9444
rect -7426 1696 -7392 1712
rect -6968 9428 -6934 9444
rect -6968 1696 -6934 1712
rect -6510 9428 -6476 9444
rect -6510 1696 -6476 1712
rect -6052 9428 -6018 9444
rect -6052 1696 -6018 1712
rect -5594 9428 -5560 9444
rect -5594 1696 -5560 1712
rect -5136 9428 -5102 9444
rect -5136 1696 -5102 1712
rect -4678 9428 -4644 9444
rect -4678 1696 -4644 1712
rect -4220 9428 -4186 9444
rect -4220 1696 -4186 1712
rect -3762 9428 -3728 9444
rect -2842 9428 -2808 9444
rect -3762 1696 -3728 1712
rect -3590 9102 -2990 9302
rect -3590 2102 -3390 9102
rect -3190 2102 -2990 9102
rect -8754 1619 -8738 1653
rect -8370 1619 -8354 1653
rect -8296 1619 -8280 1653
rect -7912 1619 -7896 1653
rect -7838 1619 -7822 1653
rect -7454 1619 -7438 1653
rect -7380 1619 -7364 1653
rect -6996 1619 -6980 1653
rect -6922 1619 -6906 1653
rect -6538 1619 -6522 1653
rect -6464 1619 -6448 1653
rect -6080 1619 -6064 1653
rect -6006 1619 -5990 1653
rect -5622 1619 -5606 1653
rect -5548 1619 -5532 1653
rect -5164 1619 -5148 1653
rect -5090 1619 -5074 1653
rect -4706 1619 -4690 1653
rect -4632 1619 -4616 1653
rect -4248 1619 -4232 1653
rect -4174 1619 -4158 1653
rect -3790 1619 -3774 1653
rect -9500 1102 -9400 1202
rect -9000 1102 -8900 1202
rect -9500 1002 -8900 1102
rect -3590 1202 -2990 2102
rect -2842 1696 -2808 1712
rect -2384 9428 -2350 9444
rect -2384 1696 -2350 1712
rect -1926 9428 -1892 9444
rect -1926 1696 -1892 1712
rect -1468 9428 -1434 9444
rect -1468 1696 -1434 1712
rect -1010 9428 -976 9444
rect -1010 1696 -976 1712
rect -552 9428 -518 9444
rect -552 1696 -518 1712
rect -94 9428 -60 9444
rect -94 1696 -60 1712
rect 364 9428 398 9444
rect 364 1696 398 1712
rect 822 9428 856 9444
rect 822 1696 856 1712
rect 1280 9428 1314 9444
rect 1280 1696 1314 1712
rect 1738 9428 1772 9444
rect 2658 9428 2692 9444
rect 1738 1696 1772 1712
rect 1910 9102 2510 9302
rect 1910 2102 2110 9102
rect 2310 2102 2510 9102
rect -2796 1619 -2780 1653
rect -2412 1619 -2396 1653
rect -2338 1619 -2322 1653
rect -1954 1619 -1938 1653
rect -1880 1619 -1864 1653
rect -1496 1619 -1480 1653
rect -1422 1619 -1406 1653
rect -1038 1619 -1022 1653
rect -964 1619 -948 1653
rect -580 1619 -564 1653
rect -506 1619 -490 1653
rect -122 1619 -106 1653
rect -48 1619 -32 1653
rect 336 1619 352 1653
rect 410 1619 426 1653
rect 794 1619 810 1653
rect 868 1619 884 1653
rect 1252 1619 1268 1653
rect 1326 1619 1342 1653
rect 1710 1619 1726 1653
rect -3590 1102 -3490 1202
rect -3090 1102 -2990 1202
rect -3590 1002 -2990 1102
rect 1910 1202 2510 2102
rect 2658 1696 2692 1712
rect 3116 9428 3150 9444
rect 3116 1696 3150 1712
rect 3574 9428 3608 9444
rect 3574 1696 3608 1712
rect 4032 9428 4066 9444
rect 4032 1696 4066 1712
rect 4490 9428 4524 9444
rect 4490 1696 4524 1712
rect 4948 9428 4982 9444
rect 4948 1696 4982 1712
rect 5406 9428 5440 9444
rect 5406 1696 5440 1712
rect 5864 9428 5898 9444
rect 5864 1696 5898 1712
rect 6322 9428 6356 9444
rect 6322 1696 6356 1712
rect 6780 9428 6814 9444
rect 6780 1696 6814 1712
rect 7238 9428 7272 9444
rect 7238 1696 7272 1712
rect 7696 9428 7730 9444
rect 7696 1696 7730 1712
rect 7866 9100 8466 9300
rect 7866 2100 8066 9100
rect 8266 2100 8466 9100
rect 2704 1619 2720 1653
rect 3088 1619 3104 1653
rect 3162 1619 3178 1653
rect 3546 1619 3562 1653
rect 3620 1619 3636 1653
rect 4004 1619 4020 1653
rect 4078 1619 4094 1653
rect 4462 1619 4478 1653
rect 4536 1619 4552 1653
rect 4920 1619 4936 1653
rect 4994 1619 5010 1653
rect 5378 1619 5394 1653
rect 5452 1619 5468 1653
rect 5836 1619 5852 1653
rect 5910 1619 5926 1653
rect 6294 1619 6310 1653
rect 6368 1619 6384 1653
rect 6752 1619 6768 1653
rect 6826 1619 6842 1653
rect 7210 1619 7226 1653
rect 7284 1619 7300 1653
rect 7668 1619 7684 1653
rect 1910 1102 2010 1202
rect 2410 1102 2510 1202
rect 1910 1002 2510 1102
rect 7866 1200 8466 2100
rect 7866 1100 7966 1200
rect 8366 1100 8466 1200
rect 7866 1000 8466 1100
<< viali >>
rect -21532 25036 -10316 25052
rect -21532 24270 -21516 25036
rect -21516 24270 -10332 25036
rect -10332 24270 -10316 25036
rect -21532 24254 -10316 24270
rect -5644 21579 -5106 21976
rect -4826 21579 -4288 21976
rect -4008 21579 -3470 21976
rect -3190 21579 -2652 21976
rect -736 21517 -198 21914
rect 82 21517 620 21914
rect 900 21517 1438 21914
rect 1718 21517 2256 21914
rect 2536 21517 3074 21914
rect 3354 21517 3892 21914
rect 4172 21517 4710 21914
rect 4990 21517 5528 21914
rect 5808 21517 6346 21914
rect 6626 21517 7164 21914
rect 7444 21517 7982 21914
rect 8262 21517 8800 21914
rect 9080 21517 9618 21914
rect 9898 21517 10436 21914
rect 10716 21517 11254 21914
rect 11534 21517 12072 21914
rect 12352 21517 12890 21914
rect -8916 20193 -8378 20590
rect -8098 20193 -7560 20590
rect -7280 20193 -6742 20590
rect -8916 16438 -8378 16835
rect -8098 16438 -7560 16835
rect -7280 16438 -6742 16835
rect -6460 16168 -5966 17234
rect -5644 16848 -5106 17245
rect -4826 16848 -4288 17245
rect -4008 16848 -3470 17245
rect -3190 16848 -2652 17245
rect -1508 16180 -996 17232
rect -736 14782 -198 15179
rect 82 14781 620 15179
rect 900 14782 1438 15179
rect 1718 14782 2256 15179
rect 2536 14781 3074 15179
rect 3354 14782 3892 15179
rect 4172 14782 4710 15179
rect 4990 14781 5528 15179
rect 5808 14782 6346 15179
rect 6626 14782 7164 15179
rect 7444 14782 7982 15179
rect 8262 14781 8800 15179
rect 9080 14782 9618 15179
rect 9898 14782 10436 15179
rect 10716 14782 11254 15179
rect 11534 14782 12072 15179
rect 12352 14782 12890 15179
rect -17888 9382 -11424 9388
rect -17888 9050 -17882 9382
rect -17882 9050 -11430 9382
rect -11430 9050 -11424 9382
rect -17888 9044 -11424 9050
rect -17164 8818 -11788 8852
rect -17248 8514 -17214 8698
rect -17164 8360 -11788 8394
rect -16728 6692 -16544 6726
rect -16156 6692 -15972 6726
rect -15584 6692 -15400 6726
rect -15012 6692 -14828 6726
rect -14440 6692 -14256 6726
rect -13868 6692 -13684 6726
rect -13296 6692 -13112 6726
rect -12724 6692 -12540 6726
rect -20906 5668 -20854 5720
rect -19990 5668 -19938 5720
rect -21658 5570 -21474 5604
rect -21200 5570 -21016 5604
rect -20742 5570 -20558 5604
rect -20284 5570 -20100 5604
rect -19826 5570 -19642 5604
rect -19368 5570 -19184 5604
rect -21812 5144 -21778 5520
rect -21354 5144 -21320 5520
rect -20896 5144 -20862 5520
rect -20438 5144 -20404 5520
rect -19980 5144 -19946 5520
rect -19522 5144 -19488 5520
rect -19064 5144 -19030 5520
rect -17434 5044 -17334 6642
rect -16882 4866 -16848 6642
rect -16424 4866 -16390 6642
rect -16310 4866 -16276 6642
rect -15852 4866 -15818 6642
rect -15738 4866 -15704 6642
rect -15280 4866 -15246 6642
rect -15166 4866 -15132 6642
rect -14708 4866 -14674 6642
rect -14594 4866 -14560 6642
rect -14136 4866 -14102 6642
rect -14022 4866 -13988 6642
rect -13564 4866 -13530 6642
rect -13450 4866 -13416 6642
rect -12992 4866 -12958 6642
rect -12878 4866 -12844 6642
rect -12420 4866 -12386 6642
rect -11934 5044 -11834 6642
rect -18454 4289 -18270 4323
rect -17882 4289 -17698 4323
rect -17310 4289 -17126 4323
rect -16738 4289 -16554 4323
rect -16166 4289 -15982 4323
rect -15594 4289 -15410 4323
rect -15022 4289 -14838 4323
rect -14450 4289 -14266 4323
rect -13878 4289 -13694 4323
rect -13306 4289 -13122 4323
rect -12734 4289 -12550 4323
rect -12162 4289 -11978 4323
rect -11590 4289 -11406 4323
rect -11018 4289 -10834 4323
rect -19250 1800 -19150 4142
rect -18608 1674 -18574 4230
rect -18150 1674 -18116 4230
rect -18036 1674 -18002 4230
rect -17578 1674 -17544 4230
rect -17464 1674 -17430 4230
rect -17006 1674 -16972 4230
rect -16892 1674 -16858 4230
rect -16434 1674 -16400 4230
rect -16320 1674 -16286 4230
rect -15862 1674 -15828 4230
rect -15748 1674 -15714 4230
rect -15290 1674 -15256 4230
rect -15176 1674 -15142 4230
rect -14718 1674 -14684 4230
rect -14604 1674 -14570 4230
rect -14146 1674 -14112 4230
rect -14032 1674 -13998 4230
rect -13574 1674 -13540 4230
rect -13460 1674 -13426 4230
rect -13002 1674 -12968 4230
rect -12888 1674 -12854 4230
rect -12430 1674 -12396 4230
rect -12316 1674 -12282 4230
rect -11858 1674 -11824 4230
rect -11744 1674 -11710 4230
rect -11286 1674 -11252 4230
rect -11172 1674 -11138 4230
rect -10714 1674 -10680 4230
rect -10122 1800 -10022 4142
rect -15668 1196 -13326 1296
rect -8800 1712 -8766 9428
rect -8342 1712 -8308 9428
rect -7884 1712 -7850 9428
rect -7426 1712 -7392 9428
rect -6968 1712 -6934 9428
rect -6510 1712 -6476 9428
rect -6052 1712 -6018 9428
rect -5594 1712 -5560 9428
rect -5136 1712 -5102 9428
rect -4678 1712 -4644 9428
rect -4220 1712 -4186 9428
rect -3762 1712 -3728 9428
rect -8646 1619 -8462 1653
rect -8188 1619 -8004 1653
rect -7730 1619 -7546 1653
rect -7272 1619 -7088 1653
rect -6814 1619 -6630 1653
rect -6356 1619 -6172 1653
rect -5898 1619 -5714 1653
rect -5440 1619 -5256 1653
rect -4982 1619 -4798 1653
rect -4524 1619 -4340 1653
rect -4066 1619 -3882 1653
rect -9400 1102 -9000 1202
rect -2842 1712 -2808 9428
rect -2384 1712 -2350 9428
rect -1926 1712 -1892 9428
rect -1468 1712 -1434 9428
rect -1010 1712 -976 9428
rect -552 1712 -518 9428
rect -94 1712 -60 9428
rect 364 1712 398 9428
rect 822 1712 856 9428
rect 1280 1712 1314 9428
rect 1738 1712 1772 9428
rect -2688 1619 -2504 1653
rect -2230 1619 -2046 1653
rect -1772 1619 -1588 1653
rect -1314 1619 -1130 1653
rect -856 1619 -672 1653
rect -398 1619 -214 1653
rect 60 1619 244 1653
rect 518 1619 702 1653
rect 976 1619 1160 1653
rect 1434 1619 1618 1653
rect -3490 1102 -3090 1202
rect 2658 1712 2692 9428
rect 3116 1712 3150 9428
rect 3574 1712 3608 9428
rect 4032 1712 4066 9428
rect 4490 1712 4524 9428
rect 4948 1712 4982 9428
rect 5406 1712 5440 9428
rect 5864 1712 5898 9428
rect 6322 1712 6356 9428
rect 6780 1712 6814 9428
rect 7238 1712 7272 9428
rect 7696 1712 7730 9428
rect 2812 1619 2996 1653
rect 3270 1619 3454 1653
rect 3728 1619 3912 1653
rect 4186 1619 4370 1653
rect 4644 1619 4828 1653
rect 5102 1619 5286 1653
rect 5560 1619 5744 1653
rect 6018 1619 6202 1653
rect 6476 1619 6660 1653
rect 6934 1619 7118 1653
rect 7392 1619 7576 1653
rect 2010 1102 2410 1202
rect 7966 1100 8366 1200
<< metal1 >>
rect -21552 25066 -10296 25072
rect -21552 24240 -21546 25066
rect -10302 24240 -10296 25066
rect -21552 24234 -10296 24240
rect 1714 23526 3908 23532
rect 1714 22968 1720 23526
rect 2278 22968 3344 23526
rect 3902 22968 3908 23526
rect 1714 22962 3908 22968
rect 7260 23526 10458 23532
rect 7260 22968 7434 23526
rect 7992 22968 9888 23526
rect 10446 22968 10458 23526
rect 7260 22962 10458 22968
rect -4842 22726 1454 22732
rect -4842 22168 -4836 22726
rect -4278 22168 890 22726
rect 1448 22168 1454 22726
rect -4842 22162 1454 22168
rect 4034 22726 7180 22732
rect 4034 22168 4162 22726
rect 4720 22168 6616 22726
rect 7174 22168 7180 22726
rect 4034 22162 7180 22168
rect 8950 22726 12088 22732
rect 8950 22168 9070 22726
rect 9628 22168 11524 22726
rect 12082 22168 12088 22726
rect 8950 22162 12088 22168
rect -4842 21988 -4272 21994
rect -5656 21976 -5094 21982
rect -5656 21579 -5644 21976
rect -5106 21579 -5094 21976
rect -5656 21573 -5094 21579
rect -4842 21568 -4836 21988
rect -4278 21568 -4272 21988
rect -4842 21562 -4272 21568
rect -4024 21988 -3454 21994
rect -4024 21568 -4018 21988
rect -3460 21568 -3454 21988
rect -3202 21976 -2640 21982
rect -3202 21579 -3190 21976
rect -2652 21579 -2640 21976
rect 66 21926 636 21932
rect -3202 21573 -2640 21579
rect -748 21914 -186 21920
rect -4024 21562 -3454 21568
rect -748 21517 -736 21914
rect -198 21517 -186 21914
rect -748 21511 -186 21517
rect 66 21506 72 21926
rect 630 21506 636 21926
rect 66 21500 636 21506
rect 884 21926 1454 21932
rect 884 21506 890 21926
rect 1448 21506 1454 21926
rect 884 21500 1454 21506
rect 1702 21926 2272 21932
rect 1702 21506 1708 21926
rect 2266 21506 2272 21926
rect 1702 21500 2272 21506
rect 2520 21926 3090 21932
rect 2520 21506 2526 21926
rect 3084 21506 3090 21926
rect 2520 21500 3090 21506
rect 3338 21926 3908 21932
rect 3338 21506 3344 21926
rect 3902 21506 3908 21926
rect 3338 21500 3908 21506
rect 4156 21926 4726 21932
rect 4156 21506 4162 21926
rect 4720 21506 4726 21926
rect 4156 21500 4726 21506
rect 4974 21926 5544 21932
rect 4974 21506 4980 21926
rect 5538 21506 5544 21926
rect 4974 21500 5544 21506
rect 5792 21926 6362 21932
rect 5792 21506 5798 21926
rect 6356 21506 6362 21926
rect 5792 21500 6362 21506
rect 6610 21926 7180 21932
rect 6610 21506 6616 21926
rect 7174 21506 7180 21926
rect 6610 21500 7180 21506
rect 7428 21926 7998 21932
rect 7428 21506 7434 21926
rect 7992 21506 7998 21926
rect 7428 21500 7998 21506
rect 8246 21926 8816 21932
rect 8246 21506 8252 21926
rect 8810 21506 8816 21926
rect 8246 21500 8816 21506
rect 9064 21926 9634 21932
rect 9064 21506 9070 21926
rect 9628 21506 9634 21926
rect 9064 21500 9634 21506
rect 9882 21926 10452 21932
rect 9882 21506 9888 21926
rect 10446 21506 10452 21926
rect 9882 21500 10452 21506
rect 10700 21926 11270 21932
rect 10700 21506 10706 21926
rect 11264 21506 11270 21926
rect 10700 21500 11270 21506
rect 11518 21926 12088 21932
rect 11518 21506 11524 21926
rect 12082 21506 12088 21926
rect 12340 21914 12902 21920
rect 12340 21517 12352 21914
rect 12890 21517 12902 21914
rect 12340 21511 12902 21517
rect 11518 21500 12088 21506
rect -4026 21264 636 21270
rect -4026 20772 -4018 21264
rect -3460 20772 72 21264
rect -4026 20706 72 20772
rect 630 20706 636 21264
rect -4026 20700 636 20706
rect 2520 21264 5544 21270
rect 2520 20706 2526 21264
rect 3084 20706 4980 21264
rect 5538 20706 5544 21264
rect 2520 20700 5544 20706
rect 8246 21264 11270 21270
rect 8246 20706 8252 21264
rect 8810 20706 10706 21264
rect 11264 20706 11270 21264
rect 8246 20700 11270 20706
rect -8928 20590 -8366 20596
rect -8928 20193 -8916 20590
rect -8378 20193 -8366 20590
rect -8928 20187 -8366 20193
rect -8110 20590 -7548 20596
rect -8110 20193 -8098 20590
rect -7560 20193 -7548 20590
rect -8110 20187 -7548 20193
rect -7292 20590 -6730 20596
rect -7292 20193 -7280 20590
rect -6742 20193 -6730 20590
rect -7292 20187 -6730 20193
rect -6482 17245 -986 17262
rect -6482 17234 -5644 17245
rect -8928 16835 -8366 16841
rect -8928 16438 -8916 16835
rect -8378 16438 -8366 16835
rect -8928 16432 -8366 16438
rect -8114 16835 -7544 16852
rect -8114 16438 -8098 16835
rect -7560 16438 -7544 16835
rect -8114 15996 -7544 16438
rect -7292 16835 -6730 16841
rect -7292 16438 -7280 16835
rect -6742 16438 -6730 16835
rect -7292 16432 -6730 16438
rect -6482 16168 -6460 17234
rect -5966 16848 -5644 17234
rect -5106 16848 -4826 17245
rect -4288 16848 -4008 17245
rect -3470 16848 -3190 17245
rect -2652 17232 -986 17245
rect -2652 16848 -1508 17232
rect -5966 16180 -1508 16848
rect -996 16180 -986 17232
rect 884 16790 4726 16796
rect 884 16232 890 16790
rect 1448 16232 4162 16790
rect 4720 16232 4726 16790
rect 884 16226 4726 16232
rect 6616 16790 9634 16796
rect 7174 16232 9070 16790
rect 9628 16232 9634 16790
rect 6616 16226 9634 16232
rect -5966 16168 -986 16180
rect -6482 16126 -986 16168
rect -8114 15990 2272 15996
rect -8114 15432 1708 15990
rect 2266 15432 2272 15990
rect -8114 15426 2272 15432
rect 3338 15990 7998 15996
rect 3338 15432 3344 15990
rect 3902 15432 7434 15990
rect 7992 15432 7998 15990
rect 3338 15426 7998 15432
rect 66 15190 636 15196
rect -748 15179 -186 15185
rect -748 14782 -736 15179
rect -198 14782 -186 15179
rect -748 14776 -186 14782
rect 66 14770 72 15190
rect 630 14770 636 15190
rect 66 14764 636 14770
rect 884 15190 1454 15196
rect 884 14770 890 15190
rect 1448 14770 1454 15190
rect 884 14764 1454 14770
rect 1702 15190 2272 15196
rect 1702 14770 1708 15190
rect 2266 14770 2272 15190
rect 1702 14764 2272 14770
rect 2520 15190 3090 15196
rect 2520 14770 2526 15190
rect 3084 14770 3090 15190
rect 2520 14764 3090 14770
rect 3338 15190 3908 15196
rect 3338 14770 3344 15190
rect 3902 14770 3908 15190
rect 3338 14764 3908 14770
rect 4156 15190 4726 15196
rect 4156 14770 4162 15190
rect 4720 14770 4726 15190
rect 4156 14764 4726 14770
rect 4974 15190 5544 15196
rect 4974 14770 4980 15190
rect 5538 14770 5544 15190
rect 4974 14764 5544 14770
rect 5714 15190 6418 15196
rect 5714 15158 5798 15190
rect 5714 14640 5720 15158
rect 6356 15158 6418 15190
rect 6412 14640 6418 15158
rect 6610 15190 7180 15196
rect 6610 14770 6616 15190
rect 7174 14770 7180 15190
rect 6610 14764 7180 14770
rect 7428 15190 7998 15196
rect 7428 14770 7434 15190
rect 7992 14770 7998 15190
rect 7428 14764 7998 14770
rect 8246 15190 8816 15196
rect 8246 14770 8252 15190
rect 8810 14770 8816 15190
rect 8246 14764 8816 14770
rect 9064 15190 9634 15196
rect 9064 14770 9070 15190
rect 9628 14770 9634 15190
rect 9064 14764 9634 14770
rect 9804 15190 10508 15196
rect 66 14528 3090 14534
rect 66 13970 72 14528
rect 630 13970 2526 14528
rect 3084 13970 3090 14528
rect 66 13964 3090 13970
rect 4974 14528 8816 14534
rect 4974 13970 4980 14528
rect 5538 13970 8252 14528
rect 8810 13970 8816 14528
rect 4974 13964 8816 13970
rect 9804 14498 9810 15190
rect 10502 14498 10508 15190
rect 9804 13500 10508 14498
rect -2890 12808 10508 13500
rect 10622 15190 11326 15196
rect 10622 14498 10628 15190
rect 11320 14498 11326 15190
rect -8390 11860 -6390 11902
rect -8390 11410 -8384 11860
rect -6396 11410 -6390 11860
rect -9908 11104 -9776 11110
rect -9908 10690 -9902 11104
rect -9782 10690 -9776 11104
rect -10364 10398 -10232 10684
rect -10364 10106 -10358 10398
rect -10238 10106 -10232 10398
rect -17900 9388 -11412 9400
rect -17900 9044 -17888 9388
rect -11424 9044 -11412 9388
rect -17900 8852 -11412 9044
rect -17900 8832 -17164 8852
rect -17176 8818 -17164 8832
rect -11788 8832 -11412 8852
rect -11788 8818 -11776 8832
rect -17176 8812 -11776 8818
rect -19254 8698 -17208 8710
rect -19254 8514 -17248 8698
rect -17214 8514 -17208 8698
rect -19254 8502 -17208 8514
rect -17176 8394 -11776 8400
rect -17894 8360 -17164 8394
rect -11788 8360 -11418 8394
rect -17894 8038 -11418 8360
rect -20918 5720 -20842 5732
rect -20918 5668 -20906 5720
rect -20854 5668 -20842 5720
rect -20918 5656 -20842 5668
rect -20002 5720 -19926 5732
rect -20002 5668 -19990 5720
rect -19938 5668 -19926 5720
rect -20002 5656 -19926 5668
rect -21670 5604 -21462 5610
rect -21224 5604 -20992 5616
rect -21670 5570 -21658 5604
rect -21474 5570 -21462 5604
rect -21670 5564 -21462 5570
rect -21360 5570 -21200 5604
rect -21016 5570 -20992 5604
rect -21360 5532 -21316 5570
rect -21224 5552 -20992 5570
rect -21818 5520 -21772 5532
rect -21818 5144 -21812 5520
rect -21778 5144 -21772 5520
rect -21818 5132 -21772 5144
rect -21360 5520 -21314 5532
rect -21360 5144 -21354 5520
rect -21320 5144 -21314 5520
rect -21360 5002 -21314 5144
rect -20902 5520 -20856 5656
rect -20754 5604 -20546 5610
rect -20754 5570 -20742 5604
rect -20558 5570 -20546 5604
rect -20754 5564 -20546 5570
rect -20296 5604 -20088 5610
rect -20296 5570 -20284 5604
rect -20100 5570 -20088 5604
rect -20296 5564 -20088 5570
rect -20902 5144 -20896 5520
rect -20862 5144 -20856 5520
rect -20902 5132 -20856 5144
rect -20444 5520 -20398 5532
rect -20444 5144 -20438 5520
rect -20404 5144 -20398 5520
rect -21370 4996 -21306 5002
rect -21370 4944 -21364 4996
rect -21312 4944 -21306 4996
rect -21370 4938 -21306 4944
rect -20444 4796 -20398 5144
rect -19986 5520 -19940 5656
rect -19860 5604 -19628 5616
rect -19380 5604 -19172 5610
rect -19860 5570 -19826 5604
rect -19642 5570 -19482 5604
rect -19860 5552 -19628 5570
rect -19986 5144 -19980 5520
rect -19946 5144 -19940 5520
rect -19986 5132 -19940 5144
rect -19528 5520 -19482 5570
rect -19380 5570 -19368 5604
rect -19184 5570 -19172 5604
rect -19380 5564 -19172 5570
rect -19528 5144 -19522 5520
rect -19488 5144 -19482 5520
rect -19528 5008 -19482 5144
rect -19070 5520 -19024 5532
rect -19070 5144 -19064 5520
rect -19030 5144 -19024 5520
rect -19070 5132 -19024 5144
rect -19536 5002 -19472 5008
rect -19536 4950 -19530 5002
rect -19478 4950 -19472 5002
rect -19536 4944 -19472 4950
rect -18930 5002 -18724 5008
rect -18930 4944 -18924 5002
rect -18730 4944 -18724 5002
rect -20452 4790 -20388 4796
rect -20452 4738 -20446 4790
rect -20394 4738 -20388 4790
rect -20452 4732 -20388 4738
rect -19266 4142 -19134 4154
rect -19266 1800 -19250 4142
rect -19150 1800 -19134 4142
rect -19266 1552 -19134 1800
rect -19266 1448 -19240 1552
rect -19188 1448 -19134 1552
rect -19266 1438 -19134 1448
rect -18930 1358 -18724 4944
rect -17894 4630 -17686 8038
rect -15584 6986 -15400 7006
rect -15584 6932 -15564 6986
rect -15420 6932 -15400 6986
rect -16156 6846 -15972 6866
rect -16156 6792 -16136 6846
rect -15992 6792 -15972 6846
rect -16156 6732 -15972 6792
rect -15584 6732 -15400 6932
rect -14440 6986 -14256 7006
rect -14440 6932 -14420 6986
rect -14276 6932 -14256 6986
rect -15012 6846 -14828 6866
rect -15012 6792 -14992 6846
rect -14848 6792 -14828 6846
rect -15012 6732 -14828 6792
rect -14440 6732 -14256 6932
rect -13296 6986 -13112 7006
rect -13296 6932 -13276 6986
rect -13132 6932 -13112 6986
rect -13868 6846 -13684 6866
rect -13868 6792 -13848 6846
rect -13704 6792 -13684 6846
rect -13868 6732 -13684 6792
rect -13296 6732 -13112 6932
rect -17440 6726 -16384 6732
rect -17440 6692 -16728 6726
rect -16544 6692 -16384 6726
rect -17440 6686 -16384 6692
rect -16168 6726 -15960 6732
rect -16168 6692 -16156 6726
rect -15972 6692 -15960 6726
rect -16168 6686 -15960 6692
rect -15596 6726 -15388 6732
rect -15596 6692 -15584 6726
rect -15400 6692 -15388 6726
rect -15596 6686 -15388 6692
rect -15024 6726 -14816 6732
rect -15024 6692 -15012 6726
rect -14828 6692 -14816 6726
rect -15024 6686 -14816 6692
rect -14452 6726 -14244 6732
rect -14452 6692 -14440 6726
rect -14256 6692 -14244 6726
rect -14452 6686 -14244 6692
rect -13880 6726 -13672 6732
rect -13880 6692 -13868 6726
rect -13684 6692 -13672 6726
rect -13880 6686 -13672 6692
rect -13308 6726 -13100 6732
rect -13308 6692 -13296 6726
rect -13112 6692 -13100 6726
rect -13308 6686 -13100 6692
rect -12884 6726 -11828 6732
rect -12884 6692 -12724 6726
rect -12540 6692 -11828 6726
rect -12884 6686 -11828 6692
rect -17440 6658 -17326 6686
rect -17450 6642 -17318 6658
rect -17450 5044 -17434 6642
rect -17334 5044 -17318 6642
rect -17450 5026 -17318 5044
rect -16888 6642 -16842 6686
rect -16888 4866 -16882 6642
rect -16848 4866 -16842 6642
rect -16888 4854 -16842 4866
rect -16430 6642 -16384 6686
rect -16430 4866 -16424 6642
rect -16390 4866 -16384 6642
rect -16430 4854 -16384 4866
rect -16316 6642 -16270 6654
rect -16316 4866 -16310 6642
rect -16276 4866 -16270 6642
rect -16316 4854 -16270 4866
rect -15858 6642 -15812 6654
rect -15858 4866 -15852 6642
rect -15818 4866 -15812 6642
rect -15858 4854 -15812 4866
rect -15744 6642 -15698 6654
rect -15744 4866 -15738 6642
rect -15704 4866 -15698 6642
rect -15744 4854 -15698 4866
rect -15286 6642 -15240 6654
rect -15286 4866 -15280 6642
rect -15246 4866 -15240 6642
rect -15286 4854 -15240 4866
rect -15172 6642 -15126 6654
rect -15172 4866 -15166 6642
rect -15132 4866 -15126 6642
rect -15172 4854 -15126 4866
rect -14714 6642 -14668 6654
rect -14714 4866 -14708 6642
rect -14674 4866 -14668 6642
rect -14714 4854 -14668 4866
rect -14600 6642 -14554 6654
rect -14600 4866 -14594 6642
rect -14560 4866 -14554 6642
rect -14600 4854 -14554 4866
rect -14142 6642 -14096 6654
rect -14142 4866 -14136 6642
rect -14102 4866 -14096 6642
rect -14142 4854 -14096 4866
rect -14028 6642 -13982 6654
rect -14028 4866 -14022 6642
rect -13988 4866 -13982 6642
rect -14028 4854 -13982 4866
rect -13570 6642 -13524 6654
rect -13570 4866 -13564 6642
rect -13530 4866 -13524 6642
rect -13570 4854 -13524 4866
rect -13456 6642 -13410 6654
rect -13456 4866 -13450 6642
rect -13416 4866 -13410 6642
rect -13456 4854 -13410 4866
rect -12998 6642 -12952 6654
rect -12998 4866 -12992 6642
rect -12958 4866 -12952 6642
rect -12998 4854 -12952 4866
rect -12884 6642 -12838 6686
rect -12884 4866 -12878 6642
rect -12844 4866 -12838 6642
rect -12884 4854 -12838 4866
rect -12426 6642 -12380 6686
rect -11942 6658 -11828 6686
rect -12426 4866 -12420 6642
rect -12386 4866 -12380 6642
rect -11950 6642 -11818 6658
rect -11950 5044 -11934 6642
rect -11834 5044 -11818 6642
rect -11950 5026 -11818 5044
rect -12426 4854 -12380 4866
rect -17894 4376 -17768 4630
rect -17716 4376 -17686 4630
rect -18614 4323 -18110 4330
rect -18614 4289 -18454 4323
rect -18270 4289 -18110 4323
rect -18614 4282 -18110 4289
rect -17894 4323 -17686 4376
rect -17894 4289 -17882 4323
rect -17698 4289 -17686 4323
rect -17894 4282 -17686 4289
rect -17334 4630 -17126 4636
rect -17334 4376 -17208 4630
rect -17156 4376 -17126 4630
rect -17334 4329 -17126 4376
rect -16774 4630 -16566 4636
rect -16774 4376 -16648 4630
rect -16596 4376 -16566 4630
rect -16774 4329 -16566 4376
rect -17334 4323 -17114 4329
rect -17334 4289 -17310 4323
rect -17126 4289 -17114 4323
rect -17334 4283 -17114 4289
rect -16774 4323 -16542 4329
rect -16774 4289 -16738 4323
rect -16554 4289 -16542 4323
rect -16774 4283 -16542 4289
rect -16312 4324 -16278 4854
rect -15852 4790 -15818 4854
rect -15878 4780 -15806 4790
rect -15878 4676 -15868 4780
rect -15816 4676 -15806 4780
rect -15878 4666 -15806 4676
rect -15740 4636 -15706 4854
rect -15280 4790 -15246 4854
rect -15306 4780 -15234 4790
rect -15306 4676 -15296 4780
rect -15244 4676 -15234 4780
rect -15306 4666 -15234 4676
rect -15754 4630 -15690 4636
rect -15754 4376 -15748 4630
rect -15696 4376 -15690 4630
rect -15754 4370 -15690 4376
rect -16176 4340 -15956 4342
rect -16176 4329 -16170 4340
rect -16178 4324 -16170 4329
rect -16312 4284 -16170 4324
rect -15962 4320 -15956 4340
rect -17334 4282 -17126 4283
rect -16774 4282 -16566 4283
rect -18614 4230 -18568 4282
rect -18614 1674 -18608 4230
rect -18574 1674 -18568 4230
rect -18614 1562 -18568 1674
rect -18156 4230 -18110 4282
rect -16312 4242 -16278 4284
rect -16178 4283 -16170 4284
rect -16176 4282 -16170 4283
rect -15962 4284 -15866 4320
rect -15962 4282 -15956 4284
rect -16176 4272 -15956 4282
rect -15740 4242 -15706 4370
rect -15604 4336 -15384 4342
rect -15604 4329 -15598 4336
rect -15606 4283 -15598 4329
rect -15604 4278 -15598 4283
rect -15390 4278 -15384 4336
rect -15604 4272 -15384 4278
rect -15168 4324 -15134 4854
rect -14708 4790 -14674 4854
rect -14734 4780 -14662 4790
rect -14734 4676 -14724 4780
rect -14672 4676 -14662 4780
rect -14734 4666 -14662 4676
rect -14596 4636 -14562 4854
rect -14136 4790 -14102 4854
rect -14162 4780 -14090 4790
rect -14162 4676 -14152 4780
rect -14100 4676 -14090 4780
rect -14162 4666 -14090 4676
rect -14610 4630 -14546 4636
rect -14610 4376 -14604 4630
rect -14552 4376 -14546 4630
rect -14610 4370 -14546 4376
rect -15032 4340 -14812 4346
rect -15032 4329 -15026 4340
rect -15034 4324 -15026 4329
rect -15168 4288 -15026 4324
rect -14818 4324 -14812 4340
rect -15168 4242 -15134 4288
rect -15034 4283 -15026 4288
rect -15032 4282 -15026 4283
rect -14818 4288 -14722 4324
rect -14818 4282 -14812 4288
rect -15032 4276 -14812 4282
rect -14596 4242 -14562 4370
rect -14460 4340 -14240 4346
rect -14460 4329 -14454 4340
rect -14462 4283 -14454 4329
rect -14460 4282 -14454 4283
rect -14246 4282 -14240 4340
rect -14460 4276 -14240 4282
rect -14024 4324 -13990 4854
rect -13564 4790 -13530 4854
rect -13590 4780 -13518 4790
rect -13590 4676 -13580 4780
rect -13528 4676 -13518 4780
rect -13590 4666 -13518 4676
rect -13452 4636 -13418 4854
rect -12992 4790 -12958 4854
rect -13018 4780 -12946 4790
rect -13018 4676 -13008 4780
rect -12956 4676 -12946 4780
rect -13018 4666 -12946 4676
rect -13466 4630 -13402 4636
rect -13466 4376 -13460 4630
rect -13408 4376 -13402 4630
rect -13466 4370 -13402 4376
rect -12746 4630 -12538 4636
rect -12746 4376 -12660 4630
rect -12608 4376 -12538 4630
rect -13888 4340 -13668 4346
rect -13888 4329 -13882 4340
rect -13890 4324 -13882 4329
rect -14024 4288 -13882 4324
rect -13674 4324 -13668 4340
rect -14024 4242 -13990 4288
rect -13890 4283 -13882 4288
rect -13888 4282 -13882 4283
rect -13674 4288 -13578 4324
rect -13674 4282 -13668 4288
rect -13888 4276 -13668 4282
rect -13452 4242 -13418 4370
rect -13316 4340 -13096 4346
rect -13316 4329 -13310 4340
rect -13318 4283 -13310 4329
rect -13316 4282 -13310 4283
rect -13102 4282 -13096 4340
rect -12746 4323 -12538 4376
rect -12746 4289 -12734 4323
rect -12550 4289 -12538 4323
rect -12746 4282 -12538 4289
rect -12186 4630 -11978 4636
rect -12186 4376 -12100 4630
rect -12048 4376 -11978 4630
rect -12186 4329 -11978 4376
rect -11626 4630 -11418 8038
rect -10364 6866 -10232 10106
rect -9908 7006 -9776 10690
rect -8390 10996 -6390 11410
rect -8390 10708 -8384 10996
rect -6396 10708 -6390 10996
rect -8390 9502 -6390 10708
rect -5690 10396 -3690 10408
rect -5690 10108 -5684 10396
rect -3696 10108 -3690 10396
rect -5690 9502 -3690 10108
rect -8350 9440 -8310 9502
rect -7430 9440 -7390 9502
rect -6510 9440 -6470 9502
rect -9908 6926 -9902 7006
rect -9782 6926 -9776 7006
rect -9908 6920 -9776 6926
rect -8806 9428 -8760 9440
rect -10364 6786 -10358 6866
rect -10248 6786 -10232 6866
rect -10364 6780 -10232 6786
rect -11626 4376 -11540 4630
rect -11488 4376 -11418 4630
rect -11626 4329 -11418 4376
rect -9496 4630 -9016 4636
rect -9496 4376 -9490 4630
rect -9022 4376 -9016 4630
rect -12186 4323 -11966 4329
rect -12186 4289 -12162 4323
rect -11978 4289 -11966 4323
rect -12186 4283 -11966 4289
rect -11626 4323 -11394 4329
rect -11626 4289 -11590 4323
rect -11406 4289 -11394 4323
rect -11626 4283 -11394 4289
rect -11178 4323 -10674 4330
rect -11178 4289 -11018 4323
rect -10834 4289 -10674 4323
rect -12186 4282 -11978 4283
rect -11626 4282 -11418 4283
rect -11178 4282 -10674 4289
rect -13316 4276 -13096 4282
rect -18156 1674 -18150 4230
rect -18116 1674 -18110 4230
rect -18156 1562 -18110 1674
rect -18042 4230 -17996 4242
rect -18042 1674 -18036 4230
rect -18002 1674 -17996 4230
rect -18042 1662 -17996 1674
rect -17584 4230 -17538 4242
rect -17584 1674 -17578 4230
rect -17544 1674 -17538 4230
rect -17584 1662 -17538 1674
rect -17470 4230 -17424 4242
rect -17470 1674 -17464 4230
rect -17430 1674 -17424 4230
rect -17470 1662 -17424 1674
rect -17012 4230 -16966 4242
rect -17012 1674 -17006 4230
rect -16972 4226 -16966 4230
rect -16898 4230 -16852 4242
rect -16972 1674 -16964 4226
rect -17012 1662 -16964 1674
rect -16898 1674 -16892 4230
rect -16858 1674 -16852 4230
rect -16898 1662 -16852 1674
rect -16440 4230 -16394 4242
rect -16440 1674 -16434 4230
rect -16400 4226 -16394 4230
rect -16326 4230 -16278 4242
rect -16400 1674 -16384 4226
rect -16440 1662 -16384 1674
rect -16326 1674 -16320 4230
rect -16286 4226 -16278 4230
rect -15868 4230 -15822 4242
rect -16286 1674 -16280 4226
rect -16326 1662 -16280 1674
rect -15868 1674 -15862 4230
rect -15828 4226 -15822 4230
rect -15754 4230 -15706 4242
rect -15296 4230 -15250 4242
rect -15828 1674 -15820 4226
rect -15868 1662 -15820 1674
rect -15754 1674 -15748 4230
rect -15714 1674 -15708 4230
rect -15754 1662 -15708 1674
rect -15296 1674 -15290 4230
rect -15256 4226 -15250 4230
rect -15182 4230 -15134 4242
rect -14724 4230 -14678 4242
rect -15256 1674 -15248 4226
rect -15296 1662 -15248 1674
rect -15182 1674 -15176 4230
rect -15142 1674 -15136 4230
rect -15182 1662 -15136 1674
rect -14724 1674 -14718 4230
rect -14684 1674 -14678 4230
rect -14724 1662 -14678 1674
rect -14610 4230 -14562 4242
rect -14152 4230 -14106 4242
rect -14610 1674 -14604 4230
rect -14570 1674 -14564 4230
rect -14610 1662 -14564 1674
rect -14152 1674 -14146 4230
rect -14112 1674 -14106 4230
rect -14152 1662 -14106 1674
rect -14038 4230 -13990 4242
rect -13580 4230 -13534 4242
rect -14038 1674 -14032 4230
rect -13998 1674 -13992 4230
rect -14038 1662 -13992 1674
rect -13580 1674 -13574 4230
rect -13540 1674 -13534 4230
rect -13580 1662 -13534 1674
rect -13466 4230 -13418 4242
rect -13008 4230 -12962 4242
rect -13466 1674 -13460 4230
rect -13426 1674 -13420 4230
rect -13466 1662 -13420 1674
rect -13008 1674 -13002 4230
rect -12968 1674 -12962 4230
rect -13008 1662 -12962 1674
rect -12894 4230 -12848 4242
rect -12894 1674 -12888 4230
rect -12854 1674 -12848 4230
rect -12894 1662 -12848 1674
rect -12436 4230 -12390 4242
rect -12436 1674 -12430 4230
rect -12396 1674 -12390 4230
rect -12436 1662 -12390 1674
rect -12322 4230 -12276 4242
rect -12322 1674 -12316 4230
rect -12282 1674 -12276 4230
rect -12322 1662 -12276 1674
rect -11864 4230 -11818 4242
rect -11864 1674 -11858 4230
rect -11824 1674 -11818 4230
rect -11864 1662 -11818 1674
rect -11750 4230 -11704 4242
rect -11750 1674 -11744 4230
rect -11710 1674 -11704 4230
rect -11750 1662 -11704 1674
rect -11292 4230 -11246 4242
rect -11292 1674 -11286 4230
rect -11252 1674 -11246 4230
rect -11292 1662 -11246 1674
rect -11178 4230 -11132 4282
rect -11178 1674 -11172 4230
rect -11138 1674 -11132 4230
rect -18628 1552 -18556 1562
rect -18628 1448 -18618 1552
rect -18566 1448 -18556 1552
rect -18628 1438 -18556 1448
rect -18170 1552 -18098 1562
rect -18170 1448 -18160 1552
rect -18108 1448 -18098 1552
rect -18170 1438 -18098 1448
rect -18040 1362 -17998 1662
rect -17578 1562 -17544 1662
rect -17594 1552 -17522 1562
rect -17594 1448 -17584 1552
rect -17532 1448 -17522 1552
rect -17594 1438 -17522 1448
rect -17468 1362 -17426 1662
rect -17006 1562 -16964 1662
rect -17022 1552 -16950 1562
rect -17022 1448 -17012 1552
rect -16960 1448 -16950 1552
rect -17022 1438 -16950 1448
rect -16896 1362 -16854 1662
rect -16434 1562 -16384 1662
rect -15862 1562 -15820 1662
rect -15290 1562 -15248 1662
rect -14718 1562 -14684 1662
rect -14146 1562 -14112 1662
rect -13574 1562 -13540 1662
rect -13002 1562 -12968 1662
rect -16450 1552 -16378 1562
rect -16450 1448 -16440 1552
rect -16388 1448 -16378 1552
rect -16450 1438 -16378 1448
rect -15878 1552 -15806 1562
rect -15878 1448 -15868 1552
rect -15816 1448 -15806 1552
rect -15878 1438 -15806 1448
rect -15306 1552 -15234 1562
rect -15306 1448 -15296 1552
rect -15244 1448 -15234 1552
rect -15306 1438 -15234 1448
rect -14734 1552 -14662 1562
rect -14734 1448 -14724 1552
rect -14672 1448 -14662 1552
rect -14734 1438 -14662 1448
rect -14162 1552 -14090 1562
rect -14162 1448 -14152 1552
rect -14100 1448 -14090 1552
rect -14162 1438 -14090 1448
rect -13590 1552 -13518 1562
rect -13590 1448 -13580 1552
rect -13528 1448 -13518 1552
rect -13590 1438 -13518 1448
rect -13018 1552 -12950 1562
rect -13018 1448 -13008 1552
rect -12956 1448 -12950 1552
rect -13018 1438 -12950 1448
rect -12892 1362 -12850 1662
rect -12430 1562 -12396 1662
rect -12446 1552 -12378 1562
rect -12446 1448 -12436 1552
rect -12384 1448 -12378 1552
rect -12446 1438 -12378 1448
rect -12320 1362 -12278 1662
rect -11858 1562 -11824 1662
rect -11874 1552 -11806 1562
rect -11874 1448 -11864 1552
rect -11812 1448 -11806 1552
rect -11874 1438 -11806 1448
rect -11748 1362 -11706 1662
rect -11286 1562 -11252 1662
rect -11178 1562 -11132 1674
rect -10720 4230 -10674 4282
rect -10720 1674 -10714 4230
rect -10680 1674 -10674 4230
rect -10720 1562 -10674 1674
rect -10138 4142 -10006 4154
rect -10138 1800 -10122 4142
rect -10022 1800 -10006 4142
rect -11302 1552 -11234 1562
rect -11302 1448 -11292 1552
rect -11240 1448 -11234 1552
rect -11302 1438 -11234 1448
rect -11192 1552 -11120 1562
rect -11192 1448 -11182 1552
rect -11130 1448 -11120 1552
rect -11192 1438 -11120 1448
rect -10734 1552 -10662 1562
rect -10734 1448 -10724 1552
rect -10672 1448 -10662 1552
rect -10734 1438 -10662 1448
rect -10138 1552 -10006 1800
rect -10138 1448 -10112 1552
rect -10060 1448 -10006 1552
rect -10138 1438 -10006 1448
rect -9496 1536 -9016 4376
rect -9496 1388 -9490 1536
rect -9022 1388 -9016 1536
rect -9496 1382 -9016 1388
rect -8806 1712 -8800 9428
rect -8766 1712 -8760 9428
rect -8350 9428 -8302 9440
rect -8350 9402 -8342 9428
rect -8806 1660 -8760 1712
rect -8348 1712 -8342 9402
rect -8308 1712 -8302 9428
rect -8348 1696 -8302 1712
rect -7890 9428 -7844 9440
rect -7890 1712 -7884 9428
rect -7850 1712 -7844 9428
rect -7890 1700 -7844 1712
rect -7432 9428 -7386 9440
rect -7432 1712 -7426 9428
rect -7392 1712 -7386 9428
rect -7432 1700 -7386 1712
rect -6974 9428 -6928 9440
rect -6974 1712 -6968 9428
rect -6934 1712 -6928 9428
rect -6974 1700 -6928 1712
rect -6516 9428 -6470 9440
rect -6516 1712 -6510 9428
rect -6476 1712 -6470 9428
rect -6516 1700 -6470 1712
rect -6058 9428 -6012 9440
rect -6058 1712 -6052 9428
rect -6018 1722 -6012 9428
rect -5610 9428 -5550 9502
rect -5610 9422 -5594 9428
rect -6018 1712 -6010 1722
rect -6058 1700 -6010 1712
rect -5600 1712 -5594 9422
rect -5560 9422 -5550 9428
rect -5142 9428 -5096 9440
rect -5560 1712 -5554 9422
rect -5142 1722 -5136 9428
rect -5600 1700 -5554 1712
rect -5150 1712 -5136 1722
rect -5102 1712 -5096 9428
rect -4690 9428 -4630 9502
rect -4690 9402 -4678 9428
rect -5150 1700 -5096 1712
rect -4684 1712 -4678 9402
rect -4644 9402 -4630 9428
rect -4226 9428 -4180 9440
rect -4644 1712 -4638 9402
rect -4226 1722 -4220 9428
rect -4684 1700 -4638 1712
rect -4230 1712 -4220 1722
rect -4186 1712 -4180 9428
rect -3770 9428 -3710 9502
rect -2890 9500 1810 12808
rect 9278 12640 10226 12646
rect 9278 12122 9286 12640
rect 10220 12122 10226 12640
rect 5310 11860 7310 11902
rect 5310 11410 5316 11860
rect 7304 11410 7310 11860
rect 5310 10996 7310 11410
rect 5310 10708 5316 10996
rect 7304 10708 7310 10996
rect 2610 10396 4610 10408
rect 2610 10108 2616 10396
rect 4604 10108 4610 10396
rect 2610 9502 4610 10108
rect 5310 9502 7310 10708
rect -3770 9402 -3762 9428
rect -4230 1700 -4180 1712
rect -3768 1712 -3762 9402
rect -3728 9402 -3710 9428
rect -2850 9440 -2810 9500
rect -1930 9440 -1890 9500
rect -1010 9440 -970 9500
rect -90 9440 -50 9500
rect -2850 9428 -2802 9440
rect -2850 9422 -2842 9428
rect -3728 1712 -3722 9402
rect -3768 1700 -3722 1712
rect -2848 1712 -2842 9422
rect -2808 1712 -2802 9428
rect -2848 1700 -2802 1712
rect -2390 9428 -2344 9440
rect -2390 1712 -2384 9428
rect -2350 1712 -2344 9428
rect -2390 1700 -2344 1712
rect -1932 9428 -1886 9440
rect -1932 1712 -1926 9428
rect -1892 1712 -1886 9428
rect -1932 1700 -1886 1712
rect -1474 9428 -1428 9440
rect -1474 1712 -1468 9428
rect -1434 1712 -1428 9428
rect -1474 1700 -1428 1712
rect -1016 9428 -970 9440
rect -1016 1712 -1010 9428
rect -976 1712 -970 9428
rect -1016 1700 -970 1712
rect -558 9428 -512 9440
rect -558 1712 -552 9428
rect -518 1722 -512 9428
rect -100 9428 -50 9440
rect -518 1712 -510 1722
rect -558 1700 -510 1712
rect -100 1712 -94 9428
rect -60 9402 -50 9428
rect 358 9428 404 9440
rect -60 1712 -54 9402
rect 358 1722 364 9428
rect -100 1700 -54 1712
rect 350 1712 364 1722
rect 398 1712 404 9428
rect 810 9428 870 9500
rect 810 9402 822 9428
rect 350 1700 404 1712
rect 816 1712 822 9402
rect 856 9402 870 9428
rect 1274 9428 1320 9440
rect 856 1712 862 9402
rect 1274 1722 1280 9428
rect 816 1700 862 1712
rect 1270 1712 1280 1722
rect 1314 1712 1320 9428
rect 1730 9428 1790 9500
rect 1730 9402 1738 9428
rect 1270 1700 1320 1712
rect 1732 1712 1738 9402
rect 1772 9402 1790 9428
rect 2650 9440 2690 9502
rect 3570 9440 3610 9502
rect 4490 9440 4530 9502
rect 2650 9428 2698 9440
rect 2650 9402 2658 9428
rect 1772 1712 1778 9402
rect 1732 1700 1778 1712
rect 2652 1712 2658 9402
rect 2692 1712 2698 9428
rect 2652 1700 2698 1712
rect 3110 9428 3156 9440
rect 3110 1712 3116 9428
rect 3150 1712 3156 9428
rect 3110 1700 3156 1712
rect 3568 9428 3614 9440
rect 3568 1712 3574 9428
rect 3608 1712 3614 9428
rect 3568 1700 3614 1712
rect 4026 9428 4072 9440
rect 4026 1712 4032 9428
rect 4066 1712 4072 9428
rect 4026 1700 4072 1712
rect 4484 9428 4530 9440
rect 4484 1712 4490 9428
rect 4524 1712 4530 9428
rect 4484 1700 4530 1712
rect 4942 9428 4988 9440
rect 4942 1712 4948 9428
rect 4982 1722 4988 9428
rect 5390 9428 5450 9502
rect 5390 9402 5406 9428
rect 4982 1712 4990 1722
rect 4942 1700 4990 1712
rect 5400 1712 5406 9402
rect 5440 9402 5450 9428
rect 5858 9428 5904 9440
rect 5440 1712 5446 9402
rect 5858 1722 5864 9428
rect 5400 1700 5446 1712
rect 5850 1712 5864 1722
rect 5898 1712 5904 9428
rect 6310 9428 6370 9502
rect 7230 9440 7270 9502
rect 6310 9422 6322 9428
rect 5850 1700 5904 1712
rect 6316 1712 6322 9422
rect 6356 9422 6370 9428
rect 6774 9428 6820 9440
rect 6356 1712 6362 9422
rect 6774 1722 6780 9428
rect 6316 1700 6362 1712
rect 6770 1712 6780 1722
rect 6814 1712 6820 9428
rect 7230 9428 7278 9440
rect 7230 9422 7238 9428
rect 6770 1700 6820 1712
rect 7232 1712 7238 9422
rect 7272 1712 7278 9428
rect -8806 1659 -8658 1660
rect -8466 1659 -8348 1660
rect -8190 1659 -8010 1662
rect -8806 1653 -8348 1659
rect -8806 1619 -8646 1653
rect -8462 1619 -8348 1653
rect -18930 1244 -18924 1358
rect -18730 1244 -18724 1358
rect -18930 1238 -18724 1244
rect -18054 1352 -17982 1362
rect -18054 1248 -18044 1352
rect -17992 1248 -17982 1352
rect -18054 1238 -17982 1248
rect -17482 1352 -17410 1362
rect -17482 1248 -17472 1352
rect -17420 1248 -17410 1352
rect -17482 1238 -17410 1248
rect -16910 1352 -16838 1362
rect -16910 1248 -16900 1352
rect -16848 1248 -16838 1352
rect -12906 1352 -12834 1362
rect -16910 1238 -16838 1248
rect -15680 1296 -13226 1312
rect -15680 1196 -15668 1296
rect -13326 1196 -13226 1296
rect -12906 1248 -12896 1352
rect -12844 1248 -12834 1352
rect -12906 1238 -12834 1248
rect -12334 1352 -12262 1362
rect -12334 1248 -12324 1352
rect -12272 1248 -12262 1352
rect -12334 1238 -12262 1248
rect -11762 1352 -11690 1362
rect -11762 1248 -11752 1352
rect -11700 1248 -11690 1352
rect -8806 1302 -8348 1619
rect -8200 1653 -7992 1659
rect -8200 1619 -8188 1653
rect -8004 1619 -7992 1653
rect -8200 1613 -7992 1619
rect -8190 1522 -8010 1613
rect -8190 1402 -8170 1522
rect -8030 1402 -8010 1522
rect -8190 1382 -8010 1402
rect -7890 1342 -7850 1700
rect -7730 1659 -7550 1662
rect -7270 1659 -7090 1662
rect -7742 1653 -7534 1659
rect -7742 1619 -7730 1653
rect -7546 1619 -7534 1653
rect -7742 1613 -7534 1619
rect -7284 1653 -7076 1659
rect -7284 1619 -7272 1653
rect -7088 1619 -7076 1653
rect -7284 1613 -7076 1619
rect -7730 1522 -7550 1613
rect -7730 1402 -7710 1522
rect -7570 1402 -7550 1522
rect -7730 1382 -7550 1402
rect -7270 1522 -7090 1613
rect -7270 1402 -7250 1522
rect -7110 1402 -7090 1522
rect -7270 1382 -7090 1402
rect -6970 1342 -6930 1700
rect -6810 1659 -6630 1662
rect -6350 1659 -6170 1662
rect -6826 1653 -6618 1659
rect -6826 1619 -6814 1653
rect -6630 1619 -6618 1653
rect -6826 1613 -6618 1619
rect -6368 1653 -6160 1659
rect -6368 1619 -6356 1653
rect -6172 1619 -6160 1653
rect -6368 1613 -6160 1619
rect -6810 1522 -6630 1613
rect -6810 1402 -6790 1522
rect -6650 1402 -6630 1522
rect -6810 1382 -6630 1402
rect -6350 1522 -6170 1613
rect -6350 1402 -6330 1522
rect -6190 1402 -6170 1522
rect -6350 1382 -6170 1402
rect -6050 1342 -6010 1700
rect -5890 1659 -5710 1662
rect -5430 1659 -5250 1662
rect -5910 1653 -5702 1659
rect -5910 1619 -5898 1653
rect -5714 1619 -5702 1653
rect -5910 1613 -5702 1619
rect -5452 1653 -5244 1659
rect -5452 1619 -5440 1653
rect -5256 1619 -5244 1653
rect -5452 1613 -5244 1619
rect -5890 1522 -5710 1613
rect -5890 1402 -5870 1522
rect -5730 1402 -5710 1522
rect -5890 1382 -5710 1402
rect -5430 1522 -5250 1613
rect -5430 1402 -5410 1522
rect -5270 1402 -5250 1522
rect -5430 1382 -5250 1402
rect -5150 1342 -5110 1700
rect -4970 1659 -4790 1662
rect -4510 1659 -4330 1662
rect -4994 1653 -4786 1659
rect -4994 1619 -4982 1653
rect -4798 1619 -4786 1653
rect -4994 1613 -4786 1619
rect -4536 1653 -4328 1659
rect -4536 1619 -4524 1653
rect -4340 1619 -4328 1653
rect -4536 1613 -4328 1619
rect -4970 1522 -4790 1613
rect -4970 1402 -4950 1522
rect -4810 1402 -4790 1522
rect -4970 1382 -4790 1402
rect -4510 1522 -4330 1613
rect -4510 1402 -4490 1522
rect -4350 1402 -4330 1522
rect -4510 1382 -4330 1402
rect -4230 1342 -4190 1700
rect -4050 1659 -3870 1662
rect -2690 1659 -2510 1662
rect -4078 1653 -3870 1659
rect -4078 1619 -4066 1653
rect -3882 1619 -3870 1653
rect -4078 1613 -3870 1619
rect -2700 1653 -2492 1659
rect -2700 1619 -2688 1653
rect -2504 1619 -2492 1653
rect -2700 1613 -2492 1619
rect -4050 1522 -3870 1613
rect -4050 1402 -4030 1522
rect -3890 1402 -3870 1522
rect -4050 1382 -3870 1402
rect -2690 1522 -2510 1613
rect -2690 1402 -2670 1522
rect -2530 1402 -2510 1522
rect -2690 1382 -2510 1402
rect -2390 1342 -2350 1700
rect -2230 1659 -2050 1662
rect -1770 1659 -1590 1662
rect -2242 1653 -2034 1659
rect -2242 1619 -2230 1653
rect -2046 1619 -2034 1653
rect -2242 1613 -2034 1619
rect -1784 1653 -1576 1659
rect -1784 1619 -1772 1653
rect -1588 1619 -1576 1653
rect -1784 1613 -1576 1619
rect -2230 1522 -2050 1613
rect -2230 1402 -2210 1522
rect -2070 1402 -2050 1522
rect -2230 1382 -2050 1402
rect -1770 1522 -1590 1613
rect -1770 1402 -1750 1522
rect -1610 1402 -1590 1522
rect -1770 1382 -1590 1402
rect -1470 1342 -1430 1700
rect -1310 1659 -1130 1662
rect -850 1659 -670 1662
rect -1326 1653 -1118 1659
rect -1326 1619 -1314 1653
rect -1130 1619 -1118 1653
rect -1326 1613 -1118 1619
rect -868 1653 -660 1659
rect -868 1619 -856 1653
rect -672 1619 -660 1653
rect -868 1613 -660 1619
rect -1310 1522 -1130 1613
rect -1310 1402 -1290 1522
rect -1150 1402 -1130 1522
rect -1310 1382 -1130 1402
rect -850 1522 -670 1613
rect -850 1402 -830 1522
rect -690 1402 -670 1522
rect -850 1382 -670 1402
rect -550 1342 -510 1700
rect -390 1659 -210 1662
rect 70 1659 250 1662
rect -410 1653 -202 1659
rect -410 1619 -398 1653
rect -214 1619 -202 1653
rect -410 1613 -202 1619
rect 48 1653 256 1659
rect 48 1619 60 1653
rect 244 1619 256 1653
rect 48 1613 256 1619
rect -390 1522 -210 1613
rect -390 1402 -370 1522
rect -230 1402 -210 1522
rect -390 1382 -210 1402
rect 70 1522 250 1613
rect 70 1402 90 1522
rect 230 1402 250 1522
rect 70 1382 250 1402
rect 350 1342 390 1700
rect 530 1659 710 1662
rect 990 1659 1170 1662
rect 506 1653 714 1659
rect 506 1619 518 1653
rect 702 1619 714 1653
rect 506 1613 714 1619
rect 964 1653 1172 1659
rect 964 1619 976 1653
rect 1160 1619 1172 1653
rect 964 1613 1172 1619
rect 530 1522 710 1613
rect 530 1402 550 1522
rect 690 1402 710 1522
rect 530 1382 710 1402
rect 990 1522 1170 1613
rect 990 1402 1010 1522
rect 1150 1402 1170 1522
rect 990 1382 1170 1402
rect 1270 1342 1310 1700
rect 1450 1659 1630 1662
rect 2810 1659 2990 1662
rect 1422 1653 1630 1659
rect 1422 1619 1434 1653
rect 1618 1619 1630 1653
rect 1422 1613 1630 1619
rect 2800 1653 3008 1659
rect 2800 1619 2812 1653
rect 2996 1619 3008 1653
rect 2800 1613 3008 1619
rect 1450 1522 1630 1613
rect 1450 1402 1470 1522
rect 1610 1402 1630 1522
rect 1450 1382 1630 1402
rect 2810 1522 2990 1613
rect 2810 1402 2830 1522
rect 2970 1402 2990 1522
rect 2810 1382 2990 1402
rect 3110 1342 3150 1700
rect 3270 1659 3450 1662
rect 3730 1659 3910 1662
rect 3258 1653 3466 1659
rect 3258 1619 3270 1653
rect 3454 1619 3466 1653
rect 3258 1613 3466 1619
rect 3716 1653 3924 1659
rect 3716 1619 3728 1653
rect 3912 1619 3924 1653
rect 3716 1613 3924 1619
rect 3270 1522 3450 1613
rect 3270 1402 3290 1522
rect 3430 1402 3450 1522
rect 3270 1382 3450 1402
rect 3730 1522 3910 1613
rect 3730 1402 3750 1522
rect 3890 1402 3910 1522
rect 3730 1382 3910 1402
rect 4030 1342 4070 1700
rect 4190 1659 4370 1662
rect 4650 1659 4830 1662
rect 4174 1653 4382 1659
rect 4174 1619 4186 1653
rect 4370 1619 4382 1653
rect 4174 1613 4382 1619
rect 4632 1653 4840 1659
rect 4632 1619 4644 1653
rect 4828 1619 4840 1653
rect 4632 1613 4840 1619
rect 4190 1522 4370 1613
rect 4190 1402 4210 1522
rect 4350 1402 4370 1522
rect 4190 1382 4370 1402
rect 4650 1522 4830 1613
rect 4650 1402 4670 1522
rect 4810 1402 4830 1522
rect 4650 1382 4830 1402
rect 4950 1342 4990 1700
rect 5110 1659 5290 1662
rect 5570 1659 5750 1662
rect 5090 1653 5298 1659
rect 5090 1619 5102 1653
rect 5286 1619 5298 1653
rect 5090 1613 5298 1619
rect 5548 1653 5756 1659
rect 5548 1619 5560 1653
rect 5744 1619 5756 1653
rect 5548 1613 5756 1619
rect 5110 1522 5290 1613
rect 5110 1402 5130 1522
rect 5270 1402 5290 1522
rect 5110 1382 5290 1402
rect 5570 1522 5750 1613
rect 5570 1402 5590 1522
rect 5730 1402 5750 1522
rect 5570 1382 5750 1402
rect 5850 1342 5890 1700
rect 6030 1659 6210 1662
rect 6490 1659 6670 1662
rect 6006 1653 6214 1659
rect 6006 1619 6018 1653
rect 6202 1619 6214 1653
rect 6006 1613 6214 1619
rect 6464 1653 6672 1659
rect 6464 1619 6476 1653
rect 6660 1619 6672 1653
rect 6464 1613 6672 1619
rect 6030 1522 6210 1613
rect 6030 1402 6050 1522
rect 6190 1402 6210 1522
rect 6030 1382 6210 1402
rect 6490 1522 6670 1613
rect 6490 1402 6510 1522
rect 6650 1402 6670 1522
rect 6490 1382 6670 1402
rect 6770 1342 6810 1700
rect 7232 1696 7278 1712
rect 7690 9428 7736 9440
rect 7690 1712 7696 9428
rect 7730 1712 7736 9428
rect 9278 3162 10226 12122
rect 10622 11860 11326 14498
rect 10622 11410 10628 11860
rect 11320 11410 11326 11860
rect 10622 8072 11326 11410
rect 11440 15190 12144 15196
rect 11440 14498 11446 15190
rect 12138 14498 12144 15190
rect 12340 15179 12902 15185
rect 12340 14782 12352 15179
rect 12890 14782 12902 15179
rect 12340 14776 12902 14782
rect 11440 10396 12144 14498
rect 11440 10108 11448 10396
rect 12138 10108 12144 10396
rect 11440 10102 12144 10108
rect 10622 7380 10628 8072
rect 11320 7380 11326 8072
rect 10622 7372 11326 7380
rect 9278 2226 9284 3162
rect 10220 2226 10226 3162
rect 9278 2220 10226 2226
rect 6950 1659 7130 1662
rect 7690 1660 7736 1712
rect 6922 1653 7130 1659
rect 6922 1619 6934 1653
rect 7118 1619 7130 1653
rect 6922 1613 7130 1619
rect 6950 1522 7130 1613
rect 6950 1402 6970 1522
rect 7110 1402 7130 1522
rect 6950 1382 7130 1402
rect 7278 1653 7736 1660
rect 7278 1619 7392 1653
rect 7576 1619 7736 1653
rect -11762 1238 -11690 1248
rect -15680 1180 -13226 1196
rect -9500 1202 -8348 1302
rect -7930 1322 -7810 1342
rect -7930 1242 -7910 1322
rect -7830 1242 -7810 1322
rect -7930 1222 -7810 1242
rect -7010 1322 -6890 1342
rect -7010 1242 -6990 1322
rect -6910 1242 -6890 1322
rect -7010 1222 -6890 1242
rect -6090 1322 -5970 1342
rect -6090 1242 -6070 1322
rect -5990 1242 -5970 1322
rect -6090 1222 -5970 1242
rect -5170 1322 -5050 1342
rect -5170 1242 -5150 1322
rect -5070 1242 -5050 1322
rect -5170 1222 -5050 1242
rect -4250 1322 -4130 1342
rect -4250 1242 -4230 1322
rect -4150 1242 -4130 1322
rect -2430 1322 -2310 1342
rect -4250 1222 -4130 1242
rect -9500 1102 -9400 1202
rect -9000 1102 -8348 1202
rect -9500 1002 -8348 1102
rect -3590 1202 -2990 1302
rect -2430 1242 -2410 1322
rect -2330 1242 -2310 1322
rect -2430 1222 -2310 1242
rect -1510 1322 -1390 1342
rect -1510 1242 -1490 1322
rect -1410 1242 -1390 1322
rect -1510 1222 -1390 1242
rect -590 1322 -470 1342
rect -590 1242 -570 1322
rect -490 1242 -470 1322
rect -590 1222 -470 1242
rect 330 1322 450 1342
rect 330 1242 350 1322
rect 430 1242 450 1322
rect 330 1222 450 1242
rect 1250 1322 1370 1342
rect 1250 1242 1270 1322
rect 1350 1242 1370 1322
rect 3070 1322 3190 1342
rect 1250 1222 1370 1242
rect -3590 1102 -3490 1202
rect -3090 1102 -2990 1202
rect -3590 1002 -2990 1102
rect 1910 1202 2510 1302
rect 3070 1242 3090 1322
rect 3170 1242 3190 1322
rect 3070 1222 3190 1242
rect 3990 1322 4110 1342
rect 3990 1242 4010 1322
rect 4090 1242 4110 1322
rect 3990 1222 4110 1242
rect 4910 1322 5030 1342
rect 4910 1242 4930 1322
rect 5010 1242 5030 1322
rect 4910 1222 5030 1242
rect 5830 1322 5950 1342
rect 5830 1242 5850 1322
rect 5930 1242 5950 1322
rect 5830 1222 5950 1242
rect 6750 1322 6870 1342
rect 6750 1242 6770 1322
rect 6850 1242 6870 1322
rect 6750 1222 6870 1242
rect 7278 1300 7736 1619
rect 1910 1102 2010 1202
rect 2410 1102 2510 1202
rect 1910 1002 2510 1102
rect 7278 1200 8466 1300
rect 7278 1100 7966 1200
rect 8366 1100 8466 1200
rect 7278 1000 8466 1100
<< via1 >>
rect -21546 25052 -10302 25066
rect -21546 24254 -21532 25052
rect -21532 24254 -10316 25052
rect -10316 24254 -10302 25052
rect -21546 24240 -10302 24254
rect 1720 22968 2278 23526
rect 3344 22968 3902 23526
rect 7434 22968 7992 23526
rect 9888 22968 10446 23526
rect -4836 22168 -4278 22726
rect 890 22168 1448 22726
rect 4162 22168 4720 22726
rect 6616 22168 7174 22726
rect 9070 22168 9628 22726
rect 11524 22168 12082 22726
rect -4836 21976 -4278 21988
rect -4836 21579 -4826 21976
rect -4826 21579 -4288 21976
rect -4288 21579 -4278 21976
rect -4836 21568 -4278 21579
rect -4018 21976 -3460 21988
rect -4018 21579 -4008 21976
rect -4008 21579 -3470 21976
rect -3470 21579 -3460 21976
rect -4018 21568 -3460 21579
rect 72 21914 630 21926
rect 72 21517 82 21914
rect 82 21517 620 21914
rect 620 21517 630 21914
rect 72 21506 630 21517
rect 890 21914 1448 21926
rect 890 21517 900 21914
rect 900 21517 1438 21914
rect 1438 21517 1448 21914
rect 890 21506 1448 21517
rect 1708 21914 2266 21926
rect 1708 21517 1718 21914
rect 1718 21517 2256 21914
rect 2256 21517 2266 21914
rect 1708 21506 2266 21517
rect 2526 21914 3084 21926
rect 2526 21517 2536 21914
rect 2536 21517 3074 21914
rect 3074 21517 3084 21914
rect 2526 21506 3084 21517
rect 3344 21914 3902 21926
rect 3344 21517 3354 21914
rect 3354 21517 3892 21914
rect 3892 21517 3902 21914
rect 3344 21506 3902 21517
rect 4162 21914 4720 21926
rect 4162 21517 4172 21914
rect 4172 21517 4710 21914
rect 4710 21517 4720 21914
rect 4162 21506 4720 21517
rect 4980 21914 5538 21926
rect 4980 21517 4990 21914
rect 4990 21517 5528 21914
rect 5528 21517 5538 21914
rect 4980 21506 5538 21517
rect 5798 21914 6356 21926
rect 5798 21517 5808 21914
rect 5808 21517 6346 21914
rect 6346 21517 6356 21914
rect 5798 21506 6356 21517
rect 6616 21914 7174 21926
rect 6616 21517 6626 21914
rect 6626 21517 7164 21914
rect 7164 21517 7174 21914
rect 6616 21506 7174 21517
rect 7434 21914 7992 21926
rect 7434 21517 7444 21914
rect 7444 21517 7982 21914
rect 7982 21517 7992 21914
rect 7434 21506 7992 21517
rect 8252 21914 8810 21926
rect 8252 21517 8262 21914
rect 8262 21517 8800 21914
rect 8800 21517 8810 21914
rect 8252 21506 8810 21517
rect 9070 21914 9628 21926
rect 9070 21517 9080 21914
rect 9080 21517 9618 21914
rect 9618 21517 9628 21914
rect 9070 21506 9628 21517
rect 9888 21914 10446 21926
rect 9888 21517 9898 21914
rect 9898 21517 10436 21914
rect 10436 21517 10446 21914
rect 9888 21506 10446 21517
rect 10706 21914 11264 21926
rect 10706 21517 10716 21914
rect 10716 21517 11254 21914
rect 11254 21517 11264 21914
rect 10706 21506 11264 21517
rect 11524 21914 12082 21926
rect 11524 21517 11534 21914
rect 11534 21517 12072 21914
rect 12072 21517 12082 21914
rect 11524 21506 12082 21517
rect -4018 20772 -3460 21264
rect 72 20706 630 21264
rect 2526 20706 3084 21264
rect 4980 20706 5538 21264
rect 8252 20706 8810 21264
rect 10706 20706 11264 21264
rect 890 16232 1448 16790
rect 4162 16232 4720 16790
rect 6616 16232 7174 16790
rect 9070 16232 9628 16790
rect 1708 15432 2266 15990
rect 3344 15432 3902 15990
rect 7434 15432 7992 15990
rect 72 15179 630 15190
rect 72 14781 82 15179
rect 82 14781 620 15179
rect 620 14781 630 15179
rect 72 14770 630 14781
rect 890 15179 1448 15190
rect 890 14782 900 15179
rect 900 14782 1438 15179
rect 1438 14782 1448 15179
rect 890 14770 1448 14782
rect 1708 15179 2266 15190
rect 1708 14782 1718 15179
rect 1718 14782 2256 15179
rect 2256 14782 2266 15179
rect 1708 14770 2266 14782
rect 2526 15179 3084 15190
rect 2526 14781 2536 15179
rect 2536 14781 3074 15179
rect 3074 14781 3084 15179
rect 2526 14770 3084 14781
rect 3344 15179 3902 15190
rect 3344 14782 3354 15179
rect 3354 14782 3892 15179
rect 3892 14782 3902 15179
rect 3344 14770 3902 14782
rect 4162 15179 4720 15190
rect 4162 14782 4172 15179
rect 4172 14782 4710 15179
rect 4710 14782 4720 15179
rect 4162 14770 4720 14782
rect 4980 15179 5538 15190
rect 4980 14781 4990 15179
rect 4990 14781 5528 15179
rect 5528 14781 5538 15179
rect 4980 14770 5538 14781
rect 5798 15179 6356 15190
rect 5798 15158 5808 15179
rect 5720 14782 5808 15158
rect 5808 14782 6346 15179
rect 6346 15158 6356 15179
rect 6346 14782 6412 15158
rect 5720 14640 6412 14782
rect 6616 15179 7174 15190
rect 6616 14782 6626 15179
rect 6626 14782 7164 15179
rect 7164 14782 7174 15179
rect 6616 14770 7174 14782
rect 7434 15179 7992 15190
rect 7434 14782 7444 15179
rect 7444 14782 7982 15179
rect 7982 14782 7992 15179
rect 7434 14770 7992 14782
rect 8252 15179 8810 15190
rect 8252 14781 8262 15179
rect 8262 14781 8800 15179
rect 8800 14781 8810 15179
rect 8252 14770 8810 14781
rect 9070 15179 9628 15190
rect 9070 14782 9080 15179
rect 9080 14782 9618 15179
rect 9618 14782 9628 15179
rect 9070 14770 9628 14782
rect 72 13970 630 14528
rect 2526 13970 3084 14528
rect 4980 13970 5538 14528
rect 8252 13970 8810 14528
rect 9810 15179 10502 15190
rect 9810 14782 9898 15179
rect 9898 14782 10436 15179
rect 10436 14782 10502 15179
rect 9810 14498 10502 14782
rect 10628 15179 11320 15190
rect 10628 14782 10716 15179
rect 10716 14782 11254 15179
rect 11254 14782 11320 15179
rect 10628 14498 11320 14782
rect -8384 11410 -6396 11860
rect -9902 10690 -9782 11104
rect -10358 10106 -10238 10398
rect -21364 4944 -21312 4996
rect -19530 4950 -19478 5002
rect -18924 4944 -18730 5002
rect -20446 4738 -20394 4790
rect -19240 1448 -19188 1552
rect -15564 6932 -15420 6986
rect -16136 6792 -15992 6846
rect -14420 6932 -14276 6986
rect -14992 6792 -14848 6846
rect -13276 6932 -13132 6986
rect -13848 6792 -13704 6846
rect -17768 4376 -17716 4630
rect -17208 4376 -17156 4630
rect -16648 4376 -16596 4630
rect -15868 4676 -15816 4780
rect -15296 4676 -15244 4780
rect -15748 4376 -15696 4630
rect -16170 4323 -15962 4340
rect -16170 4289 -16166 4323
rect -16166 4289 -15982 4323
rect -15982 4289 -15962 4323
rect -16170 4282 -15962 4289
rect -15598 4323 -15390 4336
rect -15598 4289 -15594 4323
rect -15594 4289 -15410 4323
rect -15410 4289 -15390 4323
rect -15598 4278 -15390 4289
rect -14724 4676 -14672 4780
rect -14152 4676 -14100 4780
rect -14604 4376 -14552 4630
rect -15026 4323 -14818 4340
rect -15026 4289 -15022 4323
rect -15022 4289 -14838 4323
rect -14838 4289 -14818 4323
rect -15026 4282 -14818 4289
rect -14454 4323 -14246 4340
rect -14454 4289 -14450 4323
rect -14450 4289 -14266 4323
rect -14266 4289 -14246 4323
rect -14454 4282 -14246 4289
rect -13580 4676 -13528 4780
rect -13008 4676 -12956 4780
rect -13460 4376 -13408 4630
rect -12660 4376 -12608 4630
rect -13882 4323 -13674 4340
rect -13882 4289 -13878 4323
rect -13878 4289 -13694 4323
rect -13694 4289 -13674 4323
rect -13882 4282 -13674 4289
rect -13310 4323 -13102 4340
rect -13310 4289 -13306 4323
rect -13306 4289 -13122 4323
rect -13122 4289 -13102 4323
rect -13310 4282 -13102 4289
rect -12100 4376 -12048 4630
rect -8384 10708 -6396 10996
rect -5684 10108 -3696 10396
rect -9902 6926 -9782 7006
rect -10358 6786 -10248 6866
rect -11540 4376 -11488 4630
rect -9490 4376 -9022 4630
rect -18618 1448 -18566 1552
rect -18160 1448 -18108 1552
rect -17584 1448 -17532 1552
rect -17012 1448 -16960 1552
rect -16440 1448 -16388 1552
rect -15868 1448 -15816 1552
rect -15296 1448 -15244 1552
rect -14724 1448 -14672 1552
rect -14152 1448 -14100 1552
rect -13580 1448 -13528 1552
rect -13008 1448 -12956 1552
rect -12436 1448 -12384 1552
rect -11864 1448 -11812 1552
rect -11292 1448 -11240 1552
rect -11182 1448 -11130 1552
rect -10724 1448 -10672 1552
rect -10112 1448 -10060 1552
rect -9490 1388 -9022 1536
rect 9286 12122 10220 12640
rect 5316 11410 7304 11860
rect 5316 10708 7304 10996
rect 2616 10108 4604 10396
rect -18924 1244 -18730 1358
rect -18044 1248 -17992 1352
rect -17472 1248 -17420 1352
rect -16900 1248 -16848 1352
rect -12896 1248 -12844 1352
rect -12324 1248 -12272 1352
rect -11752 1248 -11700 1352
rect -8170 1402 -8030 1522
rect -7710 1402 -7570 1522
rect -7250 1402 -7110 1522
rect -6790 1402 -6650 1522
rect -6330 1402 -6190 1522
rect -5870 1402 -5730 1522
rect -5410 1402 -5270 1522
rect -4950 1402 -4810 1522
rect -4490 1402 -4350 1522
rect -4030 1402 -3890 1522
rect -2670 1402 -2530 1522
rect -2210 1402 -2070 1522
rect -1750 1402 -1610 1522
rect -1290 1402 -1150 1522
rect -830 1402 -690 1522
rect -370 1402 -230 1522
rect 90 1402 230 1522
rect 550 1402 690 1522
rect 1010 1402 1150 1522
rect 1470 1402 1610 1522
rect 2830 1402 2970 1522
rect 3290 1402 3430 1522
rect 3750 1402 3890 1522
rect 4210 1402 4350 1522
rect 4670 1402 4810 1522
rect 5130 1402 5270 1522
rect 5590 1402 5730 1522
rect 6050 1402 6190 1522
rect 6510 1402 6650 1522
rect 10628 11410 11320 11860
rect 11446 15179 12138 15190
rect 11446 14782 11534 15179
rect 11534 14782 12072 15179
rect 12072 14782 12138 15179
rect 11446 14498 12138 14782
rect 11448 10108 12138 10396
rect 10628 7380 11320 8072
rect 9284 2226 10220 3162
rect 6970 1402 7110 1522
rect -7910 1242 -7830 1322
rect -6990 1242 -6910 1322
rect -6070 1242 -5990 1322
rect -5150 1242 -5070 1322
rect -4230 1242 -4150 1322
rect -9400 1102 -9000 1202
rect -2410 1242 -2330 1322
rect -1490 1242 -1410 1322
rect -570 1242 -490 1322
rect 350 1242 430 1322
rect 1270 1242 1350 1322
rect -3490 1102 -3090 1202
rect 3090 1242 3170 1322
rect 4010 1242 4090 1322
rect 4930 1242 5010 1322
rect 5850 1242 5930 1322
rect 6770 1242 6850 1322
rect 2010 1102 2410 1202
rect 7966 1100 8366 1200
<< metal2 >>
rect -21561 25072 -10287 25081
rect -21561 24234 -21552 25072
rect -10296 24234 -10287 25072
rect -21561 24225 -10287 24234
rect 1714 23526 2284 23532
rect 1714 22968 1720 23526
rect 2278 22968 2284 23526
rect -4842 22726 -4272 22732
rect -4842 22168 -4836 22726
rect -4278 22168 -4272 22726
rect -4842 21988 -4272 22168
rect 884 22726 1454 22732
rect 884 22168 890 22726
rect 1448 22168 1454 22726
rect -4842 21568 -4836 21988
rect -4278 21568 -4272 21988
rect -4842 21562 -4272 21568
rect -4024 21988 -3454 21994
rect -4024 21568 -4018 21988
rect -3460 21568 -3454 21988
rect -4024 21264 -3454 21568
rect -4024 20772 -4018 21264
rect -3460 20772 -3454 21264
rect -4024 20762 -3454 20772
rect 66 21926 636 21932
rect 66 21506 72 21926
rect 630 21506 636 21926
rect 66 21264 636 21506
rect 884 21926 1454 22168
rect 1714 21932 2284 22968
rect 3338 23526 3908 23532
rect 3338 22968 3344 23526
rect 3902 22968 3908 23526
rect 884 21506 890 21926
rect 1448 21506 1454 21926
rect 884 21500 1454 21506
rect 1702 21926 2284 21932
rect 1702 21506 1708 21926
rect 2266 21518 2284 21926
rect 2520 21926 3090 21932
rect 2266 21506 2272 21518
rect 1702 21500 2272 21506
rect 2520 21506 2526 21926
rect 3084 21506 3090 21926
rect 66 20706 72 21264
rect 630 20706 636 21264
rect 66 20700 636 20706
rect 2520 21264 3090 21506
rect 3338 21926 3908 22968
rect 7428 23526 7998 23532
rect 7428 22968 7434 23526
rect 7992 22968 7998 23526
rect 3338 21506 3344 21926
rect 3902 21506 3908 21926
rect 3338 21500 3908 21506
rect 4156 22726 4726 22732
rect 4156 22168 4162 22726
rect 4720 22168 4726 22726
rect 4156 21926 4726 22168
rect 6610 22726 7180 22732
rect 6610 22168 6616 22726
rect 7174 22168 7180 22726
rect 4156 21506 4162 21926
rect 4720 21506 4726 21926
rect 4156 21500 4726 21506
rect 4974 21926 5544 21932
rect 4974 21506 4980 21926
rect 5538 21506 5544 21926
rect 2520 20706 2526 21264
rect 3084 20706 3090 21264
rect 2520 20700 3090 20706
rect 4974 21264 5544 21506
rect 4974 20706 4980 21264
rect 5538 20706 5544 21264
rect 4974 20700 5544 20706
rect 5792 21926 6362 21932
rect 5792 21506 5798 21926
rect 6356 21506 6362 21926
rect 5792 19070 6362 21506
rect 6610 21926 7180 22168
rect 6610 21506 6616 21926
rect 7174 21506 7180 21926
rect 6610 21500 7180 21506
rect 7428 21926 7998 22968
rect 9888 23526 10452 23532
rect 10446 22968 10452 23526
rect 9888 22962 10452 22968
rect 9064 22726 9634 22732
rect 9064 22168 9070 22726
rect 9628 22168 9634 22726
rect 7428 21506 7434 21926
rect 7992 21506 7998 21926
rect 7428 21500 7998 21506
rect 8246 21926 8816 21932
rect 8246 21506 8252 21926
rect 8810 21506 8816 21926
rect 8246 21264 8816 21506
rect 9064 21926 9634 22168
rect 9064 21506 9070 21926
rect 9628 21506 9634 21926
rect 9064 21500 9634 21506
rect 9882 21926 10452 22962
rect 11518 22726 12088 22732
rect 11518 22168 11524 22726
rect 12082 22168 12088 22726
rect 9882 21506 9888 21926
rect 10446 21506 10452 21926
rect 9882 21500 10452 21506
rect 10700 21926 11270 21932
rect 10700 21506 10706 21926
rect 11264 21506 11270 21926
rect 8246 20706 8252 21264
rect 8810 20706 8816 21264
rect 8246 20700 8816 20706
rect 10700 21264 11270 21506
rect 11518 21926 12088 22168
rect 11518 21506 11524 21926
rect 12082 21506 12088 21926
rect 11518 21500 12088 21506
rect 10700 20706 10706 21264
rect 11264 20706 11270 21264
rect 10700 20700 11270 20706
rect 5792 18500 12076 19070
rect 884 16790 1454 16796
rect 884 16232 890 16790
rect 1448 16232 1454 16790
rect 66 15190 636 15196
rect 66 14770 72 15190
rect 630 14770 636 15190
rect 66 14528 636 14770
rect 884 15190 1454 16232
rect 4156 16790 4726 16796
rect 4156 16232 4162 16790
rect 4720 16232 4726 16790
rect 884 14770 890 15190
rect 1448 14770 1454 15190
rect 884 14764 1454 14770
rect 1702 15990 2272 15996
rect 1702 15432 1708 15990
rect 2266 15432 2272 15990
rect 1702 15190 2272 15432
rect 3338 15990 3908 15996
rect 3338 15432 3344 15990
rect 3902 15432 3908 15990
rect 1702 14770 1708 15190
rect 2266 14770 2272 15190
rect 1702 14764 2272 14770
rect 2520 15190 3090 15196
rect 2520 14770 2526 15190
rect 3084 14770 3090 15190
rect 66 13970 72 14528
rect 630 13970 636 14528
rect 2520 14528 3090 14770
rect 3338 15190 3908 15432
rect 3338 14770 3344 15190
rect 3902 14770 3908 15190
rect 3338 14764 3908 14770
rect 4156 15190 4726 16232
rect 6610 16790 7180 16796
rect 6610 16232 6616 16790
rect 7174 16232 7180 16790
rect 4156 14770 4162 15190
rect 4720 14770 4726 15190
rect 4156 14764 4726 14770
rect 4974 15190 5544 15196
rect 4974 14770 4980 15190
rect 5538 14770 5544 15190
rect 5792 15190 6362 15196
rect 5792 15158 5798 15190
rect 6356 15158 6362 15190
rect 6610 15190 7180 16232
rect 9064 16790 9634 16796
rect 9064 16232 9070 16790
rect 9628 16232 9634 16790
rect 2520 13970 2526 14528
rect 3084 13970 3090 14528
rect 4974 14528 5544 14770
rect 4974 13970 4980 14528
rect 5538 13970 5544 14528
rect 5714 14640 5720 15158
rect 6412 14640 6418 15158
rect 6610 14770 6616 15190
rect 7174 14770 7180 15190
rect 6610 14764 7180 14770
rect 7428 15990 7998 15996
rect 7428 15432 7434 15990
rect 7992 15432 7998 15990
rect 7428 15190 7998 15432
rect 7428 14770 7434 15190
rect 7992 14770 7998 15190
rect 7428 14764 7998 14770
rect 8246 15190 8816 15196
rect 8246 14770 8252 15190
rect 8810 14770 8816 15190
rect 66 13964 630 13970
rect 2520 13964 3084 13970
rect 4974 13964 5538 13970
rect 5714 13892 6418 14640
rect 8246 14528 8816 14770
rect 9064 15190 9634 16232
rect 11506 15196 12076 18500
rect 9064 14770 9070 15190
rect 9628 14770 9634 15190
rect 9064 14764 9634 14770
rect 9804 15190 10508 15196
rect 8246 13970 8252 14528
rect 8810 13970 8816 14528
rect 9804 14498 9810 15190
rect 10502 14498 10508 15190
rect 10622 15190 11326 15196
rect 10622 14498 10628 15190
rect 11320 14498 11326 15190
rect 11440 15190 12144 15196
rect 11440 14498 11446 15190
rect 12138 14498 12144 15190
rect 9804 14492 10508 14498
rect 11440 14492 12144 14498
rect 8246 13964 8816 13970
rect 5714 12646 6416 13892
rect 5714 12640 10226 12646
rect 5714 12122 9286 12640
rect 10220 12122 10226 12640
rect 5714 12116 10226 12122
rect -9906 11860 11340 11868
rect -9906 11786 -8384 11860
rect -6396 11786 5316 11860
rect 7304 11786 10628 11860
rect -9906 11110 -9252 11786
rect 11320 11410 11340 11860
rect -9908 11104 -9252 11110
rect -9908 10690 -9902 11104
rect -9782 10802 -9252 11104
rect 11070 10802 11340 11410
rect -9782 10708 -8384 10802
rect -6396 10708 5316 10802
rect 7304 10708 11340 10802
rect -9782 10690 11340 10708
rect -9908 10686 11340 10690
rect -9908 10684 -9776 10686
rect -10364 10398 12144 10402
rect -10364 10106 -10358 10398
rect -10238 10396 12144 10398
rect -10238 10108 -5684 10396
rect -3696 10108 2616 10396
rect 4604 10108 11448 10396
rect 12138 10108 12144 10396
rect -10238 10106 12144 10108
rect -10364 9802 12144 10106
rect 10622 8072 12682 8078
rect 10622 7380 10628 8072
rect 11320 7380 12682 8072
rect 10622 7374 12682 7380
rect -15584 6986 -9902 7006
rect -15584 6932 -15564 6986
rect -15420 6932 -14420 6986
rect -14276 6932 -13276 6986
rect -13132 6932 -9902 6986
rect -15584 6926 -9902 6932
rect -9782 6926 -9776 7006
rect -16156 6846 -10358 6866
rect -16156 6792 -16136 6846
rect -15992 6792 -14992 6846
rect -14848 6792 -13848 6846
rect -13704 6792 -10358 6846
rect -16156 6786 -10358 6792
rect -10248 6786 -10242 6866
rect -21370 5002 -18724 5008
rect -21370 4996 -19530 5002
rect -21370 4944 -21364 4996
rect -21312 4950 -19530 4996
rect -19478 4950 -18924 5002
rect -21312 4944 -18924 4950
rect -18730 4944 -18724 5002
rect -21370 4938 -18724 4944
rect -21317 4790 -12946 4798
rect -21317 4738 -20446 4790
rect -20394 4780 -12946 4790
rect -20394 4738 -15868 4780
rect -21317 4676 -15868 4738
rect -15816 4676 -15296 4780
rect -15244 4676 -14724 4780
rect -14672 4676 -14152 4780
rect -14100 4676 -13580 4780
rect -13528 4676 -13008 4780
rect -12956 4676 -12946 4780
rect -21317 4664 -12946 4676
rect -18620 4630 -9016 4636
rect -18620 4629 -17768 4630
rect -18620 4377 -18600 4629
rect -18000 4377 -17768 4629
rect -18620 4376 -17768 4377
rect -17716 4376 -17208 4630
rect -17156 4376 -16648 4630
rect -16596 4376 -15748 4630
rect -15696 4376 -14604 4630
rect -14552 4376 -13460 4630
rect -13408 4376 -12660 4630
rect -12608 4376 -12100 4630
rect -12048 4376 -11540 4630
rect -11488 4629 -9490 4630
rect -11488 4377 -10109 4629
rect -9509 4377 -9490 4629
rect -11488 4376 -9490 4377
rect -9022 4376 -9016 4630
rect -18620 4370 -9016 4376
rect -16176 4340 -13096 4342
rect -16176 4282 -16170 4340
rect -15962 4336 -15026 4340
rect -15962 4282 -15598 4336
rect -16176 4278 -15598 4282
rect -15390 4282 -15026 4336
rect -14818 4282 -14454 4340
rect -14246 4282 -13882 4340
rect -13674 4282 -13310 4340
rect -13102 4282 -13096 4340
rect -15390 4278 -13096 4282
rect -16176 4276 -13096 4278
rect -16176 4272 -15130 4276
rect 9278 3162 12682 3168
rect 9278 2226 9284 3162
rect 10220 2226 12682 3162
rect 9278 2220 12682 2226
rect -19268 1556 -10002 1562
rect -19268 1442 -19258 1556
rect -10012 1442 -10002 1556
rect -19268 1438 -10002 1442
rect -9496 1536 7130 1542
rect -9496 1388 -9490 1536
rect -9022 1522 7130 1536
rect -9022 1402 -8170 1522
rect -8030 1402 -7710 1522
rect -7570 1402 -7250 1522
rect -7110 1402 -6790 1522
rect -6650 1402 -6330 1522
rect -6190 1402 -5870 1522
rect -5730 1402 -5410 1522
rect -5270 1402 -4950 1522
rect -4810 1402 -4490 1522
rect -4350 1402 -4030 1522
rect -3890 1402 -2670 1522
rect -2530 1402 -2210 1522
rect -2070 1402 -1750 1522
rect -1610 1402 -1290 1522
rect -1150 1402 -830 1522
rect -690 1402 -370 1522
rect -230 1402 90 1522
rect 230 1402 550 1522
rect 690 1402 1010 1522
rect 1150 1402 1470 1522
rect 1610 1402 2830 1522
rect 2970 1402 3290 1522
rect 3430 1402 3750 1522
rect 3890 1402 4210 1522
rect 4350 1402 4670 1522
rect 4810 1402 5130 1522
rect 5270 1402 5590 1522
rect 5730 1402 6050 1522
rect 6190 1402 6510 1522
rect 6650 1402 6970 1522
rect 7110 1402 7130 1522
rect -9022 1388 7130 1402
rect -9496 1382 7130 1388
rect -18930 1362 -18724 1364
rect -18930 1358 -11690 1362
rect -18930 1244 -18924 1358
rect -18730 1352 -11690 1358
rect -18730 1248 -18044 1352
rect -17992 1248 -17472 1352
rect -17420 1248 -16900 1352
rect -16848 1248 -12896 1352
rect -12844 1248 -12324 1352
rect -12272 1248 -11752 1352
rect -11700 1248 -11690 1352
rect -7930 1334 -7810 1342
rect -7010 1334 -6890 1342
rect -6090 1334 -5970 1342
rect -5170 1334 -5050 1342
rect -4250 1334 -4130 1342
rect -2430 1334 -2310 1342
rect -1510 1334 -1390 1342
rect -590 1334 -470 1342
rect 330 1334 450 1342
rect 1250 1334 1370 1342
rect 3070 1334 3190 1342
rect 3990 1334 4110 1342
rect 4910 1334 5030 1342
rect 5830 1334 5950 1342
rect 6750 1334 6870 1342
rect -18730 1244 -11690 1248
rect -18930 1238 -11690 1244
rect -9504 1324 8454 1334
rect -9504 1006 -9494 1324
rect 8444 1300 8454 1324
rect 8444 1006 8466 1300
rect -9504 1000 8466 1006
rect -9504 998 8454 1000
<< via2 >>
rect -21552 25066 -10296 25072
rect -21552 24240 -21546 25066
rect -21546 24240 -10302 25066
rect -10302 24240 -10296 25066
rect -21552 24234 -10296 24240
rect -9252 11410 -8384 11786
rect -8384 11410 -6396 11786
rect -6396 11410 5316 11786
rect 5316 11410 7304 11786
rect 7304 11410 10628 11786
rect 10628 11410 11070 11786
rect -9252 10996 11070 11410
rect -9252 10802 -8384 10996
rect -8384 10802 -6396 10996
rect -6396 10802 5316 10996
rect 5316 10802 7304 10996
rect 7304 10802 11070 10996
rect -18600 4377 -18000 4629
rect -10109 4377 -9509 4629
rect -19258 1552 -10012 1556
rect -19258 1448 -19240 1552
rect -19240 1448 -19188 1552
rect -19188 1448 -18618 1552
rect -18618 1448 -18566 1552
rect -18566 1448 -18160 1552
rect -18160 1448 -18108 1552
rect -18108 1448 -17584 1552
rect -17584 1448 -17532 1552
rect -17532 1448 -17012 1552
rect -17012 1448 -16960 1552
rect -16960 1448 -16440 1552
rect -16440 1448 -16388 1552
rect -16388 1448 -15868 1552
rect -15868 1448 -15816 1552
rect -15816 1448 -15296 1552
rect -15296 1448 -15244 1552
rect -15244 1448 -14724 1552
rect -14724 1448 -14672 1552
rect -14672 1448 -14152 1552
rect -14152 1448 -14100 1552
rect -14100 1448 -13580 1552
rect -13580 1448 -13528 1552
rect -13528 1448 -13008 1552
rect -13008 1448 -12956 1552
rect -12956 1448 -12436 1552
rect -12436 1448 -12384 1552
rect -12384 1448 -11864 1552
rect -11864 1448 -11812 1552
rect -11812 1448 -11292 1552
rect -11292 1448 -11240 1552
rect -11240 1448 -11182 1552
rect -11182 1448 -11130 1552
rect -11130 1448 -10724 1552
rect -10724 1448 -10672 1552
rect -10672 1448 -10112 1552
rect -10112 1448 -10060 1552
rect -10060 1448 -10012 1552
rect -19258 1442 -10012 1448
rect -9494 1322 8444 1324
rect -9494 1242 -7910 1322
rect -7910 1242 -7830 1322
rect -7830 1242 -6990 1322
rect -6990 1242 -6910 1322
rect -6910 1242 -6070 1322
rect -6070 1242 -5990 1322
rect -5990 1242 -5150 1322
rect -5150 1242 -5070 1322
rect -5070 1242 -4230 1322
rect -4230 1242 -4150 1322
rect -4150 1242 -2410 1322
rect -2410 1242 -2330 1322
rect -2330 1242 -1490 1322
rect -1490 1242 -1410 1322
rect -1410 1242 -570 1322
rect -570 1242 -490 1322
rect -490 1242 350 1322
rect 350 1242 430 1322
rect 430 1242 1270 1322
rect 1270 1242 1350 1322
rect 1350 1242 3090 1322
rect 3090 1242 3170 1322
rect 3170 1242 4010 1322
rect 4010 1242 4090 1322
rect 4090 1242 4930 1322
rect 4930 1242 5010 1322
rect 5010 1242 5850 1322
rect 5850 1242 5930 1322
rect 5930 1242 6770 1322
rect 6770 1242 6850 1322
rect 6850 1242 8444 1322
rect -9494 1202 8444 1242
rect -9494 1102 -9400 1202
rect -9400 1102 -9000 1202
rect -9000 1102 -3490 1202
rect -3490 1102 -3090 1202
rect -3090 1102 2010 1202
rect 2010 1102 2410 1202
rect 2410 1200 8444 1202
rect 2410 1102 7966 1200
rect -9494 1100 7966 1102
rect 7966 1100 8366 1200
rect 8366 1100 8444 1200
rect -9494 1006 8444 1100
<< metal3 >>
rect -21567 25081 -10281 25087
rect -21567 24225 -21561 25081
rect -10287 24225 -10281 25081
rect -21567 24219 -10281 24225
rect -17888 16638 -10718 16666
rect -17888 16094 -17273 16638
rect -17209 16094 -16554 16638
rect -16490 16094 -15835 16638
rect -15771 16094 -15116 16638
rect -15052 16094 -14397 16638
rect -14333 16094 -13678 16638
rect -13614 16094 -12959 16638
rect -12895 16094 -12240 16638
rect -12176 16094 -11521 16638
rect -11457 16094 -10802 16638
rect -10738 16094 -10718 16638
rect -17888 15938 -10718 16094
rect -17888 15394 -17273 15938
rect -17209 15394 -16554 15938
rect -16490 15394 -15835 15938
rect -15771 15394 -15116 15938
rect -15052 15394 -14397 15938
rect -14333 15394 -13678 15938
rect -13614 15394 -12959 15938
rect -12895 15394 -12240 15938
rect -12176 15394 -11521 15938
rect -11457 15394 -10802 15938
rect -10738 15394 -10718 15938
rect -17888 15238 -10718 15394
rect -17888 14694 -17273 15238
rect -17209 14694 -16554 15238
rect -16490 14694 -15835 15238
rect -15771 14694 -15116 15238
rect -15052 14694 -14397 15238
rect -14333 14694 -13678 15238
rect -13614 14694 -12959 15238
rect -12895 14694 -12240 15238
rect -12176 14694 -11521 15238
rect -11457 14694 -10802 15238
rect -10738 14694 -10718 15238
rect -17888 14538 -10718 14694
rect -17888 13994 -17273 14538
rect -17209 13994 -16554 14538
rect -16490 13994 -15835 14538
rect -15771 13994 -15116 14538
rect -15052 13994 -14397 14538
rect -14333 13994 -13678 14538
rect -13614 13994 -12959 14538
rect -12895 13994 -12240 14538
rect -12176 13994 -11521 14538
rect -11457 13994 -10802 14538
rect -10738 13994 -10718 14538
rect -17888 13838 -10718 13994
rect -17888 13294 -17273 13838
rect -17209 13294 -16554 13838
rect -16490 13294 -15835 13838
rect -15771 13294 -15116 13838
rect -15052 13294 -14397 13838
rect -14333 13294 -13678 13838
rect -13614 13294 -12959 13838
rect -12895 13294 -12240 13838
rect -12176 13294 -11521 13838
rect -11457 13294 -10802 13838
rect -10738 13294 -10718 13838
rect -17888 13138 -10718 13294
rect -17888 12594 -17273 13138
rect -17209 12594 -16554 13138
rect -16490 12594 -15835 13138
rect -15771 12594 -15116 13138
rect -15052 12594 -14397 13138
rect -14333 12594 -13678 13138
rect -13614 12594 -12959 13138
rect -12895 12594 -12240 13138
rect -12176 12594 -11521 13138
rect -11457 12594 -10802 13138
rect -10738 12594 -10718 13138
rect -17888 12438 -10718 12594
rect -17888 11894 -17273 12438
rect -17209 11894 -16554 12438
rect -16490 11894 -15835 12438
rect -15771 11894 -15116 12438
rect -15052 11894 -14397 12438
rect -14333 11894 -13678 12438
rect -13614 11894 -12959 12438
rect -12895 11894 -12240 12438
rect -12176 11894 -11521 12438
rect -11457 11894 -10802 12438
rect -10738 11894 -10718 12438
rect -17888 11738 -10718 11894
rect -17888 11194 -17273 11738
rect -17209 11194 -16554 11738
rect -16490 11194 -15835 11738
rect -15771 11194 -15116 11738
rect -15052 11194 -14397 11738
rect -14333 11194 -13678 11738
rect -13614 11194 -12959 11738
rect -12895 11194 -12240 11738
rect -12176 11194 -11521 11738
rect -11457 11194 -10802 11738
rect -10738 11194 -10718 11738
rect -17888 11038 -10718 11194
rect -17888 10494 -17273 11038
rect -17209 10494 -16554 11038
rect -16490 10494 -15835 11038
rect -15771 10494 -15116 11038
rect -15052 10494 -14397 11038
rect -14333 10494 -13678 11038
rect -13614 10494 -12959 11038
rect -12895 10494 -12240 11038
rect -12176 10494 -11521 11038
rect -11457 10494 -10802 11038
rect -10738 10494 -10718 11038
rect -9257 11786 11075 11791
rect -9257 10802 -9252 11786
rect 11070 10802 11075 11786
rect -9257 10797 11075 10802
rect -17888 10338 -10718 10494
rect -17888 9794 -17273 10338
rect -17209 9794 -16554 10338
rect -16490 9794 -15835 10338
rect -15771 9794 -15116 10338
rect -15052 9794 -14397 10338
rect -14333 9794 -13678 10338
rect -13614 9794 -12959 10338
rect -12895 9794 -12240 10338
rect -12176 9794 -11521 10338
rect -11457 9794 -10802 10338
rect -10738 9794 -10718 10338
rect -18620 4643 -17980 4649
rect -18620 4363 -18614 4643
rect -17986 4363 -17980 4643
rect -18620 4357 -17980 4363
rect -17888 1562 -10718 9794
rect -10129 4643 -9489 4649
rect -10129 4363 -10123 4643
rect -9495 4363 -9489 4643
rect -10129 4357 -9489 4363
rect -19266 1556 8465 1562
rect -19266 1442 -19258 1556
rect -10012 1442 8465 1556
rect -20266 1340 8465 1442
rect -20266 1324 8466 1340
rect -20266 1006 -9494 1324
rect 8444 1006 8466 1324
rect -20266 1000 8466 1006
rect -17888 966 -10718 1000
<< via3 >>
rect -21561 25072 -10287 25081
rect -21561 24234 -21552 25072
rect -21552 24234 -10296 25072
rect -10296 24234 -10287 25072
rect -21561 24225 -10287 24234
rect -17273 16094 -17209 16638
rect -16554 16094 -16490 16638
rect -15835 16094 -15771 16638
rect -15116 16094 -15052 16638
rect -14397 16094 -14333 16638
rect -13678 16094 -13614 16638
rect -12959 16094 -12895 16638
rect -12240 16094 -12176 16638
rect -11521 16094 -11457 16638
rect -10802 16094 -10738 16638
rect -17273 15394 -17209 15938
rect -16554 15394 -16490 15938
rect -15835 15394 -15771 15938
rect -15116 15394 -15052 15938
rect -14397 15394 -14333 15938
rect -13678 15394 -13614 15938
rect -12959 15394 -12895 15938
rect -12240 15394 -12176 15938
rect -11521 15394 -11457 15938
rect -10802 15394 -10738 15938
rect -17273 14694 -17209 15238
rect -16554 14694 -16490 15238
rect -15835 14694 -15771 15238
rect -15116 14694 -15052 15238
rect -14397 14694 -14333 15238
rect -13678 14694 -13614 15238
rect -12959 14694 -12895 15238
rect -12240 14694 -12176 15238
rect -11521 14694 -11457 15238
rect -10802 14694 -10738 15238
rect -17273 13994 -17209 14538
rect -16554 13994 -16490 14538
rect -15835 13994 -15771 14538
rect -15116 13994 -15052 14538
rect -14397 13994 -14333 14538
rect -13678 13994 -13614 14538
rect -12959 13994 -12895 14538
rect -12240 13994 -12176 14538
rect -11521 13994 -11457 14538
rect -10802 13994 -10738 14538
rect -17273 13294 -17209 13838
rect -16554 13294 -16490 13838
rect -15835 13294 -15771 13838
rect -15116 13294 -15052 13838
rect -14397 13294 -14333 13838
rect -13678 13294 -13614 13838
rect -12959 13294 -12895 13838
rect -12240 13294 -12176 13838
rect -11521 13294 -11457 13838
rect -10802 13294 -10738 13838
rect -17273 12594 -17209 13138
rect -16554 12594 -16490 13138
rect -15835 12594 -15771 13138
rect -15116 12594 -15052 13138
rect -14397 12594 -14333 13138
rect -13678 12594 -13614 13138
rect -12959 12594 -12895 13138
rect -12240 12594 -12176 13138
rect -11521 12594 -11457 13138
rect -10802 12594 -10738 13138
rect -17273 11894 -17209 12438
rect -16554 11894 -16490 12438
rect -15835 11894 -15771 12438
rect -15116 11894 -15052 12438
rect -14397 11894 -14333 12438
rect -13678 11894 -13614 12438
rect -12959 11894 -12895 12438
rect -12240 11894 -12176 12438
rect -11521 11894 -11457 12438
rect -10802 11894 -10738 12438
rect -17273 11194 -17209 11738
rect -16554 11194 -16490 11738
rect -15835 11194 -15771 11738
rect -15116 11194 -15052 11738
rect -14397 11194 -14333 11738
rect -13678 11194 -13614 11738
rect -12959 11194 -12895 11738
rect -12240 11194 -12176 11738
rect -11521 11194 -11457 11738
rect -10802 11194 -10738 11738
rect -17273 10494 -17209 11038
rect -16554 10494 -16490 11038
rect -15835 10494 -15771 11038
rect -15116 10494 -15052 11038
rect -14397 10494 -14333 11038
rect -13678 10494 -13614 11038
rect -12959 10494 -12895 11038
rect -12240 10494 -12176 11038
rect -11521 10494 -11457 11038
rect -10802 10494 -10738 11038
rect -9246 10808 11064 11780
rect -17273 9794 -17209 10338
rect -16554 9794 -16490 10338
rect -15835 9794 -15771 10338
rect -15116 9794 -15052 10338
rect -14397 9794 -14333 10338
rect -13678 9794 -13614 10338
rect -12959 9794 -12895 10338
rect -12240 9794 -12176 10338
rect -11521 9794 -11457 10338
rect -10802 9794 -10738 10338
rect -18614 4629 -17986 4643
rect -18614 4377 -18600 4629
rect -18600 4377 -18000 4629
rect -18000 4377 -17986 4629
rect -18614 4363 -17986 4377
rect -10123 4629 -9495 4643
rect -10123 4377 -10109 4629
rect -10109 4377 -9509 4629
rect -9509 4377 -9495 4629
rect -10123 4363 -9495 4377
<< mimcap >>
rect -17788 16526 -17388 16566
rect -17788 16206 -17748 16526
rect -17428 16206 -17388 16526
rect -17788 16166 -17388 16206
rect -17069 16526 -16669 16566
rect -17069 16206 -17029 16526
rect -16709 16206 -16669 16526
rect -17069 16166 -16669 16206
rect -16350 16526 -15950 16566
rect -16350 16206 -16310 16526
rect -15990 16206 -15950 16526
rect -16350 16166 -15950 16206
rect -15631 16526 -15231 16566
rect -15631 16206 -15591 16526
rect -15271 16206 -15231 16526
rect -15631 16166 -15231 16206
rect -14912 16526 -14512 16566
rect -14912 16206 -14872 16526
rect -14552 16206 -14512 16526
rect -14912 16166 -14512 16206
rect -14193 16526 -13793 16566
rect -14193 16206 -14153 16526
rect -13833 16206 -13793 16526
rect -14193 16166 -13793 16206
rect -13474 16526 -13074 16566
rect -13474 16206 -13434 16526
rect -13114 16206 -13074 16526
rect -13474 16166 -13074 16206
rect -12755 16526 -12355 16566
rect -12755 16206 -12715 16526
rect -12395 16206 -12355 16526
rect -12755 16166 -12355 16206
rect -12036 16526 -11636 16566
rect -12036 16206 -11996 16526
rect -11676 16206 -11636 16526
rect -12036 16166 -11636 16206
rect -11317 16526 -10917 16566
rect -11317 16206 -11277 16526
rect -10957 16206 -10917 16526
rect -11317 16166 -10917 16206
rect -17788 15826 -17388 15866
rect -17788 15506 -17748 15826
rect -17428 15506 -17388 15826
rect -17788 15466 -17388 15506
rect -17069 15826 -16669 15866
rect -17069 15506 -17029 15826
rect -16709 15506 -16669 15826
rect -17069 15466 -16669 15506
rect -16350 15826 -15950 15866
rect -16350 15506 -16310 15826
rect -15990 15506 -15950 15826
rect -16350 15466 -15950 15506
rect -15631 15826 -15231 15866
rect -15631 15506 -15591 15826
rect -15271 15506 -15231 15826
rect -15631 15466 -15231 15506
rect -14912 15826 -14512 15866
rect -14912 15506 -14872 15826
rect -14552 15506 -14512 15826
rect -14912 15466 -14512 15506
rect -14193 15826 -13793 15866
rect -14193 15506 -14153 15826
rect -13833 15506 -13793 15826
rect -14193 15466 -13793 15506
rect -13474 15826 -13074 15866
rect -13474 15506 -13434 15826
rect -13114 15506 -13074 15826
rect -13474 15466 -13074 15506
rect -12755 15826 -12355 15866
rect -12755 15506 -12715 15826
rect -12395 15506 -12355 15826
rect -12755 15466 -12355 15506
rect -12036 15826 -11636 15866
rect -12036 15506 -11996 15826
rect -11676 15506 -11636 15826
rect -12036 15466 -11636 15506
rect -11317 15826 -10917 15866
rect -11317 15506 -11277 15826
rect -10957 15506 -10917 15826
rect -11317 15466 -10917 15506
rect -17788 15126 -17388 15166
rect -17788 14806 -17748 15126
rect -17428 14806 -17388 15126
rect -17788 14766 -17388 14806
rect -17069 15126 -16669 15166
rect -17069 14806 -17029 15126
rect -16709 14806 -16669 15126
rect -17069 14766 -16669 14806
rect -16350 15126 -15950 15166
rect -16350 14806 -16310 15126
rect -15990 14806 -15950 15126
rect -16350 14766 -15950 14806
rect -15631 15126 -15231 15166
rect -15631 14806 -15591 15126
rect -15271 14806 -15231 15126
rect -15631 14766 -15231 14806
rect -14912 15126 -14512 15166
rect -14912 14806 -14872 15126
rect -14552 14806 -14512 15126
rect -14912 14766 -14512 14806
rect -14193 15126 -13793 15166
rect -14193 14806 -14153 15126
rect -13833 14806 -13793 15126
rect -14193 14766 -13793 14806
rect -13474 15126 -13074 15166
rect -13474 14806 -13434 15126
rect -13114 14806 -13074 15126
rect -13474 14766 -13074 14806
rect -12755 15126 -12355 15166
rect -12755 14806 -12715 15126
rect -12395 14806 -12355 15126
rect -12755 14766 -12355 14806
rect -12036 15126 -11636 15166
rect -12036 14806 -11996 15126
rect -11676 14806 -11636 15126
rect -12036 14766 -11636 14806
rect -11317 15126 -10917 15166
rect -11317 14806 -11277 15126
rect -10957 14806 -10917 15126
rect -11317 14766 -10917 14806
rect -17788 14426 -17388 14466
rect -17788 14106 -17748 14426
rect -17428 14106 -17388 14426
rect -17788 14066 -17388 14106
rect -17069 14426 -16669 14466
rect -17069 14106 -17029 14426
rect -16709 14106 -16669 14426
rect -17069 14066 -16669 14106
rect -16350 14426 -15950 14466
rect -16350 14106 -16310 14426
rect -15990 14106 -15950 14426
rect -16350 14066 -15950 14106
rect -15631 14426 -15231 14466
rect -15631 14106 -15591 14426
rect -15271 14106 -15231 14426
rect -15631 14066 -15231 14106
rect -14912 14426 -14512 14466
rect -14912 14106 -14872 14426
rect -14552 14106 -14512 14426
rect -14912 14066 -14512 14106
rect -14193 14426 -13793 14466
rect -14193 14106 -14153 14426
rect -13833 14106 -13793 14426
rect -14193 14066 -13793 14106
rect -13474 14426 -13074 14466
rect -13474 14106 -13434 14426
rect -13114 14106 -13074 14426
rect -13474 14066 -13074 14106
rect -12755 14426 -12355 14466
rect -12755 14106 -12715 14426
rect -12395 14106 -12355 14426
rect -12755 14066 -12355 14106
rect -12036 14426 -11636 14466
rect -12036 14106 -11996 14426
rect -11676 14106 -11636 14426
rect -12036 14066 -11636 14106
rect -11317 14426 -10917 14466
rect -11317 14106 -11277 14426
rect -10957 14106 -10917 14426
rect -11317 14066 -10917 14106
rect -17788 13726 -17388 13766
rect -17788 13406 -17748 13726
rect -17428 13406 -17388 13726
rect -17788 13366 -17388 13406
rect -17069 13726 -16669 13766
rect -17069 13406 -17029 13726
rect -16709 13406 -16669 13726
rect -17069 13366 -16669 13406
rect -16350 13726 -15950 13766
rect -16350 13406 -16310 13726
rect -15990 13406 -15950 13726
rect -16350 13366 -15950 13406
rect -15631 13726 -15231 13766
rect -15631 13406 -15591 13726
rect -15271 13406 -15231 13726
rect -15631 13366 -15231 13406
rect -14912 13726 -14512 13766
rect -14912 13406 -14872 13726
rect -14552 13406 -14512 13726
rect -14912 13366 -14512 13406
rect -14193 13726 -13793 13766
rect -14193 13406 -14153 13726
rect -13833 13406 -13793 13726
rect -14193 13366 -13793 13406
rect -13474 13726 -13074 13766
rect -13474 13406 -13434 13726
rect -13114 13406 -13074 13726
rect -13474 13366 -13074 13406
rect -12755 13726 -12355 13766
rect -12755 13406 -12715 13726
rect -12395 13406 -12355 13726
rect -12755 13366 -12355 13406
rect -12036 13726 -11636 13766
rect -12036 13406 -11996 13726
rect -11676 13406 -11636 13726
rect -12036 13366 -11636 13406
rect -11317 13726 -10917 13766
rect -11317 13406 -11277 13726
rect -10957 13406 -10917 13726
rect -11317 13366 -10917 13406
rect -17788 13026 -17388 13066
rect -17788 12706 -17748 13026
rect -17428 12706 -17388 13026
rect -17788 12666 -17388 12706
rect -17069 13026 -16669 13066
rect -17069 12706 -17029 13026
rect -16709 12706 -16669 13026
rect -17069 12666 -16669 12706
rect -16350 13026 -15950 13066
rect -16350 12706 -16310 13026
rect -15990 12706 -15950 13026
rect -16350 12666 -15950 12706
rect -15631 13026 -15231 13066
rect -15631 12706 -15591 13026
rect -15271 12706 -15231 13026
rect -15631 12666 -15231 12706
rect -14912 13026 -14512 13066
rect -14912 12706 -14872 13026
rect -14552 12706 -14512 13026
rect -14912 12666 -14512 12706
rect -14193 13026 -13793 13066
rect -14193 12706 -14153 13026
rect -13833 12706 -13793 13026
rect -14193 12666 -13793 12706
rect -13474 13026 -13074 13066
rect -13474 12706 -13434 13026
rect -13114 12706 -13074 13026
rect -13474 12666 -13074 12706
rect -12755 13026 -12355 13066
rect -12755 12706 -12715 13026
rect -12395 12706 -12355 13026
rect -12755 12666 -12355 12706
rect -12036 13026 -11636 13066
rect -12036 12706 -11996 13026
rect -11676 12706 -11636 13026
rect -12036 12666 -11636 12706
rect -11317 13026 -10917 13066
rect -11317 12706 -11277 13026
rect -10957 12706 -10917 13026
rect -11317 12666 -10917 12706
rect -17788 12326 -17388 12366
rect -17788 12006 -17748 12326
rect -17428 12006 -17388 12326
rect -17788 11966 -17388 12006
rect -17069 12326 -16669 12366
rect -17069 12006 -17029 12326
rect -16709 12006 -16669 12326
rect -17069 11966 -16669 12006
rect -16350 12326 -15950 12366
rect -16350 12006 -16310 12326
rect -15990 12006 -15950 12326
rect -16350 11966 -15950 12006
rect -15631 12326 -15231 12366
rect -15631 12006 -15591 12326
rect -15271 12006 -15231 12326
rect -15631 11966 -15231 12006
rect -14912 12326 -14512 12366
rect -14912 12006 -14872 12326
rect -14552 12006 -14512 12326
rect -14912 11966 -14512 12006
rect -14193 12326 -13793 12366
rect -14193 12006 -14153 12326
rect -13833 12006 -13793 12326
rect -14193 11966 -13793 12006
rect -13474 12326 -13074 12366
rect -13474 12006 -13434 12326
rect -13114 12006 -13074 12326
rect -13474 11966 -13074 12006
rect -12755 12326 -12355 12366
rect -12755 12006 -12715 12326
rect -12395 12006 -12355 12326
rect -12755 11966 -12355 12006
rect -12036 12326 -11636 12366
rect -12036 12006 -11996 12326
rect -11676 12006 -11636 12326
rect -12036 11966 -11636 12006
rect -11317 12326 -10917 12366
rect -11317 12006 -11277 12326
rect -10957 12006 -10917 12326
rect -11317 11966 -10917 12006
rect -17788 11626 -17388 11666
rect -17788 11306 -17748 11626
rect -17428 11306 -17388 11626
rect -17788 11266 -17388 11306
rect -17069 11626 -16669 11666
rect -17069 11306 -17029 11626
rect -16709 11306 -16669 11626
rect -17069 11266 -16669 11306
rect -16350 11626 -15950 11666
rect -16350 11306 -16310 11626
rect -15990 11306 -15950 11626
rect -16350 11266 -15950 11306
rect -15631 11626 -15231 11666
rect -15631 11306 -15591 11626
rect -15271 11306 -15231 11626
rect -15631 11266 -15231 11306
rect -14912 11626 -14512 11666
rect -14912 11306 -14872 11626
rect -14552 11306 -14512 11626
rect -14912 11266 -14512 11306
rect -14193 11626 -13793 11666
rect -14193 11306 -14153 11626
rect -13833 11306 -13793 11626
rect -14193 11266 -13793 11306
rect -13474 11626 -13074 11666
rect -13474 11306 -13434 11626
rect -13114 11306 -13074 11626
rect -13474 11266 -13074 11306
rect -12755 11626 -12355 11666
rect -12755 11306 -12715 11626
rect -12395 11306 -12355 11626
rect -12755 11266 -12355 11306
rect -12036 11626 -11636 11666
rect -12036 11306 -11996 11626
rect -11676 11306 -11636 11626
rect -12036 11266 -11636 11306
rect -11317 11626 -10917 11666
rect -11317 11306 -11277 11626
rect -10957 11306 -10917 11626
rect -11317 11266 -10917 11306
rect -17788 10926 -17388 10966
rect -17788 10606 -17748 10926
rect -17428 10606 -17388 10926
rect -17788 10566 -17388 10606
rect -17069 10926 -16669 10966
rect -17069 10606 -17029 10926
rect -16709 10606 -16669 10926
rect -17069 10566 -16669 10606
rect -16350 10926 -15950 10966
rect -16350 10606 -16310 10926
rect -15990 10606 -15950 10926
rect -16350 10566 -15950 10606
rect -15631 10926 -15231 10966
rect -15631 10606 -15591 10926
rect -15271 10606 -15231 10926
rect -15631 10566 -15231 10606
rect -14912 10926 -14512 10966
rect -14912 10606 -14872 10926
rect -14552 10606 -14512 10926
rect -14912 10566 -14512 10606
rect -14193 10926 -13793 10966
rect -14193 10606 -14153 10926
rect -13833 10606 -13793 10926
rect -14193 10566 -13793 10606
rect -13474 10926 -13074 10966
rect -13474 10606 -13434 10926
rect -13114 10606 -13074 10926
rect -13474 10566 -13074 10606
rect -12755 10926 -12355 10966
rect -12755 10606 -12715 10926
rect -12395 10606 -12355 10926
rect -12755 10566 -12355 10606
rect -12036 10926 -11636 10966
rect -12036 10606 -11996 10926
rect -11676 10606 -11636 10926
rect -12036 10566 -11636 10606
rect -11317 10926 -10917 10966
rect -11317 10606 -11277 10926
rect -10957 10606 -10917 10926
rect -11317 10566 -10917 10606
rect -17788 10226 -17388 10266
rect -17788 9906 -17748 10226
rect -17428 9906 -17388 10226
rect -17788 9866 -17388 9906
rect -17069 10226 -16669 10266
rect -17069 9906 -17029 10226
rect -16709 9906 -16669 10226
rect -17069 9866 -16669 9906
rect -16350 10226 -15950 10266
rect -16350 9906 -16310 10226
rect -15990 9906 -15950 10226
rect -16350 9866 -15950 9906
rect -15631 10226 -15231 10266
rect -15631 9906 -15591 10226
rect -15271 9906 -15231 10226
rect -15631 9866 -15231 9906
rect -14912 10226 -14512 10266
rect -14912 9906 -14872 10226
rect -14552 9906 -14512 10226
rect -14912 9866 -14512 9906
rect -14193 10226 -13793 10266
rect -14193 9906 -14153 10226
rect -13833 9906 -13793 10226
rect -14193 9866 -13793 9906
rect -13474 10226 -13074 10266
rect -13474 9906 -13434 10226
rect -13114 9906 -13074 10226
rect -13474 9866 -13074 9906
rect -12755 10226 -12355 10266
rect -12755 9906 -12715 10226
rect -12395 9906 -12355 10226
rect -12755 9866 -12355 9906
rect -12036 10226 -11636 10266
rect -12036 9906 -11996 10226
rect -11676 9906 -11636 10226
rect -12036 9866 -11636 9906
rect -11317 10226 -10917 10266
rect -11317 9906 -11277 10226
rect -10957 9906 -10917 10226
rect -11317 9866 -10917 9906
<< mimcapcontact >>
rect -17748 16206 -17428 16526
rect -17029 16206 -16709 16526
rect -16310 16206 -15990 16526
rect -15591 16206 -15271 16526
rect -14872 16206 -14552 16526
rect -14153 16206 -13833 16526
rect -13434 16206 -13114 16526
rect -12715 16206 -12395 16526
rect -11996 16206 -11676 16526
rect -11277 16206 -10957 16526
rect -17748 15506 -17428 15826
rect -17029 15506 -16709 15826
rect -16310 15506 -15990 15826
rect -15591 15506 -15271 15826
rect -14872 15506 -14552 15826
rect -14153 15506 -13833 15826
rect -13434 15506 -13114 15826
rect -12715 15506 -12395 15826
rect -11996 15506 -11676 15826
rect -11277 15506 -10957 15826
rect -17748 14806 -17428 15126
rect -17029 14806 -16709 15126
rect -16310 14806 -15990 15126
rect -15591 14806 -15271 15126
rect -14872 14806 -14552 15126
rect -14153 14806 -13833 15126
rect -13434 14806 -13114 15126
rect -12715 14806 -12395 15126
rect -11996 14806 -11676 15126
rect -11277 14806 -10957 15126
rect -17748 14106 -17428 14426
rect -17029 14106 -16709 14426
rect -16310 14106 -15990 14426
rect -15591 14106 -15271 14426
rect -14872 14106 -14552 14426
rect -14153 14106 -13833 14426
rect -13434 14106 -13114 14426
rect -12715 14106 -12395 14426
rect -11996 14106 -11676 14426
rect -11277 14106 -10957 14426
rect -17748 13406 -17428 13726
rect -17029 13406 -16709 13726
rect -16310 13406 -15990 13726
rect -15591 13406 -15271 13726
rect -14872 13406 -14552 13726
rect -14153 13406 -13833 13726
rect -13434 13406 -13114 13726
rect -12715 13406 -12395 13726
rect -11996 13406 -11676 13726
rect -11277 13406 -10957 13726
rect -17748 12706 -17428 13026
rect -17029 12706 -16709 13026
rect -16310 12706 -15990 13026
rect -15591 12706 -15271 13026
rect -14872 12706 -14552 13026
rect -14153 12706 -13833 13026
rect -13434 12706 -13114 13026
rect -12715 12706 -12395 13026
rect -11996 12706 -11676 13026
rect -11277 12706 -10957 13026
rect -17748 12006 -17428 12326
rect -17029 12006 -16709 12326
rect -16310 12006 -15990 12326
rect -15591 12006 -15271 12326
rect -14872 12006 -14552 12326
rect -14153 12006 -13833 12326
rect -13434 12006 -13114 12326
rect -12715 12006 -12395 12326
rect -11996 12006 -11676 12326
rect -11277 12006 -10957 12326
rect -17748 11306 -17428 11626
rect -17029 11306 -16709 11626
rect -16310 11306 -15990 11626
rect -15591 11306 -15271 11626
rect -14872 11306 -14552 11626
rect -14153 11306 -13833 11626
rect -13434 11306 -13114 11626
rect -12715 11306 -12395 11626
rect -11996 11306 -11676 11626
rect -11277 11306 -10957 11626
rect -17748 10606 -17428 10926
rect -17029 10606 -16709 10926
rect -16310 10606 -15990 10926
rect -15591 10606 -15271 10926
rect -14872 10606 -14552 10926
rect -14153 10606 -13833 10926
rect -13434 10606 -13114 10926
rect -12715 10606 -12395 10926
rect -11996 10606 -11676 10926
rect -11277 10606 -10957 10926
rect -17748 9906 -17428 10226
rect -17029 9906 -16709 10226
rect -16310 9906 -15990 10226
rect -15591 9906 -15271 10226
rect -14872 9906 -14552 10226
rect -14153 9906 -13833 10226
rect -13434 9906 -13114 10226
rect -12715 9906 -12395 10226
rect -11996 9906 -11676 10226
rect -11277 9906 -10957 10226
<< metal4 >>
rect -21578 25081 -10252 25118
rect -21578 24225 -21561 25081
rect -10287 24225 -10252 25081
rect -21578 16956 -10252 24225
rect -21532 16950 -10252 16956
rect -17289 16638 -17193 16654
rect -17788 16526 -17388 16566
rect -17788 16206 -17748 16526
rect -17428 16206 -17388 16526
rect -17788 15826 -17388 16206
rect -17289 16094 -17273 16638
rect -17209 16094 -17193 16638
rect -16570 16638 -16474 16654
rect -17289 16078 -17193 16094
rect -17068 16526 -16668 16566
rect -17068 16206 -17029 16526
rect -16709 16206 -16668 16526
rect -17788 15506 -17748 15826
rect -17428 15506 -17388 15826
rect -17788 15126 -17388 15506
rect -17289 15938 -17193 15954
rect -17289 15394 -17273 15938
rect -17209 15394 -17193 15938
rect -17289 15378 -17193 15394
rect -17068 15826 -16668 16206
rect -16570 16094 -16554 16638
rect -16490 16094 -16474 16638
rect -15851 16638 -15755 16654
rect -16570 16078 -16474 16094
rect -16348 16526 -15948 16566
rect -16348 16206 -16310 16526
rect -15990 16206 -15948 16526
rect -17068 15506 -17029 15826
rect -16709 15506 -16668 15826
rect -17788 14806 -17748 15126
rect -17428 14806 -17388 15126
rect -17788 14426 -17388 14806
rect -17289 15238 -17193 15254
rect -17289 14694 -17273 15238
rect -17209 14694 -17193 15238
rect -17289 14678 -17193 14694
rect -17068 15126 -16668 15506
rect -16570 15938 -16474 15954
rect -16570 15394 -16554 15938
rect -16490 15394 -16474 15938
rect -16570 15378 -16474 15394
rect -16348 15826 -15948 16206
rect -15851 16094 -15835 16638
rect -15771 16094 -15755 16638
rect -15132 16638 -15036 16654
rect -15851 16078 -15755 16094
rect -15628 16526 -15228 16566
rect -15628 16206 -15591 16526
rect -15271 16206 -15228 16526
rect -16348 15506 -16310 15826
rect -15990 15506 -15948 15826
rect -17068 14806 -17029 15126
rect -16709 14806 -16668 15126
rect -17788 14106 -17748 14426
rect -17428 14106 -17388 14426
rect -17788 13726 -17388 14106
rect -17289 14538 -17193 14554
rect -17289 13994 -17273 14538
rect -17209 13994 -17193 14538
rect -17289 13978 -17193 13994
rect -17068 14426 -16668 14806
rect -16570 15238 -16474 15254
rect -16570 14694 -16554 15238
rect -16490 14694 -16474 15238
rect -16570 14678 -16474 14694
rect -16348 15126 -15948 15506
rect -15851 15938 -15755 15954
rect -15851 15394 -15835 15938
rect -15771 15394 -15755 15938
rect -15851 15378 -15755 15394
rect -15628 15826 -15228 16206
rect -15132 16094 -15116 16638
rect -15052 16094 -15036 16638
rect -14413 16638 -14317 16654
rect -15132 16078 -15036 16094
rect -14908 16526 -14508 16566
rect -14908 16206 -14872 16526
rect -14552 16206 -14508 16526
rect -15628 15506 -15591 15826
rect -15271 15506 -15228 15826
rect -16348 14806 -16310 15126
rect -15990 14806 -15948 15126
rect -17068 14106 -17029 14426
rect -16709 14106 -16668 14426
rect -17788 13406 -17748 13726
rect -17428 13406 -17388 13726
rect -17788 13026 -17388 13406
rect -17289 13838 -17193 13854
rect -17289 13294 -17273 13838
rect -17209 13294 -17193 13838
rect -17289 13278 -17193 13294
rect -17068 13726 -16668 14106
rect -16570 14538 -16474 14554
rect -16570 13994 -16554 14538
rect -16490 13994 -16474 14538
rect -16570 13978 -16474 13994
rect -16348 14426 -15948 14806
rect -15851 15238 -15755 15254
rect -15851 14694 -15835 15238
rect -15771 14694 -15755 15238
rect -15851 14678 -15755 14694
rect -15628 15126 -15228 15506
rect -15132 15938 -15036 15954
rect -15132 15394 -15116 15938
rect -15052 15394 -15036 15938
rect -15132 15378 -15036 15394
rect -14908 15826 -14508 16206
rect -14413 16094 -14397 16638
rect -14333 16094 -14317 16638
rect -13694 16638 -13598 16654
rect -14413 16078 -14317 16094
rect -14188 16526 -13788 16566
rect -14188 16206 -14153 16526
rect -13833 16206 -13788 16526
rect -14908 15506 -14872 15826
rect -14552 15506 -14508 15826
rect -15628 14806 -15591 15126
rect -15271 14806 -15228 15126
rect -16348 14106 -16310 14426
rect -15990 14106 -15948 14426
rect -17068 13406 -17029 13726
rect -16709 13406 -16668 13726
rect -17788 12706 -17748 13026
rect -17428 12706 -17388 13026
rect -17788 12326 -17388 12706
rect -17289 13138 -17193 13154
rect -17289 12594 -17273 13138
rect -17209 12594 -17193 13138
rect -17289 12578 -17193 12594
rect -17068 13026 -16668 13406
rect -16570 13838 -16474 13854
rect -16570 13294 -16554 13838
rect -16490 13294 -16474 13838
rect -16570 13278 -16474 13294
rect -16348 13726 -15948 14106
rect -15851 14538 -15755 14554
rect -15851 13994 -15835 14538
rect -15771 13994 -15755 14538
rect -15851 13978 -15755 13994
rect -15628 14426 -15228 14806
rect -15132 15238 -15036 15254
rect -15132 14694 -15116 15238
rect -15052 14694 -15036 15238
rect -15132 14678 -15036 14694
rect -14908 15126 -14508 15506
rect -14413 15938 -14317 15954
rect -14413 15394 -14397 15938
rect -14333 15394 -14317 15938
rect -14413 15378 -14317 15394
rect -14188 15826 -13788 16206
rect -13694 16094 -13678 16638
rect -13614 16094 -13598 16638
rect -12975 16638 -12879 16654
rect -13694 16078 -13598 16094
rect -13468 16526 -13068 16566
rect -13468 16206 -13434 16526
rect -13114 16206 -13068 16526
rect -14188 15506 -14153 15826
rect -13833 15506 -13788 15826
rect -14908 14806 -14872 15126
rect -14552 14806 -14508 15126
rect -15628 14106 -15591 14426
rect -15271 14106 -15228 14426
rect -16348 13406 -16310 13726
rect -15990 13406 -15948 13726
rect -17068 12706 -17029 13026
rect -16709 12706 -16668 13026
rect -17788 12006 -17748 12326
rect -17428 12006 -17388 12326
rect -17788 11626 -17388 12006
rect -17289 12438 -17193 12454
rect -17289 11894 -17273 12438
rect -17209 11894 -17193 12438
rect -17289 11878 -17193 11894
rect -17068 12326 -16668 12706
rect -16570 13138 -16474 13154
rect -16570 12594 -16554 13138
rect -16490 12594 -16474 13138
rect -16570 12578 -16474 12594
rect -16348 13026 -15948 13406
rect -15851 13838 -15755 13854
rect -15851 13294 -15835 13838
rect -15771 13294 -15755 13838
rect -15851 13278 -15755 13294
rect -15628 13726 -15228 14106
rect -15132 14538 -15036 14554
rect -15132 13994 -15116 14538
rect -15052 13994 -15036 14538
rect -15132 13978 -15036 13994
rect -14908 14426 -14508 14806
rect -14413 15238 -14317 15254
rect -14413 14694 -14397 15238
rect -14333 14694 -14317 15238
rect -14413 14678 -14317 14694
rect -14188 15126 -13788 15506
rect -13694 15938 -13598 15954
rect -13694 15394 -13678 15938
rect -13614 15394 -13598 15938
rect -13694 15378 -13598 15394
rect -13468 15826 -13068 16206
rect -12975 16094 -12959 16638
rect -12895 16094 -12879 16638
rect -12256 16638 -12160 16654
rect -12975 16078 -12879 16094
rect -12748 16526 -12348 16566
rect -12748 16206 -12715 16526
rect -12395 16206 -12348 16526
rect -13468 15506 -13434 15826
rect -13114 15506 -13068 15826
rect -14188 14806 -14153 15126
rect -13833 14806 -13788 15126
rect -14908 14106 -14872 14426
rect -14552 14106 -14508 14426
rect -15628 13406 -15591 13726
rect -15271 13406 -15228 13726
rect -16348 12706 -16310 13026
rect -15990 12706 -15948 13026
rect -17068 12006 -17029 12326
rect -16709 12006 -16668 12326
rect -17788 11306 -17748 11626
rect -17428 11306 -17388 11626
rect -17788 10926 -17388 11306
rect -17289 11738 -17193 11754
rect -17289 11194 -17273 11738
rect -17209 11194 -17193 11738
rect -17289 11178 -17193 11194
rect -17068 11626 -16668 12006
rect -16570 12438 -16474 12454
rect -16570 11894 -16554 12438
rect -16490 11894 -16474 12438
rect -16570 11878 -16474 11894
rect -16348 12326 -15948 12706
rect -15851 13138 -15755 13154
rect -15851 12594 -15835 13138
rect -15771 12594 -15755 13138
rect -15851 12578 -15755 12594
rect -15628 13026 -15228 13406
rect -15132 13838 -15036 13854
rect -15132 13294 -15116 13838
rect -15052 13294 -15036 13838
rect -15132 13278 -15036 13294
rect -14908 13726 -14508 14106
rect -14413 14538 -14317 14554
rect -14413 13994 -14397 14538
rect -14333 13994 -14317 14538
rect -14413 13978 -14317 13994
rect -14188 14426 -13788 14806
rect -13694 15238 -13598 15254
rect -13694 14694 -13678 15238
rect -13614 14694 -13598 15238
rect -13694 14678 -13598 14694
rect -13468 15126 -13068 15506
rect -12975 15938 -12879 15954
rect -12975 15394 -12959 15938
rect -12895 15394 -12879 15938
rect -12975 15378 -12879 15394
rect -12748 15826 -12348 16206
rect -12256 16094 -12240 16638
rect -12176 16094 -12160 16638
rect -11537 16638 -11441 16654
rect -12256 16078 -12160 16094
rect -12028 16526 -11628 16566
rect -12028 16206 -11996 16526
rect -11676 16206 -11628 16526
rect -12748 15506 -12715 15826
rect -12395 15506 -12348 15826
rect -13468 14806 -13434 15126
rect -13114 14806 -13068 15126
rect -14188 14106 -14153 14426
rect -13833 14106 -13788 14426
rect -14908 13406 -14872 13726
rect -14552 13406 -14508 13726
rect -15628 12706 -15591 13026
rect -15271 12706 -15228 13026
rect -16348 12006 -16310 12326
rect -15990 12006 -15948 12326
rect -17068 11306 -17029 11626
rect -16709 11306 -16668 11626
rect -17788 10606 -17748 10926
rect -17428 10606 -17388 10926
rect -17788 10226 -17388 10606
rect -17289 11038 -17193 11054
rect -17289 10494 -17273 11038
rect -17209 10494 -17193 11038
rect -17289 10478 -17193 10494
rect -17068 10926 -16668 11306
rect -16570 11738 -16474 11754
rect -16570 11194 -16554 11738
rect -16490 11194 -16474 11738
rect -16570 11178 -16474 11194
rect -16348 11626 -15948 12006
rect -15851 12438 -15755 12454
rect -15851 11894 -15835 12438
rect -15771 11894 -15755 12438
rect -15851 11878 -15755 11894
rect -15628 12326 -15228 12706
rect -15132 13138 -15036 13154
rect -15132 12594 -15116 13138
rect -15052 12594 -15036 13138
rect -15132 12578 -15036 12594
rect -14908 13026 -14508 13406
rect -14413 13838 -14317 13854
rect -14413 13294 -14397 13838
rect -14333 13294 -14317 13838
rect -14413 13278 -14317 13294
rect -14188 13726 -13788 14106
rect -13694 14538 -13598 14554
rect -13694 13994 -13678 14538
rect -13614 13994 -13598 14538
rect -13694 13978 -13598 13994
rect -13468 14426 -13068 14806
rect -12975 15238 -12879 15254
rect -12975 14694 -12959 15238
rect -12895 14694 -12879 15238
rect -12975 14678 -12879 14694
rect -12748 15126 -12348 15506
rect -12256 15938 -12160 15954
rect -12256 15394 -12240 15938
rect -12176 15394 -12160 15938
rect -12256 15378 -12160 15394
rect -12028 15826 -11628 16206
rect -11537 16094 -11521 16638
rect -11457 16094 -11441 16638
rect -10818 16638 -10722 16654
rect -11317 16526 -10908 16566
rect -11317 16206 -11277 16526
rect -10957 16206 -10908 16526
rect -11317 16166 -10908 16206
rect -11537 16078 -11441 16094
rect -12028 15506 -11996 15826
rect -11676 15506 -11628 15826
rect -12748 14806 -12715 15126
rect -12395 14806 -12348 15126
rect -13468 14106 -13434 14426
rect -13114 14106 -13068 14426
rect -14188 13406 -14153 13726
rect -13833 13406 -13788 13726
rect -14908 12706 -14872 13026
rect -14552 12706 -14508 13026
rect -15628 12006 -15591 12326
rect -15271 12006 -15228 12326
rect -16348 11306 -16310 11626
rect -15990 11306 -15948 11626
rect -17068 10606 -17029 10926
rect -16709 10606 -16668 10926
rect -17788 9906 -17748 10226
rect -17428 9906 -17388 10226
rect -17788 9698 -17388 9906
rect -17289 10338 -17193 10354
rect -17289 9794 -17273 10338
rect -17209 9794 -17193 10338
rect -17289 9778 -17193 9794
rect -17068 10226 -16668 10606
rect -16570 11038 -16474 11054
rect -16570 10494 -16554 11038
rect -16490 10494 -16474 11038
rect -16570 10478 -16474 10494
rect -16348 10926 -15948 11306
rect -15851 11738 -15755 11754
rect -15851 11194 -15835 11738
rect -15771 11194 -15755 11738
rect -15851 11178 -15755 11194
rect -15628 11626 -15228 12006
rect -15132 12438 -15036 12454
rect -15132 11894 -15116 12438
rect -15052 11894 -15036 12438
rect -15132 11878 -15036 11894
rect -14908 12326 -14508 12706
rect -14413 13138 -14317 13154
rect -14413 12594 -14397 13138
rect -14333 12594 -14317 13138
rect -14413 12578 -14317 12594
rect -14188 13026 -13788 13406
rect -13694 13838 -13598 13854
rect -13694 13294 -13678 13838
rect -13614 13294 -13598 13838
rect -13694 13278 -13598 13294
rect -13468 13726 -13068 14106
rect -12975 14538 -12879 14554
rect -12975 13994 -12959 14538
rect -12895 13994 -12879 14538
rect -12975 13978 -12879 13994
rect -12748 14426 -12348 14806
rect -12256 15238 -12160 15254
rect -12256 14694 -12240 15238
rect -12176 14694 -12160 15238
rect -12256 14678 -12160 14694
rect -12028 15126 -11628 15506
rect -11537 15938 -11441 15954
rect -11537 15394 -11521 15938
rect -11457 15394 -11441 15938
rect -11537 15378 -11441 15394
rect -11308 15826 -10908 16166
rect -10818 16094 -10802 16638
rect -10738 16094 -10722 16638
rect -10818 16078 -10722 16094
rect -11308 15506 -11277 15826
rect -10957 15506 -10908 15826
rect -12028 14806 -11996 15126
rect -11676 14806 -11628 15126
rect -12748 14106 -12715 14426
rect -12395 14106 -12348 14426
rect -13468 13406 -13434 13726
rect -13114 13406 -13068 13726
rect -14188 12706 -14153 13026
rect -13833 12706 -13788 13026
rect -14908 12006 -14872 12326
rect -14552 12006 -14508 12326
rect -15628 11306 -15591 11626
rect -15271 11306 -15228 11626
rect -16348 10606 -16310 10926
rect -15990 10606 -15948 10926
rect -17068 9906 -17029 10226
rect -16709 9906 -16668 10226
rect -17068 9698 -16668 9906
rect -16570 10338 -16474 10354
rect -16570 9794 -16554 10338
rect -16490 9794 -16474 10338
rect -16570 9778 -16474 9794
rect -16348 10226 -15948 10606
rect -15851 11038 -15755 11054
rect -15851 10494 -15835 11038
rect -15771 10494 -15755 11038
rect -15851 10478 -15755 10494
rect -15628 10926 -15228 11306
rect -15132 11738 -15036 11754
rect -15132 11194 -15116 11738
rect -15052 11194 -15036 11738
rect -15132 11178 -15036 11194
rect -14908 11626 -14508 12006
rect -14413 12438 -14317 12454
rect -14413 11894 -14397 12438
rect -14333 11894 -14317 12438
rect -14413 11878 -14317 11894
rect -14188 12326 -13788 12706
rect -13694 13138 -13598 13154
rect -13694 12594 -13678 13138
rect -13614 12594 -13598 13138
rect -13694 12578 -13598 12594
rect -13468 13026 -13068 13406
rect -12975 13838 -12879 13854
rect -12975 13294 -12959 13838
rect -12895 13294 -12879 13838
rect -12975 13278 -12879 13294
rect -12748 13726 -12348 14106
rect -12256 14538 -12160 14554
rect -12256 13994 -12240 14538
rect -12176 13994 -12160 14538
rect -12256 13978 -12160 13994
rect -12028 14426 -11628 14806
rect -11537 15238 -11441 15254
rect -11537 14694 -11521 15238
rect -11457 14694 -11441 15238
rect -11537 14678 -11441 14694
rect -11308 15126 -10908 15506
rect -10818 15938 -10722 15954
rect -10818 15394 -10802 15938
rect -10738 15394 -10722 15938
rect -10818 15378 -10722 15394
rect -11308 14806 -11277 15126
rect -10957 14806 -10908 15126
rect -12028 14106 -11996 14426
rect -11676 14106 -11628 14426
rect -12748 13406 -12715 13726
rect -12395 13406 -12348 13726
rect -13468 12706 -13434 13026
rect -13114 12706 -13068 13026
rect -14188 12006 -14153 12326
rect -13833 12006 -13788 12326
rect -14908 11306 -14872 11626
rect -14552 11306 -14508 11626
rect -15628 10606 -15591 10926
rect -15271 10606 -15228 10926
rect -16348 9906 -16310 10226
rect -15990 9906 -15948 10226
rect -16348 9698 -15948 9906
rect -15851 10338 -15755 10354
rect -15851 9794 -15835 10338
rect -15771 9794 -15755 10338
rect -15851 9778 -15755 9794
rect -15628 10226 -15228 10606
rect -15132 11038 -15036 11054
rect -15132 10494 -15116 11038
rect -15052 10494 -15036 11038
rect -15132 10478 -15036 10494
rect -14908 10926 -14508 11306
rect -14413 11738 -14317 11754
rect -14413 11194 -14397 11738
rect -14333 11194 -14317 11738
rect -14413 11178 -14317 11194
rect -14188 11626 -13788 12006
rect -13694 12438 -13598 12454
rect -13694 11894 -13678 12438
rect -13614 11894 -13598 12438
rect -13694 11878 -13598 11894
rect -13468 12326 -13068 12706
rect -12975 13138 -12879 13154
rect -12975 12594 -12959 13138
rect -12895 12594 -12879 13138
rect -12975 12578 -12879 12594
rect -12748 13026 -12348 13406
rect -12256 13838 -12160 13854
rect -12256 13294 -12240 13838
rect -12176 13294 -12160 13838
rect -12256 13278 -12160 13294
rect -12028 13726 -11628 14106
rect -11537 14538 -11441 14554
rect -11537 13994 -11521 14538
rect -11457 13994 -11441 14538
rect -11537 13978 -11441 13994
rect -11308 14426 -10908 14806
rect -10818 15238 -10722 15254
rect -10818 14694 -10802 15238
rect -10738 14694 -10722 15238
rect -10818 14678 -10722 14694
rect -11308 14106 -11277 14426
rect -10957 14106 -10908 14426
rect -12028 13406 -11996 13726
rect -11676 13406 -11628 13726
rect -12748 12706 -12715 13026
rect -12395 12706 -12348 13026
rect -13468 12006 -13434 12326
rect -13114 12006 -13068 12326
rect -14188 11306 -14153 11626
rect -13833 11306 -13788 11626
rect -14908 10606 -14872 10926
rect -14552 10606 -14508 10926
rect -15628 9906 -15591 10226
rect -15271 9906 -15228 10226
rect -15628 9698 -15228 9906
rect -15132 10338 -15036 10354
rect -15132 9794 -15116 10338
rect -15052 9794 -15036 10338
rect -15132 9778 -15036 9794
rect -14908 10226 -14508 10606
rect -14413 11038 -14317 11054
rect -14413 10494 -14397 11038
rect -14333 10494 -14317 11038
rect -14413 10478 -14317 10494
rect -14188 10926 -13788 11306
rect -13694 11738 -13598 11754
rect -13694 11194 -13678 11738
rect -13614 11194 -13598 11738
rect -13694 11178 -13598 11194
rect -13468 11626 -13068 12006
rect -12975 12438 -12879 12454
rect -12975 11894 -12959 12438
rect -12895 11894 -12879 12438
rect -12975 11878 -12879 11894
rect -12748 12326 -12348 12706
rect -12256 13138 -12160 13154
rect -12256 12594 -12240 13138
rect -12176 12594 -12160 13138
rect -12256 12578 -12160 12594
rect -12028 13026 -11628 13406
rect -11537 13838 -11441 13854
rect -11537 13294 -11521 13838
rect -11457 13294 -11441 13838
rect -11537 13278 -11441 13294
rect -11308 13726 -10908 14106
rect -10818 14538 -10722 14554
rect -10818 13994 -10802 14538
rect -10738 13994 -10722 14538
rect -10818 13978 -10722 13994
rect -11308 13406 -11277 13726
rect -10957 13406 -10908 13726
rect -12028 12706 -11996 13026
rect -11676 12706 -11628 13026
rect -12748 12006 -12715 12326
rect -12395 12006 -12348 12326
rect -13468 11306 -13434 11626
rect -13114 11306 -13068 11626
rect -14188 10606 -14153 10926
rect -13833 10606 -13788 10926
rect -14908 9906 -14872 10226
rect -14552 9906 -14508 10226
rect -14908 9698 -14508 9906
rect -14413 10338 -14317 10354
rect -14413 9794 -14397 10338
rect -14333 9794 -14317 10338
rect -14413 9778 -14317 9794
rect -14188 10226 -13788 10606
rect -13694 11038 -13598 11054
rect -13694 10494 -13678 11038
rect -13614 10494 -13598 11038
rect -13694 10478 -13598 10494
rect -13468 10926 -13068 11306
rect -12975 11738 -12879 11754
rect -12975 11194 -12959 11738
rect -12895 11194 -12879 11738
rect -12975 11178 -12879 11194
rect -12748 11626 -12348 12006
rect -12256 12438 -12160 12454
rect -12256 11894 -12240 12438
rect -12176 11894 -12160 12438
rect -12256 11878 -12160 11894
rect -12028 12326 -11628 12706
rect -11537 13138 -11441 13154
rect -11537 12594 -11521 13138
rect -11457 12594 -11441 13138
rect -11537 12578 -11441 12594
rect -11308 13026 -10908 13406
rect -10818 13838 -10722 13854
rect -10818 13294 -10802 13838
rect -10738 13294 -10722 13838
rect -10818 13278 -10722 13294
rect -11308 12706 -11277 13026
rect -10957 12706 -10908 13026
rect -12028 12006 -11996 12326
rect -11676 12006 -11628 12326
rect -12748 11306 -12715 11626
rect -12395 11306 -12348 11626
rect -13468 10606 -13434 10926
rect -13114 10606 -13068 10926
rect -14188 9906 -14153 10226
rect -13833 9906 -13788 10226
rect -14188 9698 -13788 9906
rect -13694 10338 -13598 10354
rect -13694 9794 -13678 10338
rect -13614 9794 -13598 10338
rect -13694 9778 -13598 9794
rect -13468 10226 -13068 10606
rect -12975 11038 -12879 11054
rect -12975 10494 -12959 11038
rect -12895 10494 -12879 11038
rect -12975 10478 -12879 10494
rect -12748 10926 -12348 11306
rect -12256 11738 -12160 11754
rect -12256 11194 -12240 11738
rect -12176 11194 -12160 11738
rect -12256 11178 -12160 11194
rect -12028 11626 -11628 12006
rect -11537 12438 -11441 12454
rect -11537 11894 -11521 12438
rect -11457 11894 -11441 12438
rect -11537 11878 -11441 11894
rect -11308 12326 -10908 12706
rect -10818 13138 -10722 13154
rect -10818 12594 -10802 13138
rect -10738 12594 -10722 13138
rect -10818 12578 -10722 12594
rect -11308 12006 -11277 12326
rect -10957 12006 -10908 12326
rect -12028 11306 -11996 11626
rect -11676 11306 -11628 11626
rect -12748 10606 -12715 10926
rect -12395 10606 -12348 10926
rect -13468 9906 -13434 10226
rect -13114 9906 -13068 10226
rect -13468 9698 -13068 9906
rect -12975 10338 -12879 10354
rect -12975 9794 -12959 10338
rect -12895 9794 -12879 10338
rect -12975 9778 -12879 9794
rect -12748 10226 -12348 10606
rect -12256 11038 -12160 11054
rect -12256 10494 -12240 11038
rect -12176 10494 -12160 11038
rect -12256 10478 -12160 10494
rect -12028 10926 -11628 11306
rect -11537 11738 -11441 11754
rect -11537 11194 -11521 11738
rect -11457 11194 -11441 11738
rect -11537 11178 -11441 11194
rect -11308 11626 -10908 12006
rect -10818 12438 -10722 12454
rect -10818 11894 -10802 12438
rect -10738 11894 -10722 12438
rect -10818 11878 -10722 11894
rect -9247 11780 11065 11781
rect -11308 11306 -11277 11626
rect -10957 11306 -10908 11626
rect -12028 10606 -11996 10926
rect -11676 10606 -11628 10926
rect -12748 9906 -12715 10226
rect -12395 9906 -12348 10226
rect -12748 9698 -12348 9906
rect -12256 10338 -12160 10354
rect -12256 9794 -12240 10338
rect -12176 9794 -12160 10338
rect -12256 9778 -12160 9794
rect -12028 10226 -11628 10606
rect -11537 11038 -11441 11054
rect -11537 10494 -11521 11038
rect -11457 10494 -11441 11038
rect -11537 10478 -11441 10494
rect -11308 10926 -10908 11306
rect -10818 11738 -10722 11754
rect -10818 11194 -10802 11738
rect -10738 11194 -10722 11738
rect -10818 11178 -10722 11194
rect -11308 10606 -11277 10926
rect -10957 10606 -10908 10926
rect -12028 9906 -11996 10226
rect -11676 9906 -11628 10226
rect -12028 9698 -11628 9906
rect -11537 10338 -11441 10354
rect -11537 9794 -11521 10338
rect -11457 9794 -11441 10338
rect -11537 9778 -11441 9794
rect -11308 10226 -10908 10606
rect -10818 11038 -10722 11054
rect -10818 10494 -10802 11038
rect -10738 10494 -10722 11038
rect -9247 10808 -9246 11780
rect 11064 10808 11065 11780
rect -9247 10807 11065 10808
rect -10818 10478 -10722 10494
rect -11308 9906 -11277 10226
rect -10957 9906 -10908 10226
rect -11308 9706 -10908 9906
rect -10818 10338 -10722 10354
rect -10818 9794 -10802 10338
rect -10738 9794 -10722 10338
rect -10818 9778 -10722 9794
rect -11308 9698 -10888 9706
rect -17788 9691 -10888 9698
rect -18614 4645 -9482 9691
rect -18616 4643 -9482 4645
rect -18616 4363 -18614 4643
rect -17986 4363 -10123 4643
rect -9495 4363 -9482 4643
rect -18616 4361 -9482 4363
rect -18614 4360 -9482 4361
<< via4 >>
rect -9246 10808 11064 11780
<< mimcap2 >>
rect -21478 23766 -21078 23806
rect -21478 23446 -21438 23766
rect -21118 23446 -21078 23766
rect -21478 23406 -21078 23446
rect -20356 23766 -19956 23806
rect -20356 23446 -20316 23766
rect -19996 23446 -19956 23766
rect -20356 23406 -19956 23446
rect -19234 23766 -18834 23806
rect -19234 23446 -19194 23766
rect -18874 23446 -18834 23766
rect -19234 23406 -18834 23446
rect -18112 23766 -17712 23806
rect -18112 23446 -18072 23766
rect -17752 23446 -17712 23766
rect -18112 23406 -17712 23446
rect -16990 23766 -16590 23806
rect -16990 23446 -16950 23766
rect -16630 23446 -16590 23766
rect -16990 23406 -16590 23446
rect -15868 23766 -15468 23806
rect -15868 23446 -15828 23766
rect -15508 23446 -15468 23766
rect -15868 23406 -15468 23446
rect -14746 23766 -14346 23806
rect -14746 23446 -14706 23766
rect -14386 23446 -14346 23766
rect -14746 23406 -14346 23446
rect -13624 23766 -13224 23806
rect -13624 23446 -13584 23766
rect -13264 23446 -13224 23766
rect -13624 23406 -13224 23446
rect -12502 23766 -12102 23806
rect -12502 23446 -12462 23766
rect -12142 23446 -12102 23766
rect -12502 23406 -12102 23446
rect -11380 23766 -10980 23806
rect -11380 23446 -11340 23766
rect -11020 23446 -10980 23766
rect -11380 23406 -10980 23446
rect -21478 23066 -21078 23106
rect -21478 22746 -21438 23066
rect -21118 22746 -21078 23066
rect -21478 22706 -21078 22746
rect -20356 23066 -19956 23106
rect -20356 22746 -20316 23066
rect -19996 22746 -19956 23066
rect -20356 22706 -19956 22746
rect -19234 23066 -18834 23106
rect -19234 22746 -19194 23066
rect -18874 22746 -18834 23066
rect -19234 22706 -18834 22746
rect -18112 23066 -17712 23106
rect -18112 22746 -18072 23066
rect -17752 22746 -17712 23066
rect -18112 22706 -17712 22746
rect -16990 23066 -16590 23106
rect -16990 22746 -16950 23066
rect -16630 22746 -16590 23066
rect -16990 22706 -16590 22746
rect -15868 23066 -15468 23106
rect -15868 22746 -15828 23066
rect -15508 22746 -15468 23066
rect -15868 22706 -15468 22746
rect -14746 23066 -14346 23106
rect -14746 22746 -14706 23066
rect -14386 22746 -14346 23066
rect -14746 22706 -14346 22746
rect -13624 23066 -13224 23106
rect -13624 22746 -13584 23066
rect -13264 22746 -13224 23066
rect -13624 22706 -13224 22746
rect -12502 23066 -12102 23106
rect -12502 22746 -12462 23066
rect -12142 22746 -12102 23066
rect -12502 22706 -12102 22746
rect -11380 23066 -10980 23106
rect -11380 22746 -11340 23066
rect -11020 22746 -10980 23066
rect -11380 22706 -10980 22746
rect -21478 22366 -21078 22406
rect -21478 22046 -21438 22366
rect -21118 22046 -21078 22366
rect -21478 22006 -21078 22046
rect -20356 22366 -19956 22406
rect -20356 22046 -20316 22366
rect -19996 22046 -19956 22366
rect -20356 22006 -19956 22046
rect -19234 22366 -18834 22406
rect -19234 22046 -19194 22366
rect -18874 22046 -18834 22366
rect -19234 22006 -18834 22046
rect -18112 22366 -17712 22406
rect -18112 22046 -18072 22366
rect -17752 22046 -17712 22366
rect -18112 22006 -17712 22046
rect -16990 22366 -16590 22406
rect -16990 22046 -16950 22366
rect -16630 22046 -16590 22366
rect -16990 22006 -16590 22046
rect -15868 22366 -15468 22406
rect -15868 22046 -15828 22366
rect -15508 22046 -15468 22366
rect -15868 22006 -15468 22046
rect -14746 22366 -14346 22406
rect -14746 22046 -14706 22366
rect -14386 22046 -14346 22366
rect -14746 22006 -14346 22046
rect -13624 22366 -13224 22406
rect -13624 22046 -13584 22366
rect -13264 22046 -13224 22366
rect -13624 22006 -13224 22046
rect -12502 22366 -12102 22406
rect -12502 22046 -12462 22366
rect -12142 22046 -12102 22366
rect -12502 22006 -12102 22046
rect -11380 22366 -10980 22406
rect -11380 22046 -11340 22366
rect -11020 22046 -10980 22366
rect -11380 22006 -10980 22046
rect -21478 21666 -21078 21706
rect -21478 21346 -21438 21666
rect -21118 21346 -21078 21666
rect -21478 21306 -21078 21346
rect -20356 21666 -19956 21706
rect -20356 21346 -20316 21666
rect -19996 21346 -19956 21666
rect -20356 21306 -19956 21346
rect -19234 21666 -18834 21706
rect -19234 21346 -19194 21666
rect -18874 21346 -18834 21666
rect -19234 21306 -18834 21346
rect -18112 21666 -17712 21706
rect -18112 21346 -18072 21666
rect -17752 21346 -17712 21666
rect -18112 21306 -17712 21346
rect -16990 21666 -16590 21706
rect -16990 21346 -16950 21666
rect -16630 21346 -16590 21666
rect -16990 21306 -16590 21346
rect -15868 21666 -15468 21706
rect -15868 21346 -15828 21666
rect -15508 21346 -15468 21666
rect -15868 21306 -15468 21346
rect -14746 21666 -14346 21706
rect -14746 21346 -14706 21666
rect -14386 21346 -14346 21666
rect -14746 21306 -14346 21346
rect -13624 21666 -13224 21706
rect -13624 21346 -13584 21666
rect -13264 21346 -13224 21666
rect -13624 21306 -13224 21346
rect -12502 21666 -12102 21706
rect -12502 21346 -12462 21666
rect -12142 21346 -12102 21666
rect -12502 21306 -12102 21346
rect -11380 21666 -10980 21706
rect -11380 21346 -11340 21666
rect -11020 21346 -10980 21666
rect -11380 21306 -10980 21346
rect -21478 20966 -21078 21006
rect -21478 20646 -21438 20966
rect -21118 20646 -21078 20966
rect -21478 20606 -21078 20646
rect -20356 20966 -19956 21006
rect -20356 20646 -20316 20966
rect -19996 20646 -19956 20966
rect -20356 20606 -19956 20646
rect -19234 20966 -18834 21006
rect -19234 20646 -19194 20966
rect -18874 20646 -18834 20966
rect -19234 20606 -18834 20646
rect -18112 20966 -17712 21006
rect -18112 20646 -18072 20966
rect -17752 20646 -17712 20966
rect -18112 20606 -17712 20646
rect -16990 20966 -16590 21006
rect -16990 20646 -16950 20966
rect -16630 20646 -16590 20966
rect -16990 20606 -16590 20646
rect -15868 20966 -15468 21006
rect -15868 20646 -15828 20966
rect -15508 20646 -15468 20966
rect -15868 20606 -15468 20646
rect -14746 20966 -14346 21006
rect -14746 20646 -14706 20966
rect -14386 20646 -14346 20966
rect -14746 20606 -14346 20646
rect -13624 20966 -13224 21006
rect -13624 20646 -13584 20966
rect -13264 20646 -13224 20966
rect -13624 20606 -13224 20646
rect -12502 20966 -12102 21006
rect -12502 20646 -12462 20966
rect -12142 20646 -12102 20966
rect -12502 20606 -12102 20646
rect -11380 20966 -10980 21006
rect -11380 20646 -11340 20966
rect -11020 20646 -10980 20966
rect -11380 20606 -10980 20646
rect -21478 20266 -21078 20306
rect -21478 19946 -21438 20266
rect -21118 19946 -21078 20266
rect -21478 19906 -21078 19946
rect -20356 20266 -19956 20306
rect -20356 19946 -20316 20266
rect -19996 19946 -19956 20266
rect -20356 19906 -19956 19946
rect -19234 20266 -18834 20306
rect -19234 19946 -19194 20266
rect -18874 19946 -18834 20266
rect -19234 19906 -18834 19946
rect -18112 20266 -17712 20306
rect -18112 19946 -18072 20266
rect -17752 19946 -17712 20266
rect -18112 19906 -17712 19946
rect -16990 20266 -16590 20306
rect -16990 19946 -16950 20266
rect -16630 19946 -16590 20266
rect -16990 19906 -16590 19946
rect -15868 20266 -15468 20306
rect -15868 19946 -15828 20266
rect -15508 19946 -15468 20266
rect -15868 19906 -15468 19946
rect -14746 20266 -14346 20306
rect -14746 19946 -14706 20266
rect -14386 19946 -14346 20266
rect -14746 19906 -14346 19946
rect -13624 20266 -13224 20306
rect -13624 19946 -13584 20266
rect -13264 19946 -13224 20266
rect -13624 19906 -13224 19946
rect -12502 20266 -12102 20306
rect -12502 19946 -12462 20266
rect -12142 19946 -12102 20266
rect -12502 19906 -12102 19946
rect -11380 20266 -10980 20306
rect -11380 19946 -11340 20266
rect -11020 19946 -10980 20266
rect -11380 19906 -10980 19946
rect -21478 19566 -21078 19606
rect -21478 19246 -21438 19566
rect -21118 19246 -21078 19566
rect -21478 19206 -21078 19246
rect -20356 19566 -19956 19606
rect -20356 19246 -20316 19566
rect -19996 19246 -19956 19566
rect -20356 19206 -19956 19246
rect -19234 19566 -18834 19606
rect -19234 19246 -19194 19566
rect -18874 19246 -18834 19566
rect -19234 19206 -18834 19246
rect -18112 19566 -17712 19606
rect -18112 19246 -18072 19566
rect -17752 19246 -17712 19566
rect -18112 19206 -17712 19246
rect -16990 19566 -16590 19606
rect -16990 19246 -16950 19566
rect -16630 19246 -16590 19566
rect -16990 19206 -16590 19246
rect -15868 19566 -15468 19606
rect -15868 19246 -15828 19566
rect -15508 19246 -15468 19566
rect -15868 19206 -15468 19246
rect -14746 19566 -14346 19606
rect -14746 19246 -14706 19566
rect -14386 19246 -14346 19566
rect -14746 19206 -14346 19246
rect -13624 19566 -13224 19606
rect -13624 19246 -13584 19566
rect -13264 19246 -13224 19566
rect -13624 19206 -13224 19246
rect -12502 19566 -12102 19606
rect -12502 19246 -12462 19566
rect -12142 19246 -12102 19566
rect -12502 19206 -12102 19246
rect -11380 19566 -10980 19606
rect -11380 19246 -11340 19566
rect -11020 19246 -10980 19566
rect -11380 19206 -10980 19246
rect -21478 18866 -21078 18906
rect -21478 18546 -21438 18866
rect -21118 18546 -21078 18866
rect -21478 18506 -21078 18546
rect -20356 18866 -19956 18906
rect -20356 18546 -20316 18866
rect -19996 18546 -19956 18866
rect -20356 18506 -19956 18546
rect -19234 18866 -18834 18906
rect -19234 18546 -19194 18866
rect -18874 18546 -18834 18866
rect -19234 18506 -18834 18546
rect -18112 18866 -17712 18906
rect -18112 18546 -18072 18866
rect -17752 18546 -17712 18866
rect -18112 18506 -17712 18546
rect -16990 18866 -16590 18906
rect -16990 18546 -16950 18866
rect -16630 18546 -16590 18866
rect -16990 18506 -16590 18546
rect -15868 18866 -15468 18906
rect -15868 18546 -15828 18866
rect -15508 18546 -15468 18866
rect -15868 18506 -15468 18546
rect -14746 18866 -14346 18906
rect -14746 18546 -14706 18866
rect -14386 18546 -14346 18866
rect -14746 18506 -14346 18546
rect -13624 18866 -13224 18906
rect -13624 18546 -13584 18866
rect -13264 18546 -13224 18866
rect -13624 18506 -13224 18546
rect -12502 18866 -12102 18906
rect -12502 18546 -12462 18866
rect -12142 18546 -12102 18866
rect -12502 18506 -12102 18546
rect -11380 18866 -10980 18906
rect -11380 18546 -11340 18866
rect -11020 18546 -10980 18866
rect -11380 18506 -10980 18546
rect -21478 18166 -21078 18206
rect -21478 17846 -21438 18166
rect -21118 17846 -21078 18166
rect -21478 17806 -21078 17846
rect -20356 18166 -19956 18206
rect -20356 17846 -20316 18166
rect -19996 17846 -19956 18166
rect -20356 17806 -19956 17846
rect -19234 18166 -18834 18206
rect -19234 17846 -19194 18166
rect -18874 17846 -18834 18166
rect -19234 17806 -18834 17846
rect -18112 18166 -17712 18206
rect -18112 17846 -18072 18166
rect -17752 17846 -17712 18166
rect -18112 17806 -17712 17846
rect -16990 18166 -16590 18206
rect -16990 17846 -16950 18166
rect -16630 17846 -16590 18166
rect -16990 17806 -16590 17846
rect -15868 18166 -15468 18206
rect -15868 17846 -15828 18166
rect -15508 17846 -15468 18166
rect -15868 17806 -15468 17846
rect -14746 18166 -14346 18206
rect -14746 17846 -14706 18166
rect -14386 17846 -14346 18166
rect -14746 17806 -14346 17846
rect -13624 18166 -13224 18206
rect -13624 17846 -13584 18166
rect -13264 17846 -13224 18166
rect -13624 17806 -13224 17846
rect -12502 18166 -12102 18206
rect -12502 17846 -12462 18166
rect -12142 17846 -12102 18166
rect -12502 17806 -12102 17846
rect -11380 18166 -10980 18206
rect -11380 17846 -11340 18166
rect -11020 17846 -10980 18166
rect -11380 17806 -10980 17846
rect -21478 17466 -21078 17506
rect -21478 17146 -21438 17466
rect -21118 17146 -21078 17466
rect -21478 17106 -21078 17146
rect -20356 17466 -19956 17506
rect -20356 17146 -20316 17466
rect -19996 17146 -19956 17466
rect -20356 17106 -19956 17146
rect -19234 17466 -18834 17506
rect -19234 17146 -19194 17466
rect -18874 17146 -18834 17466
rect -19234 17106 -18834 17146
rect -18112 17466 -17712 17506
rect -18112 17146 -18072 17466
rect -17752 17146 -17712 17466
rect -18112 17106 -17712 17146
rect -16990 17466 -16590 17506
rect -16990 17146 -16950 17466
rect -16630 17146 -16590 17466
rect -16990 17106 -16590 17146
rect -15868 17466 -15468 17506
rect -15868 17146 -15828 17466
rect -15508 17146 -15468 17466
rect -15868 17106 -15468 17146
rect -14746 17466 -14346 17506
rect -14746 17146 -14706 17466
rect -14386 17146 -14346 17466
rect -14746 17106 -14346 17146
rect -13624 17466 -13224 17506
rect -13624 17146 -13584 17466
rect -13264 17146 -13224 17466
rect -13624 17106 -13224 17146
rect -12502 17466 -12102 17506
rect -12502 17146 -12462 17466
rect -12142 17146 -12102 17466
rect -12502 17106 -12102 17146
rect -11380 17466 -10980 17506
rect -11380 17146 -11340 17466
rect -11020 17146 -10980 17466
rect -11380 17106 -10980 17146
<< mimcap2contact >>
rect -21438 23446 -21118 23766
rect -20316 23446 -19996 23766
rect -19194 23446 -18874 23766
rect -18072 23446 -17752 23766
rect -16950 23446 -16630 23766
rect -15828 23446 -15508 23766
rect -14706 23446 -14386 23766
rect -13584 23446 -13264 23766
rect -12462 23446 -12142 23766
rect -11340 23446 -11020 23766
rect -21438 22746 -21118 23066
rect -20316 22746 -19996 23066
rect -19194 22746 -18874 23066
rect -18072 22746 -17752 23066
rect -16950 22746 -16630 23066
rect -15828 22746 -15508 23066
rect -14706 22746 -14386 23066
rect -13584 22746 -13264 23066
rect -12462 22746 -12142 23066
rect -11340 22746 -11020 23066
rect -21438 22046 -21118 22366
rect -20316 22046 -19996 22366
rect -19194 22046 -18874 22366
rect -18072 22046 -17752 22366
rect -16950 22046 -16630 22366
rect -15828 22046 -15508 22366
rect -14706 22046 -14386 22366
rect -13584 22046 -13264 22366
rect -12462 22046 -12142 22366
rect -11340 22046 -11020 22366
rect -21438 21346 -21118 21666
rect -20316 21346 -19996 21666
rect -19194 21346 -18874 21666
rect -18072 21346 -17752 21666
rect -16950 21346 -16630 21666
rect -15828 21346 -15508 21666
rect -14706 21346 -14386 21666
rect -13584 21346 -13264 21666
rect -12462 21346 -12142 21666
rect -11340 21346 -11020 21666
rect -21438 20646 -21118 20966
rect -20316 20646 -19996 20966
rect -19194 20646 -18874 20966
rect -18072 20646 -17752 20966
rect -16950 20646 -16630 20966
rect -15828 20646 -15508 20966
rect -14706 20646 -14386 20966
rect -13584 20646 -13264 20966
rect -12462 20646 -12142 20966
rect -11340 20646 -11020 20966
rect -21438 19946 -21118 20266
rect -20316 19946 -19996 20266
rect -19194 19946 -18874 20266
rect -18072 19946 -17752 20266
rect -16950 19946 -16630 20266
rect -15828 19946 -15508 20266
rect -14706 19946 -14386 20266
rect -13584 19946 -13264 20266
rect -12462 19946 -12142 20266
rect -11340 19946 -11020 20266
rect -21438 19246 -21118 19566
rect -20316 19246 -19996 19566
rect -19194 19246 -18874 19566
rect -18072 19246 -17752 19566
rect -16950 19246 -16630 19566
rect -15828 19246 -15508 19566
rect -14706 19246 -14386 19566
rect -13584 19246 -13264 19566
rect -12462 19246 -12142 19566
rect -11340 19246 -11020 19566
rect -21438 18546 -21118 18866
rect -20316 18546 -19996 18866
rect -19194 18546 -18874 18866
rect -18072 18546 -17752 18866
rect -16950 18546 -16630 18866
rect -15828 18546 -15508 18866
rect -14706 18546 -14386 18866
rect -13584 18546 -13264 18866
rect -12462 18546 -12142 18866
rect -11340 18546 -11020 18866
rect -21438 17846 -21118 18166
rect -20316 17846 -19996 18166
rect -19194 17846 -18874 18166
rect -18072 17846 -17752 18166
rect -16950 17846 -16630 18166
rect -15828 17846 -15508 18166
rect -14706 17846 -14386 18166
rect -13584 17846 -13264 18166
rect -12462 17846 -12142 18166
rect -11340 17846 -11020 18166
rect -21438 17146 -21118 17466
rect -20316 17146 -19996 17466
rect -19194 17146 -18874 17466
rect -18072 17146 -17752 17466
rect -16950 17146 -16630 17466
rect -15828 17146 -15508 17466
rect -14706 17146 -14386 17466
rect -13584 17146 -13264 17466
rect -12462 17146 -12142 17466
rect -11340 17146 -11020 17466
<< metal5 >>
rect -21532 23950 11082 24225
rect -21532 23766 11238 23950
rect -21532 23446 -21438 23766
rect -21118 23446 -20316 23766
rect -19996 23446 -19194 23766
rect -18874 23446 -18072 23766
rect -17752 23446 -16950 23766
rect -16630 23446 -15828 23766
rect -15508 23446 -14706 23766
rect -14386 23446 -13584 23766
rect -13264 23446 -12462 23766
rect -12142 23446 -11340 23766
rect -11020 23446 11238 23766
rect -21532 23066 11238 23446
rect -21532 22746 -21438 23066
rect -21118 22746 -20316 23066
rect -19996 22746 -19194 23066
rect -18874 22746 -18072 23066
rect -17752 22746 -16950 23066
rect -16630 22746 -15828 23066
rect -15508 22746 -14706 23066
rect -14386 22746 -13584 23066
rect -13264 22746 -12462 23066
rect -12142 22746 -11340 23066
rect -11020 22746 11238 23066
rect -21532 22366 11238 22746
rect -21532 22046 -21438 22366
rect -21118 22046 -20316 22366
rect -19996 22046 -19194 22366
rect -18874 22046 -18072 22366
rect -17752 22046 -16950 22366
rect -16630 22046 -15828 22366
rect -15508 22046 -14706 22366
rect -14386 22046 -13584 22366
rect -13264 22046 -12462 22366
rect -12142 22046 -11340 22366
rect -11020 22046 11238 22366
rect -21532 21666 11238 22046
rect -21532 21346 -21438 21666
rect -21118 21346 -20316 21666
rect -19996 21346 -19194 21666
rect -18874 21346 -18072 21666
rect -17752 21346 -16950 21666
rect -16630 21346 -15828 21666
rect -15508 21346 -14706 21666
rect -14386 21346 -13584 21666
rect -13264 21346 -12462 21666
rect -12142 21346 -11340 21666
rect -11020 21346 11238 21666
rect -21532 20966 11238 21346
rect -21532 20646 -21438 20966
rect -21118 20646 -20316 20966
rect -19996 20646 -19194 20966
rect -18874 20646 -18072 20966
rect -17752 20646 -16950 20966
rect -16630 20646 -15828 20966
rect -15508 20646 -14706 20966
rect -14386 20646 -13584 20966
rect -13264 20646 -12462 20966
rect -12142 20646 -11340 20966
rect -11020 20646 11238 20966
rect -21532 20266 11238 20646
rect -21532 19946 -21438 20266
rect -21118 19946 -20316 20266
rect -19996 19946 -19194 20266
rect -18874 19946 -18072 20266
rect -17752 19946 -16950 20266
rect -16630 19946 -15828 20266
rect -15508 19946 -14706 20266
rect -14386 19946 -13584 20266
rect -13264 19946 -12462 20266
rect -12142 19946 -11340 20266
rect -11020 19946 11238 20266
rect -21532 19566 11238 19946
rect -21532 19246 -21438 19566
rect -21118 19246 -20316 19566
rect -19996 19246 -19194 19566
rect -18874 19246 -18072 19566
rect -17752 19246 -16950 19566
rect -16630 19246 -15828 19566
rect -15508 19246 -14706 19566
rect -14386 19246 -13584 19566
rect -13264 19246 -12462 19566
rect -12142 19246 -11340 19566
rect -11020 19246 11238 19566
rect -21532 18866 11238 19246
rect -21532 18546 -21438 18866
rect -21118 18546 -20316 18866
rect -19996 18546 -19194 18866
rect -18874 18546 -18072 18866
rect -17752 18546 -16950 18866
rect -16630 18546 -15828 18866
rect -15508 18546 -14706 18866
rect -14386 18546 -13584 18866
rect -13264 18546 -12462 18866
rect -12142 18546 -11340 18866
rect -11020 18546 11238 18866
rect -21532 18166 11238 18546
rect -21532 17846 -21438 18166
rect -21118 17846 -20316 18166
rect -19996 17846 -19194 18166
rect -18874 17846 -18072 18166
rect -17752 17846 -16950 18166
rect -16630 17846 -15828 18166
rect -15508 17846 -14706 18166
rect -14386 17846 -13584 18166
rect -13264 17846 -12462 18166
rect -12142 17846 -11340 18166
rect -11020 17846 11238 18166
rect -21532 17466 11238 17846
rect -21532 17146 -21438 17466
rect -21118 17146 -20316 17466
rect -19996 17146 -19194 17466
rect -18874 17146 -18072 17466
rect -17752 17146 -16950 17466
rect -16630 17146 -15828 17466
rect -15508 17146 -14706 17466
rect -14386 17146 -13584 17466
rect -13264 17146 -12462 17466
rect -12142 17146 -11340 17466
rect -11020 17146 11238 17466
rect -21532 11780 11238 17146
rect -21532 10808 -9246 11780
rect 11064 10808 11238 11780
rect -21532 10748 11238 10808
rect -9246 10710 11238 10748
<< res2p85 >>
rect -8934 16850 -8360 20178
rect -8116 16850 -7542 20178
rect -7298 16850 -6724 20178
rect -5662 17260 -5088 21564
rect -4844 17260 -4270 21564
rect -4026 17260 -3452 21564
rect -3208 17260 -2634 21564
rect -754 15194 -180 21502
rect 64 15194 638 21502
rect 882 15194 1456 21502
rect 1700 15194 2274 21502
rect 2518 15194 3092 21502
rect 3336 15194 3910 21502
rect 4154 15194 4728 21502
rect 4972 15194 5546 21502
rect 5790 15194 6364 21502
rect 6608 15194 7182 21502
rect 7426 15194 8000 21502
rect 8244 15194 8818 21502
rect 9062 15194 9636 21502
rect 9880 15194 10454 21502
rect 10698 15194 11272 21502
rect 11516 15194 12090 21502
rect 12334 15194 12908 21502
use pnps  pnps_0
timestamp 1621317379
transform 0 1 30178 -1 0 28812
box 16166 -20906 26884 -11302
<< labels >>
flabel metal1 -19254 8502 -18792 8700 1 FreeSans 1600 0 0 0 porst
port 2 n
flabel metal1 -2858 12824 1810 13500 1 FreeSans 1600 0 0 0 Vbg
port 1 n
flabel metal3 -20266 1000 -19556 1422 1 FreeSans 1600 0 0 0 VDD!
flabel metal2 -21312 4728 -19530 4798 1 FreeSans 800 0 0 0 ampcurrentsource_0/Vq
flabel metal2 -21312 4938 -19530 5008 1 FreeSans 800 0 0 0 ampcurrentsource_0/Vx
flabel locali -20452 5698 -20370 5726 1 FreeSans 800 0 0 0 ampcurrentsource_0/GND!
rlabel via1 -8118 1418 -8072 1462 5 currentmirror_0/Vgate
rlabel metal3 -7396 1062 -7262 1180 5 currentmirror_0/VDD!
flabel metal1 -590 9602 -290 9702 5 FreeSans 1600 0 0 0 currentmirror_0/Vbg
flabel metal2 -590 10202 -390 10302 5 FreeSans 1600 0 0 0 currentmirror_0/Vb
flabel metal2 -590 10802 -390 10902 5 FreeSans 1600 0 0 0 currentmirror_0/Va
flabel metal2 -14560 1438 -14544 1562 5 FreeSans 800 0 0 0 amplifier_0/VDD!
flabel metal2 -13906 4666 -13890 4790 5 FreeSans 800 0 0 0 amplifier_0/Vq
flabel metal2 -13964 6926 -13948 7006 5 FreeSans 800 0 0 0 amplifier_0/Va
flabel metal2 -14736 6786 -14720 6866 5 FreeSans 800 0 0 0 amplifier_0/Vb
flabel metal2 -13230 4370 -13136 4636 5 FreeSans 800 0 0 0 amplifier_0/Vgate
flabel metal2 -14954 4370 -14860 4636 5 FreeSans 800 0 0 0 amplifier_0/Vgate
flabel metal1 -16312 4384 -16278 4476 5 FreeSans 800 0 0 0 amplifier_0/vg
flabel metal2 -12212 1238 -12190 1362 5 FreeSans 800 0 0 0 amplifier_0/Vx
flabel psubdiffcont -17434 5042 -17334 6642 5 FreeSans 800 0 0 0 amplifier_0/GND!
flabel psubdiff -11984 6642 -11784 6742 5 FreeSans 800 180 0 0 amplifier_0/GND!
flabel metal2 884 21500 1454 21932 1 FreeSans 800 90 0 0 bandgapcorev3_0/VbEnd
flabel metal2 1702 14764 2272 15196 1 FreeSans 800 90 0 0 bandgapcorev3_0/VbgEnd
flabel metal2 66 20700 636 21932 1 FreeSans 800 90 0 0 bandgapcorev3_0/VaEnd
flabel metal2 9810 14498 10502 15190 1 FreeSans 1600 90 0 0 bandgapcorev3_0/Vbg
flabel metal2 11440 14492 12144 15196 1 FreeSans 1600 90 0 0 bandgapcorev3_0/Vb
flabel metal1 10622 13926 11326 14498 3 FreeSans 1600 0 0 0 bandgapcorev3_0/Va
flabel metal1 -4846 16332 -3380 16774 3 FreeSans 1600 0 0 0 bandgapcorev3_0/GND!
flabel space 11606 2220 12742 3168 7 FreeSans 1600 0 0 0 bandgapcorev3_0/Vbneg
<< end >>
