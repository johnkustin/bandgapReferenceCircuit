magic
tech sky130A
magscale 1 2
timestamp 1620883575
<< xpolycontact >>
rect -35 376 35 808
rect -35 -808 35 -376
<< xpolyres >>
rect -35 -376 35 376
<< viali >>
rect -19 393 19 790
rect -19 -790 19 -393
<< metal1 >>
rect -25 790 25 802
rect -25 393 -19 790
rect 19 393 25 790
rect -25 381 25 393
rect -25 -393 25 -381
rect -25 -790 -19 -393
rect 19 -790 25 -393
rect -25 -802 25 -790
<< res0p35 >>
rect -37 -378 37 378
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 3.763 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 22.188k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
