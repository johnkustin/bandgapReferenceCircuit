magic
tech sky130A
magscale 1 2
timestamp 1621208350
<< xpolycontact >>
rect -65316 570 -64746 1002
rect -65316 -1002 -64746 -570
rect -64498 570 -63928 1002
rect -64498 -1002 -63928 -570
rect -63680 570 -63110 1002
rect -63680 -1002 -63110 -570
rect -62862 570 -62292 1002
rect -62862 -1002 -62292 -570
rect -62044 570 -61474 1002
rect -62044 -1002 -61474 -570
rect -61226 570 -60656 1002
rect -61226 -1002 -60656 -570
rect -60408 570 -59838 1002
rect -60408 -1002 -59838 -570
rect -59590 570 -59020 1002
rect -59590 -1002 -59020 -570
rect -58772 570 -58202 1002
rect -58772 -1002 -58202 -570
rect -57954 570 -57384 1002
rect -57954 -1002 -57384 -570
rect -57136 570 -56566 1002
rect -57136 -1002 -56566 -570
rect -56318 570 -55748 1002
rect -56318 -1002 -55748 -570
rect -55500 570 -54930 1002
rect -55500 -1002 -54930 -570
rect -54682 570 -54112 1002
rect -54682 -1002 -54112 -570
rect -53864 570 -53294 1002
rect -53864 -1002 -53294 -570
rect -53046 570 -52476 1002
rect -53046 -1002 -52476 -570
rect -52228 570 -51658 1002
rect -52228 -1002 -51658 -570
rect -51410 570 -50840 1002
rect -51410 -1002 -50840 -570
rect -50592 570 -50022 1002
rect -50592 -1002 -50022 -570
rect -49774 570 -49204 1002
rect -49774 -1002 -49204 -570
rect -48956 570 -48386 1002
rect -48956 -1002 -48386 -570
rect -48138 570 -47568 1002
rect -48138 -1002 -47568 -570
rect -47320 570 -46750 1002
rect -47320 -1002 -46750 -570
rect -46502 570 -45932 1002
rect -46502 -1002 -45932 -570
rect -45684 570 -45114 1002
rect -45684 -1002 -45114 -570
rect -44866 570 -44296 1002
rect -44866 -1002 -44296 -570
rect -44048 570 -43478 1002
rect -44048 -1002 -43478 -570
rect -43230 570 -42660 1002
rect -43230 -1002 -42660 -570
rect -42412 570 -41842 1002
rect -42412 -1002 -41842 -570
rect -41594 570 -41024 1002
rect -41594 -1002 -41024 -570
rect -40776 570 -40206 1002
rect -40776 -1002 -40206 -570
rect -39958 570 -39388 1002
rect -39958 -1002 -39388 -570
rect -39140 570 -38570 1002
rect -39140 -1002 -38570 -570
rect -38322 570 -37752 1002
rect -38322 -1002 -37752 -570
rect -37504 570 -36934 1002
rect -37504 -1002 -36934 -570
rect -36686 570 -36116 1002
rect -36686 -1002 -36116 -570
rect -35868 570 -35298 1002
rect -35868 -1002 -35298 -570
rect -35050 570 -34480 1002
rect -35050 -1002 -34480 -570
rect -34232 570 -33662 1002
rect -34232 -1002 -33662 -570
rect -33414 570 -32844 1002
rect -33414 -1002 -32844 -570
rect -32596 570 -32026 1002
rect -32596 -1002 -32026 -570
rect -31778 570 -31208 1002
rect -31778 -1002 -31208 -570
rect -30960 570 -30390 1002
rect -30960 -1002 -30390 -570
rect -30142 570 -29572 1002
rect -30142 -1002 -29572 -570
rect -29324 570 -28754 1002
rect -29324 -1002 -28754 -570
rect -28506 570 -27936 1002
rect -28506 -1002 -27936 -570
rect -27688 570 -27118 1002
rect -27688 -1002 -27118 -570
rect -26870 570 -26300 1002
rect -26870 -1002 -26300 -570
rect -26052 570 -25482 1002
rect -26052 -1002 -25482 -570
rect -25234 570 -24664 1002
rect -25234 -1002 -24664 -570
rect -24416 570 -23846 1002
rect -24416 -1002 -23846 -570
rect -23598 570 -23028 1002
rect -23598 -1002 -23028 -570
rect -22780 570 -22210 1002
rect -22780 -1002 -22210 -570
rect -21962 570 -21392 1002
rect -21962 -1002 -21392 -570
rect -21144 570 -20574 1002
rect -21144 -1002 -20574 -570
rect -20326 570 -19756 1002
rect -20326 -1002 -19756 -570
rect -19508 570 -18938 1002
rect -19508 -1002 -18938 -570
rect -18690 570 -18120 1002
rect -18690 -1002 -18120 -570
rect -17872 570 -17302 1002
rect -17872 -1002 -17302 -570
rect -17054 570 -16484 1002
rect -17054 -1002 -16484 -570
rect -16236 570 -15666 1002
rect -16236 -1002 -15666 -570
rect -15418 570 -14848 1002
rect -15418 -1002 -14848 -570
rect -14600 570 -14030 1002
rect -14600 -1002 -14030 -570
rect -13782 570 -13212 1002
rect -13782 -1002 -13212 -570
rect -12964 570 -12394 1002
rect -12964 -1002 -12394 -570
rect -12146 570 -11576 1002
rect -12146 -1002 -11576 -570
rect -11328 570 -10758 1002
rect -11328 -1002 -10758 -570
rect -10510 570 -9940 1002
rect -10510 -1002 -9940 -570
rect -9692 570 -9122 1002
rect -9692 -1002 -9122 -570
rect -8874 570 -8304 1002
rect -8874 -1002 -8304 -570
rect -8056 570 -7486 1002
rect -8056 -1002 -7486 -570
rect -7238 570 -6668 1002
rect -7238 -1002 -6668 -570
rect -6420 570 -5850 1002
rect -6420 -1002 -5850 -570
rect -5602 570 -5032 1002
rect -5602 -1002 -5032 -570
rect -4784 570 -4214 1002
rect -4784 -1002 -4214 -570
rect -3966 570 -3396 1002
rect -3966 -1002 -3396 -570
rect -3148 570 -2578 1002
rect -3148 -1002 -2578 -570
rect -2330 570 -1760 1002
rect -2330 -1002 -1760 -570
rect -1512 570 -942 1002
rect -1512 -1002 -942 -570
rect -694 570 -124 1002
rect -694 -1002 -124 -570
rect 124 570 694 1002
rect 124 -1002 694 -570
rect 942 570 1512 1002
rect 942 -1002 1512 -570
rect 1760 570 2330 1002
rect 1760 -1002 2330 -570
rect 2578 570 3148 1002
rect 2578 -1002 3148 -570
rect 3396 570 3966 1002
rect 3396 -1002 3966 -570
rect 4214 570 4784 1002
rect 4214 -1002 4784 -570
rect 5032 570 5602 1002
rect 5032 -1002 5602 -570
rect 5850 570 6420 1002
rect 5850 -1002 6420 -570
rect 6668 570 7238 1002
rect 6668 -1002 7238 -570
rect 7486 570 8056 1002
rect 7486 -1002 8056 -570
rect 8304 570 8874 1002
rect 8304 -1002 8874 -570
rect 9122 570 9692 1002
rect 9122 -1002 9692 -570
rect 9940 570 10510 1002
rect 9940 -1002 10510 -570
rect 10758 570 11328 1002
rect 10758 -1002 11328 -570
rect 11576 570 12146 1002
rect 11576 -1002 12146 -570
rect 12394 570 12964 1002
rect 12394 -1002 12964 -570
rect 13212 570 13782 1002
rect 13212 -1002 13782 -570
rect 14030 570 14600 1002
rect 14030 -1002 14600 -570
rect 14848 570 15418 1002
rect 14848 -1002 15418 -570
rect 15666 570 16236 1002
rect 15666 -1002 16236 -570
rect 16484 570 17054 1002
rect 16484 -1002 17054 -570
rect 17302 570 17872 1002
rect 17302 -1002 17872 -570
rect 18120 570 18690 1002
rect 18120 -1002 18690 -570
rect 18938 570 19508 1002
rect 18938 -1002 19508 -570
rect 19756 570 20326 1002
rect 19756 -1002 20326 -570
rect 20574 570 21144 1002
rect 20574 -1002 21144 -570
rect 21392 570 21962 1002
rect 21392 -1002 21962 -570
rect 22210 570 22780 1002
rect 22210 -1002 22780 -570
rect 23028 570 23598 1002
rect 23028 -1002 23598 -570
rect 23846 570 24416 1002
rect 23846 -1002 24416 -570
rect 24664 570 25234 1002
rect 24664 -1002 25234 -570
rect 25482 570 26052 1002
rect 25482 -1002 26052 -570
rect 26300 570 26870 1002
rect 26300 -1002 26870 -570
rect 27118 570 27688 1002
rect 27118 -1002 27688 -570
rect 27936 570 28506 1002
rect 27936 -1002 28506 -570
rect 28754 570 29324 1002
rect 28754 -1002 29324 -570
rect 29572 570 30142 1002
rect 29572 -1002 30142 -570
rect 30390 570 30960 1002
rect 30390 -1002 30960 -570
rect 31208 570 31778 1002
rect 31208 -1002 31778 -570
rect 32026 570 32596 1002
rect 32026 -1002 32596 -570
rect 32844 570 33414 1002
rect 32844 -1002 33414 -570
rect 33662 570 34232 1002
rect 33662 -1002 34232 -570
rect 34480 570 35050 1002
rect 34480 -1002 35050 -570
rect 35298 570 35868 1002
rect 35298 -1002 35868 -570
rect 36116 570 36686 1002
rect 36116 -1002 36686 -570
rect 36934 570 37504 1002
rect 36934 -1002 37504 -570
rect 37752 570 38322 1002
rect 37752 -1002 38322 -570
rect 38570 570 39140 1002
rect 38570 -1002 39140 -570
rect 39388 570 39958 1002
rect 39388 -1002 39958 -570
rect 40206 570 40776 1002
rect 40206 -1002 40776 -570
rect 41024 570 41594 1002
rect 41024 -1002 41594 -570
rect 41842 570 42412 1002
rect 41842 -1002 42412 -570
rect 42660 570 43230 1002
rect 42660 -1002 43230 -570
rect 43478 570 44048 1002
rect 43478 -1002 44048 -570
rect 44296 570 44866 1002
rect 44296 -1002 44866 -570
rect 45114 570 45684 1002
rect 45114 -1002 45684 -570
rect 45932 570 46502 1002
rect 45932 -1002 46502 -570
rect 46750 570 47320 1002
rect 46750 -1002 47320 -570
rect 47568 570 48138 1002
rect 47568 -1002 48138 -570
rect 48386 570 48956 1002
rect 48386 -1002 48956 -570
rect 49204 570 49774 1002
rect 49204 -1002 49774 -570
rect 50022 570 50592 1002
rect 50022 -1002 50592 -570
rect 50840 570 51410 1002
rect 50840 -1002 51410 -570
rect 51658 570 52228 1002
rect 51658 -1002 52228 -570
rect 52476 570 53046 1002
rect 52476 -1002 53046 -570
rect 53294 570 53864 1002
rect 53294 -1002 53864 -570
rect 54112 570 54682 1002
rect 54112 -1002 54682 -570
rect 54930 570 55500 1002
rect 54930 -1002 55500 -570
rect 55748 570 56318 1002
rect 55748 -1002 56318 -570
rect 56566 570 57136 1002
rect 56566 -1002 57136 -570
rect 57384 570 57954 1002
rect 57384 -1002 57954 -570
rect 58202 570 58772 1002
rect 58202 -1002 58772 -570
rect 59020 570 59590 1002
rect 59020 -1002 59590 -570
rect 59838 570 60408 1002
rect 59838 -1002 60408 -570
rect 60656 570 61226 1002
rect 60656 -1002 61226 -570
rect 61474 570 62044 1002
rect 61474 -1002 62044 -570
rect 62292 570 62862 1002
rect 62292 -1002 62862 -570
rect 63110 570 63680 1002
rect 63110 -1002 63680 -570
rect 63928 570 64498 1002
rect 63928 -1002 64498 -570
rect 64746 570 65316 1002
rect 64746 -1002 65316 -570
<< xpolyres >>
rect -65316 -570 -64746 570
rect -64498 -570 -63928 570
rect -63680 -570 -63110 570
rect -62862 -570 -62292 570
rect -62044 -570 -61474 570
rect -61226 -570 -60656 570
rect -60408 -570 -59838 570
rect -59590 -570 -59020 570
rect -58772 -570 -58202 570
rect -57954 -570 -57384 570
rect -57136 -570 -56566 570
rect -56318 -570 -55748 570
rect -55500 -570 -54930 570
rect -54682 -570 -54112 570
rect -53864 -570 -53294 570
rect -53046 -570 -52476 570
rect -52228 -570 -51658 570
rect -51410 -570 -50840 570
rect -50592 -570 -50022 570
rect -49774 -570 -49204 570
rect -48956 -570 -48386 570
rect -48138 -570 -47568 570
rect -47320 -570 -46750 570
rect -46502 -570 -45932 570
rect -45684 -570 -45114 570
rect -44866 -570 -44296 570
rect -44048 -570 -43478 570
rect -43230 -570 -42660 570
rect -42412 -570 -41842 570
rect -41594 -570 -41024 570
rect -40776 -570 -40206 570
rect -39958 -570 -39388 570
rect -39140 -570 -38570 570
rect -38322 -570 -37752 570
rect -37504 -570 -36934 570
rect -36686 -570 -36116 570
rect -35868 -570 -35298 570
rect -35050 -570 -34480 570
rect -34232 -570 -33662 570
rect -33414 -570 -32844 570
rect -32596 -570 -32026 570
rect -31778 -570 -31208 570
rect -30960 -570 -30390 570
rect -30142 -570 -29572 570
rect -29324 -570 -28754 570
rect -28506 -570 -27936 570
rect -27688 -570 -27118 570
rect -26870 -570 -26300 570
rect -26052 -570 -25482 570
rect -25234 -570 -24664 570
rect -24416 -570 -23846 570
rect -23598 -570 -23028 570
rect -22780 -570 -22210 570
rect -21962 -570 -21392 570
rect -21144 -570 -20574 570
rect -20326 -570 -19756 570
rect -19508 -570 -18938 570
rect -18690 -570 -18120 570
rect -17872 -570 -17302 570
rect -17054 -570 -16484 570
rect -16236 -570 -15666 570
rect -15418 -570 -14848 570
rect -14600 -570 -14030 570
rect -13782 -570 -13212 570
rect -12964 -570 -12394 570
rect -12146 -570 -11576 570
rect -11328 -570 -10758 570
rect -10510 -570 -9940 570
rect -9692 -570 -9122 570
rect -8874 -570 -8304 570
rect -8056 -570 -7486 570
rect -7238 -570 -6668 570
rect -6420 -570 -5850 570
rect -5602 -570 -5032 570
rect -4784 -570 -4214 570
rect -3966 -570 -3396 570
rect -3148 -570 -2578 570
rect -2330 -570 -1760 570
rect -1512 -570 -942 570
rect -694 -570 -124 570
rect 124 -570 694 570
rect 942 -570 1512 570
rect 1760 -570 2330 570
rect 2578 -570 3148 570
rect 3396 -570 3966 570
rect 4214 -570 4784 570
rect 5032 -570 5602 570
rect 5850 -570 6420 570
rect 6668 -570 7238 570
rect 7486 -570 8056 570
rect 8304 -570 8874 570
rect 9122 -570 9692 570
rect 9940 -570 10510 570
rect 10758 -570 11328 570
rect 11576 -570 12146 570
rect 12394 -570 12964 570
rect 13212 -570 13782 570
rect 14030 -570 14600 570
rect 14848 -570 15418 570
rect 15666 -570 16236 570
rect 16484 -570 17054 570
rect 17302 -570 17872 570
rect 18120 -570 18690 570
rect 18938 -570 19508 570
rect 19756 -570 20326 570
rect 20574 -570 21144 570
rect 21392 -570 21962 570
rect 22210 -570 22780 570
rect 23028 -570 23598 570
rect 23846 -570 24416 570
rect 24664 -570 25234 570
rect 25482 -570 26052 570
rect 26300 -570 26870 570
rect 27118 -570 27688 570
rect 27936 -570 28506 570
rect 28754 -570 29324 570
rect 29572 -570 30142 570
rect 30390 -570 30960 570
rect 31208 -570 31778 570
rect 32026 -570 32596 570
rect 32844 -570 33414 570
rect 33662 -570 34232 570
rect 34480 -570 35050 570
rect 35298 -570 35868 570
rect 36116 -570 36686 570
rect 36934 -570 37504 570
rect 37752 -570 38322 570
rect 38570 -570 39140 570
rect 39388 -570 39958 570
rect 40206 -570 40776 570
rect 41024 -570 41594 570
rect 41842 -570 42412 570
rect 42660 -570 43230 570
rect 43478 -570 44048 570
rect 44296 -570 44866 570
rect 45114 -570 45684 570
rect 45932 -570 46502 570
rect 46750 -570 47320 570
rect 47568 -570 48138 570
rect 48386 -570 48956 570
rect 49204 -570 49774 570
rect 50022 -570 50592 570
rect 50840 -570 51410 570
rect 51658 -570 52228 570
rect 52476 -570 53046 570
rect 53294 -570 53864 570
rect 54112 -570 54682 570
rect 54930 -570 55500 570
rect 55748 -570 56318 570
rect 56566 -570 57136 570
rect 57384 -570 57954 570
rect 58202 -570 58772 570
rect 59020 -570 59590 570
rect 59838 -570 60408 570
rect 60656 -570 61226 570
rect 61474 -570 62044 570
rect 62292 -570 62862 570
rect 63110 -570 63680 570
rect 63928 -570 64498 570
rect 64746 -570 65316 570
<< viali >>
rect -65300 587 -64762 984
rect -64482 587 -63944 984
rect -63664 587 -63126 984
rect -62846 587 -62308 984
rect -62028 587 -61490 984
rect -61210 587 -60672 984
rect -60392 587 -59854 984
rect -59574 587 -59036 984
rect -58756 587 -58218 984
rect -57938 587 -57400 984
rect -57120 587 -56582 984
rect -56302 587 -55764 984
rect -55484 587 -54946 984
rect -54666 587 -54128 984
rect -53848 587 -53310 984
rect -53030 587 -52492 984
rect -52212 587 -51674 984
rect -51394 587 -50856 984
rect -50576 587 -50038 984
rect -49758 587 -49220 984
rect -48940 587 -48402 984
rect -48122 587 -47584 984
rect -47304 587 -46766 984
rect -46486 587 -45948 984
rect -45668 587 -45130 984
rect -44850 587 -44312 984
rect -44032 587 -43494 984
rect -43214 587 -42676 984
rect -42396 587 -41858 984
rect -41578 587 -41040 984
rect -40760 587 -40222 984
rect -39942 587 -39404 984
rect -39124 587 -38586 984
rect -38306 587 -37768 984
rect -37488 587 -36950 984
rect -36670 587 -36132 984
rect -35852 587 -35314 984
rect -35034 587 -34496 984
rect -34216 587 -33678 984
rect -33398 587 -32860 984
rect -32580 587 -32042 984
rect -31762 587 -31224 984
rect -30944 587 -30406 984
rect -30126 587 -29588 984
rect -29308 587 -28770 984
rect -28490 587 -27952 984
rect -27672 587 -27134 984
rect -26854 587 -26316 984
rect -26036 587 -25498 984
rect -25218 587 -24680 984
rect -24400 587 -23862 984
rect -23582 587 -23044 984
rect -22764 587 -22226 984
rect -21946 587 -21408 984
rect -21128 587 -20590 984
rect -20310 587 -19772 984
rect -19492 587 -18954 984
rect -18674 587 -18136 984
rect -17856 587 -17318 984
rect -17038 587 -16500 984
rect -16220 587 -15682 984
rect -15402 587 -14864 984
rect -14584 587 -14046 984
rect -13766 587 -13228 984
rect -12948 587 -12410 984
rect -12130 587 -11592 984
rect -11312 587 -10774 984
rect -10494 587 -9956 984
rect -9676 587 -9138 984
rect -8858 587 -8320 984
rect -8040 587 -7502 984
rect -7222 587 -6684 984
rect -6404 587 -5866 984
rect -5586 587 -5048 984
rect -4768 587 -4230 984
rect -3950 587 -3412 984
rect -3132 587 -2594 984
rect -2314 587 -1776 984
rect -1496 587 -958 984
rect -678 587 -140 984
rect 140 587 678 984
rect 958 587 1496 984
rect 1776 587 2314 984
rect 2594 587 3132 984
rect 3412 587 3950 984
rect 4230 587 4768 984
rect 5048 587 5586 984
rect 5866 587 6404 984
rect 6684 587 7222 984
rect 7502 587 8040 984
rect 8320 587 8858 984
rect 9138 587 9676 984
rect 9956 587 10494 984
rect 10774 587 11312 984
rect 11592 587 12130 984
rect 12410 587 12948 984
rect 13228 587 13766 984
rect 14046 587 14584 984
rect 14864 587 15402 984
rect 15682 587 16220 984
rect 16500 587 17038 984
rect 17318 587 17856 984
rect 18136 587 18674 984
rect 18954 587 19492 984
rect 19772 587 20310 984
rect 20590 587 21128 984
rect 21408 587 21946 984
rect 22226 587 22764 984
rect 23044 587 23582 984
rect 23862 587 24400 984
rect 24680 587 25218 984
rect 25498 587 26036 984
rect 26316 587 26854 984
rect 27134 587 27672 984
rect 27952 587 28490 984
rect 28770 587 29308 984
rect 29588 587 30126 984
rect 30406 587 30944 984
rect 31224 587 31762 984
rect 32042 587 32580 984
rect 32860 587 33398 984
rect 33678 587 34216 984
rect 34496 587 35034 984
rect 35314 587 35852 984
rect 36132 587 36670 984
rect 36950 587 37488 984
rect 37768 587 38306 984
rect 38586 587 39124 984
rect 39404 587 39942 984
rect 40222 587 40760 984
rect 41040 587 41578 984
rect 41858 587 42396 984
rect 42676 587 43214 984
rect 43494 587 44032 984
rect 44312 587 44850 984
rect 45130 587 45668 984
rect 45948 587 46486 984
rect 46766 587 47304 984
rect 47584 587 48122 984
rect 48402 587 48940 984
rect 49220 587 49758 984
rect 50038 587 50576 984
rect 50856 587 51394 984
rect 51674 587 52212 984
rect 52492 587 53030 984
rect 53310 587 53848 984
rect 54128 587 54666 984
rect 54946 587 55484 984
rect 55764 587 56302 984
rect 56582 587 57120 984
rect 57400 587 57938 984
rect 58218 587 58756 984
rect 59036 587 59574 984
rect 59854 587 60392 984
rect 60672 587 61210 984
rect 61490 587 62028 984
rect 62308 587 62846 984
rect 63126 587 63664 984
rect 63944 587 64482 984
rect 64762 587 65300 984
rect -65300 -984 -64762 -587
rect -64482 -984 -63944 -587
rect -63664 -984 -63126 -587
rect -62846 -984 -62308 -587
rect -62028 -984 -61490 -587
rect -61210 -984 -60672 -587
rect -60392 -984 -59854 -587
rect -59574 -984 -59036 -587
rect -58756 -984 -58218 -587
rect -57938 -984 -57400 -587
rect -57120 -984 -56582 -587
rect -56302 -984 -55764 -587
rect -55484 -984 -54946 -587
rect -54666 -984 -54128 -587
rect -53848 -984 -53310 -587
rect -53030 -984 -52492 -587
rect -52212 -984 -51674 -587
rect -51394 -984 -50856 -587
rect -50576 -984 -50038 -587
rect -49758 -984 -49220 -587
rect -48940 -984 -48402 -587
rect -48122 -984 -47584 -587
rect -47304 -984 -46766 -587
rect -46486 -984 -45948 -587
rect -45668 -984 -45130 -587
rect -44850 -984 -44312 -587
rect -44032 -984 -43494 -587
rect -43214 -984 -42676 -587
rect -42396 -984 -41858 -587
rect -41578 -984 -41040 -587
rect -40760 -984 -40222 -587
rect -39942 -984 -39404 -587
rect -39124 -984 -38586 -587
rect -38306 -984 -37768 -587
rect -37488 -984 -36950 -587
rect -36670 -984 -36132 -587
rect -35852 -984 -35314 -587
rect -35034 -984 -34496 -587
rect -34216 -984 -33678 -587
rect -33398 -984 -32860 -587
rect -32580 -984 -32042 -587
rect -31762 -984 -31224 -587
rect -30944 -984 -30406 -587
rect -30126 -984 -29588 -587
rect -29308 -984 -28770 -587
rect -28490 -984 -27952 -587
rect -27672 -984 -27134 -587
rect -26854 -984 -26316 -587
rect -26036 -984 -25498 -587
rect -25218 -984 -24680 -587
rect -24400 -984 -23862 -587
rect -23582 -984 -23044 -587
rect -22764 -984 -22226 -587
rect -21946 -984 -21408 -587
rect -21128 -984 -20590 -587
rect -20310 -984 -19772 -587
rect -19492 -984 -18954 -587
rect -18674 -984 -18136 -587
rect -17856 -984 -17318 -587
rect -17038 -984 -16500 -587
rect -16220 -984 -15682 -587
rect -15402 -984 -14864 -587
rect -14584 -984 -14046 -587
rect -13766 -984 -13228 -587
rect -12948 -984 -12410 -587
rect -12130 -984 -11592 -587
rect -11312 -984 -10774 -587
rect -10494 -984 -9956 -587
rect -9676 -984 -9138 -587
rect -8858 -984 -8320 -587
rect -8040 -984 -7502 -587
rect -7222 -984 -6684 -587
rect -6404 -984 -5866 -587
rect -5586 -984 -5048 -587
rect -4768 -984 -4230 -587
rect -3950 -984 -3412 -587
rect -3132 -984 -2594 -587
rect -2314 -984 -1776 -587
rect -1496 -984 -958 -587
rect -678 -984 -140 -587
rect 140 -984 678 -587
rect 958 -984 1496 -587
rect 1776 -984 2314 -587
rect 2594 -984 3132 -587
rect 3412 -984 3950 -587
rect 4230 -984 4768 -587
rect 5048 -984 5586 -587
rect 5866 -984 6404 -587
rect 6684 -984 7222 -587
rect 7502 -984 8040 -587
rect 8320 -984 8858 -587
rect 9138 -984 9676 -587
rect 9956 -984 10494 -587
rect 10774 -984 11312 -587
rect 11592 -984 12130 -587
rect 12410 -984 12948 -587
rect 13228 -984 13766 -587
rect 14046 -984 14584 -587
rect 14864 -984 15402 -587
rect 15682 -984 16220 -587
rect 16500 -984 17038 -587
rect 17318 -984 17856 -587
rect 18136 -984 18674 -587
rect 18954 -984 19492 -587
rect 19772 -984 20310 -587
rect 20590 -984 21128 -587
rect 21408 -984 21946 -587
rect 22226 -984 22764 -587
rect 23044 -984 23582 -587
rect 23862 -984 24400 -587
rect 24680 -984 25218 -587
rect 25498 -984 26036 -587
rect 26316 -984 26854 -587
rect 27134 -984 27672 -587
rect 27952 -984 28490 -587
rect 28770 -984 29308 -587
rect 29588 -984 30126 -587
rect 30406 -984 30944 -587
rect 31224 -984 31762 -587
rect 32042 -984 32580 -587
rect 32860 -984 33398 -587
rect 33678 -984 34216 -587
rect 34496 -984 35034 -587
rect 35314 -984 35852 -587
rect 36132 -984 36670 -587
rect 36950 -984 37488 -587
rect 37768 -984 38306 -587
rect 38586 -984 39124 -587
rect 39404 -984 39942 -587
rect 40222 -984 40760 -587
rect 41040 -984 41578 -587
rect 41858 -984 42396 -587
rect 42676 -984 43214 -587
rect 43494 -984 44032 -587
rect 44312 -984 44850 -587
rect 45130 -984 45668 -587
rect 45948 -984 46486 -587
rect 46766 -984 47304 -587
rect 47584 -984 48122 -587
rect 48402 -984 48940 -587
rect 49220 -984 49758 -587
rect 50038 -984 50576 -587
rect 50856 -984 51394 -587
rect 51674 -984 52212 -587
rect 52492 -984 53030 -587
rect 53310 -984 53848 -587
rect 54128 -984 54666 -587
rect 54946 -984 55484 -587
rect 55764 -984 56302 -587
rect 56582 -984 57120 -587
rect 57400 -984 57938 -587
rect 58218 -984 58756 -587
rect 59036 -984 59574 -587
rect 59854 -984 60392 -587
rect 60672 -984 61210 -587
rect 61490 -984 62028 -587
rect 62308 -984 62846 -587
rect 63126 -984 63664 -587
rect 63944 -984 64482 -587
rect 64762 -984 65300 -587
<< metal1 >>
rect -65312 984 -64750 990
rect -65312 587 -65300 984
rect -64762 587 -64750 984
rect -65312 581 -64750 587
rect -64494 984 -63932 990
rect -64494 587 -64482 984
rect -63944 587 -63932 984
rect -64494 581 -63932 587
rect -63676 984 -63114 990
rect -63676 587 -63664 984
rect -63126 587 -63114 984
rect -63676 581 -63114 587
rect -62858 984 -62296 990
rect -62858 587 -62846 984
rect -62308 587 -62296 984
rect -62858 581 -62296 587
rect -62040 984 -61478 990
rect -62040 587 -62028 984
rect -61490 587 -61478 984
rect -62040 581 -61478 587
rect -61222 984 -60660 990
rect -61222 587 -61210 984
rect -60672 587 -60660 984
rect -61222 581 -60660 587
rect -60404 984 -59842 990
rect -60404 587 -60392 984
rect -59854 587 -59842 984
rect -60404 581 -59842 587
rect -59586 984 -59024 990
rect -59586 587 -59574 984
rect -59036 587 -59024 984
rect -59586 581 -59024 587
rect -58768 984 -58206 990
rect -58768 587 -58756 984
rect -58218 587 -58206 984
rect -58768 581 -58206 587
rect -57950 984 -57388 990
rect -57950 587 -57938 984
rect -57400 587 -57388 984
rect -57950 581 -57388 587
rect -57132 984 -56570 990
rect -57132 587 -57120 984
rect -56582 587 -56570 984
rect -57132 581 -56570 587
rect -56314 984 -55752 990
rect -56314 587 -56302 984
rect -55764 587 -55752 984
rect -56314 581 -55752 587
rect -55496 984 -54934 990
rect -55496 587 -55484 984
rect -54946 587 -54934 984
rect -55496 581 -54934 587
rect -54678 984 -54116 990
rect -54678 587 -54666 984
rect -54128 587 -54116 984
rect -54678 581 -54116 587
rect -53860 984 -53298 990
rect -53860 587 -53848 984
rect -53310 587 -53298 984
rect -53860 581 -53298 587
rect -53042 984 -52480 990
rect -53042 587 -53030 984
rect -52492 587 -52480 984
rect -53042 581 -52480 587
rect -52224 984 -51662 990
rect -52224 587 -52212 984
rect -51674 587 -51662 984
rect -52224 581 -51662 587
rect -51406 984 -50844 990
rect -51406 587 -51394 984
rect -50856 587 -50844 984
rect -51406 581 -50844 587
rect -50588 984 -50026 990
rect -50588 587 -50576 984
rect -50038 587 -50026 984
rect -50588 581 -50026 587
rect -49770 984 -49208 990
rect -49770 587 -49758 984
rect -49220 587 -49208 984
rect -49770 581 -49208 587
rect -48952 984 -48390 990
rect -48952 587 -48940 984
rect -48402 587 -48390 984
rect -48952 581 -48390 587
rect -48134 984 -47572 990
rect -48134 587 -48122 984
rect -47584 587 -47572 984
rect -48134 581 -47572 587
rect -47316 984 -46754 990
rect -47316 587 -47304 984
rect -46766 587 -46754 984
rect -47316 581 -46754 587
rect -46498 984 -45936 990
rect -46498 587 -46486 984
rect -45948 587 -45936 984
rect -46498 581 -45936 587
rect -45680 984 -45118 990
rect -45680 587 -45668 984
rect -45130 587 -45118 984
rect -45680 581 -45118 587
rect -44862 984 -44300 990
rect -44862 587 -44850 984
rect -44312 587 -44300 984
rect -44862 581 -44300 587
rect -44044 984 -43482 990
rect -44044 587 -44032 984
rect -43494 587 -43482 984
rect -44044 581 -43482 587
rect -43226 984 -42664 990
rect -43226 587 -43214 984
rect -42676 587 -42664 984
rect -43226 581 -42664 587
rect -42408 984 -41846 990
rect -42408 587 -42396 984
rect -41858 587 -41846 984
rect -42408 581 -41846 587
rect -41590 984 -41028 990
rect -41590 587 -41578 984
rect -41040 587 -41028 984
rect -41590 581 -41028 587
rect -40772 984 -40210 990
rect -40772 587 -40760 984
rect -40222 587 -40210 984
rect -40772 581 -40210 587
rect -39954 984 -39392 990
rect -39954 587 -39942 984
rect -39404 587 -39392 984
rect -39954 581 -39392 587
rect -39136 984 -38574 990
rect -39136 587 -39124 984
rect -38586 587 -38574 984
rect -39136 581 -38574 587
rect -38318 984 -37756 990
rect -38318 587 -38306 984
rect -37768 587 -37756 984
rect -38318 581 -37756 587
rect -37500 984 -36938 990
rect -37500 587 -37488 984
rect -36950 587 -36938 984
rect -37500 581 -36938 587
rect -36682 984 -36120 990
rect -36682 587 -36670 984
rect -36132 587 -36120 984
rect -36682 581 -36120 587
rect -35864 984 -35302 990
rect -35864 587 -35852 984
rect -35314 587 -35302 984
rect -35864 581 -35302 587
rect -35046 984 -34484 990
rect -35046 587 -35034 984
rect -34496 587 -34484 984
rect -35046 581 -34484 587
rect -34228 984 -33666 990
rect -34228 587 -34216 984
rect -33678 587 -33666 984
rect -34228 581 -33666 587
rect -33410 984 -32848 990
rect -33410 587 -33398 984
rect -32860 587 -32848 984
rect -33410 581 -32848 587
rect -32592 984 -32030 990
rect -32592 587 -32580 984
rect -32042 587 -32030 984
rect -32592 581 -32030 587
rect -31774 984 -31212 990
rect -31774 587 -31762 984
rect -31224 587 -31212 984
rect -31774 581 -31212 587
rect -30956 984 -30394 990
rect -30956 587 -30944 984
rect -30406 587 -30394 984
rect -30956 581 -30394 587
rect -30138 984 -29576 990
rect -30138 587 -30126 984
rect -29588 587 -29576 984
rect -30138 581 -29576 587
rect -29320 984 -28758 990
rect -29320 587 -29308 984
rect -28770 587 -28758 984
rect -29320 581 -28758 587
rect -28502 984 -27940 990
rect -28502 587 -28490 984
rect -27952 587 -27940 984
rect -28502 581 -27940 587
rect -27684 984 -27122 990
rect -27684 587 -27672 984
rect -27134 587 -27122 984
rect -27684 581 -27122 587
rect -26866 984 -26304 990
rect -26866 587 -26854 984
rect -26316 587 -26304 984
rect -26866 581 -26304 587
rect -26048 984 -25486 990
rect -26048 587 -26036 984
rect -25498 587 -25486 984
rect -26048 581 -25486 587
rect -25230 984 -24668 990
rect -25230 587 -25218 984
rect -24680 587 -24668 984
rect -25230 581 -24668 587
rect -24412 984 -23850 990
rect -24412 587 -24400 984
rect -23862 587 -23850 984
rect -24412 581 -23850 587
rect -23594 984 -23032 990
rect -23594 587 -23582 984
rect -23044 587 -23032 984
rect -23594 581 -23032 587
rect -22776 984 -22214 990
rect -22776 587 -22764 984
rect -22226 587 -22214 984
rect -22776 581 -22214 587
rect -21958 984 -21396 990
rect -21958 587 -21946 984
rect -21408 587 -21396 984
rect -21958 581 -21396 587
rect -21140 984 -20578 990
rect -21140 587 -21128 984
rect -20590 587 -20578 984
rect -21140 581 -20578 587
rect -20322 984 -19760 990
rect -20322 587 -20310 984
rect -19772 587 -19760 984
rect -20322 581 -19760 587
rect -19504 984 -18942 990
rect -19504 587 -19492 984
rect -18954 587 -18942 984
rect -19504 581 -18942 587
rect -18686 984 -18124 990
rect -18686 587 -18674 984
rect -18136 587 -18124 984
rect -18686 581 -18124 587
rect -17868 984 -17306 990
rect -17868 587 -17856 984
rect -17318 587 -17306 984
rect -17868 581 -17306 587
rect -17050 984 -16488 990
rect -17050 587 -17038 984
rect -16500 587 -16488 984
rect -17050 581 -16488 587
rect -16232 984 -15670 990
rect -16232 587 -16220 984
rect -15682 587 -15670 984
rect -16232 581 -15670 587
rect -15414 984 -14852 990
rect -15414 587 -15402 984
rect -14864 587 -14852 984
rect -15414 581 -14852 587
rect -14596 984 -14034 990
rect -14596 587 -14584 984
rect -14046 587 -14034 984
rect -14596 581 -14034 587
rect -13778 984 -13216 990
rect -13778 587 -13766 984
rect -13228 587 -13216 984
rect -13778 581 -13216 587
rect -12960 984 -12398 990
rect -12960 587 -12948 984
rect -12410 587 -12398 984
rect -12960 581 -12398 587
rect -12142 984 -11580 990
rect -12142 587 -12130 984
rect -11592 587 -11580 984
rect -12142 581 -11580 587
rect -11324 984 -10762 990
rect -11324 587 -11312 984
rect -10774 587 -10762 984
rect -11324 581 -10762 587
rect -10506 984 -9944 990
rect -10506 587 -10494 984
rect -9956 587 -9944 984
rect -10506 581 -9944 587
rect -9688 984 -9126 990
rect -9688 587 -9676 984
rect -9138 587 -9126 984
rect -9688 581 -9126 587
rect -8870 984 -8308 990
rect -8870 587 -8858 984
rect -8320 587 -8308 984
rect -8870 581 -8308 587
rect -8052 984 -7490 990
rect -8052 587 -8040 984
rect -7502 587 -7490 984
rect -8052 581 -7490 587
rect -7234 984 -6672 990
rect -7234 587 -7222 984
rect -6684 587 -6672 984
rect -7234 581 -6672 587
rect -6416 984 -5854 990
rect -6416 587 -6404 984
rect -5866 587 -5854 984
rect -6416 581 -5854 587
rect -5598 984 -5036 990
rect -5598 587 -5586 984
rect -5048 587 -5036 984
rect -5598 581 -5036 587
rect -4780 984 -4218 990
rect -4780 587 -4768 984
rect -4230 587 -4218 984
rect -4780 581 -4218 587
rect -3962 984 -3400 990
rect -3962 587 -3950 984
rect -3412 587 -3400 984
rect -3962 581 -3400 587
rect -3144 984 -2582 990
rect -3144 587 -3132 984
rect -2594 587 -2582 984
rect -3144 581 -2582 587
rect -2326 984 -1764 990
rect -2326 587 -2314 984
rect -1776 587 -1764 984
rect -2326 581 -1764 587
rect -1508 984 -946 990
rect -1508 587 -1496 984
rect -958 587 -946 984
rect -1508 581 -946 587
rect -690 984 -128 990
rect -690 587 -678 984
rect -140 587 -128 984
rect -690 581 -128 587
rect 128 984 690 990
rect 128 587 140 984
rect 678 587 690 984
rect 128 581 690 587
rect 946 984 1508 990
rect 946 587 958 984
rect 1496 587 1508 984
rect 946 581 1508 587
rect 1764 984 2326 990
rect 1764 587 1776 984
rect 2314 587 2326 984
rect 1764 581 2326 587
rect 2582 984 3144 990
rect 2582 587 2594 984
rect 3132 587 3144 984
rect 2582 581 3144 587
rect 3400 984 3962 990
rect 3400 587 3412 984
rect 3950 587 3962 984
rect 3400 581 3962 587
rect 4218 984 4780 990
rect 4218 587 4230 984
rect 4768 587 4780 984
rect 4218 581 4780 587
rect 5036 984 5598 990
rect 5036 587 5048 984
rect 5586 587 5598 984
rect 5036 581 5598 587
rect 5854 984 6416 990
rect 5854 587 5866 984
rect 6404 587 6416 984
rect 5854 581 6416 587
rect 6672 984 7234 990
rect 6672 587 6684 984
rect 7222 587 7234 984
rect 6672 581 7234 587
rect 7490 984 8052 990
rect 7490 587 7502 984
rect 8040 587 8052 984
rect 7490 581 8052 587
rect 8308 984 8870 990
rect 8308 587 8320 984
rect 8858 587 8870 984
rect 8308 581 8870 587
rect 9126 984 9688 990
rect 9126 587 9138 984
rect 9676 587 9688 984
rect 9126 581 9688 587
rect 9944 984 10506 990
rect 9944 587 9956 984
rect 10494 587 10506 984
rect 9944 581 10506 587
rect 10762 984 11324 990
rect 10762 587 10774 984
rect 11312 587 11324 984
rect 10762 581 11324 587
rect 11580 984 12142 990
rect 11580 587 11592 984
rect 12130 587 12142 984
rect 11580 581 12142 587
rect 12398 984 12960 990
rect 12398 587 12410 984
rect 12948 587 12960 984
rect 12398 581 12960 587
rect 13216 984 13778 990
rect 13216 587 13228 984
rect 13766 587 13778 984
rect 13216 581 13778 587
rect 14034 984 14596 990
rect 14034 587 14046 984
rect 14584 587 14596 984
rect 14034 581 14596 587
rect 14852 984 15414 990
rect 14852 587 14864 984
rect 15402 587 15414 984
rect 14852 581 15414 587
rect 15670 984 16232 990
rect 15670 587 15682 984
rect 16220 587 16232 984
rect 15670 581 16232 587
rect 16488 984 17050 990
rect 16488 587 16500 984
rect 17038 587 17050 984
rect 16488 581 17050 587
rect 17306 984 17868 990
rect 17306 587 17318 984
rect 17856 587 17868 984
rect 17306 581 17868 587
rect 18124 984 18686 990
rect 18124 587 18136 984
rect 18674 587 18686 984
rect 18124 581 18686 587
rect 18942 984 19504 990
rect 18942 587 18954 984
rect 19492 587 19504 984
rect 18942 581 19504 587
rect 19760 984 20322 990
rect 19760 587 19772 984
rect 20310 587 20322 984
rect 19760 581 20322 587
rect 20578 984 21140 990
rect 20578 587 20590 984
rect 21128 587 21140 984
rect 20578 581 21140 587
rect 21396 984 21958 990
rect 21396 587 21408 984
rect 21946 587 21958 984
rect 21396 581 21958 587
rect 22214 984 22776 990
rect 22214 587 22226 984
rect 22764 587 22776 984
rect 22214 581 22776 587
rect 23032 984 23594 990
rect 23032 587 23044 984
rect 23582 587 23594 984
rect 23032 581 23594 587
rect 23850 984 24412 990
rect 23850 587 23862 984
rect 24400 587 24412 984
rect 23850 581 24412 587
rect 24668 984 25230 990
rect 24668 587 24680 984
rect 25218 587 25230 984
rect 24668 581 25230 587
rect 25486 984 26048 990
rect 25486 587 25498 984
rect 26036 587 26048 984
rect 25486 581 26048 587
rect 26304 984 26866 990
rect 26304 587 26316 984
rect 26854 587 26866 984
rect 26304 581 26866 587
rect 27122 984 27684 990
rect 27122 587 27134 984
rect 27672 587 27684 984
rect 27122 581 27684 587
rect 27940 984 28502 990
rect 27940 587 27952 984
rect 28490 587 28502 984
rect 27940 581 28502 587
rect 28758 984 29320 990
rect 28758 587 28770 984
rect 29308 587 29320 984
rect 28758 581 29320 587
rect 29576 984 30138 990
rect 29576 587 29588 984
rect 30126 587 30138 984
rect 29576 581 30138 587
rect 30394 984 30956 990
rect 30394 587 30406 984
rect 30944 587 30956 984
rect 30394 581 30956 587
rect 31212 984 31774 990
rect 31212 587 31224 984
rect 31762 587 31774 984
rect 31212 581 31774 587
rect 32030 984 32592 990
rect 32030 587 32042 984
rect 32580 587 32592 984
rect 32030 581 32592 587
rect 32848 984 33410 990
rect 32848 587 32860 984
rect 33398 587 33410 984
rect 32848 581 33410 587
rect 33666 984 34228 990
rect 33666 587 33678 984
rect 34216 587 34228 984
rect 33666 581 34228 587
rect 34484 984 35046 990
rect 34484 587 34496 984
rect 35034 587 35046 984
rect 34484 581 35046 587
rect 35302 984 35864 990
rect 35302 587 35314 984
rect 35852 587 35864 984
rect 35302 581 35864 587
rect 36120 984 36682 990
rect 36120 587 36132 984
rect 36670 587 36682 984
rect 36120 581 36682 587
rect 36938 984 37500 990
rect 36938 587 36950 984
rect 37488 587 37500 984
rect 36938 581 37500 587
rect 37756 984 38318 990
rect 37756 587 37768 984
rect 38306 587 38318 984
rect 37756 581 38318 587
rect 38574 984 39136 990
rect 38574 587 38586 984
rect 39124 587 39136 984
rect 38574 581 39136 587
rect 39392 984 39954 990
rect 39392 587 39404 984
rect 39942 587 39954 984
rect 39392 581 39954 587
rect 40210 984 40772 990
rect 40210 587 40222 984
rect 40760 587 40772 984
rect 40210 581 40772 587
rect 41028 984 41590 990
rect 41028 587 41040 984
rect 41578 587 41590 984
rect 41028 581 41590 587
rect 41846 984 42408 990
rect 41846 587 41858 984
rect 42396 587 42408 984
rect 41846 581 42408 587
rect 42664 984 43226 990
rect 42664 587 42676 984
rect 43214 587 43226 984
rect 42664 581 43226 587
rect 43482 984 44044 990
rect 43482 587 43494 984
rect 44032 587 44044 984
rect 43482 581 44044 587
rect 44300 984 44862 990
rect 44300 587 44312 984
rect 44850 587 44862 984
rect 44300 581 44862 587
rect 45118 984 45680 990
rect 45118 587 45130 984
rect 45668 587 45680 984
rect 45118 581 45680 587
rect 45936 984 46498 990
rect 45936 587 45948 984
rect 46486 587 46498 984
rect 45936 581 46498 587
rect 46754 984 47316 990
rect 46754 587 46766 984
rect 47304 587 47316 984
rect 46754 581 47316 587
rect 47572 984 48134 990
rect 47572 587 47584 984
rect 48122 587 48134 984
rect 47572 581 48134 587
rect 48390 984 48952 990
rect 48390 587 48402 984
rect 48940 587 48952 984
rect 48390 581 48952 587
rect 49208 984 49770 990
rect 49208 587 49220 984
rect 49758 587 49770 984
rect 49208 581 49770 587
rect 50026 984 50588 990
rect 50026 587 50038 984
rect 50576 587 50588 984
rect 50026 581 50588 587
rect 50844 984 51406 990
rect 50844 587 50856 984
rect 51394 587 51406 984
rect 50844 581 51406 587
rect 51662 984 52224 990
rect 51662 587 51674 984
rect 52212 587 52224 984
rect 51662 581 52224 587
rect 52480 984 53042 990
rect 52480 587 52492 984
rect 53030 587 53042 984
rect 52480 581 53042 587
rect 53298 984 53860 990
rect 53298 587 53310 984
rect 53848 587 53860 984
rect 53298 581 53860 587
rect 54116 984 54678 990
rect 54116 587 54128 984
rect 54666 587 54678 984
rect 54116 581 54678 587
rect 54934 984 55496 990
rect 54934 587 54946 984
rect 55484 587 55496 984
rect 54934 581 55496 587
rect 55752 984 56314 990
rect 55752 587 55764 984
rect 56302 587 56314 984
rect 55752 581 56314 587
rect 56570 984 57132 990
rect 56570 587 56582 984
rect 57120 587 57132 984
rect 56570 581 57132 587
rect 57388 984 57950 990
rect 57388 587 57400 984
rect 57938 587 57950 984
rect 57388 581 57950 587
rect 58206 984 58768 990
rect 58206 587 58218 984
rect 58756 587 58768 984
rect 58206 581 58768 587
rect 59024 984 59586 990
rect 59024 587 59036 984
rect 59574 587 59586 984
rect 59024 581 59586 587
rect 59842 984 60404 990
rect 59842 587 59854 984
rect 60392 587 60404 984
rect 59842 581 60404 587
rect 60660 984 61222 990
rect 60660 587 60672 984
rect 61210 587 61222 984
rect 60660 581 61222 587
rect 61478 984 62040 990
rect 61478 587 61490 984
rect 62028 587 62040 984
rect 61478 581 62040 587
rect 62296 984 62858 990
rect 62296 587 62308 984
rect 62846 587 62858 984
rect 62296 581 62858 587
rect 63114 984 63676 990
rect 63114 587 63126 984
rect 63664 587 63676 984
rect 63114 581 63676 587
rect 63932 984 64494 990
rect 63932 587 63944 984
rect 64482 587 64494 984
rect 63932 581 64494 587
rect 64750 984 65312 990
rect 64750 587 64762 984
rect 65300 587 65312 984
rect 64750 581 65312 587
rect -65312 -587 -64750 -581
rect -65312 -984 -65300 -587
rect -64762 -984 -64750 -587
rect -65312 -990 -64750 -984
rect -64494 -587 -63932 -581
rect -64494 -984 -64482 -587
rect -63944 -984 -63932 -587
rect -64494 -990 -63932 -984
rect -63676 -587 -63114 -581
rect -63676 -984 -63664 -587
rect -63126 -984 -63114 -587
rect -63676 -990 -63114 -984
rect -62858 -587 -62296 -581
rect -62858 -984 -62846 -587
rect -62308 -984 -62296 -587
rect -62858 -990 -62296 -984
rect -62040 -587 -61478 -581
rect -62040 -984 -62028 -587
rect -61490 -984 -61478 -587
rect -62040 -990 -61478 -984
rect -61222 -587 -60660 -581
rect -61222 -984 -61210 -587
rect -60672 -984 -60660 -587
rect -61222 -990 -60660 -984
rect -60404 -587 -59842 -581
rect -60404 -984 -60392 -587
rect -59854 -984 -59842 -587
rect -60404 -990 -59842 -984
rect -59586 -587 -59024 -581
rect -59586 -984 -59574 -587
rect -59036 -984 -59024 -587
rect -59586 -990 -59024 -984
rect -58768 -587 -58206 -581
rect -58768 -984 -58756 -587
rect -58218 -984 -58206 -587
rect -58768 -990 -58206 -984
rect -57950 -587 -57388 -581
rect -57950 -984 -57938 -587
rect -57400 -984 -57388 -587
rect -57950 -990 -57388 -984
rect -57132 -587 -56570 -581
rect -57132 -984 -57120 -587
rect -56582 -984 -56570 -587
rect -57132 -990 -56570 -984
rect -56314 -587 -55752 -581
rect -56314 -984 -56302 -587
rect -55764 -984 -55752 -587
rect -56314 -990 -55752 -984
rect -55496 -587 -54934 -581
rect -55496 -984 -55484 -587
rect -54946 -984 -54934 -587
rect -55496 -990 -54934 -984
rect -54678 -587 -54116 -581
rect -54678 -984 -54666 -587
rect -54128 -984 -54116 -587
rect -54678 -990 -54116 -984
rect -53860 -587 -53298 -581
rect -53860 -984 -53848 -587
rect -53310 -984 -53298 -587
rect -53860 -990 -53298 -984
rect -53042 -587 -52480 -581
rect -53042 -984 -53030 -587
rect -52492 -984 -52480 -587
rect -53042 -990 -52480 -984
rect -52224 -587 -51662 -581
rect -52224 -984 -52212 -587
rect -51674 -984 -51662 -587
rect -52224 -990 -51662 -984
rect -51406 -587 -50844 -581
rect -51406 -984 -51394 -587
rect -50856 -984 -50844 -587
rect -51406 -990 -50844 -984
rect -50588 -587 -50026 -581
rect -50588 -984 -50576 -587
rect -50038 -984 -50026 -587
rect -50588 -990 -50026 -984
rect -49770 -587 -49208 -581
rect -49770 -984 -49758 -587
rect -49220 -984 -49208 -587
rect -49770 -990 -49208 -984
rect -48952 -587 -48390 -581
rect -48952 -984 -48940 -587
rect -48402 -984 -48390 -587
rect -48952 -990 -48390 -984
rect -48134 -587 -47572 -581
rect -48134 -984 -48122 -587
rect -47584 -984 -47572 -587
rect -48134 -990 -47572 -984
rect -47316 -587 -46754 -581
rect -47316 -984 -47304 -587
rect -46766 -984 -46754 -587
rect -47316 -990 -46754 -984
rect -46498 -587 -45936 -581
rect -46498 -984 -46486 -587
rect -45948 -984 -45936 -587
rect -46498 -990 -45936 -984
rect -45680 -587 -45118 -581
rect -45680 -984 -45668 -587
rect -45130 -984 -45118 -587
rect -45680 -990 -45118 -984
rect -44862 -587 -44300 -581
rect -44862 -984 -44850 -587
rect -44312 -984 -44300 -587
rect -44862 -990 -44300 -984
rect -44044 -587 -43482 -581
rect -44044 -984 -44032 -587
rect -43494 -984 -43482 -587
rect -44044 -990 -43482 -984
rect -43226 -587 -42664 -581
rect -43226 -984 -43214 -587
rect -42676 -984 -42664 -587
rect -43226 -990 -42664 -984
rect -42408 -587 -41846 -581
rect -42408 -984 -42396 -587
rect -41858 -984 -41846 -587
rect -42408 -990 -41846 -984
rect -41590 -587 -41028 -581
rect -41590 -984 -41578 -587
rect -41040 -984 -41028 -587
rect -41590 -990 -41028 -984
rect -40772 -587 -40210 -581
rect -40772 -984 -40760 -587
rect -40222 -984 -40210 -587
rect -40772 -990 -40210 -984
rect -39954 -587 -39392 -581
rect -39954 -984 -39942 -587
rect -39404 -984 -39392 -587
rect -39954 -990 -39392 -984
rect -39136 -587 -38574 -581
rect -39136 -984 -39124 -587
rect -38586 -984 -38574 -587
rect -39136 -990 -38574 -984
rect -38318 -587 -37756 -581
rect -38318 -984 -38306 -587
rect -37768 -984 -37756 -587
rect -38318 -990 -37756 -984
rect -37500 -587 -36938 -581
rect -37500 -984 -37488 -587
rect -36950 -984 -36938 -587
rect -37500 -990 -36938 -984
rect -36682 -587 -36120 -581
rect -36682 -984 -36670 -587
rect -36132 -984 -36120 -587
rect -36682 -990 -36120 -984
rect -35864 -587 -35302 -581
rect -35864 -984 -35852 -587
rect -35314 -984 -35302 -587
rect -35864 -990 -35302 -984
rect -35046 -587 -34484 -581
rect -35046 -984 -35034 -587
rect -34496 -984 -34484 -587
rect -35046 -990 -34484 -984
rect -34228 -587 -33666 -581
rect -34228 -984 -34216 -587
rect -33678 -984 -33666 -587
rect -34228 -990 -33666 -984
rect -33410 -587 -32848 -581
rect -33410 -984 -33398 -587
rect -32860 -984 -32848 -587
rect -33410 -990 -32848 -984
rect -32592 -587 -32030 -581
rect -32592 -984 -32580 -587
rect -32042 -984 -32030 -587
rect -32592 -990 -32030 -984
rect -31774 -587 -31212 -581
rect -31774 -984 -31762 -587
rect -31224 -984 -31212 -587
rect -31774 -990 -31212 -984
rect -30956 -587 -30394 -581
rect -30956 -984 -30944 -587
rect -30406 -984 -30394 -587
rect -30956 -990 -30394 -984
rect -30138 -587 -29576 -581
rect -30138 -984 -30126 -587
rect -29588 -984 -29576 -587
rect -30138 -990 -29576 -984
rect -29320 -587 -28758 -581
rect -29320 -984 -29308 -587
rect -28770 -984 -28758 -587
rect -29320 -990 -28758 -984
rect -28502 -587 -27940 -581
rect -28502 -984 -28490 -587
rect -27952 -984 -27940 -587
rect -28502 -990 -27940 -984
rect -27684 -587 -27122 -581
rect -27684 -984 -27672 -587
rect -27134 -984 -27122 -587
rect -27684 -990 -27122 -984
rect -26866 -587 -26304 -581
rect -26866 -984 -26854 -587
rect -26316 -984 -26304 -587
rect -26866 -990 -26304 -984
rect -26048 -587 -25486 -581
rect -26048 -984 -26036 -587
rect -25498 -984 -25486 -587
rect -26048 -990 -25486 -984
rect -25230 -587 -24668 -581
rect -25230 -984 -25218 -587
rect -24680 -984 -24668 -587
rect -25230 -990 -24668 -984
rect -24412 -587 -23850 -581
rect -24412 -984 -24400 -587
rect -23862 -984 -23850 -587
rect -24412 -990 -23850 -984
rect -23594 -587 -23032 -581
rect -23594 -984 -23582 -587
rect -23044 -984 -23032 -587
rect -23594 -990 -23032 -984
rect -22776 -587 -22214 -581
rect -22776 -984 -22764 -587
rect -22226 -984 -22214 -587
rect -22776 -990 -22214 -984
rect -21958 -587 -21396 -581
rect -21958 -984 -21946 -587
rect -21408 -984 -21396 -587
rect -21958 -990 -21396 -984
rect -21140 -587 -20578 -581
rect -21140 -984 -21128 -587
rect -20590 -984 -20578 -587
rect -21140 -990 -20578 -984
rect -20322 -587 -19760 -581
rect -20322 -984 -20310 -587
rect -19772 -984 -19760 -587
rect -20322 -990 -19760 -984
rect -19504 -587 -18942 -581
rect -19504 -984 -19492 -587
rect -18954 -984 -18942 -587
rect -19504 -990 -18942 -984
rect -18686 -587 -18124 -581
rect -18686 -984 -18674 -587
rect -18136 -984 -18124 -587
rect -18686 -990 -18124 -984
rect -17868 -587 -17306 -581
rect -17868 -984 -17856 -587
rect -17318 -984 -17306 -587
rect -17868 -990 -17306 -984
rect -17050 -587 -16488 -581
rect -17050 -984 -17038 -587
rect -16500 -984 -16488 -587
rect -17050 -990 -16488 -984
rect -16232 -587 -15670 -581
rect -16232 -984 -16220 -587
rect -15682 -984 -15670 -587
rect -16232 -990 -15670 -984
rect -15414 -587 -14852 -581
rect -15414 -984 -15402 -587
rect -14864 -984 -14852 -587
rect -15414 -990 -14852 -984
rect -14596 -587 -14034 -581
rect -14596 -984 -14584 -587
rect -14046 -984 -14034 -587
rect -14596 -990 -14034 -984
rect -13778 -587 -13216 -581
rect -13778 -984 -13766 -587
rect -13228 -984 -13216 -587
rect -13778 -990 -13216 -984
rect -12960 -587 -12398 -581
rect -12960 -984 -12948 -587
rect -12410 -984 -12398 -587
rect -12960 -990 -12398 -984
rect -12142 -587 -11580 -581
rect -12142 -984 -12130 -587
rect -11592 -984 -11580 -587
rect -12142 -990 -11580 -984
rect -11324 -587 -10762 -581
rect -11324 -984 -11312 -587
rect -10774 -984 -10762 -587
rect -11324 -990 -10762 -984
rect -10506 -587 -9944 -581
rect -10506 -984 -10494 -587
rect -9956 -984 -9944 -587
rect -10506 -990 -9944 -984
rect -9688 -587 -9126 -581
rect -9688 -984 -9676 -587
rect -9138 -984 -9126 -587
rect -9688 -990 -9126 -984
rect -8870 -587 -8308 -581
rect -8870 -984 -8858 -587
rect -8320 -984 -8308 -587
rect -8870 -990 -8308 -984
rect -8052 -587 -7490 -581
rect -8052 -984 -8040 -587
rect -7502 -984 -7490 -587
rect -8052 -990 -7490 -984
rect -7234 -587 -6672 -581
rect -7234 -984 -7222 -587
rect -6684 -984 -6672 -587
rect -7234 -990 -6672 -984
rect -6416 -587 -5854 -581
rect -6416 -984 -6404 -587
rect -5866 -984 -5854 -587
rect -6416 -990 -5854 -984
rect -5598 -587 -5036 -581
rect -5598 -984 -5586 -587
rect -5048 -984 -5036 -587
rect -5598 -990 -5036 -984
rect -4780 -587 -4218 -581
rect -4780 -984 -4768 -587
rect -4230 -984 -4218 -587
rect -4780 -990 -4218 -984
rect -3962 -587 -3400 -581
rect -3962 -984 -3950 -587
rect -3412 -984 -3400 -587
rect -3962 -990 -3400 -984
rect -3144 -587 -2582 -581
rect -3144 -984 -3132 -587
rect -2594 -984 -2582 -587
rect -3144 -990 -2582 -984
rect -2326 -587 -1764 -581
rect -2326 -984 -2314 -587
rect -1776 -984 -1764 -587
rect -2326 -990 -1764 -984
rect -1508 -587 -946 -581
rect -1508 -984 -1496 -587
rect -958 -984 -946 -587
rect -1508 -990 -946 -984
rect -690 -587 -128 -581
rect -690 -984 -678 -587
rect -140 -984 -128 -587
rect -690 -990 -128 -984
rect 128 -587 690 -581
rect 128 -984 140 -587
rect 678 -984 690 -587
rect 128 -990 690 -984
rect 946 -587 1508 -581
rect 946 -984 958 -587
rect 1496 -984 1508 -587
rect 946 -990 1508 -984
rect 1764 -587 2326 -581
rect 1764 -984 1776 -587
rect 2314 -984 2326 -587
rect 1764 -990 2326 -984
rect 2582 -587 3144 -581
rect 2582 -984 2594 -587
rect 3132 -984 3144 -587
rect 2582 -990 3144 -984
rect 3400 -587 3962 -581
rect 3400 -984 3412 -587
rect 3950 -984 3962 -587
rect 3400 -990 3962 -984
rect 4218 -587 4780 -581
rect 4218 -984 4230 -587
rect 4768 -984 4780 -587
rect 4218 -990 4780 -984
rect 5036 -587 5598 -581
rect 5036 -984 5048 -587
rect 5586 -984 5598 -587
rect 5036 -990 5598 -984
rect 5854 -587 6416 -581
rect 5854 -984 5866 -587
rect 6404 -984 6416 -587
rect 5854 -990 6416 -984
rect 6672 -587 7234 -581
rect 6672 -984 6684 -587
rect 7222 -984 7234 -587
rect 6672 -990 7234 -984
rect 7490 -587 8052 -581
rect 7490 -984 7502 -587
rect 8040 -984 8052 -587
rect 7490 -990 8052 -984
rect 8308 -587 8870 -581
rect 8308 -984 8320 -587
rect 8858 -984 8870 -587
rect 8308 -990 8870 -984
rect 9126 -587 9688 -581
rect 9126 -984 9138 -587
rect 9676 -984 9688 -587
rect 9126 -990 9688 -984
rect 9944 -587 10506 -581
rect 9944 -984 9956 -587
rect 10494 -984 10506 -587
rect 9944 -990 10506 -984
rect 10762 -587 11324 -581
rect 10762 -984 10774 -587
rect 11312 -984 11324 -587
rect 10762 -990 11324 -984
rect 11580 -587 12142 -581
rect 11580 -984 11592 -587
rect 12130 -984 12142 -587
rect 11580 -990 12142 -984
rect 12398 -587 12960 -581
rect 12398 -984 12410 -587
rect 12948 -984 12960 -587
rect 12398 -990 12960 -984
rect 13216 -587 13778 -581
rect 13216 -984 13228 -587
rect 13766 -984 13778 -587
rect 13216 -990 13778 -984
rect 14034 -587 14596 -581
rect 14034 -984 14046 -587
rect 14584 -984 14596 -587
rect 14034 -990 14596 -984
rect 14852 -587 15414 -581
rect 14852 -984 14864 -587
rect 15402 -984 15414 -587
rect 14852 -990 15414 -984
rect 15670 -587 16232 -581
rect 15670 -984 15682 -587
rect 16220 -984 16232 -587
rect 15670 -990 16232 -984
rect 16488 -587 17050 -581
rect 16488 -984 16500 -587
rect 17038 -984 17050 -587
rect 16488 -990 17050 -984
rect 17306 -587 17868 -581
rect 17306 -984 17318 -587
rect 17856 -984 17868 -587
rect 17306 -990 17868 -984
rect 18124 -587 18686 -581
rect 18124 -984 18136 -587
rect 18674 -984 18686 -587
rect 18124 -990 18686 -984
rect 18942 -587 19504 -581
rect 18942 -984 18954 -587
rect 19492 -984 19504 -587
rect 18942 -990 19504 -984
rect 19760 -587 20322 -581
rect 19760 -984 19772 -587
rect 20310 -984 20322 -587
rect 19760 -990 20322 -984
rect 20578 -587 21140 -581
rect 20578 -984 20590 -587
rect 21128 -984 21140 -587
rect 20578 -990 21140 -984
rect 21396 -587 21958 -581
rect 21396 -984 21408 -587
rect 21946 -984 21958 -587
rect 21396 -990 21958 -984
rect 22214 -587 22776 -581
rect 22214 -984 22226 -587
rect 22764 -984 22776 -587
rect 22214 -990 22776 -984
rect 23032 -587 23594 -581
rect 23032 -984 23044 -587
rect 23582 -984 23594 -587
rect 23032 -990 23594 -984
rect 23850 -587 24412 -581
rect 23850 -984 23862 -587
rect 24400 -984 24412 -587
rect 23850 -990 24412 -984
rect 24668 -587 25230 -581
rect 24668 -984 24680 -587
rect 25218 -984 25230 -587
rect 24668 -990 25230 -984
rect 25486 -587 26048 -581
rect 25486 -984 25498 -587
rect 26036 -984 26048 -587
rect 25486 -990 26048 -984
rect 26304 -587 26866 -581
rect 26304 -984 26316 -587
rect 26854 -984 26866 -587
rect 26304 -990 26866 -984
rect 27122 -587 27684 -581
rect 27122 -984 27134 -587
rect 27672 -984 27684 -587
rect 27122 -990 27684 -984
rect 27940 -587 28502 -581
rect 27940 -984 27952 -587
rect 28490 -984 28502 -587
rect 27940 -990 28502 -984
rect 28758 -587 29320 -581
rect 28758 -984 28770 -587
rect 29308 -984 29320 -587
rect 28758 -990 29320 -984
rect 29576 -587 30138 -581
rect 29576 -984 29588 -587
rect 30126 -984 30138 -587
rect 29576 -990 30138 -984
rect 30394 -587 30956 -581
rect 30394 -984 30406 -587
rect 30944 -984 30956 -587
rect 30394 -990 30956 -984
rect 31212 -587 31774 -581
rect 31212 -984 31224 -587
rect 31762 -984 31774 -587
rect 31212 -990 31774 -984
rect 32030 -587 32592 -581
rect 32030 -984 32042 -587
rect 32580 -984 32592 -587
rect 32030 -990 32592 -984
rect 32848 -587 33410 -581
rect 32848 -984 32860 -587
rect 33398 -984 33410 -587
rect 32848 -990 33410 -984
rect 33666 -587 34228 -581
rect 33666 -984 33678 -587
rect 34216 -984 34228 -587
rect 33666 -990 34228 -984
rect 34484 -587 35046 -581
rect 34484 -984 34496 -587
rect 35034 -984 35046 -587
rect 34484 -990 35046 -984
rect 35302 -587 35864 -581
rect 35302 -984 35314 -587
rect 35852 -984 35864 -587
rect 35302 -990 35864 -984
rect 36120 -587 36682 -581
rect 36120 -984 36132 -587
rect 36670 -984 36682 -587
rect 36120 -990 36682 -984
rect 36938 -587 37500 -581
rect 36938 -984 36950 -587
rect 37488 -984 37500 -587
rect 36938 -990 37500 -984
rect 37756 -587 38318 -581
rect 37756 -984 37768 -587
rect 38306 -984 38318 -587
rect 37756 -990 38318 -984
rect 38574 -587 39136 -581
rect 38574 -984 38586 -587
rect 39124 -984 39136 -587
rect 38574 -990 39136 -984
rect 39392 -587 39954 -581
rect 39392 -984 39404 -587
rect 39942 -984 39954 -587
rect 39392 -990 39954 -984
rect 40210 -587 40772 -581
rect 40210 -984 40222 -587
rect 40760 -984 40772 -587
rect 40210 -990 40772 -984
rect 41028 -587 41590 -581
rect 41028 -984 41040 -587
rect 41578 -984 41590 -587
rect 41028 -990 41590 -984
rect 41846 -587 42408 -581
rect 41846 -984 41858 -587
rect 42396 -984 42408 -587
rect 41846 -990 42408 -984
rect 42664 -587 43226 -581
rect 42664 -984 42676 -587
rect 43214 -984 43226 -587
rect 42664 -990 43226 -984
rect 43482 -587 44044 -581
rect 43482 -984 43494 -587
rect 44032 -984 44044 -587
rect 43482 -990 44044 -984
rect 44300 -587 44862 -581
rect 44300 -984 44312 -587
rect 44850 -984 44862 -587
rect 44300 -990 44862 -984
rect 45118 -587 45680 -581
rect 45118 -984 45130 -587
rect 45668 -984 45680 -587
rect 45118 -990 45680 -984
rect 45936 -587 46498 -581
rect 45936 -984 45948 -587
rect 46486 -984 46498 -587
rect 45936 -990 46498 -984
rect 46754 -587 47316 -581
rect 46754 -984 46766 -587
rect 47304 -984 47316 -587
rect 46754 -990 47316 -984
rect 47572 -587 48134 -581
rect 47572 -984 47584 -587
rect 48122 -984 48134 -587
rect 47572 -990 48134 -984
rect 48390 -587 48952 -581
rect 48390 -984 48402 -587
rect 48940 -984 48952 -587
rect 48390 -990 48952 -984
rect 49208 -587 49770 -581
rect 49208 -984 49220 -587
rect 49758 -984 49770 -587
rect 49208 -990 49770 -984
rect 50026 -587 50588 -581
rect 50026 -984 50038 -587
rect 50576 -984 50588 -587
rect 50026 -990 50588 -984
rect 50844 -587 51406 -581
rect 50844 -984 50856 -587
rect 51394 -984 51406 -587
rect 50844 -990 51406 -984
rect 51662 -587 52224 -581
rect 51662 -984 51674 -587
rect 52212 -984 52224 -587
rect 51662 -990 52224 -984
rect 52480 -587 53042 -581
rect 52480 -984 52492 -587
rect 53030 -984 53042 -587
rect 52480 -990 53042 -984
rect 53298 -587 53860 -581
rect 53298 -984 53310 -587
rect 53848 -984 53860 -587
rect 53298 -990 53860 -984
rect 54116 -587 54678 -581
rect 54116 -984 54128 -587
rect 54666 -984 54678 -587
rect 54116 -990 54678 -984
rect 54934 -587 55496 -581
rect 54934 -984 54946 -587
rect 55484 -984 55496 -587
rect 54934 -990 55496 -984
rect 55752 -587 56314 -581
rect 55752 -984 55764 -587
rect 56302 -984 56314 -587
rect 55752 -990 56314 -984
rect 56570 -587 57132 -581
rect 56570 -984 56582 -587
rect 57120 -984 57132 -587
rect 56570 -990 57132 -984
rect 57388 -587 57950 -581
rect 57388 -984 57400 -587
rect 57938 -984 57950 -587
rect 57388 -990 57950 -984
rect 58206 -587 58768 -581
rect 58206 -984 58218 -587
rect 58756 -984 58768 -587
rect 58206 -990 58768 -984
rect 59024 -587 59586 -581
rect 59024 -984 59036 -587
rect 59574 -984 59586 -587
rect 59024 -990 59586 -984
rect 59842 -587 60404 -581
rect 59842 -984 59854 -587
rect 60392 -984 60404 -587
rect 59842 -990 60404 -984
rect 60660 -587 61222 -581
rect 60660 -984 60672 -587
rect 61210 -984 61222 -587
rect 60660 -990 61222 -984
rect 61478 -587 62040 -581
rect 61478 -984 61490 -587
rect 62028 -984 62040 -587
rect 61478 -990 62040 -984
rect 62296 -587 62858 -581
rect 62296 -984 62308 -587
rect 62846 -984 62858 -587
rect 62296 -990 62858 -984
rect 63114 -587 63676 -581
rect 63114 -984 63126 -587
rect 63664 -984 63676 -587
rect 63114 -990 63676 -984
rect 63932 -587 64494 -581
rect 63932 -984 63944 -587
rect 64482 -984 64494 -587
rect 63932 -990 64494 -984
rect 64750 -587 65312 -581
rect 64750 -984 64762 -587
rect 65300 -984 65312 -587
rect 64750 -990 65312 -984
<< res2p85 >>
rect -65318 -572 -64744 572
rect -64500 -572 -63926 572
rect -63682 -572 -63108 572
rect -62864 -572 -62290 572
rect -62046 -572 -61472 572
rect -61228 -572 -60654 572
rect -60410 -572 -59836 572
rect -59592 -572 -59018 572
rect -58774 -572 -58200 572
rect -57956 -572 -57382 572
rect -57138 -572 -56564 572
rect -56320 -572 -55746 572
rect -55502 -572 -54928 572
rect -54684 -572 -54110 572
rect -53866 -572 -53292 572
rect -53048 -572 -52474 572
rect -52230 -572 -51656 572
rect -51412 -572 -50838 572
rect -50594 -572 -50020 572
rect -49776 -572 -49202 572
rect -48958 -572 -48384 572
rect -48140 -572 -47566 572
rect -47322 -572 -46748 572
rect -46504 -572 -45930 572
rect -45686 -572 -45112 572
rect -44868 -572 -44294 572
rect -44050 -572 -43476 572
rect -43232 -572 -42658 572
rect -42414 -572 -41840 572
rect -41596 -572 -41022 572
rect -40778 -572 -40204 572
rect -39960 -572 -39386 572
rect -39142 -572 -38568 572
rect -38324 -572 -37750 572
rect -37506 -572 -36932 572
rect -36688 -572 -36114 572
rect -35870 -572 -35296 572
rect -35052 -572 -34478 572
rect -34234 -572 -33660 572
rect -33416 -572 -32842 572
rect -32598 -572 -32024 572
rect -31780 -572 -31206 572
rect -30962 -572 -30388 572
rect -30144 -572 -29570 572
rect -29326 -572 -28752 572
rect -28508 -572 -27934 572
rect -27690 -572 -27116 572
rect -26872 -572 -26298 572
rect -26054 -572 -25480 572
rect -25236 -572 -24662 572
rect -24418 -572 -23844 572
rect -23600 -572 -23026 572
rect -22782 -572 -22208 572
rect -21964 -572 -21390 572
rect -21146 -572 -20572 572
rect -20328 -572 -19754 572
rect -19510 -572 -18936 572
rect -18692 -572 -18118 572
rect -17874 -572 -17300 572
rect -17056 -572 -16482 572
rect -16238 -572 -15664 572
rect -15420 -572 -14846 572
rect -14602 -572 -14028 572
rect -13784 -572 -13210 572
rect -12966 -572 -12392 572
rect -12148 -572 -11574 572
rect -11330 -572 -10756 572
rect -10512 -572 -9938 572
rect -9694 -572 -9120 572
rect -8876 -572 -8302 572
rect -8058 -572 -7484 572
rect -7240 -572 -6666 572
rect -6422 -572 -5848 572
rect -5604 -572 -5030 572
rect -4786 -572 -4212 572
rect -3968 -572 -3394 572
rect -3150 -572 -2576 572
rect -2332 -572 -1758 572
rect -1514 -572 -940 572
rect -696 -572 -122 572
rect 122 -572 696 572
rect 940 -572 1514 572
rect 1758 -572 2332 572
rect 2576 -572 3150 572
rect 3394 -572 3968 572
rect 4212 -572 4786 572
rect 5030 -572 5604 572
rect 5848 -572 6422 572
rect 6666 -572 7240 572
rect 7484 -572 8058 572
rect 8302 -572 8876 572
rect 9120 -572 9694 572
rect 9938 -572 10512 572
rect 10756 -572 11330 572
rect 11574 -572 12148 572
rect 12392 -572 12966 572
rect 13210 -572 13784 572
rect 14028 -572 14602 572
rect 14846 -572 15420 572
rect 15664 -572 16238 572
rect 16482 -572 17056 572
rect 17300 -572 17874 572
rect 18118 -572 18692 572
rect 18936 -572 19510 572
rect 19754 -572 20328 572
rect 20572 -572 21146 572
rect 21390 -572 21964 572
rect 22208 -572 22782 572
rect 23026 -572 23600 572
rect 23844 -572 24418 572
rect 24662 -572 25236 572
rect 25480 -572 26054 572
rect 26298 -572 26872 572
rect 27116 -572 27690 572
rect 27934 -572 28508 572
rect 28752 -572 29326 572
rect 29570 -572 30144 572
rect 30388 -572 30962 572
rect 31206 -572 31780 572
rect 32024 -572 32598 572
rect 32842 -572 33416 572
rect 33660 -572 34234 572
rect 34478 -572 35052 572
rect 35296 -572 35870 572
rect 36114 -572 36688 572
rect 36932 -572 37506 572
rect 37750 -572 38324 572
rect 38568 -572 39142 572
rect 39386 -572 39960 572
rect 40204 -572 40778 572
rect 41022 -572 41596 572
rect 41840 -572 42414 572
rect 42658 -572 43232 572
rect 43476 -572 44050 572
rect 44294 -572 44868 572
rect 45112 -572 45686 572
rect 45930 -572 46504 572
rect 46748 -572 47322 572
rect 47566 -572 48140 572
rect 48384 -572 48958 572
rect 49202 -572 49776 572
rect 50020 -572 50594 572
rect 50838 -572 51412 572
rect 51656 -572 52230 572
rect 52474 -572 53048 572
rect 53292 -572 53866 572
rect 54110 -572 54684 572
rect 54928 -572 55502 572
rect 55746 -572 56320 572
rect 56564 -572 57138 572
rect 57382 -572 57956 572
rect 58200 -572 58774 572
rect 59018 -572 59592 572
rect 59836 -572 60410 572
rect 60654 -572 61228 572
rect 61472 -572 62046 572
rect 62290 -572 62864 572
rect 63108 -572 63682 572
rect 63926 -572 64500 572
rect 64744 -572 65318 572
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_2p85
string parameters w 2.850 l 5.7 m 1 nx 160 wmin 2.850 lmin 0.50 rho 2000 val 4.013k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 2.850 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
