magic
tech sky130A
magscale 1 2
timestamp 1620853902
<< nwell >>
rect -3440 -1354 3440 1388
<< pmoslvt >>
rect -3346 -1254 -2946 1326
rect -2774 -1254 -2374 1326
rect -2202 -1254 -1802 1326
rect -1630 -1254 -1230 1326
rect -1058 -1254 -658 1326
rect -486 -1254 -86 1326
rect 86 -1254 486 1326
rect 658 -1254 1058 1326
rect 1230 -1254 1630 1326
rect 1802 -1254 2202 1326
rect 2374 -1254 2774 1326
rect 2946 -1254 3346 1326
<< pdiff >>
rect -3404 1314 -3346 1326
rect -3404 -1242 -3392 1314
rect -3358 -1242 -3346 1314
rect -3404 -1254 -3346 -1242
rect -2946 1314 -2888 1326
rect -2946 -1242 -2934 1314
rect -2900 -1242 -2888 1314
rect -2946 -1254 -2888 -1242
rect -2832 1314 -2774 1326
rect -2832 -1242 -2820 1314
rect -2786 -1242 -2774 1314
rect -2832 -1254 -2774 -1242
rect -2374 1314 -2316 1326
rect -2374 -1242 -2362 1314
rect -2328 -1242 -2316 1314
rect -2374 -1254 -2316 -1242
rect -2260 1314 -2202 1326
rect -2260 -1242 -2248 1314
rect -2214 -1242 -2202 1314
rect -2260 -1254 -2202 -1242
rect -1802 1314 -1744 1326
rect -1802 -1242 -1790 1314
rect -1756 -1242 -1744 1314
rect -1802 -1254 -1744 -1242
rect -1688 1314 -1630 1326
rect -1688 -1242 -1676 1314
rect -1642 -1242 -1630 1314
rect -1688 -1254 -1630 -1242
rect -1230 1314 -1172 1326
rect -1230 -1242 -1218 1314
rect -1184 -1242 -1172 1314
rect -1230 -1254 -1172 -1242
rect -1116 1314 -1058 1326
rect -1116 -1242 -1104 1314
rect -1070 -1242 -1058 1314
rect -1116 -1254 -1058 -1242
rect -658 1314 -600 1326
rect -658 -1242 -646 1314
rect -612 -1242 -600 1314
rect -658 -1254 -600 -1242
rect -544 1314 -486 1326
rect -544 -1242 -532 1314
rect -498 -1242 -486 1314
rect -544 -1254 -486 -1242
rect -86 1314 -28 1326
rect -86 -1242 -74 1314
rect -40 -1242 -28 1314
rect -86 -1254 -28 -1242
rect 28 1314 86 1326
rect 28 -1242 40 1314
rect 74 -1242 86 1314
rect 28 -1254 86 -1242
rect 486 1314 544 1326
rect 486 -1242 498 1314
rect 532 -1242 544 1314
rect 486 -1254 544 -1242
rect 600 1314 658 1326
rect 600 -1242 612 1314
rect 646 -1242 658 1314
rect 600 -1254 658 -1242
rect 1058 1314 1116 1326
rect 1058 -1242 1070 1314
rect 1104 -1242 1116 1314
rect 1058 -1254 1116 -1242
rect 1172 1314 1230 1326
rect 1172 -1242 1184 1314
rect 1218 -1242 1230 1314
rect 1172 -1254 1230 -1242
rect 1630 1314 1688 1326
rect 1630 -1242 1642 1314
rect 1676 -1242 1688 1314
rect 1630 -1254 1688 -1242
rect 1744 1314 1802 1326
rect 1744 -1242 1756 1314
rect 1790 -1242 1802 1314
rect 1744 -1254 1802 -1242
rect 2202 1314 2260 1326
rect 2202 -1242 2214 1314
rect 2248 -1242 2260 1314
rect 2202 -1254 2260 -1242
rect 2316 1314 2374 1326
rect 2316 -1242 2328 1314
rect 2362 -1242 2374 1314
rect 2316 -1254 2374 -1242
rect 2774 1314 2832 1326
rect 2774 -1242 2786 1314
rect 2820 -1242 2832 1314
rect 2774 -1254 2832 -1242
rect 2888 1314 2946 1326
rect 2888 -1242 2900 1314
rect 2934 -1242 2946 1314
rect 2888 -1254 2946 -1242
rect 3346 1314 3404 1326
rect 3346 -1242 3358 1314
rect 3392 -1242 3404 1314
rect 3346 -1254 3404 -1242
<< pdiffc >>
rect -3392 -1242 -3358 1314
rect -2934 -1242 -2900 1314
rect -2820 -1242 -2786 1314
rect -2362 -1242 -2328 1314
rect -2248 -1242 -2214 1314
rect -1790 -1242 -1756 1314
rect -1676 -1242 -1642 1314
rect -1218 -1242 -1184 1314
rect -1104 -1242 -1070 1314
rect -646 -1242 -612 1314
rect -532 -1242 -498 1314
rect -74 -1242 -40 1314
rect 40 -1242 74 1314
rect 498 -1242 532 1314
rect 612 -1242 646 1314
rect 1070 -1242 1104 1314
rect 1184 -1242 1218 1314
rect 1642 -1242 1676 1314
rect 1756 -1242 1790 1314
rect 2214 -1242 2248 1314
rect 2328 -1242 2362 1314
rect 2786 -1242 2820 1314
rect 2900 -1242 2934 1314
rect 3358 -1242 3392 1314
<< poly >>
rect -3346 1326 -2946 1352
rect -2774 1326 -2374 1352
rect -2202 1326 -1802 1352
rect -1630 1326 -1230 1352
rect -1058 1326 -658 1352
rect -486 1326 -86 1352
rect 86 1326 486 1352
rect 658 1326 1058 1352
rect 1230 1326 1630 1352
rect 1802 1326 2202 1352
rect 2374 1326 2774 1352
rect 2946 1326 3346 1352
rect -3346 -1301 -2946 -1254
rect -3346 -1335 -3330 -1301
rect -2962 -1335 -2946 -1301
rect -3346 -1351 -2946 -1335
rect -2774 -1301 -2374 -1254
rect -2774 -1335 -2758 -1301
rect -2390 -1335 -2374 -1301
rect -2774 -1351 -2374 -1335
rect -2202 -1301 -1802 -1254
rect -2202 -1335 -2186 -1301
rect -1818 -1335 -1802 -1301
rect -2202 -1351 -1802 -1335
rect -1630 -1301 -1230 -1254
rect -1630 -1335 -1614 -1301
rect -1246 -1335 -1230 -1301
rect -1630 -1351 -1230 -1335
rect -1058 -1301 -658 -1254
rect -1058 -1335 -1042 -1301
rect -674 -1335 -658 -1301
rect -1058 -1351 -658 -1335
rect -486 -1301 -86 -1254
rect -486 -1335 -470 -1301
rect -102 -1335 -86 -1301
rect -486 -1351 -86 -1335
rect 86 -1301 486 -1254
rect 86 -1335 102 -1301
rect 470 -1335 486 -1301
rect 86 -1351 486 -1335
rect 658 -1301 1058 -1254
rect 658 -1335 674 -1301
rect 1042 -1335 1058 -1301
rect 658 -1351 1058 -1335
rect 1230 -1301 1630 -1254
rect 1230 -1335 1246 -1301
rect 1614 -1335 1630 -1301
rect 1230 -1351 1630 -1335
rect 1802 -1301 2202 -1254
rect 1802 -1335 1818 -1301
rect 2186 -1335 2202 -1301
rect 1802 -1351 2202 -1335
rect 2374 -1301 2774 -1254
rect 2374 -1335 2390 -1301
rect 2758 -1335 2774 -1301
rect 2374 -1351 2774 -1335
rect 2946 -1301 3346 -1254
rect 2946 -1335 2962 -1301
rect 3330 -1335 3346 -1301
rect 2946 -1351 3346 -1335
<< polycont >>
rect -3330 -1335 -2962 -1301
rect -2758 -1335 -2390 -1301
rect -2186 -1335 -1818 -1301
rect -1614 -1335 -1246 -1301
rect -1042 -1335 -674 -1301
rect -470 -1335 -102 -1301
rect 102 -1335 470 -1301
rect 674 -1335 1042 -1301
rect 1246 -1335 1614 -1301
rect 1818 -1335 2186 -1301
rect 2390 -1335 2758 -1301
rect 2962 -1335 3330 -1301
<< locali >>
rect -3392 1314 -3358 1330
rect -3392 -1258 -3358 -1242
rect -2934 1314 -2900 1330
rect -2934 -1258 -2900 -1242
rect -2820 1314 -2786 1330
rect -2820 -1258 -2786 -1242
rect -2362 1314 -2328 1330
rect -2362 -1258 -2328 -1242
rect -2248 1314 -2214 1330
rect -2248 -1258 -2214 -1242
rect -1790 1314 -1756 1330
rect -1790 -1258 -1756 -1242
rect -1676 1314 -1642 1330
rect -1676 -1258 -1642 -1242
rect -1218 1314 -1184 1330
rect -1218 -1258 -1184 -1242
rect -1104 1314 -1070 1330
rect -1104 -1258 -1070 -1242
rect -646 1314 -612 1330
rect -646 -1258 -612 -1242
rect -532 1314 -498 1330
rect -532 -1258 -498 -1242
rect -74 1314 -40 1330
rect -74 -1258 -40 -1242
rect 40 1314 74 1330
rect 40 -1258 74 -1242
rect 498 1314 532 1330
rect 498 -1258 532 -1242
rect 612 1314 646 1330
rect 612 -1258 646 -1242
rect 1070 1314 1104 1330
rect 1070 -1258 1104 -1242
rect 1184 1314 1218 1330
rect 1184 -1258 1218 -1242
rect 1642 1314 1676 1330
rect 1642 -1258 1676 -1242
rect 1756 1314 1790 1330
rect 1756 -1258 1790 -1242
rect 2214 1314 2248 1330
rect 2214 -1258 2248 -1242
rect 2328 1314 2362 1330
rect 2328 -1258 2362 -1242
rect 2786 1314 2820 1330
rect 2786 -1258 2820 -1242
rect 2900 1314 2934 1330
rect 2900 -1258 2934 -1242
rect 3358 1314 3392 1330
rect 3358 -1258 3392 -1242
rect -3346 -1335 -3330 -1301
rect -2962 -1335 -2946 -1301
rect -2774 -1335 -2758 -1301
rect -2390 -1335 -2374 -1301
rect -2202 -1335 -2186 -1301
rect -1818 -1335 -1802 -1301
rect -1630 -1335 -1614 -1301
rect -1246 -1335 -1230 -1301
rect -1058 -1335 -1042 -1301
rect -674 -1335 -658 -1301
rect -486 -1335 -470 -1301
rect -102 -1335 -86 -1301
rect 86 -1335 102 -1301
rect 470 -1335 486 -1301
rect 658 -1335 674 -1301
rect 1042 -1335 1058 -1301
rect 1230 -1335 1246 -1301
rect 1614 -1335 1630 -1301
rect 1802 -1335 1818 -1301
rect 2186 -1335 2202 -1301
rect 2374 -1335 2390 -1301
rect 2758 -1335 2774 -1301
rect 2946 -1335 2962 -1301
rect 3330 -1335 3346 -1301
<< viali >>
rect -3392 -1242 -3358 1314
rect -2934 -1242 -2900 1314
rect -2820 -1242 -2786 1314
rect -2362 -1242 -2328 1314
rect -2248 -1242 -2214 1314
rect -1790 -1242 -1756 1314
rect -1676 -1242 -1642 1314
rect -1218 -1242 -1184 1314
rect -1104 -1242 -1070 1314
rect -646 -1242 -612 1314
rect -532 -1242 -498 1314
rect -74 -1242 -40 1314
rect 40 -1242 74 1314
rect 498 -1242 532 1314
rect 612 -1242 646 1314
rect 1070 -1242 1104 1314
rect 1184 -1242 1218 1314
rect 1642 -1242 1676 1314
rect 1756 -1242 1790 1314
rect 2214 -1242 2248 1314
rect 2328 -1242 2362 1314
rect 2786 -1242 2820 1314
rect 2900 -1242 2934 1314
rect 3358 -1242 3392 1314
rect -3238 -1335 -3054 -1301
rect -2666 -1335 -2482 -1301
rect -2094 -1335 -1910 -1301
rect -1522 -1335 -1338 -1301
rect -950 -1335 -766 -1301
rect -378 -1335 -194 -1301
rect 194 -1335 378 -1301
rect 766 -1335 950 -1301
rect 1338 -1335 1522 -1301
rect 1910 -1335 2094 -1301
rect 2482 -1335 2666 -1301
rect 3054 -1335 3238 -1301
<< metal1 >>
rect -3398 1314 -3352 1326
rect -3398 -1242 -3392 1314
rect -3358 -1242 -3352 1314
rect -3398 -1254 -3352 -1242
rect -2940 1314 -2894 1326
rect -2940 -1242 -2934 1314
rect -2900 -1242 -2894 1314
rect -2940 -1254 -2894 -1242
rect -2826 1314 -2780 1326
rect -2826 -1242 -2820 1314
rect -2786 -1242 -2780 1314
rect -2826 -1254 -2780 -1242
rect -2368 1314 -2322 1326
rect -2368 -1242 -2362 1314
rect -2328 -1242 -2322 1314
rect -2368 -1254 -2322 -1242
rect -2254 1314 -2208 1326
rect -2254 -1242 -2248 1314
rect -2214 -1242 -2208 1314
rect -2254 -1254 -2208 -1242
rect -1796 1314 -1750 1326
rect -1796 -1242 -1790 1314
rect -1756 -1242 -1750 1314
rect -1796 -1254 -1750 -1242
rect -1682 1314 -1636 1326
rect -1682 -1242 -1676 1314
rect -1642 -1242 -1636 1314
rect -1682 -1254 -1636 -1242
rect -1224 1314 -1178 1326
rect -1224 -1242 -1218 1314
rect -1184 -1242 -1178 1314
rect -1224 -1254 -1178 -1242
rect -1110 1314 -1064 1326
rect -1110 -1242 -1104 1314
rect -1070 -1242 -1064 1314
rect -1110 -1254 -1064 -1242
rect -652 1314 -606 1326
rect -652 -1242 -646 1314
rect -612 -1242 -606 1314
rect -652 -1254 -606 -1242
rect -538 1314 -492 1326
rect -538 -1242 -532 1314
rect -498 -1242 -492 1314
rect -538 -1254 -492 -1242
rect -80 1314 -34 1326
rect -80 -1242 -74 1314
rect -40 -1242 -34 1314
rect -80 -1254 -34 -1242
rect 34 1314 80 1326
rect 34 -1242 40 1314
rect 74 -1242 80 1314
rect 34 -1254 80 -1242
rect 492 1314 538 1326
rect 492 -1242 498 1314
rect 532 -1242 538 1314
rect 492 -1254 538 -1242
rect 606 1314 652 1326
rect 606 -1242 612 1314
rect 646 -1242 652 1314
rect 606 -1254 652 -1242
rect 1064 1314 1110 1326
rect 1064 -1242 1070 1314
rect 1104 -1242 1110 1314
rect 1064 -1254 1110 -1242
rect 1178 1314 1224 1326
rect 1178 -1242 1184 1314
rect 1218 -1242 1224 1314
rect 1178 -1254 1224 -1242
rect 1636 1314 1682 1326
rect 1636 -1242 1642 1314
rect 1676 -1242 1682 1314
rect 1636 -1254 1682 -1242
rect 1750 1314 1796 1326
rect 1750 -1242 1756 1314
rect 1790 -1242 1796 1314
rect 1750 -1254 1796 -1242
rect 2208 1314 2254 1326
rect 2208 -1242 2214 1314
rect 2248 -1242 2254 1314
rect 2208 -1254 2254 -1242
rect 2322 1314 2368 1326
rect 2322 -1242 2328 1314
rect 2362 -1242 2368 1314
rect 2322 -1254 2368 -1242
rect 2780 1314 2826 1326
rect 2780 -1242 2786 1314
rect 2820 -1242 2826 1314
rect 2780 -1254 2826 -1242
rect 2894 1314 2940 1326
rect 2894 -1242 2900 1314
rect 2934 -1242 2940 1314
rect 2894 -1254 2940 -1242
rect 3352 1314 3398 1326
rect 3352 -1242 3358 1314
rect 3392 -1242 3398 1314
rect 3352 -1254 3398 -1242
rect -3250 -1301 -3042 -1295
rect -3250 -1335 -3238 -1301
rect -3054 -1335 -3042 -1301
rect -3250 -1341 -3042 -1335
rect -2678 -1301 -2470 -1295
rect -2678 -1335 -2666 -1301
rect -2482 -1335 -2470 -1301
rect -2678 -1341 -2470 -1335
rect -2106 -1301 -1898 -1295
rect -2106 -1335 -2094 -1301
rect -1910 -1335 -1898 -1301
rect -2106 -1341 -1898 -1335
rect -1534 -1301 -1326 -1295
rect -1534 -1335 -1522 -1301
rect -1338 -1335 -1326 -1301
rect -1534 -1341 -1326 -1335
rect -962 -1301 -754 -1295
rect -962 -1335 -950 -1301
rect -766 -1335 -754 -1301
rect -962 -1341 -754 -1335
rect -390 -1301 -182 -1295
rect -390 -1335 -378 -1301
rect -194 -1335 -182 -1301
rect -390 -1341 -182 -1335
rect 182 -1301 390 -1295
rect 182 -1335 194 -1301
rect 378 -1335 390 -1301
rect 182 -1341 390 -1335
rect 754 -1301 962 -1295
rect 754 -1335 766 -1301
rect 950 -1335 962 -1301
rect 754 -1341 962 -1335
rect 1326 -1301 1534 -1295
rect 1326 -1335 1338 -1301
rect 1522 -1335 1534 -1301
rect 1326 -1341 1534 -1335
rect 1898 -1301 2106 -1295
rect 1898 -1335 1910 -1301
rect 2094 -1335 2106 -1301
rect 1898 -1341 2106 -1335
rect 2470 -1301 2678 -1295
rect 2470 -1335 2482 -1301
rect 2666 -1335 2678 -1301
rect 2470 -1341 2678 -1335
rect 3042 -1301 3250 -1295
rect 3042 -1335 3054 -1301
rect 3238 -1335 3250 -1301
rect 3042 -1341 3250 -1335
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 12.9 l 2 m 1 nf 12 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
