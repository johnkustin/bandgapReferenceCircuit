.option SEED=random
.ic v(x0.amplifier_0/Vgate)=0 v(x0.amplifier_0/vg)=0 
+ v(x0.amplifier_0/Vx)=0 v(x0.amplifier_0/vq)=0 v(Vbg)=0 
+ v(x0.amplifier_0/va)=0 v(x0.amplifier_0/vb)=0
.param mc_mm_switch=1
.param VDD=1.8

V1 VDD GND {VDD} pwl 0us 0 1us {VDD}
V2 porst GND 0 pulse(0V 1.8V 2us 1us 1us 1us)
V3 VSUBS GND 0

X0 Vbg porst VDD GND bandgaptop_flat

.option RSHUNT=1e20

.control

let run=1
option temp=27

  dowhile run <= 400
    if run > 1
      reset
      set appendwrite
    end
    save all

    let randomseed = $rndseed
    tran 1n 11u

    write TESTTYPENAMEHERE_mc_1_27degc_run_{$&run}.raw vbg
    write TESTTYPENAMEHERE_mc_1_27degc_run_{$&run}_randomseed.raw randomseed
    let run = run + 1
  end

.endc

.GLOBAL VDD
.GLOBAL GND
.GLOBAL VSUBS
.end

