magic
tech sky130A
magscale 1 2
timestamp 1621270775
<< error_p >>
rect -5116 2990 -4820 3500
rect -4796 3450 -4476 3451
rect -4796 3334 -4258 3450
rect -4796 2990 -4156 3334
rect -3994 2990 -3698 3500
rect -3674 3450 -3354 3451
rect -3674 3334 -3136 3450
rect -3674 2990 -3034 3334
rect -2872 2990 -2576 3500
rect -2552 3450 -2232 3451
rect -2552 3334 -2014 3450
rect -2552 2990 -1912 3334
rect -1750 2990 -1454 3500
rect -1430 3450 -1110 3451
rect -1430 3334 -892 3450
rect -1430 2990 -790 3334
rect -628 2990 -332 3500
rect -308 3450 12 3451
rect -308 3334 230 3450
rect -308 2990 332 3334
rect 494 2990 790 3500
rect 814 3450 1134 3451
rect 814 3334 1352 3450
rect 814 2990 1454 3334
rect 1616 2990 1912 3500
rect 1936 3450 2256 3451
rect 1936 3334 2474 3450
rect 1936 2990 2576 3334
rect 2738 2990 3034 3500
rect 3058 3450 3378 3451
rect 3058 3334 3596 3450
rect 3058 2990 3698 3334
rect 3860 2990 4156 3500
rect 4180 3450 4500 3451
rect 4180 3334 4718 3450
rect 4180 2990 4820 3334
rect 4982 2990 5278 3500
rect 5302 3071 5598 3451
rect 5302 2990 5622 3071
rect -5600 2850 5622 2990
rect -5116 2750 -4820 2850
rect -4796 2849 -4476 2850
rect -4796 2750 -4476 2751
rect -3994 2750 -3698 2850
rect -3674 2849 -3354 2850
rect -3674 2750 -3354 2751
rect -2872 2750 -2576 2850
rect -2552 2849 -2232 2850
rect -2552 2750 -2232 2751
rect -1750 2750 -1454 2850
rect -1430 2849 -1110 2850
rect -1430 2750 -1110 2751
rect -628 2750 -332 2850
rect -308 2849 12 2850
rect -308 2750 12 2751
rect 494 2750 790 2850
rect 814 2849 1134 2850
rect 814 2750 1134 2751
rect 1616 2750 1912 2850
rect 1936 2849 2256 2850
rect 1936 2750 2256 2751
rect 2738 2750 3034 2850
rect 3058 2849 3378 2850
rect 3058 2750 3378 2751
rect 3860 2750 4156 2850
rect 4180 2849 4500 2850
rect 4180 2750 4500 2751
rect 4982 2750 5278 2850
rect 5302 2849 5622 2850
rect 5302 2750 5622 2751
rect -5600 2610 5622 2750
rect -5116 2290 -4820 2610
rect -4796 2290 -4156 2610
rect -3994 2290 -3698 2610
rect -3674 2290 -3034 2610
rect -2872 2290 -2576 2610
rect -2552 2290 -1912 2610
rect -1750 2290 -1454 2610
rect -1430 2290 -790 2610
rect -628 2290 -332 2610
rect -308 2290 332 2610
rect 494 2290 790 2610
rect 814 2290 1454 2610
rect 1616 2290 1912 2610
rect 1936 2290 2576 2610
rect 2738 2290 3034 2610
rect 3058 2290 3698 2610
rect 3860 2290 4156 2610
rect 4180 2290 4820 2610
rect 4982 2290 5278 2610
rect 5302 2529 5622 2610
rect 5302 2371 5598 2529
rect 5302 2290 5622 2371
rect -5600 2150 5622 2290
rect -5116 2050 -4820 2150
rect -4796 2149 -4476 2150
rect -4796 2050 -4476 2051
rect -3994 2050 -3698 2150
rect -3674 2149 -3354 2150
rect -3674 2050 -3354 2051
rect -2872 2050 -2576 2150
rect -2552 2149 -2232 2150
rect -2552 2050 -2232 2051
rect -1750 2050 -1454 2150
rect -1430 2149 -1110 2150
rect -1430 2050 -1110 2051
rect -628 2050 -332 2150
rect -308 2149 12 2150
rect -308 2050 12 2051
rect 494 2050 790 2150
rect 814 2149 1134 2150
rect 814 2050 1134 2051
rect 1616 2050 1912 2150
rect 1936 2149 2256 2150
rect 1936 2050 2256 2051
rect 2738 2050 3034 2150
rect 3058 2149 3378 2150
rect 3058 2050 3378 2051
rect 3860 2050 4156 2150
rect 4180 2149 4500 2150
rect 4180 2050 4500 2051
rect 4982 2050 5278 2150
rect 5302 2149 5622 2150
rect 5302 2050 5622 2051
rect -5600 1910 5622 2050
rect -5116 1590 -4820 1910
rect -4796 1590 -4156 1910
rect -3994 1590 -3698 1910
rect -3674 1590 -3034 1910
rect -2872 1590 -2576 1910
rect -2552 1590 -1912 1910
rect -1750 1590 -1454 1910
rect -1430 1590 -790 1910
rect -628 1590 -332 1910
rect -308 1590 332 1910
rect 494 1590 790 1910
rect 814 1590 1454 1910
rect 1616 1590 1912 1910
rect 1936 1590 2576 1910
rect 2738 1590 3034 1910
rect 3058 1590 3698 1910
rect 3860 1590 4156 1910
rect 4180 1590 4820 1910
rect 4982 1590 5278 1910
rect 5302 1829 5622 1910
rect 5302 1671 5598 1829
rect 5302 1590 5622 1671
rect -5600 1450 5622 1590
rect -5116 1350 -4820 1450
rect -4796 1449 -4476 1450
rect -4796 1350 -4476 1351
rect -3994 1350 -3698 1450
rect -3674 1449 -3354 1450
rect -3674 1350 -3354 1351
rect -2872 1350 -2576 1450
rect -2552 1449 -2232 1450
rect -2552 1350 -2232 1351
rect -1750 1350 -1454 1450
rect -1430 1449 -1110 1450
rect -1430 1350 -1110 1351
rect -628 1350 -332 1450
rect -308 1449 12 1450
rect -308 1350 12 1351
rect 494 1350 790 1450
rect 814 1449 1134 1450
rect 814 1350 1134 1351
rect 1616 1350 1912 1450
rect 1936 1449 2256 1450
rect 1936 1350 2256 1351
rect 2738 1350 3034 1450
rect 3058 1449 3378 1450
rect 3058 1350 3378 1351
rect 3860 1350 4156 1450
rect 4180 1449 4500 1450
rect 4180 1350 4500 1351
rect 4982 1350 5278 1450
rect 5302 1449 5622 1450
rect 5302 1350 5622 1351
rect -5600 1210 5622 1350
rect -5116 890 -4820 1210
rect -4796 890 -4156 1210
rect -3994 890 -3698 1210
rect -3674 890 -3034 1210
rect -2872 890 -2576 1210
rect -2552 890 -1912 1210
rect -1750 890 -1454 1210
rect -1430 890 -790 1210
rect -628 890 -332 1210
rect -308 890 332 1210
rect 494 890 790 1210
rect 814 890 1454 1210
rect 1616 890 1912 1210
rect 1936 890 2576 1210
rect 2738 890 3034 1210
rect 3058 890 3698 1210
rect 3860 890 4156 1210
rect 4180 890 4820 1210
rect 4982 890 5278 1210
rect 5302 1129 5622 1210
rect 5302 971 5598 1129
rect 5302 890 5622 971
rect -5600 750 5622 890
rect -5116 650 -4820 750
rect -4796 749 -4476 750
rect -4796 650 -4476 651
rect -3994 650 -3698 750
rect -3674 749 -3354 750
rect -3674 650 -3354 651
rect -2872 650 -2576 750
rect -2552 749 -2232 750
rect -2552 650 -2232 651
rect -1750 650 -1454 750
rect -1430 749 -1110 750
rect -1430 650 -1110 651
rect -628 650 -332 750
rect -308 749 12 750
rect -308 650 12 651
rect 494 650 790 750
rect 814 749 1134 750
rect 814 650 1134 651
rect 1616 650 1912 750
rect 1936 749 2256 750
rect 1936 650 2256 651
rect 2738 650 3034 750
rect 3058 749 3378 750
rect 3058 650 3378 651
rect 3860 650 4156 750
rect 4180 749 4500 750
rect 4180 650 4500 651
rect 4982 650 5278 750
rect 5302 749 5622 750
rect 5302 650 5622 651
rect -5600 510 5622 650
rect -5116 190 -4820 510
rect -4796 190 -4156 510
rect -3994 190 -3698 510
rect -3674 190 -3034 510
rect -2872 190 -2576 510
rect -2552 190 -1912 510
rect -1750 190 -1454 510
rect -1430 190 -790 510
rect -628 190 -332 510
rect -308 190 332 510
rect 494 190 790 510
rect 814 190 1454 510
rect 1616 190 1912 510
rect 1936 190 2576 510
rect 2738 190 3034 510
rect 3058 190 3698 510
rect 3860 190 4156 510
rect 4180 190 4820 510
rect 4982 190 5278 510
rect 5302 429 5622 510
rect 5302 271 5598 429
rect 5302 190 5622 271
rect -5600 50 5622 190
rect -5116 -50 -4820 50
rect -4796 49 -4476 50
rect -4796 -50 -4476 -49
rect -3994 -50 -3698 50
rect -3674 49 -3354 50
rect -3674 -50 -3354 -49
rect -2872 -50 -2576 50
rect -2552 49 -2232 50
rect -2552 -50 -2232 -49
rect -1750 -50 -1454 50
rect -1430 49 -1110 50
rect -1430 -50 -1110 -49
rect -628 -50 -332 50
rect -308 49 12 50
rect -308 -50 12 -49
rect 494 -50 790 50
rect 814 49 1134 50
rect 814 -50 1134 -49
rect 1616 -50 1912 50
rect 1936 49 2256 50
rect 1936 -50 2256 -49
rect 2738 -50 3034 50
rect 3058 49 3378 50
rect 3058 -50 3378 -49
rect 3860 -50 4156 50
rect 4180 49 4500 50
rect 4180 -50 4500 -49
rect 4982 -50 5278 50
rect 5302 49 5622 50
rect 5302 -50 5622 -49
rect -5600 -190 5622 -50
rect -5116 -510 -4820 -190
rect -4796 -510 -4156 -190
rect -3994 -510 -3698 -190
rect -3674 -510 -3034 -190
rect -2872 -510 -2576 -190
rect -2552 -510 -1912 -190
rect -1750 -510 -1454 -190
rect -1430 -510 -790 -190
rect -628 -510 -332 -190
rect -308 -510 332 -190
rect 494 -510 790 -190
rect 814 -510 1454 -190
rect 1616 -510 1912 -190
rect 1936 -510 2576 -190
rect 2738 -510 3034 -190
rect 3058 -510 3698 -190
rect 3860 -510 4156 -190
rect 4180 -510 4820 -190
rect 4982 -510 5278 -190
rect 5302 -271 5622 -190
rect 5302 -429 5598 -271
rect 5302 -510 5622 -429
rect -5600 -650 5622 -510
rect -5116 -750 -4820 -650
rect -4796 -651 -4476 -650
rect -4796 -750 -4476 -749
rect -3994 -750 -3698 -650
rect -3674 -651 -3354 -650
rect -3674 -750 -3354 -749
rect -2872 -750 -2576 -650
rect -2552 -651 -2232 -650
rect -2552 -750 -2232 -749
rect -1750 -750 -1454 -650
rect -1430 -651 -1110 -650
rect -1430 -750 -1110 -749
rect -628 -750 -332 -650
rect -308 -651 12 -650
rect -308 -750 12 -749
rect 494 -750 790 -650
rect 814 -651 1134 -650
rect 814 -750 1134 -749
rect 1616 -750 1912 -650
rect 1936 -651 2256 -650
rect 1936 -750 2256 -749
rect 2738 -750 3034 -650
rect 3058 -651 3378 -650
rect 3058 -750 3378 -749
rect 3860 -750 4156 -650
rect 4180 -651 4500 -650
rect 4180 -750 4500 -749
rect 4982 -750 5278 -650
rect 5302 -651 5622 -650
rect 5302 -750 5622 -749
rect -5600 -890 5622 -750
rect -5116 -1210 -4820 -890
rect -4796 -1210 -4156 -890
rect -3994 -1210 -3698 -890
rect -3674 -1210 -3034 -890
rect -2872 -1210 -2576 -890
rect -2552 -1210 -1912 -890
rect -1750 -1210 -1454 -890
rect -1430 -1210 -790 -890
rect -628 -1210 -332 -890
rect -308 -1210 332 -890
rect 494 -1210 790 -890
rect 814 -1210 1454 -890
rect 1616 -1210 1912 -890
rect 1936 -1210 2576 -890
rect 2738 -1210 3034 -890
rect 3058 -1210 3698 -890
rect 3860 -1210 4156 -890
rect 4180 -1210 4820 -890
rect 4982 -1210 5278 -890
rect 5302 -971 5622 -890
rect 5302 -1129 5598 -971
rect 5302 -1210 5622 -1129
rect -5600 -1350 5622 -1210
rect -5116 -1450 -4820 -1350
rect -4796 -1351 -4476 -1350
rect -4796 -1450 -4476 -1449
rect -3994 -1450 -3698 -1350
rect -3674 -1351 -3354 -1350
rect -3674 -1450 -3354 -1449
rect -2872 -1450 -2576 -1350
rect -2552 -1351 -2232 -1350
rect -2552 -1450 -2232 -1449
rect -1750 -1450 -1454 -1350
rect -1430 -1351 -1110 -1350
rect -1430 -1450 -1110 -1449
rect -628 -1450 -332 -1350
rect -308 -1351 12 -1350
rect -308 -1450 12 -1449
rect 494 -1450 790 -1350
rect 814 -1351 1134 -1350
rect 814 -1450 1134 -1449
rect 1616 -1450 1912 -1350
rect 1936 -1351 2256 -1350
rect 1936 -1450 2256 -1449
rect 2738 -1450 3034 -1350
rect 3058 -1351 3378 -1350
rect 3058 -1450 3378 -1449
rect 3860 -1450 4156 -1350
rect 4180 -1351 4500 -1350
rect 4180 -1450 4500 -1449
rect 4982 -1450 5278 -1350
rect 5302 -1351 5622 -1350
rect 5302 -1450 5622 -1449
rect -5600 -1590 5622 -1450
rect -5116 -1910 -4820 -1590
rect -4796 -1910 -4156 -1590
rect -3994 -1910 -3698 -1590
rect -3674 -1910 -3034 -1590
rect -2872 -1910 -2576 -1590
rect -2552 -1910 -1912 -1590
rect -1750 -1910 -1454 -1590
rect -1430 -1910 -790 -1590
rect -628 -1910 -332 -1590
rect -308 -1910 332 -1590
rect 494 -1910 790 -1590
rect 814 -1910 1454 -1590
rect 1616 -1910 1912 -1590
rect 1936 -1910 2576 -1590
rect 2738 -1910 3034 -1590
rect 3058 -1910 3698 -1590
rect 3860 -1910 4156 -1590
rect 4180 -1910 4820 -1590
rect 4982 -1910 5278 -1590
rect 5302 -1671 5622 -1590
rect 5302 -1829 5598 -1671
rect 5302 -1910 5622 -1829
rect -5600 -2050 5622 -1910
rect -5116 -2150 -4820 -2050
rect -4796 -2051 -4476 -2050
rect -4796 -2150 -4476 -2149
rect -3994 -2150 -3698 -2050
rect -3674 -2051 -3354 -2050
rect -3674 -2150 -3354 -2149
rect -2872 -2150 -2576 -2050
rect -2552 -2051 -2232 -2050
rect -2552 -2150 -2232 -2149
rect -1750 -2150 -1454 -2050
rect -1430 -2051 -1110 -2050
rect -1430 -2150 -1110 -2149
rect -628 -2150 -332 -2050
rect -308 -2051 12 -2050
rect -308 -2150 12 -2149
rect 494 -2150 790 -2050
rect 814 -2051 1134 -2050
rect 814 -2150 1134 -2149
rect 1616 -2150 1912 -2050
rect 1936 -2051 2256 -2050
rect 1936 -2150 2256 -2149
rect 2738 -2150 3034 -2050
rect 3058 -2051 3378 -2050
rect 3058 -2150 3378 -2149
rect 3860 -2150 4156 -2050
rect 4180 -2051 4500 -2050
rect 4180 -2150 4500 -2149
rect 4982 -2150 5278 -2050
rect 5302 -2051 5622 -2050
rect 5302 -2150 5622 -2149
rect -5600 -2290 5622 -2150
rect -5116 -2610 -4820 -2290
rect -4796 -2610 -4156 -2290
rect -3994 -2610 -3698 -2290
rect -3674 -2610 -3034 -2290
rect -2872 -2610 -2576 -2290
rect -2552 -2610 -1912 -2290
rect -1750 -2610 -1454 -2290
rect -1430 -2610 -790 -2290
rect -628 -2610 -332 -2290
rect -308 -2610 332 -2290
rect 494 -2610 790 -2290
rect 814 -2610 1454 -2290
rect 1616 -2610 1912 -2290
rect 1936 -2610 2576 -2290
rect 2738 -2610 3034 -2290
rect 3058 -2610 3698 -2290
rect 3860 -2610 4156 -2290
rect 4180 -2610 4820 -2290
rect 4982 -2610 5278 -2290
rect 5302 -2371 5622 -2290
rect 5302 -2529 5598 -2371
rect 5302 -2610 5622 -2529
rect -5600 -2750 5622 -2610
rect -5116 -2850 -4820 -2750
rect -4796 -2751 -4476 -2750
rect -4796 -2850 -4476 -2849
rect -3994 -2850 -3698 -2750
rect -3674 -2751 -3354 -2750
rect -3674 -2850 -3354 -2849
rect -2872 -2850 -2576 -2750
rect -2552 -2751 -2232 -2750
rect -2552 -2850 -2232 -2849
rect -1750 -2850 -1454 -2750
rect -1430 -2751 -1110 -2750
rect -1430 -2850 -1110 -2849
rect -628 -2850 -332 -2750
rect -308 -2751 12 -2750
rect -308 -2850 12 -2849
rect 494 -2850 790 -2750
rect 814 -2751 1134 -2750
rect 814 -2850 1134 -2849
rect 1616 -2850 1912 -2750
rect 1936 -2751 2256 -2750
rect 1936 -2850 2256 -2849
rect 2738 -2850 3034 -2750
rect 3058 -2751 3378 -2750
rect 3058 -2850 3378 -2849
rect 3860 -2850 4156 -2750
rect 4180 -2751 4500 -2750
rect 4180 -2850 4500 -2849
rect 4982 -2850 5278 -2750
rect 5302 -2751 5622 -2750
rect 5302 -2850 5622 -2849
rect -5600 -2990 5622 -2850
rect -5116 -3500 -4820 -2990
rect -4796 -3334 -4156 -2990
rect -4796 -3450 -4258 -3334
rect -4796 -3451 -4476 -3450
rect -3994 -3500 -3698 -2990
rect -3674 -3334 -3034 -2990
rect -3674 -3450 -3136 -3334
rect -3674 -3451 -3354 -3450
rect -2872 -3500 -2576 -2990
rect -2552 -3334 -1912 -2990
rect -2552 -3450 -2014 -3334
rect -2552 -3451 -2232 -3450
rect -1750 -3500 -1454 -2990
rect -1430 -3334 -790 -2990
rect -1430 -3450 -892 -3334
rect -1430 -3451 -1110 -3450
rect -628 -3500 -332 -2990
rect -308 -3334 332 -2990
rect -308 -3450 230 -3334
rect -308 -3451 12 -3450
rect 494 -3500 790 -2990
rect 814 -3334 1454 -2990
rect 814 -3450 1352 -3334
rect 814 -3451 1134 -3450
rect 1616 -3500 1912 -2990
rect 1936 -3334 2576 -2990
rect 1936 -3450 2474 -3334
rect 1936 -3451 2256 -3450
rect 2738 -3500 3034 -2990
rect 3058 -3334 3698 -2990
rect 3058 -3450 3596 -3334
rect 3058 -3451 3378 -3450
rect 3860 -3500 4156 -2990
rect 4180 -3334 4820 -2990
rect 4180 -3450 4718 -3334
rect 4180 -3451 4500 -3450
rect 4982 -3500 5278 -2990
rect 5302 -3071 5622 -2990
rect 5302 -3451 5598 -3071
<< metal4 >>
rect -5600 3409 -4498 3450
rect -5600 2891 -4754 3409
rect -4518 2891 -4498 3409
rect -5600 2850 -4498 2891
rect -4478 3409 -3376 3450
rect -4478 2891 -3632 3409
rect -3396 2891 -3376 3409
rect -4478 2850 -3376 2891
rect -3356 3409 -2254 3450
rect -3356 2891 -2510 3409
rect -2274 2891 -2254 3409
rect -3356 2850 -2254 2891
rect -2234 3409 -1132 3450
rect -2234 2891 -1388 3409
rect -1152 2891 -1132 3409
rect -2234 2850 -1132 2891
rect -1112 3409 -10 3450
rect -1112 2891 -266 3409
rect -30 2891 -10 3409
rect -1112 2850 -10 2891
rect 10 3409 1112 3450
rect 10 2891 856 3409
rect 1092 2891 1112 3409
rect 10 2850 1112 2891
rect 1132 3409 2234 3450
rect 1132 2891 1978 3409
rect 2214 2891 2234 3409
rect 1132 2850 2234 2891
rect 2254 3409 3356 3450
rect 2254 2891 3100 3409
rect 3336 2891 3356 3409
rect 2254 2850 3356 2891
rect 3376 3409 4478 3450
rect 3376 2891 4222 3409
rect 4458 2891 4478 3409
rect 3376 2850 4478 2891
rect 4498 3409 5600 3450
rect 4498 2891 5344 3409
rect 5580 2891 5600 3409
rect 4498 2850 5600 2891
rect -5600 2709 -4498 2750
rect -5600 2191 -4754 2709
rect -4518 2191 -4498 2709
rect -5600 2150 -4498 2191
rect -4478 2709 -3376 2750
rect -4478 2191 -3632 2709
rect -3396 2191 -3376 2709
rect -4478 2150 -3376 2191
rect -3356 2709 -2254 2750
rect -3356 2191 -2510 2709
rect -2274 2191 -2254 2709
rect -3356 2150 -2254 2191
rect -2234 2709 -1132 2750
rect -2234 2191 -1388 2709
rect -1152 2191 -1132 2709
rect -2234 2150 -1132 2191
rect -1112 2709 -10 2750
rect -1112 2191 -266 2709
rect -30 2191 -10 2709
rect -1112 2150 -10 2191
rect 10 2709 1112 2750
rect 10 2191 856 2709
rect 1092 2191 1112 2709
rect 10 2150 1112 2191
rect 1132 2709 2234 2750
rect 1132 2191 1978 2709
rect 2214 2191 2234 2709
rect 1132 2150 2234 2191
rect 2254 2709 3356 2750
rect 2254 2191 3100 2709
rect 3336 2191 3356 2709
rect 2254 2150 3356 2191
rect 3376 2709 4478 2750
rect 3376 2191 4222 2709
rect 4458 2191 4478 2709
rect 3376 2150 4478 2191
rect 4498 2709 5600 2750
rect 4498 2191 5344 2709
rect 5580 2191 5600 2709
rect 4498 2150 5600 2191
rect -5600 2009 -4498 2050
rect -5600 1491 -4754 2009
rect -4518 1491 -4498 2009
rect -5600 1450 -4498 1491
rect -4478 2009 -3376 2050
rect -4478 1491 -3632 2009
rect -3396 1491 -3376 2009
rect -4478 1450 -3376 1491
rect -3356 2009 -2254 2050
rect -3356 1491 -2510 2009
rect -2274 1491 -2254 2009
rect -3356 1450 -2254 1491
rect -2234 2009 -1132 2050
rect -2234 1491 -1388 2009
rect -1152 1491 -1132 2009
rect -2234 1450 -1132 1491
rect -1112 2009 -10 2050
rect -1112 1491 -266 2009
rect -30 1491 -10 2009
rect -1112 1450 -10 1491
rect 10 2009 1112 2050
rect 10 1491 856 2009
rect 1092 1491 1112 2009
rect 10 1450 1112 1491
rect 1132 2009 2234 2050
rect 1132 1491 1978 2009
rect 2214 1491 2234 2009
rect 1132 1450 2234 1491
rect 2254 2009 3356 2050
rect 2254 1491 3100 2009
rect 3336 1491 3356 2009
rect 2254 1450 3356 1491
rect 3376 2009 4478 2050
rect 3376 1491 4222 2009
rect 4458 1491 4478 2009
rect 3376 1450 4478 1491
rect 4498 2009 5600 2050
rect 4498 1491 5344 2009
rect 5580 1491 5600 2009
rect 4498 1450 5600 1491
rect -5600 1309 -4498 1350
rect -5600 791 -4754 1309
rect -4518 791 -4498 1309
rect -5600 750 -4498 791
rect -4478 1309 -3376 1350
rect -4478 791 -3632 1309
rect -3396 791 -3376 1309
rect -4478 750 -3376 791
rect -3356 1309 -2254 1350
rect -3356 791 -2510 1309
rect -2274 791 -2254 1309
rect -3356 750 -2254 791
rect -2234 1309 -1132 1350
rect -2234 791 -1388 1309
rect -1152 791 -1132 1309
rect -2234 750 -1132 791
rect -1112 1309 -10 1350
rect -1112 791 -266 1309
rect -30 791 -10 1309
rect -1112 750 -10 791
rect 10 1309 1112 1350
rect 10 791 856 1309
rect 1092 791 1112 1309
rect 10 750 1112 791
rect 1132 1309 2234 1350
rect 1132 791 1978 1309
rect 2214 791 2234 1309
rect 1132 750 2234 791
rect 2254 1309 3356 1350
rect 2254 791 3100 1309
rect 3336 791 3356 1309
rect 2254 750 3356 791
rect 3376 1309 4478 1350
rect 3376 791 4222 1309
rect 4458 791 4478 1309
rect 3376 750 4478 791
rect 4498 1309 5600 1350
rect 4498 791 5344 1309
rect 5580 791 5600 1309
rect 4498 750 5600 791
rect -5600 609 -4498 650
rect -5600 91 -4754 609
rect -4518 91 -4498 609
rect -5600 50 -4498 91
rect -4478 609 -3376 650
rect -4478 91 -3632 609
rect -3396 91 -3376 609
rect -4478 50 -3376 91
rect -3356 609 -2254 650
rect -3356 91 -2510 609
rect -2274 91 -2254 609
rect -3356 50 -2254 91
rect -2234 609 -1132 650
rect -2234 91 -1388 609
rect -1152 91 -1132 609
rect -2234 50 -1132 91
rect -1112 609 -10 650
rect -1112 91 -266 609
rect -30 91 -10 609
rect -1112 50 -10 91
rect 10 609 1112 650
rect 10 91 856 609
rect 1092 91 1112 609
rect 10 50 1112 91
rect 1132 609 2234 650
rect 1132 91 1978 609
rect 2214 91 2234 609
rect 1132 50 2234 91
rect 2254 609 3356 650
rect 2254 91 3100 609
rect 3336 91 3356 609
rect 2254 50 3356 91
rect 3376 609 4478 650
rect 3376 91 4222 609
rect 4458 91 4478 609
rect 3376 50 4478 91
rect 4498 609 5600 650
rect 4498 91 5344 609
rect 5580 91 5600 609
rect 4498 50 5600 91
rect -5600 -91 -4498 -50
rect -5600 -609 -4754 -91
rect -4518 -609 -4498 -91
rect -5600 -650 -4498 -609
rect -4478 -91 -3376 -50
rect -4478 -609 -3632 -91
rect -3396 -609 -3376 -91
rect -4478 -650 -3376 -609
rect -3356 -91 -2254 -50
rect -3356 -609 -2510 -91
rect -2274 -609 -2254 -91
rect -3356 -650 -2254 -609
rect -2234 -91 -1132 -50
rect -2234 -609 -1388 -91
rect -1152 -609 -1132 -91
rect -2234 -650 -1132 -609
rect -1112 -91 -10 -50
rect -1112 -609 -266 -91
rect -30 -609 -10 -91
rect -1112 -650 -10 -609
rect 10 -91 1112 -50
rect 10 -609 856 -91
rect 1092 -609 1112 -91
rect 10 -650 1112 -609
rect 1132 -91 2234 -50
rect 1132 -609 1978 -91
rect 2214 -609 2234 -91
rect 1132 -650 2234 -609
rect 2254 -91 3356 -50
rect 2254 -609 3100 -91
rect 3336 -609 3356 -91
rect 2254 -650 3356 -609
rect 3376 -91 4478 -50
rect 3376 -609 4222 -91
rect 4458 -609 4478 -91
rect 3376 -650 4478 -609
rect 4498 -91 5600 -50
rect 4498 -609 5344 -91
rect 5580 -609 5600 -91
rect 4498 -650 5600 -609
rect -5600 -791 -4498 -750
rect -5600 -1309 -4754 -791
rect -4518 -1309 -4498 -791
rect -5600 -1350 -4498 -1309
rect -4478 -791 -3376 -750
rect -4478 -1309 -3632 -791
rect -3396 -1309 -3376 -791
rect -4478 -1350 -3376 -1309
rect -3356 -791 -2254 -750
rect -3356 -1309 -2510 -791
rect -2274 -1309 -2254 -791
rect -3356 -1350 -2254 -1309
rect -2234 -791 -1132 -750
rect -2234 -1309 -1388 -791
rect -1152 -1309 -1132 -791
rect -2234 -1350 -1132 -1309
rect -1112 -791 -10 -750
rect -1112 -1309 -266 -791
rect -30 -1309 -10 -791
rect -1112 -1350 -10 -1309
rect 10 -791 1112 -750
rect 10 -1309 856 -791
rect 1092 -1309 1112 -791
rect 10 -1350 1112 -1309
rect 1132 -791 2234 -750
rect 1132 -1309 1978 -791
rect 2214 -1309 2234 -791
rect 1132 -1350 2234 -1309
rect 2254 -791 3356 -750
rect 2254 -1309 3100 -791
rect 3336 -1309 3356 -791
rect 2254 -1350 3356 -1309
rect 3376 -791 4478 -750
rect 3376 -1309 4222 -791
rect 4458 -1309 4478 -791
rect 3376 -1350 4478 -1309
rect 4498 -791 5600 -750
rect 4498 -1309 5344 -791
rect 5580 -1309 5600 -791
rect 4498 -1350 5600 -1309
rect -5600 -1491 -4498 -1450
rect -5600 -2009 -4754 -1491
rect -4518 -2009 -4498 -1491
rect -5600 -2050 -4498 -2009
rect -4478 -1491 -3376 -1450
rect -4478 -2009 -3632 -1491
rect -3396 -2009 -3376 -1491
rect -4478 -2050 -3376 -2009
rect -3356 -1491 -2254 -1450
rect -3356 -2009 -2510 -1491
rect -2274 -2009 -2254 -1491
rect -3356 -2050 -2254 -2009
rect -2234 -1491 -1132 -1450
rect -2234 -2009 -1388 -1491
rect -1152 -2009 -1132 -1491
rect -2234 -2050 -1132 -2009
rect -1112 -1491 -10 -1450
rect -1112 -2009 -266 -1491
rect -30 -2009 -10 -1491
rect -1112 -2050 -10 -2009
rect 10 -1491 1112 -1450
rect 10 -2009 856 -1491
rect 1092 -2009 1112 -1491
rect 10 -2050 1112 -2009
rect 1132 -1491 2234 -1450
rect 1132 -2009 1978 -1491
rect 2214 -2009 2234 -1491
rect 1132 -2050 2234 -2009
rect 2254 -1491 3356 -1450
rect 2254 -2009 3100 -1491
rect 3336 -2009 3356 -1491
rect 2254 -2050 3356 -2009
rect 3376 -1491 4478 -1450
rect 3376 -2009 4222 -1491
rect 4458 -2009 4478 -1491
rect 3376 -2050 4478 -2009
rect 4498 -1491 5600 -1450
rect 4498 -2009 5344 -1491
rect 5580 -2009 5600 -1491
rect 4498 -2050 5600 -2009
rect -5600 -2191 -4498 -2150
rect -5600 -2709 -4754 -2191
rect -4518 -2709 -4498 -2191
rect -5600 -2750 -4498 -2709
rect -4478 -2191 -3376 -2150
rect -4478 -2709 -3632 -2191
rect -3396 -2709 -3376 -2191
rect -4478 -2750 -3376 -2709
rect -3356 -2191 -2254 -2150
rect -3356 -2709 -2510 -2191
rect -2274 -2709 -2254 -2191
rect -3356 -2750 -2254 -2709
rect -2234 -2191 -1132 -2150
rect -2234 -2709 -1388 -2191
rect -1152 -2709 -1132 -2191
rect -2234 -2750 -1132 -2709
rect -1112 -2191 -10 -2150
rect -1112 -2709 -266 -2191
rect -30 -2709 -10 -2191
rect -1112 -2750 -10 -2709
rect 10 -2191 1112 -2150
rect 10 -2709 856 -2191
rect 1092 -2709 1112 -2191
rect 10 -2750 1112 -2709
rect 1132 -2191 2234 -2150
rect 1132 -2709 1978 -2191
rect 2214 -2709 2234 -2191
rect 1132 -2750 2234 -2709
rect 2254 -2191 3356 -2150
rect 2254 -2709 3100 -2191
rect 3336 -2709 3356 -2191
rect 2254 -2750 3356 -2709
rect 3376 -2191 4478 -2150
rect 3376 -2709 4222 -2191
rect 4458 -2709 4478 -2191
rect 3376 -2750 4478 -2709
rect 4498 -2191 5600 -2150
rect 4498 -2709 5344 -2191
rect 5580 -2709 5600 -2191
rect 4498 -2750 5600 -2709
rect -5600 -2891 -4498 -2850
rect -5600 -3409 -4754 -2891
rect -4518 -3409 -4498 -2891
rect -5600 -3450 -4498 -3409
rect -4478 -2891 -3376 -2850
rect -4478 -3409 -3632 -2891
rect -3396 -3409 -3376 -2891
rect -4478 -3450 -3376 -3409
rect -3356 -2891 -2254 -2850
rect -3356 -3409 -2510 -2891
rect -2274 -3409 -2254 -2891
rect -3356 -3450 -2254 -3409
rect -2234 -2891 -1132 -2850
rect -2234 -3409 -1388 -2891
rect -1152 -3409 -1132 -2891
rect -2234 -3450 -1132 -3409
rect -1112 -2891 -10 -2850
rect -1112 -3409 -266 -2891
rect -30 -3409 -10 -2891
rect -1112 -3450 -10 -3409
rect 10 -2891 1112 -2850
rect 10 -3409 856 -2891
rect 1092 -3409 1112 -2891
rect 10 -3450 1112 -3409
rect 1132 -2891 2234 -2850
rect 1132 -3409 1978 -2891
rect 2214 -3409 2234 -2891
rect 1132 -3450 2234 -3409
rect 2254 -2891 3356 -2850
rect 2254 -3409 3100 -2891
rect 3336 -3409 3356 -2891
rect 2254 -3450 3356 -3409
rect 3376 -2891 4478 -2850
rect 3376 -3409 4222 -2891
rect 4458 -3409 4478 -2891
rect 3376 -3450 4478 -3409
rect 4498 -2891 5600 -2850
rect 4498 -3409 5344 -2891
rect 5580 -3409 5600 -2891
rect 4498 -3450 5600 -3409
<< via4 >>
rect -4754 2891 -4518 3409
rect -3632 2891 -3396 3409
rect -2510 2891 -2274 3409
rect -1388 2891 -1152 3409
rect -266 2891 -30 3409
rect 856 2891 1092 3409
rect 1978 2891 2214 3409
rect 3100 2891 3336 3409
rect 4222 2891 4458 3409
rect 5344 2891 5580 3409
rect -4754 2191 -4518 2709
rect -3632 2191 -3396 2709
rect -2510 2191 -2274 2709
rect -1388 2191 -1152 2709
rect -266 2191 -30 2709
rect 856 2191 1092 2709
rect 1978 2191 2214 2709
rect 3100 2191 3336 2709
rect 4222 2191 4458 2709
rect 5344 2191 5580 2709
rect -4754 1491 -4518 2009
rect -3632 1491 -3396 2009
rect -2510 1491 -2274 2009
rect -1388 1491 -1152 2009
rect -266 1491 -30 2009
rect 856 1491 1092 2009
rect 1978 1491 2214 2009
rect 3100 1491 3336 2009
rect 4222 1491 4458 2009
rect 5344 1491 5580 2009
rect -4754 791 -4518 1309
rect -3632 791 -3396 1309
rect -2510 791 -2274 1309
rect -1388 791 -1152 1309
rect -266 791 -30 1309
rect 856 791 1092 1309
rect 1978 791 2214 1309
rect 3100 791 3336 1309
rect 4222 791 4458 1309
rect 5344 791 5580 1309
rect -4754 91 -4518 609
rect -3632 91 -3396 609
rect -2510 91 -2274 609
rect -1388 91 -1152 609
rect -266 91 -30 609
rect 856 91 1092 609
rect 1978 91 2214 609
rect 3100 91 3336 609
rect 4222 91 4458 609
rect 5344 91 5580 609
rect -4754 -609 -4518 -91
rect -3632 -609 -3396 -91
rect -2510 -609 -2274 -91
rect -1388 -609 -1152 -91
rect -266 -609 -30 -91
rect 856 -609 1092 -91
rect 1978 -609 2214 -91
rect 3100 -609 3336 -91
rect 4222 -609 4458 -91
rect 5344 -609 5580 -91
rect -4754 -1309 -4518 -791
rect -3632 -1309 -3396 -791
rect -2510 -1309 -2274 -791
rect -1388 -1309 -1152 -791
rect -266 -1309 -30 -791
rect 856 -1309 1092 -791
rect 1978 -1309 2214 -791
rect 3100 -1309 3336 -791
rect 4222 -1309 4458 -791
rect 5344 -1309 5580 -791
rect -4754 -2009 -4518 -1491
rect -3632 -2009 -3396 -1491
rect -2510 -2009 -2274 -1491
rect -1388 -2009 -1152 -1491
rect -266 -2009 -30 -1491
rect 856 -2009 1092 -1491
rect 1978 -2009 2214 -1491
rect 3100 -2009 3336 -1491
rect 4222 -2009 4458 -1491
rect 5344 -2009 5580 -1491
rect -4754 -2709 -4518 -2191
rect -3632 -2709 -3396 -2191
rect -2510 -2709 -2274 -2191
rect -1388 -2709 -1152 -2191
rect -266 -2709 -30 -2191
rect 856 -2709 1092 -2191
rect 1978 -2709 2214 -2191
rect 3100 -2709 3336 -2191
rect 4222 -2709 4458 -2191
rect 5344 -2709 5580 -2191
rect -4754 -3409 -4518 -2891
rect -3632 -3409 -3396 -2891
rect -2510 -3409 -2274 -2891
rect -1388 -3409 -1152 -2891
rect -266 -3409 -30 -2891
rect 856 -3409 1092 -2891
rect 1978 -3409 2214 -2891
rect 3100 -3409 3336 -2891
rect 4222 -3409 4458 -2891
rect 5344 -3409 5580 -2891
<< mimcap2 >>
rect -5500 3310 -5100 3350
rect -5500 2990 -5460 3310
rect -5140 2990 -5100 3310
rect -5500 2950 -5100 2990
rect -4378 3310 -3978 3350
rect -4378 2990 -4338 3310
rect -4018 2990 -3978 3310
rect -4378 2950 -3978 2990
rect -3256 3310 -2856 3350
rect -3256 2990 -3216 3310
rect -2896 2990 -2856 3310
rect -3256 2950 -2856 2990
rect -2134 3310 -1734 3350
rect -2134 2990 -2094 3310
rect -1774 2990 -1734 3310
rect -2134 2950 -1734 2990
rect -1012 3310 -612 3350
rect -1012 2990 -972 3310
rect -652 2990 -612 3310
rect -1012 2950 -612 2990
rect 110 3310 510 3350
rect 110 2990 150 3310
rect 470 2990 510 3310
rect 110 2950 510 2990
rect 1232 3310 1632 3350
rect 1232 2990 1272 3310
rect 1592 2990 1632 3310
rect 1232 2950 1632 2990
rect 2354 3310 2754 3350
rect 2354 2990 2394 3310
rect 2714 2990 2754 3310
rect 2354 2950 2754 2990
rect 3476 3310 3876 3350
rect 3476 2990 3516 3310
rect 3836 2990 3876 3310
rect 3476 2950 3876 2990
rect 4598 3310 4998 3350
rect 4598 2990 4638 3310
rect 4958 2990 4998 3310
rect 4598 2950 4998 2990
rect -5500 2610 -5100 2650
rect -5500 2290 -5460 2610
rect -5140 2290 -5100 2610
rect -5500 2250 -5100 2290
rect -4378 2610 -3978 2650
rect -4378 2290 -4338 2610
rect -4018 2290 -3978 2610
rect -4378 2250 -3978 2290
rect -3256 2610 -2856 2650
rect -3256 2290 -3216 2610
rect -2896 2290 -2856 2610
rect -3256 2250 -2856 2290
rect -2134 2610 -1734 2650
rect -2134 2290 -2094 2610
rect -1774 2290 -1734 2610
rect -2134 2250 -1734 2290
rect -1012 2610 -612 2650
rect -1012 2290 -972 2610
rect -652 2290 -612 2610
rect -1012 2250 -612 2290
rect 110 2610 510 2650
rect 110 2290 150 2610
rect 470 2290 510 2610
rect 110 2250 510 2290
rect 1232 2610 1632 2650
rect 1232 2290 1272 2610
rect 1592 2290 1632 2610
rect 1232 2250 1632 2290
rect 2354 2610 2754 2650
rect 2354 2290 2394 2610
rect 2714 2290 2754 2610
rect 2354 2250 2754 2290
rect 3476 2610 3876 2650
rect 3476 2290 3516 2610
rect 3836 2290 3876 2610
rect 3476 2250 3876 2290
rect 4598 2610 4998 2650
rect 4598 2290 4638 2610
rect 4958 2290 4998 2610
rect 4598 2250 4998 2290
rect -5500 1910 -5100 1950
rect -5500 1590 -5460 1910
rect -5140 1590 -5100 1910
rect -5500 1550 -5100 1590
rect -4378 1910 -3978 1950
rect -4378 1590 -4338 1910
rect -4018 1590 -3978 1910
rect -4378 1550 -3978 1590
rect -3256 1910 -2856 1950
rect -3256 1590 -3216 1910
rect -2896 1590 -2856 1910
rect -3256 1550 -2856 1590
rect -2134 1910 -1734 1950
rect -2134 1590 -2094 1910
rect -1774 1590 -1734 1910
rect -2134 1550 -1734 1590
rect -1012 1910 -612 1950
rect -1012 1590 -972 1910
rect -652 1590 -612 1910
rect -1012 1550 -612 1590
rect 110 1910 510 1950
rect 110 1590 150 1910
rect 470 1590 510 1910
rect 110 1550 510 1590
rect 1232 1910 1632 1950
rect 1232 1590 1272 1910
rect 1592 1590 1632 1910
rect 1232 1550 1632 1590
rect 2354 1910 2754 1950
rect 2354 1590 2394 1910
rect 2714 1590 2754 1910
rect 2354 1550 2754 1590
rect 3476 1910 3876 1950
rect 3476 1590 3516 1910
rect 3836 1590 3876 1910
rect 3476 1550 3876 1590
rect 4598 1910 4998 1950
rect 4598 1590 4638 1910
rect 4958 1590 4998 1910
rect 4598 1550 4998 1590
rect -5500 1210 -5100 1250
rect -5500 890 -5460 1210
rect -5140 890 -5100 1210
rect -5500 850 -5100 890
rect -4378 1210 -3978 1250
rect -4378 890 -4338 1210
rect -4018 890 -3978 1210
rect -4378 850 -3978 890
rect -3256 1210 -2856 1250
rect -3256 890 -3216 1210
rect -2896 890 -2856 1210
rect -3256 850 -2856 890
rect -2134 1210 -1734 1250
rect -2134 890 -2094 1210
rect -1774 890 -1734 1210
rect -2134 850 -1734 890
rect -1012 1210 -612 1250
rect -1012 890 -972 1210
rect -652 890 -612 1210
rect -1012 850 -612 890
rect 110 1210 510 1250
rect 110 890 150 1210
rect 470 890 510 1210
rect 110 850 510 890
rect 1232 1210 1632 1250
rect 1232 890 1272 1210
rect 1592 890 1632 1210
rect 1232 850 1632 890
rect 2354 1210 2754 1250
rect 2354 890 2394 1210
rect 2714 890 2754 1210
rect 2354 850 2754 890
rect 3476 1210 3876 1250
rect 3476 890 3516 1210
rect 3836 890 3876 1210
rect 3476 850 3876 890
rect 4598 1210 4998 1250
rect 4598 890 4638 1210
rect 4958 890 4998 1210
rect 4598 850 4998 890
rect -5500 510 -5100 550
rect -5500 190 -5460 510
rect -5140 190 -5100 510
rect -5500 150 -5100 190
rect -4378 510 -3978 550
rect -4378 190 -4338 510
rect -4018 190 -3978 510
rect -4378 150 -3978 190
rect -3256 510 -2856 550
rect -3256 190 -3216 510
rect -2896 190 -2856 510
rect -3256 150 -2856 190
rect -2134 510 -1734 550
rect -2134 190 -2094 510
rect -1774 190 -1734 510
rect -2134 150 -1734 190
rect -1012 510 -612 550
rect -1012 190 -972 510
rect -652 190 -612 510
rect -1012 150 -612 190
rect 110 510 510 550
rect 110 190 150 510
rect 470 190 510 510
rect 110 150 510 190
rect 1232 510 1632 550
rect 1232 190 1272 510
rect 1592 190 1632 510
rect 1232 150 1632 190
rect 2354 510 2754 550
rect 2354 190 2394 510
rect 2714 190 2754 510
rect 2354 150 2754 190
rect 3476 510 3876 550
rect 3476 190 3516 510
rect 3836 190 3876 510
rect 3476 150 3876 190
rect 4598 510 4998 550
rect 4598 190 4638 510
rect 4958 190 4998 510
rect 4598 150 4998 190
rect -5500 -190 -5100 -150
rect -5500 -510 -5460 -190
rect -5140 -510 -5100 -190
rect -5500 -550 -5100 -510
rect -4378 -190 -3978 -150
rect -4378 -510 -4338 -190
rect -4018 -510 -3978 -190
rect -4378 -550 -3978 -510
rect -3256 -190 -2856 -150
rect -3256 -510 -3216 -190
rect -2896 -510 -2856 -190
rect -3256 -550 -2856 -510
rect -2134 -190 -1734 -150
rect -2134 -510 -2094 -190
rect -1774 -510 -1734 -190
rect -2134 -550 -1734 -510
rect -1012 -190 -612 -150
rect -1012 -510 -972 -190
rect -652 -510 -612 -190
rect -1012 -550 -612 -510
rect 110 -190 510 -150
rect 110 -510 150 -190
rect 470 -510 510 -190
rect 110 -550 510 -510
rect 1232 -190 1632 -150
rect 1232 -510 1272 -190
rect 1592 -510 1632 -190
rect 1232 -550 1632 -510
rect 2354 -190 2754 -150
rect 2354 -510 2394 -190
rect 2714 -510 2754 -190
rect 2354 -550 2754 -510
rect 3476 -190 3876 -150
rect 3476 -510 3516 -190
rect 3836 -510 3876 -190
rect 3476 -550 3876 -510
rect 4598 -190 4998 -150
rect 4598 -510 4638 -190
rect 4958 -510 4998 -190
rect 4598 -550 4998 -510
rect -5500 -890 -5100 -850
rect -5500 -1210 -5460 -890
rect -5140 -1210 -5100 -890
rect -5500 -1250 -5100 -1210
rect -4378 -890 -3978 -850
rect -4378 -1210 -4338 -890
rect -4018 -1210 -3978 -890
rect -4378 -1250 -3978 -1210
rect -3256 -890 -2856 -850
rect -3256 -1210 -3216 -890
rect -2896 -1210 -2856 -890
rect -3256 -1250 -2856 -1210
rect -2134 -890 -1734 -850
rect -2134 -1210 -2094 -890
rect -1774 -1210 -1734 -890
rect -2134 -1250 -1734 -1210
rect -1012 -890 -612 -850
rect -1012 -1210 -972 -890
rect -652 -1210 -612 -890
rect -1012 -1250 -612 -1210
rect 110 -890 510 -850
rect 110 -1210 150 -890
rect 470 -1210 510 -890
rect 110 -1250 510 -1210
rect 1232 -890 1632 -850
rect 1232 -1210 1272 -890
rect 1592 -1210 1632 -890
rect 1232 -1250 1632 -1210
rect 2354 -890 2754 -850
rect 2354 -1210 2394 -890
rect 2714 -1210 2754 -890
rect 2354 -1250 2754 -1210
rect 3476 -890 3876 -850
rect 3476 -1210 3516 -890
rect 3836 -1210 3876 -890
rect 3476 -1250 3876 -1210
rect 4598 -890 4998 -850
rect 4598 -1210 4638 -890
rect 4958 -1210 4998 -890
rect 4598 -1250 4998 -1210
rect -5500 -1590 -5100 -1550
rect -5500 -1910 -5460 -1590
rect -5140 -1910 -5100 -1590
rect -5500 -1950 -5100 -1910
rect -4378 -1590 -3978 -1550
rect -4378 -1910 -4338 -1590
rect -4018 -1910 -3978 -1590
rect -4378 -1950 -3978 -1910
rect -3256 -1590 -2856 -1550
rect -3256 -1910 -3216 -1590
rect -2896 -1910 -2856 -1590
rect -3256 -1950 -2856 -1910
rect -2134 -1590 -1734 -1550
rect -2134 -1910 -2094 -1590
rect -1774 -1910 -1734 -1590
rect -2134 -1950 -1734 -1910
rect -1012 -1590 -612 -1550
rect -1012 -1910 -972 -1590
rect -652 -1910 -612 -1590
rect -1012 -1950 -612 -1910
rect 110 -1590 510 -1550
rect 110 -1910 150 -1590
rect 470 -1910 510 -1590
rect 110 -1950 510 -1910
rect 1232 -1590 1632 -1550
rect 1232 -1910 1272 -1590
rect 1592 -1910 1632 -1590
rect 1232 -1950 1632 -1910
rect 2354 -1590 2754 -1550
rect 2354 -1910 2394 -1590
rect 2714 -1910 2754 -1590
rect 2354 -1950 2754 -1910
rect 3476 -1590 3876 -1550
rect 3476 -1910 3516 -1590
rect 3836 -1910 3876 -1590
rect 3476 -1950 3876 -1910
rect 4598 -1590 4998 -1550
rect 4598 -1910 4638 -1590
rect 4958 -1910 4998 -1590
rect 4598 -1950 4998 -1910
rect -5500 -2290 -5100 -2250
rect -5500 -2610 -5460 -2290
rect -5140 -2610 -5100 -2290
rect -5500 -2650 -5100 -2610
rect -4378 -2290 -3978 -2250
rect -4378 -2610 -4338 -2290
rect -4018 -2610 -3978 -2290
rect -4378 -2650 -3978 -2610
rect -3256 -2290 -2856 -2250
rect -3256 -2610 -3216 -2290
rect -2896 -2610 -2856 -2290
rect -3256 -2650 -2856 -2610
rect -2134 -2290 -1734 -2250
rect -2134 -2610 -2094 -2290
rect -1774 -2610 -1734 -2290
rect -2134 -2650 -1734 -2610
rect -1012 -2290 -612 -2250
rect -1012 -2610 -972 -2290
rect -652 -2610 -612 -2290
rect -1012 -2650 -612 -2610
rect 110 -2290 510 -2250
rect 110 -2610 150 -2290
rect 470 -2610 510 -2290
rect 110 -2650 510 -2610
rect 1232 -2290 1632 -2250
rect 1232 -2610 1272 -2290
rect 1592 -2610 1632 -2290
rect 1232 -2650 1632 -2610
rect 2354 -2290 2754 -2250
rect 2354 -2610 2394 -2290
rect 2714 -2610 2754 -2290
rect 2354 -2650 2754 -2610
rect 3476 -2290 3876 -2250
rect 3476 -2610 3516 -2290
rect 3836 -2610 3876 -2290
rect 3476 -2650 3876 -2610
rect 4598 -2290 4998 -2250
rect 4598 -2610 4638 -2290
rect 4958 -2610 4998 -2290
rect 4598 -2650 4998 -2610
rect -5500 -2990 -5100 -2950
rect -5500 -3310 -5460 -2990
rect -5140 -3310 -5100 -2990
rect -5500 -3350 -5100 -3310
rect -4378 -2990 -3978 -2950
rect -4378 -3310 -4338 -2990
rect -4018 -3310 -3978 -2990
rect -4378 -3350 -3978 -3310
rect -3256 -2990 -2856 -2950
rect -3256 -3310 -3216 -2990
rect -2896 -3310 -2856 -2990
rect -3256 -3350 -2856 -3310
rect -2134 -2990 -1734 -2950
rect -2134 -3310 -2094 -2990
rect -1774 -3310 -1734 -2990
rect -2134 -3350 -1734 -3310
rect -1012 -2990 -612 -2950
rect -1012 -3310 -972 -2990
rect -652 -3310 -612 -2990
rect -1012 -3350 -612 -3310
rect 110 -2990 510 -2950
rect 110 -3310 150 -2990
rect 470 -3310 510 -2990
rect 110 -3350 510 -3310
rect 1232 -2990 1632 -2950
rect 1232 -3310 1272 -2990
rect 1592 -3310 1632 -2990
rect 1232 -3350 1632 -3310
rect 2354 -2990 2754 -2950
rect 2354 -3310 2394 -2990
rect 2714 -3310 2754 -2990
rect 2354 -3350 2754 -3310
rect 3476 -2990 3876 -2950
rect 3476 -3310 3516 -2990
rect 3836 -3310 3876 -2990
rect 3476 -3350 3876 -3310
rect 4598 -2990 4998 -2950
rect 4598 -3310 4638 -2990
rect 4958 -3310 4998 -2990
rect 4598 -3350 4998 -3310
<< mimcap2contact >>
rect -5460 2990 -5140 3310
rect -4338 2990 -4018 3310
rect -3216 2990 -2896 3310
rect -2094 2990 -1774 3310
rect -972 2990 -652 3310
rect 150 2990 470 3310
rect 1272 2990 1592 3310
rect 2394 2990 2714 3310
rect 3516 2990 3836 3310
rect 4638 2990 4958 3310
rect -5460 2290 -5140 2610
rect -4338 2290 -4018 2610
rect -3216 2290 -2896 2610
rect -2094 2290 -1774 2610
rect -972 2290 -652 2610
rect 150 2290 470 2610
rect 1272 2290 1592 2610
rect 2394 2290 2714 2610
rect 3516 2290 3836 2610
rect 4638 2290 4958 2610
rect -5460 1590 -5140 1910
rect -4338 1590 -4018 1910
rect -3216 1590 -2896 1910
rect -2094 1590 -1774 1910
rect -972 1590 -652 1910
rect 150 1590 470 1910
rect 1272 1590 1592 1910
rect 2394 1590 2714 1910
rect 3516 1590 3836 1910
rect 4638 1590 4958 1910
rect -5460 890 -5140 1210
rect -4338 890 -4018 1210
rect -3216 890 -2896 1210
rect -2094 890 -1774 1210
rect -972 890 -652 1210
rect 150 890 470 1210
rect 1272 890 1592 1210
rect 2394 890 2714 1210
rect 3516 890 3836 1210
rect 4638 890 4958 1210
rect -5460 190 -5140 510
rect -4338 190 -4018 510
rect -3216 190 -2896 510
rect -2094 190 -1774 510
rect -972 190 -652 510
rect 150 190 470 510
rect 1272 190 1592 510
rect 2394 190 2714 510
rect 3516 190 3836 510
rect 4638 190 4958 510
rect -5460 -510 -5140 -190
rect -4338 -510 -4018 -190
rect -3216 -510 -2896 -190
rect -2094 -510 -1774 -190
rect -972 -510 -652 -190
rect 150 -510 470 -190
rect 1272 -510 1592 -190
rect 2394 -510 2714 -190
rect 3516 -510 3836 -190
rect 4638 -510 4958 -190
rect -5460 -1210 -5140 -890
rect -4338 -1210 -4018 -890
rect -3216 -1210 -2896 -890
rect -2094 -1210 -1774 -890
rect -972 -1210 -652 -890
rect 150 -1210 470 -890
rect 1272 -1210 1592 -890
rect 2394 -1210 2714 -890
rect 3516 -1210 3836 -890
rect 4638 -1210 4958 -890
rect -5460 -1910 -5140 -1590
rect -4338 -1910 -4018 -1590
rect -3216 -1910 -2896 -1590
rect -2094 -1910 -1774 -1590
rect -972 -1910 -652 -1590
rect 150 -1910 470 -1590
rect 1272 -1910 1592 -1590
rect 2394 -1910 2714 -1590
rect 3516 -1910 3836 -1590
rect 4638 -1910 4958 -1590
rect -5460 -2610 -5140 -2290
rect -4338 -2610 -4018 -2290
rect -3216 -2610 -2896 -2290
rect -2094 -2610 -1774 -2290
rect -972 -2610 -652 -2290
rect 150 -2610 470 -2290
rect 1272 -2610 1592 -2290
rect 2394 -2610 2714 -2290
rect 3516 -2610 3836 -2290
rect 4638 -2610 4958 -2290
rect -5460 -3310 -5140 -2990
rect -4338 -3310 -4018 -2990
rect -3216 -3310 -2896 -2990
rect -2094 -3310 -1774 -2990
rect -972 -3310 -652 -2990
rect 150 -3310 470 -2990
rect 1272 -3310 1592 -2990
rect 2394 -3310 2714 -2990
rect 3516 -3310 3836 -2990
rect 4638 -3310 4958 -2990
<< metal5 >>
rect -5140 3334 -4820 3500
rect -5484 3310 -4820 3334
rect -5484 2990 -5460 3310
rect -5140 2990 -4820 3310
rect -5484 2966 -4820 2990
rect -5140 2634 -4820 2966
rect -4796 3409 -4476 3451
rect -4796 2891 -4754 3409
rect -4518 2891 -4476 3409
rect -4018 3334 -3698 3500
rect -4362 3310 -3698 3334
rect -4362 2990 -4338 3310
rect -4018 2990 -3698 3310
rect -4362 2966 -3698 2990
rect -4796 2849 -4476 2891
rect -5484 2610 -4820 2634
rect -5484 2290 -5460 2610
rect -5140 2290 -4820 2610
rect -5484 2266 -4820 2290
rect -5140 1934 -4820 2266
rect -4796 2709 -4476 2751
rect -4796 2191 -4754 2709
rect -4518 2191 -4476 2709
rect -4018 2634 -3698 2966
rect -3674 3409 -3354 3451
rect -3674 2891 -3632 3409
rect -3396 2891 -3354 3409
rect -2896 3334 -2576 3500
rect -3240 3310 -2576 3334
rect -3240 2990 -3216 3310
rect -2896 2990 -2576 3310
rect -3240 2966 -2576 2990
rect -3674 2849 -3354 2891
rect -4362 2610 -3698 2634
rect -4362 2290 -4338 2610
rect -4018 2290 -3698 2610
rect -4362 2266 -3698 2290
rect -4796 2149 -4476 2191
rect -5484 1910 -4820 1934
rect -5484 1590 -5460 1910
rect -5140 1590 -4820 1910
rect -5484 1566 -4820 1590
rect -5140 1234 -4820 1566
rect -4796 2009 -4476 2051
rect -4796 1491 -4754 2009
rect -4518 1491 -4476 2009
rect -4018 1934 -3698 2266
rect -3674 2709 -3354 2751
rect -3674 2191 -3632 2709
rect -3396 2191 -3354 2709
rect -2896 2634 -2576 2966
rect -2552 3409 -2232 3451
rect -2552 2891 -2510 3409
rect -2274 2891 -2232 3409
rect -1774 3334 -1454 3500
rect -2118 3310 -1454 3334
rect -2118 2990 -2094 3310
rect -1774 2990 -1454 3310
rect -2118 2966 -1454 2990
rect -2552 2849 -2232 2891
rect -3240 2610 -2576 2634
rect -3240 2290 -3216 2610
rect -2896 2290 -2576 2610
rect -3240 2266 -2576 2290
rect -3674 2149 -3354 2191
rect -4362 1910 -3698 1934
rect -4362 1590 -4338 1910
rect -4018 1590 -3698 1910
rect -4362 1566 -3698 1590
rect -4796 1449 -4476 1491
rect -5484 1210 -4820 1234
rect -5484 890 -5460 1210
rect -5140 890 -4820 1210
rect -5484 866 -4820 890
rect -5140 534 -4820 866
rect -4796 1309 -4476 1351
rect -4796 791 -4754 1309
rect -4518 791 -4476 1309
rect -4018 1234 -3698 1566
rect -3674 2009 -3354 2051
rect -3674 1491 -3632 2009
rect -3396 1491 -3354 2009
rect -2896 1934 -2576 2266
rect -2552 2709 -2232 2751
rect -2552 2191 -2510 2709
rect -2274 2191 -2232 2709
rect -1774 2634 -1454 2966
rect -1430 3409 -1110 3451
rect -1430 2891 -1388 3409
rect -1152 2891 -1110 3409
rect -652 3334 -332 3500
rect -996 3310 -332 3334
rect -996 2990 -972 3310
rect -652 2990 -332 3310
rect -996 2966 -332 2990
rect -1430 2849 -1110 2891
rect -2118 2610 -1454 2634
rect -2118 2290 -2094 2610
rect -1774 2290 -1454 2610
rect -2118 2266 -1454 2290
rect -2552 2149 -2232 2191
rect -3240 1910 -2576 1934
rect -3240 1590 -3216 1910
rect -2896 1590 -2576 1910
rect -3240 1566 -2576 1590
rect -3674 1449 -3354 1491
rect -4362 1210 -3698 1234
rect -4362 890 -4338 1210
rect -4018 890 -3698 1210
rect -4362 866 -3698 890
rect -4796 749 -4476 791
rect -5484 510 -4820 534
rect -5484 190 -5460 510
rect -5140 190 -4820 510
rect -5484 166 -4820 190
rect -5140 -166 -4820 166
rect -4796 609 -4476 651
rect -4796 91 -4754 609
rect -4518 91 -4476 609
rect -4018 534 -3698 866
rect -3674 1309 -3354 1351
rect -3674 791 -3632 1309
rect -3396 791 -3354 1309
rect -2896 1234 -2576 1566
rect -2552 2009 -2232 2051
rect -2552 1491 -2510 2009
rect -2274 1491 -2232 2009
rect -1774 1934 -1454 2266
rect -1430 2709 -1110 2751
rect -1430 2191 -1388 2709
rect -1152 2191 -1110 2709
rect -652 2634 -332 2966
rect -308 3409 12 3451
rect -308 2891 -266 3409
rect -30 2891 12 3409
rect 470 3334 790 3500
rect 126 3310 790 3334
rect 126 2990 150 3310
rect 470 2990 790 3310
rect 126 2966 790 2990
rect -308 2849 12 2891
rect -996 2610 -332 2634
rect -996 2290 -972 2610
rect -652 2290 -332 2610
rect -996 2266 -332 2290
rect -1430 2149 -1110 2191
rect -2118 1910 -1454 1934
rect -2118 1590 -2094 1910
rect -1774 1590 -1454 1910
rect -2118 1566 -1454 1590
rect -2552 1449 -2232 1491
rect -3240 1210 -2576 1234
rect -3240 890 -3216 1210
rect -2896 890 -2576 1210
rect -3240 866 -2576 890
rect -3674 749 -3354 791
rect -4362 510 -3698 534
rect -4362 190 -4338 510
rect -4018 190 -3698 510
rect -4362 166 -3698 190
rect -4796 49 -4476 91
rect -5484 -190 -4820 -166
rect -5484 -510 -5460 -190
rect -5140 -510 -4820 -190
rect -5484 -534 -4820 -510
rect -5140 -866 -4820 -534
rect -4796 -91 -4476 -49
rect -4796 -609 -4754 -91
rect -4518 -609 -4476 -91
rect -4018 -166 -3698 166
rect -3674 609 -3354 651
rect -3674 91 -3632 609
rect -3396 91 -3354 609
rect -2896 534 -2576 866
rect -2552 1309 -2232 1351
rect -2552 791 -2510 1309
rect -2274 791 -2232 1309
rect -1774 1234 -1454 1566
rect -1430 2009 -1110 2051
rect -1430 1491 -1388 2009
rect -1152 1491 -1110 2009
rect -652 1934 -332 2266
rect -308 2709 12 2751
rect -308 2191 -266 2709
rect -30 2191 12 2709
rect 470 2634 790 2966
rect 814 3409 1134 3451
rect 814 2891 856 3409
rect 1092 2891 1134 3409
rect 1592 3334 1912 3500
rect 1248 3310 1912 3334
rect 1248 2990 1272 3310
rect 1592 2990 1912 3310
rect 1248 2966 1912 2990
rect 814 2849 1134 2891
rect 126 2610 790 2634
rect 126 2290 150 2610
rect 470 2290 790 2610
rect 126 2266 790 2290
rect -308 2149 12 2191
rect -996 1910 -332 1934
rect -996 1590 -972 1910
rect -652 1590 -332 1910
rect -996 1566 -332 1590
rect -1430 1449 -1110 1491
rect -2118 1210 -1454 1234
rect -2118 890 -2094 1210
rect -1774 890 -1454 1210
rect -2118 866 -1454 890
rect -2552 749 -2232 791
rect -3240 510 -2576 534
rect -3240 190 -3216 510
rect -2896 190 -2576 510
rect -3240 166 -2576 190
rect -3674 49 -3354 91
rect -4362 -190 -3698 -166
rect -4362 -510 -4338 -190
rect -4018 -510 -3698 -190
rect -4362 -534 -3698 -510
rect -4796 -651 -4476 -609
rect -5484 -890 -4820 -866
rect -5484 -1210 -5460 -890
rect -5140 -1210 -4820 -890
rect -5484 -1234 -4820 -1210
rect -5140 -1566 -4820 -1234
rect -4796 -791 -4476 -749
rect -4796 -1309 -4754 -791
rect -4518 -1309 -4476 -791
rect -4018 -866 -3698 -534
rect -3674 -91 -3354 -49
rect -3674 -609 -3632 -91
rect -3396 -609 -3354 -91
rect -2896 -166 -2576 166
rect -2552 609 -2232 651
rect -2552 91 -2510 609
rect -2274 91 -2232 609
rect -1774 534 -1454 866
rect -1430 1309 -1110 1351
rect -1430 791 -1388 1309
rect -1152 791 -1110 1309
rect -652 1234 -332 1566
rect -308 2009 12 2051
rect -308 1491 -266 2009
rect -30 1491 12 2009
rect 470 1934 790 2266
rect 814 2709 1134 2751
rect 814 2191 856 2709
rect 1092 2191 1134 2709
rect 1592 2634 1912 2966
rect 1936 3409 2256 3451
rect 1936 2891 1978 3409
rect 2214 2891 2256 3409
rect 2714 3334 3034 3500
rect 2370 3310 3034 3334
rect 2370 2990 2394 3310
rect 2714 2990 3034 3310
rect 2370 2966 3034 2990
rect 1936 2849 2256 2891
rect 1248 2610 1912 2634
rect 1248 2290 1272 2610
rect 1592 2290 1912 2610
rect 1248 2266 1912 2290
rect 814 2149 1134 2191
rect 126 1910 790 1934
rect 126 1590 150 1910
rect 470 1590 790 1910
rect 126 1566 790 1590
rect -308 1449 12 1491
rect -996 1210 -332 1234
rect -996 890 -972 1210
rect -652 890 -332 1210
rect -996 866 -332 890
rect -1430 749 -1110 791
rect -2118 510 -1454 534
rect -2118 190 -2094 510
rect -1774 190 -1454 510
rect -2118 166 -1454 190
rect -2552 49 -2232 91
rect -3240 -190 -2576 -166
rect -3240 -510 -3216 -190
rect -2896 -510 -2576 -190
rect -3240 -534 -2576 -510
rect -3674 -651 -3354 -609
rect -4362 -890 -3698 -866
rect -4362 -1210 -4338 -890
rect -4018 -1210 -3698 -890
rect -4362 -1234 -3698 -1210
rect -4796 -1351 -4476 -1309
rect -5484 -1590 -4820 -1566
rect -5484 -1910 -5460 -1590
rect -5140 -1910 -4820 -1590
rect -5484 -1934 -4820 -1910
rect -5140 -2266 -4820 -1934
rect -4796 -1491 -4476 -1449
rect -4796 -2009 -4754 -1491
rect -4518 -2009 -4476 -1491
rect -4018 -1566 -3698 -1234
rect -3674 -791 -3354 -749
rect -3674 -1309 -3632 -791
rect -3396 -1309 -3354 -791
rect -2896 -866 -2576 -534
rect -2552 -91 -2232 -49
rect -2552 -609 -2510 -91
rect -2274 -609 -2232 -91
rect -1774 -166 -1454 166
rect -1430 609 -1110 651
rect -1430 91 -1388 609
rect -1152 91 -1110 609
rect -652 534 -332 866
rect -308 1309 12 1351
rect -308 791 -266 1309
rect -30 791 12 1309
rect 470 1234 790 1566
rect 814 2009 1134 2051
rect 814 1491 856 2009
rect 1092 1491 1134 2009
rect 1592 1934 1912 2266
rect 1936 2709 2256 2751
rect 1936 2191 1978 2709
rect 2214 2191 2256 2709
rect 2714 2634 3034 2966
rect 3058 3409 3378 3451
rect 3058 2891 3100 3409
rect 3336 2891 3378 3409
rect 3836 3334 4156 3500
rect 3492 3310 4156 3334
rect 3492 2990 3516 3310
rect 3836 2990 4156 3310
rect 3492 2966 4156 2990
rect 3058 2849 3378 2891
rect 2370 2610 3034 2634
rect 2370 2290 2394 2610
rect 2714 2290 3034 2610
rect 2370 2266 3034 2290
rect 1936 2149 2256 2191
rect 1248 1910 1912 1934
rect 1248 1590 1272 1910
rect 1592 1590 1912 1910
rect 1248 1566 1912 1590
rect 814 1449 1134 1491
rect 126 1210 790 1234
rect 126 890 150 1210
rect 470 890 790 1210
rect 126 866 790 890
rect -308 749 12 791
rect -996 510 -332 534
rect -996 190 -972 510
rect -652 190 -332 510
rect -996 166 -332 190
rect -1430 49 -1110 91
rect -2118 -190 -1454 -166
rect -2118 -510 -2094 -190
rect -1774 -510 -1454 -190
rect -2118 -534 -1454 -510
rect -2552 -651 -2232 -609
rect -3240 -890 -2576 -866
rect -3240 -1210 -3216 -890
rect -2896 -1210 -2576 -890
rect -3240 -1234 -2576 -1210
rect -3674 -1351 -3354 -1309
rect -4362 -1590 -3698 -1566
rect -4362 -1910 -4338 -1590
rect -4018 -1910 -3698 -1590
rect -4362 -1934 -3698 -1910
rect -4796 -2051 -4476 -2009
rect -5484 -2290 -4820 -2266
rect -5484 -2610 -5460 -2290
rect -5140 -2610 -4820 -2290
rect -5484 -2634 -4820 -2610
rect -5140 -2966 -4820 -2634
rect -4796 -2191 -4476 -2149
rect -4796 -2709 -4754 -2191
rect -4518 -2709 -4476 -2191
rect -4018 -2266 -3698 -1934
rect -3674 -1491 -3354 -1449
rect -3674 -2009 -3632 -1491
rect -3396 -2009 -3354 -1491
rect -2896 -1566 -2576 -1234
rect -2552 -791 -2232 -749
rect -2552 -1309 -2510 -791
rect -2274 -1309 -2232 -791
rect -1774 -866 -1454 -534
rect -1430 -91 -1110 -49
rect -1430 -609 -1388 -91
rect -1152 -609 -1110 -91
rect -652 -166 -332 166
rect -308 609 12 651
rect -308 91 -266 609
rect -30 91 12 609
rect 470 534 790 866
rect 814 1309 1134 1351
rect 814 791 856 1309
rect 1092 791 1134 1309
rect 1592 1234 1912 1566
rect 1936 2009 2256 2051
rect 1936 1491 1978 2009
rect 2214 1491 2256 2009
rect 2714 1934 3034 2266
rect 3058 2709 3378 2751
rect 3058 2191 3100 2709
rect 3336 2191 3378 2709
rect 3836 2634 4156 2966
rect 4180 3409 4500 3451
rect 4180 2891 4222 3409
rect 4458 2891 4500 3409
rect 4958 3334 5278 3500
rect 4614 3310 5278 3334
rect 4614 2990 4638 3310
rect 4958 2990 5278 3310
rect 4614 2966 5278 2990
rect 4180 2849 4500 2891
rect 3492 2610 4156 2634
rect 3492 2290 3516 2610
rect 3836 2290 4156 2610
rect 3492 2266 4156 2290
rect 3058 2149 3378 2191
rect 2370 1910 3034 1934
rect 2370 1590 2394 1910
rect 2714 1590 3034 1910
rect 2370 1566 3034 1590
rect 1936 1449 2256 1491
rect 1248 1210 1912 1234
rect 1248 890 1272 1210
rect 1592 890 1912 1210
rect 1248 866 1912 890
rect 814 749 1134 791
rect 126 510 790 534
rect 126 190 150 510
rect 470 190 790 510
rect 126 166 790 190
rect -308 49 12 91
rect -996 -190 -332 -166
rect -996 -510 -972 -190
rect -652 -510 -332 -190
rect -996 -534 -332 -510
rect -1430 -651 -1110 -609
rect -2118 -890 -1454 -866
rect -2118 -1210 -2094 -890
rect -1774 -1210 -1454 -890
rect -2118 -1234 -1454 -1210
rect -2552 -1351 -2232 -1309
rect -3240 -1590 -2576 -1566
rect -3240 -1910 -3216 -1590
rect -2896 -1910 -2576 -1590
rect -3240 -1934 -2576 -1910
rect -3674 -2051 -3354 -2009
rect -4362 -2290 -3698 -2266
rect -4362 -2610 -4338 -2290
rect -4018 -2610 -3698 -2290
rect -4362 -2634 -3698 -2610
rect -4796 -2751 -4476 -2709
rect -5484 -2990 -4820 -2966
rect -5484 -3310 -5460 -2990
rect -5140 -3310 -4820 -2990
rect -5484 -3334 -4820 -3310
rect -5140 -3500 -4820 -3334
rect -4796 -2891 -4476 -2849
rect -4796 -3409 -4754 -2891
rect -4518 -3409 -4476 -2891
rect -4018 -2966 -3698 -2634
rect -3674 -2191 -3354 -2149
rect -3674 -2709 -3632 -2191
rect -3396 -2709 -3354 -2191
rect -2896 -2266 -2576 -1934
rect -2552 -1491 -2232 -1449
rect -2552 -2009 -2510 -1491
rect -2274 -2009 -2232 -1491
rect -1774 -1566 -1454 -1234
rect -1430 -791 -1110 -749
rect -1430 -1309 -1388 -791
rect -1152 -1309 -1110 -791
rect -652 -866 -332 -534
rect -308 -91 12 -49
rect -308 -609 -266 -91
rect -30 -609 12 -91
rect 470 -166 790 166
rect 814 609 1134 651
rect 814 91 856 609
rect 1092 91 1134 609
rect 1592 534 1912 866
rect 1936 1309 2256 1351
rect 1936 791 1978 1309
rect 2214 791 2256 1309
rect 2714 1234 3034 1566
rect 3058 2009 3378 2051
rect 3058 1491 3100 2009
rect 3336 1491 3378 2009
rect 3836 1934 4156 2266
rect 4180 2709 4500 2751
rect 4180 2191 4222 2709
rect 4458 2191 4500 2709
rect 4958 2634 5278 2966
rect 5302 3409 5622 3451
rect 5302 2891 5344 3409
rect 5580 2891 5622 3409
rect 5302 2849 5622 2891
rect 4614 2610 5278 2634
rect 4614 2290 4638 2610
rect 4958 2290 5278 2610
rect 4614 2266 5278 2290
rect 4180 2149 4500 2191
rect 3492 1910 4156 1934
rect 3492 1590 3516 1910
rect 3836 1590 4156 1910
rect 3492 1566 4156 1590
rect 3058 1449 3378 1491
rect 2370 1210 3034 1234
rect 2370 890 2394 1210
rect 2714 890 3034 1210
rect 2370 866 3034 890
rect 1936 749 2256 791
rect 1248 510 1912 534
rect 1248 190 1272 510
rect 1592 190 1912 510
rect 1248 166 1912 190
rect 814 49 1134 91
rect 126 -190 790 -166
rect 126 -510 150 -190
rect 470 -510 790 -190
rect 126 -534 790 -510
rect -308 -651 12 -609
rect -996 -890 -332 -866
rect -996 -1210 -972 -890
rect -652 -1210 -332 -890
rect -996 -1234 -332 -1210
rect -1430 -1351 -1110 -1309
rect -2118 -1590 -1454 -1566
rect -2118 -1910 -2094 -1590
rect -1774 -1910 -1454 -1590
rect -2118 -1934 -1454 -1910
rect -2552 -2051 -2232 -2009
rect -3240 -2290 -2576 -2266
rect -3240 -2610 -3216 -2290
rect -2896 -2610 -2576 -2290
rect -3240 -2634 -2576 -2610
rect -3674 -2751 -3354 -2709
rect -4362 -2990 -3698 -2966
rect -4362 -3310 -4338 -2990
rect -4018 -3310 -3698 -2990
rect -4362 -3334 -3698 -3310
rect -4796 -3451 -4476 -3409
rect -4018 -3500 -3698 -3334
rect -3674 -2891 -3354 -2849
rect -3674 -3409 -3632 -2891
rect -3396 -3409 -3354 -2891
rect -2896 -2966 -2576 -2634
rect -2552 -2191 -2232 -2149
rect -2552 -2709 -2510 -2191
rect -2274 -2709 -2232 -2191
rect -1774 -2266 -1454 -1934
rect -1430 -1491 -1110 -1449
rect -1430 -2009 -1388 -1491
rect -1152 -2009 -1110 -1491
rect -652 -1566 -332 -1234
rect -308 -791 12 -749
rect -308 -1309 -266 -791
rect -30 -1309 12 -791
rect 470 -866 790 -534
rect 814 -91 1134 -49
rect 814 -609 856 -91
rect 1092 -609 1134 -91
rect 1592 -166 1912 166
rect 1936 609 2256 651
rect 1936 91 1978 609
rect 2214 91 2256 609
rect 2714 534 3034 866
rect 3058 1309 3378 1351
rect 3058 791 3100 1309
rect 3336 791 3378 1309
rect 3836 1234 4156 1566
rect 4180 2009 4500 2051
rect 4180 1491 4222 2009
rect 4458 1491 4500 2009
rect 4958 1934 5278 2266
rect 5302 2709 5622 2751
rect 5302 2191 5344 2709
rect 5580 2191 5622 2709
rect 5302 2149 5622 2191
rect 4614 1910 5278 1934
rect 4614 1590 4638 1910
rect 4958 1590 5278 1910
rect 4614 1566 5278 1590
rect 4180 1449 4500 1491
rect 3492 1210 4156 1234
rect 3492 890 3516 1210
rect 3836 890 4156 1210
rect 3492 866 4156 890
rect 3058 749 3378 791
rect 2370 510 3034 534
rect 2370 190 2394 510
rect 2714 190 3034 510
rect 2370 166 3034 190
rect 1936 49 2256 91
rect 1248 -190 1912 -166
rect 1248 -510 1272 -190
rect 1592 -510 1912 -190
rect 1248 -534 1912 -510
rect 814 -651 1134 -609
rect 126 -890 790 -866
rect 126 -1210 150 -890
rect 470 -1210 790 -890
rect 126 -1234 790 -1210
rect -308 -1351 12 -1309
rect -996 -1590 -332 -1566
rect -996 -1910 -972 -1590
rect -652 -1910 -332 -1590
rect -996 -1934 -332 -1910
rect -1430 -2051 -1110 -2009
rect -2118 -2290 -1454 -2266
rect -2118 -2610 -2094 -2290
rect -1774 -2610 -1454 -2290
rect -2118 -2634 -1454 -2610
rect -2552 -2751 -2232 -2709
rect -3240 -2990 -2576 -2966
rect -3240 -3310 -3216 -2990
rect -2896 -3310 -2576 -2990
rect -3240 -3334 -2576 -3310
rect -3674 -3451 -3354 -3409
rect -2896 -3500 -2576 -3334
rect -2552 -2891 -2232 -2849
rect -2552 -3409 -2510 -2891
rect -2274 -3409 -2232 -2891
rect -1774 -2966 -1454 -2634
rect -1430 -2191 -1110 -2149
rect -1430 -2709 -1388 -2191
rect -1152 -2709 -1110 -2191
rect -652 -2266 -332 -1934
rect -308 -1491 12 -1449
rect -308 -2009 -266 -1491
rect -30 -2009 12 -1491
rect 470 -1566 790 -1234
rect 814 -791 1134 -749
rect 814 -1309 856 -791
rect 1092 -1309 1134 -791
rect 1592 -866 1912 -534
rect 1936 -91 2256 -49
rect 1936 -609 1978 -91
rect 2214 -609 2256 -91
rect 2714 -166 3034 166
rect 3058 609 3378 651
rect 3058 91 3100 609
rect 3336 91 3378 609
rect 3836 534 4156 866
rect 4180 1309 4500 1351
rect 4180 791 4222 1309
rect 4458 791 4500 1309
rect 4958 1234 5278 1566
rect 5302 2009 5622 2051
rect 5302 1491 5344 2009
rect 5580 1491 5622 2009
rect 5302 1449 5622 1491
rect 4614 1210 5278 1234
rect 4614 890 4638 1210
rect 4958 890 5278 1210
rect 4614 866 5278 890
rect 4180 749 4500 791
rect 3492 510 4156 534
rect 3492 190 3516 510
rect 3836 190 4156 510
rect 3492 166 4156 190
rect 3058 49 3378 91
rect 2370 -190 3034 -166
rect 2370 -510 2394 -190
rect 2714 -510 3034 -190
rect 2370 -534 3034 -510
rect 1936 -651 2256 -609
rect 1248 -890 1912 -866
rect 1248 -1210 1272 -890
rect 1592 -1210 1912 -890
rect 1248 -1234 1912 -1210
rect 814 -1351 1134 -1309
rect 126 -1590 790 -1566
rect 126 -1910 150 -1590
rect 470 -1910 790 -1590
rect 126 -1934 790 -1910
rect -308 -2051 12 -2009
rect -996 -2290 -332 -2266
rect -996 -2610 -972 -2290
rect -652 -2610 -332 -2290
rect -996 -2634 -332 -2610
rect -1430 -2751 -1110 -2709
rect -2118 -2990 -1454 -2966
rect -2118 -3310 -2094 -2990
rect -1774 -3310 -1454 -2990
rect -2118 -3334 -1454 -3310
rect -2552 -3451 -2232 -3409
rect -1774 -3500 -1454 -3334
rect -1430 -2891 -1110 -2849
rect -1430 -3409 -1388 -2891
rect -1152 -3409 -1110 -2891
rect -652 -2966 -332 -2634
rect -308 -2191 12 -2149
rect -308 -2709 -266 -2191
rect -30 -2709 12 -2191
rect 470 -2266 790 -1934
rect 814 -1491 1134 -1449
rect 814 -2009 856 -1491
rect 1092 -2009 1134 -1491
rect 1592 -1566 1912 -1234
rect 1936 -791 2256 -749
rect 1936 -1309 1978 -791
rect 2214 -1309 2256 -791
rect 2714 -866 3034 -534
rect 3058 -91 3378 -49
rect 3058 -609 3100 -91
rect 3336 -609 3378 -91
rect 3836 -166 4156 166
rect 4180 609 4500 651
rect 4180 91 4222 609
rect 4458 91 4500 609
rect 4958 534 5278 866
rect 5302 1309 5622 1351
rect 5302 791 5344 1309
rect 5580 791 5622 1309
rect 5302 749 5622 791
rect 4614 510 5278 534
rect 4614 190 4638 510
rect 4958 190 5278 510
rect 4614 166 5278 190
rect 4180 49 4500 91
rect 3492 -190 4156 -166
rect 3492 -510 3516 -190
rect 3836 -510 4156 -190
rect 3492 -534 4156 -510
rect 3058 -651 3378 -609
rect 2370 -890 3034 -866
rect 2370 -1210 2394 -890
rect 2714 -1210 3034 -890
rect 2370 -1234 3034 -1210
rect 1936 -1351 2256 -1309
rect 1248 -1590 1912 -1566
rect 1248 -1910 1272 -1590
rect 1592 -1910 1912 -1590
rect 1248 -1934 1912 -1910
rect 814 -2051 1134 -2009
rect 126 -2290 790 -2266
rect 126 -2610 150 -2290
rect 470 -2610 790 -2290
rect 126 -2634 790 -2610
rect -308 -2751 12 -2709
rect -996 -2990 -332 -2966
rect -996 -3310 -972 -2990
rect -652 -3310 -332 -2990
rect -996 -3334 -332 -3310
rect -1430 -3451 -1110 -3409
rect -652 -3500 -332 -3334
rect -308 -2891 12 -2849
rect -308 -3409 -266 -2891
rect -30 -3409 12 -2891
rect 470 -2966 790 -2634
rect 814 -2191 1134 -2149
rect 814 -2709 856 -2191
rect 1092 -2709 1134 -2191
rect 1592 -2266 1912 -1934
rect 1936 -1491 2256 -1449
rect 1936 -2009 1978 -1491
rect 2214 -2009 2256 -1491
rect 2714 -1566 3034 -1234
rect 3058 -791 3378 -749
rect 3058 -1309 3100 -791
rect 3336 -1309 3378 -791
rect 3836 -866 4156 -534
rect 4180 -91 4500 -49
rect 4180 -609 4222 -91
rect 4458 -609 4500 -91
rect 4958 -166 5278 166
rect 5302 609 5622 651
rect 5302 91 5344 609
rect 5580 91 5622 609
rect 5302 49 5622 91
rect 4614 -190 5278 -166
rect 4614 -510 4638 -190
rect 4958 -510 5278 -190
rect 4614 -534 5278 -510
rect 4180 -651 4500 -609
rect 3492 -890 4156 -866
rect 3492 -1210 3516 -890
rect 3836 -1210 4156 -890
rect 3492 -1234 4156 -1210
rect 3058 -1351 3378 -1309
rect 2370 -1590 3034 -1566
rect 2370 -1910 2394 -1590
rect 2714 -1910 3034 -1590
rect 2370 -1934 3034 -1910
rect 1936 -2051 2256 -2009
rect 1248 -2290 1912 -2266
rect 1248 -2610 1272 -2290
rect 1592 -2610 1912 -2290
rect 1248 -2634 1912 -2610
rect 814 -2751 1134 -2709
rect 126 -2990 790 -2966
rect 126 -3310 150 -2990
rect 470 -3310 790 -2990
rect 126 -3334 790 -3310
rect -308 -3451 12 -3409
rect 470 -3500 790 -3334
rect 814 -2891 1134 -2849
rect 814 -3409 856 -2891
rect 1092 -3409 1134 -2891
rect 1592 -2966 1912 -2634
rect 1936 -2191 2256 -2149
rect 1936 -2709 1978 -2191
rect 2214 -2709 2256 -2191
rect 2714 -2266 3034 -1934
rect 3058 -1491 3378 -1449
rect 3058 -2009 3100 -1491
rect 3336 -2009 3378 -1491
rect 3836 -1566 4156 -1234
rect 4180 -791 4500 -749
rect 4180 -1309 4222 -791
rect 4458 -1309 4500 -791
rect 4958 -866 5278 -534
rect 5302 -91 5622 -49
rect 5302 -609 5344 -91
rect 5580 -609 5622 -91
rect 5302 -651 5622 -609
rect 4614 -890 5278 -866
rect 4614 -1210 4638 -890
rect 4958 -1210 5278 -890
rect 4614 -1234 5278 -1210
rect 4180 -1351 4500 -1309
rect 3492 -1590 4156 -1566
rect 3492 -1910 3516 -1590
rect 3836 -1910 4156 -1590
rect 3492 -1934 4156 -1910
rect 3058 -2051 3378 -2009
rect 2370 -2290 3034 -2266
rect 2370 -2610 2394 -2290
rect 2714 -2610 3034 -2290
rect 2370 -2634 3034 -2610
rect 1936 -2751 2256 -2709
rect 1248 -2990 1912 -2966
rect 1248 -3310 1272 -2990
rect 1592 -3310 1912 -2990
rect 1248 -3334 1912 -3310
rect 814 -3451 1134 -3409
rect 1592 -3500 1912 -3334
rect 1936 -2891 2256 -2849
rect 1936 -3409 1978 -2891
rect 2214 -3409 2256 -2891
rect 2714 -2966 3034 -2634
rect 3058 -2191 3378 -2149
rect 3058 -2709 3100 -2191
rect 3336 -2709 3378 -2191
rect 3836 -2266 4156 -1934
rect 4180 -1491 4500 -1449
rect 4180 -2009 4222 -1491
rect 4458 -2009 4500 -1491
rect 4958 -1566 5278 -1234
rect 5302 -791 5622 -749
rect 5302 -1309 5344 -791
rect 5580 -1309 5622 -791
rect 5302 -1351 5622 -1309
rect 4614 -1590 5278 -1566
rect 4614 -1910 4638 -1590
rect 4958 -1910 5278 -1590
rect 4614 -1934 5278 -1910
rect 4180 -2051 4500 -2009
rect 3492 -2290 4156 -2266
rect 3492 -2610 3516 -2290
rect 3836 -2610 4156 -2290
rect 3492 -2634 4156 -2610
rect 3058 -2751 3378 -2709
rect 2370 -2990 3034 -2966
rect 2370 -3310 2394 -2990
rect 2714 -3310 3034 -2990
rect 2370 -3334 3034 -3310
rect 1936 -3451 2256 -3409
rect 2714 -3500 3034 -3334
rect 3058 -2891 3378 -2849
rect 3058 -3409 3100 -2891
rect 3336 -3409 3378 -2891
rect 3836 -2966 4156 -2634
rect 4180 -2191 4500 -2149
rect 4180 -2709 4222 -2191
rect 4458 -2709 4500 -2191
rect 4958 -2266 5278 -1934
rect 5302 -1491 5622 -1449
rect 5302 -2009 5344 -1491
rect 5580 -2009 5622 -1491
rect 5302 -2051 5622 -2009
rect 4614 -2290 5278 -2266
rect 4614 -2610 4638 -2290
rect 4958 -2610 5278 -2290
rect 4614 -2634 5278 -2610
rect 4180 -2751 4500 -2709
rect 3492 -2990 4156 -2966
rect 3492 -3310 3516 -2990
rect 3836 -3310 4156 -2990
rect 3492 -3334 4156 -3310
rect 3058 -3451 3378 -3409
rect 3836 -3500 4156 -3334
rect 4180 -2891 4500 -2849
rect 4180 -3409 4222 -2891
rect 4458 -3409 4500 -2891
rect 4958 -2966 5278 -2634
rect 5302 -2191 5622 -2149
rect 5302 -2709 5344 -2191
rect 5580 -2709 5622 -2191
rect 5302 -2751 5622 -2709
rect 4614 -2990 5278 -2966
rect 4614 -3310 4638 -2990
rect 4958 -3310 5278 -2990
rect 4614 -3334 5278 -3310
rect 4180 -3451 4500 -3409
rect 4958 -3500 5278 -3334
rect 5302 -2891 5622 -2849
rect 5302 -3409 5344 -2891
rect 5580 -3409 5622 -2891
rect 5302 -3451 5622 -3409
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX 4498 2850 5098 3450
string parameters w 2.00 l 2.00 val 5.36 carea 1.00 cperi 0.17 nx 10 ny 10 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 0 ccov 100
string library sky130
<< end >>
