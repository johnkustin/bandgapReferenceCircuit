magic
tech sky130A
magscale 1 2
timestamp 1620340193
<< nwell >>
rect -752 -4398 752 4364
<< pmoslvt >>
rect -658 -4336 -258 4264
rect -200 -4336 200 4264
rect 258 -4336 658 4264
<< pdiff >>
rect -716 4252 -658 4264
rect -716 -4324 -704 4252
rect -670 -4324 -658 4252
rect -716 -4336 -658 -4324
rect -258 4252 -200 4264
rect -258 -4324 -246 4252
rect -212 -4324 -200 4252
rect -258 -4336 -200 -4324
rect 200 4252 258 4264
rect 200 -4324 212 4252
rect 246 -4324 258 4252
rect 200 -4336 258 -4324
rect 658 4252 716 4264
rect 658 -4324 670 4252
rect 704 -4324 716 4252
rect 658 -4336 716 -4324
<< pdiffc >>
rect -704 -4324 -670 4252
rect -246 -4324 -212 4252
rect 212 -4324 246 4252
rect 670 -4324 704 4252
<< poly >>
rect -658 4345 -258 4361
rect -658 4311 -642 4345
rect -274 4311 -258 4345
rect -658 4264 -258 4311
rect -200 4345 200 4361
rect -200 4311 -184 4345
rect 184 4311 200 4345
rect -200 4264 200 4311
rect 258 4345 658 4361
rect 258 4311 274 4345
rect 642 4311 658 4345
rect 258 4264 658 4311
rect -658 -4362 -258 -4336
rect -200 -4362 200 -4336
rect 258 -4362 658 -4336
<< polycont >>
rect -642 4311 -274 4345
rect -184 4311 184 4345
rect 274 4311 642 4345
<< locali >>
rect -658 4311 -642 4345
rect -274 4311 -258 4345
rect -200 4311 -184 4345
rect 184 4311 200 4345
rect 258 4311 274 4345
rect 642 4311 658 4345
rect -704 4252 -670 4268
rect -704 -4340 -670 -4324
rect -246 4252 -212 4268
rect -246 -4340 -212 -4324
rect 212 4252 246 4268
rect 212 -4340 246 -4324
rect 670 4252 704 4268
rect 670 -4340 704 -4324
<< viali >>
rect -550 4311 -366 4345
rect -92 4311 92 4345
rect 366 4311 550 4345
rect -704 -4324 -670 4252
rect -246 -4324 -212 4252
rect 212 -4324 246 4252
rect 670 -4324 704 4252
<< metal1 >>
rect -562 4345 -354 4351
rect -562 4311 -550 4345
rect -366 4311 -354 4345
rect -562 4305 -354 4311
rect -104 4345 104 4351
rect -104 4311 -92 4345
rect 92 4311 104 4345
rect -104 4305 104 4311
rect 354 4345 562 4351
rect 354 4311 366 4345
rect 550 4311 562 4345
rect 354 4305 562 4311
rect -710 4252 -664 4264
rect -710 -4324 -704 4252
rect -670 -4324 -664 4252
rect -710 -4336 -664 -4324
rect -252 4252 -206 4264
rect -252 -4324 -246 4252
rect -212 -4324 -206 4252
rect -252 -4336 -206 -4324
rect 206 4252 252 4264
rect 206 -4324 212 4252
rect 246 -4324 252 4252
rect 206 -4336 252 -4324
rect 664 4252 710 4264
rect 664 -4324 670 4252
rect 704 -4324 710 4252
rect 664 -4336 710 -4324
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 43 l 2 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 50 viadrn 100 viasrc 100
string library sky130
<< end >>
