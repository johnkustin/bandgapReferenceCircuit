magic
tech sky130A
magscale 1 2
timestamp 1620886664
<< xpolycontact >>
rect -35 487 35 919
rect -35 -919 35 -487
<< xpolyres >>
rect -35 -487 35 487
<< viali >>
rect -19 504 19 901
rect -19 -901 19 -504
<< metal1 >>
rect -25 901 25 913
rect -25 504 -19 901
rect 19 504 25 901
rect -25 492 25 504
rect -25 -504 25 -492
rect -25 -901 -19 -504
rect 19 -901 25 -504
rect -25 -913 25 -901
<< res0p69 >>
rect -37 -489 37 489
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p69
string parameters w 0.350 l 4.87 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 27.938k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
