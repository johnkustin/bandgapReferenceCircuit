magic
tech sky130A
magscale 1 2
timestamp 1620594042
<< error_p >>
rect -2355 -3968 2355 3934
<< nwell >>
rect -2355 -3968 2355 3934
<< pmoslvt >>
rect -2261 -3906 -1861 3834
rect -1803 -3906 -1403 3834
rect -1345 -3906 -945 3834
rect -887 -3906 -487 3834
rect -429 -3906 -29 3834
rect 29 -3906 429 3834
rect 487 -3906 887 3834
rect 945 -3906 1345 3834
rect 1403 -3906 1803 3834
rect 1861 -3906 2261 3834
<< pdiff >>
rect -2319 3822 -2261 3834
rect -2319 -3894 -2307 3822
rect -2273 -3894 -2261 3822
rect -2319 -3906 -2261 -3894
rect -1861 3822 -1803 3834
rect -1861 -3894 -1849 3822
rect -1815 -3894 -1803 3822
rect -1861 -3906 -1803 -3894
rect -1403 3822 -1345 3834
rect -1403 -3894 -1391 3822
rect -1357 -3894 -1345 3822
rect -1403 -3906 -1345 -3894
rect -945 3822 -887 3834
rect -945 -3894 -933 3822
rect -899 -3894 -887 3822
rect -945 -3906 -887 -3894
rect -487 3822 -429 3834
rect -487 -3894 -475 3822
rect -441 -3894 -429 3822
rect -487 -3906 -429 -3894
rect -29 3822 29 3834
rect -29 -3894 -17 3822
rect 17 -3894 29 3822
rect -29 -3906 29 -3894
rect 429 3822 487 3834
rect 429 -3894 441 3822
rect 475 -3894 487 3822
rect 429 -3906 487 -3894
rect 887 3822 945 3834
rect 887 -3894 899 3822
rect 933 -3894 945 3822
rect 887 -3906 945 -3894
rect 1345 3822 1403 3834
rect 1345 -3894 1357 3822
rect 1391 -3894 1403 3822
rect 1345 -3906 1403 -3894
rect 1803 3822 1861 3834
rect 1803 -3894 1815 3822
rect 1849 -3894 1861 3822
rect 1803 -3906 1861 -3894
rect 2261 3822 2319 3834
rect 2261 -3894 2273 3822
rect 2307 -3894 2319 3822
rect 2261 -3906 2319 -3894
<< pdiffc >>
rect -2307 -3894 -2273 3822
rect -1849 -3894 -1815 3822
rect -1391 -3894 -1357 3822
rect -933 -3894 -899 3822
rect -475 -3894 -441 3822
rect -17 -3894 17 3822
rect 441 -3894 475 3822
rect 899 -3894 933 3822
rect 1357 -3894 1391 3822
rect 1815 -3894 1849 3822
rect 2273 -3894 2307 3822
<< poly >>
rect -2261 3915 -1861 3931
rect -2261 3881 -2245 3915
rect -1877 3881 -1861 3915
rect -2261 3834 -1861 3881
rect -1803 3915 -1403 3931
rect -1803 3881 -1787 3915
rect -1419 3881 -1403 3915
rect -1803 3834 -1403 3881
rect -1345 3915 -945 3931
rect -1345 3881 -1329 3915
rect -961 3881 -945 3915
rect -1345 3834 -945 3881
rect -887 3915 -487 3931
rect -887 3881 -871 3915
rect -503 3881 -487 3915
rect -887 3834 -487 3881
rect -429 3915 -29 3931
rect -429 3881 -413 3915
rect -45 3881 -29 3915
rect -429 3834 -29 3881
rect 29 3915 429 3931
rect 29 3881 45 3915
rect 413 3881 429 3915
rect 29 3834 429 3881
rect 487 3915 887 3931
rect 487 3881 503 3915
rect 871 3881 887 3915
rect 487 3834 887 3881
rect 945 3915 1345 3931
rect 945 3881 961 3915
rect 1329 3881 1345 3915
rect 945 3834 1345 3881
rect 1403 3915 1803 3931
rect 1403 3881 1419 3915
rect 1787 3881 1803 3915
rect 1403 3834 1803 3881
rect 1861 3915 2261 3931
rect 1861 3881 1877 3915
rect 2245 3881 2261 3915
rect 1861 3834 2261 3881
rect -2261 -3932 -1861 -3906
rect -1803 -3932 -1403 -3906
rect -1345 -3932 -945 -3906
rect -887 -3932 -487 -3906
rect -429 -3932 -29 -3906
rect 29 -3932 429 -3906
rect 487 -3932 887 -3906
rect 945 -3932 1345 -3906
rect 1403 -3932 1803 -3906
rect 1861 -3932 2261 -3906
<< polycont >>
rect -2245 3881 -1877 3915
rect -1787 3881 -1419 3915
rect -1329 3881 -961 3915
rect -871 3881 -503 3915
rect -413 3881 -45 3915
rect 45 3881 413 3915
rect 503 3881 871 3915
rect 961 3881 1329 3915
rect 1419 3881 1787 3915
rect 1877 3881 2245 3915
<< locali >>
rect -2261 3881 -2245 3915
rect -1877 3881 -1861 3915
rect -1803 3881 -1787 3915
rect -1419 3881 -1403 3915
rect -1345 3881 -1329 3915
rect -961 3881 -945 3915
rect -887 3881 -871 3915
rect -503 3881 -487 3915
rect -429 3881 -413 3915
rect -45 3881 -29 3915
rect 29 3881 45 3915
rect 413 3881 429 3915
rect 487 3881 503 3915
rect 871 3881 887 3915
rect 945 3881 961 3915
rect 1329 3881 1345 3915
rect 1403 3881 1419 3915
rect 1787 3881 1803 3915
rect 1861 3881 1877 3915
rect 2245 3881 2261 3915
rect -2307 3822 -2273 3838
rect -2307 -3910 -2273 -3894
rect -1849 3822 -1815 3838
rect -1849 -3910 -1815 -3894
rect -1391 3822 -1357 3838
rect -1391 -3910 -1357 -3894
rect -933 3822 -899 3838
rect -933 -3910 -899 -3894
rect -475 3822 -441 3838
rect -475 -3910 -441 -3894
rect -17 3822 17 3838
rect -17 -3910 17 -3894
rect 441 3822 475 3838
rect 441 -3910 475 -3894
rect 899 3822 933 3838
rect 899 -3910 933 -3894
rect 1357 3822 1391 3838
rect 1357 -3910 1391 -3894
rect 1815 3822 1849 3838
rect 1815 -3910 1849 -3894
rect 2273 3822 2307 3838
rect 2273 -3910 2307 -3894
<< viali >>
rect -2153 3881 -1969 3915
rect -1695 3881 -1511 3915
rect -1237 3881 -1053 3915
rect -779 3881 -595 3915
rect -321 3881 -137 3915
rect 137 3881 321 3915
rect 595 3881 779 3915
rect 1053 3881 1237 3915
rect 1511 3881 1695 3915
rect 1969 3881 2153 3915
rect -2307 -3894 -2273 3822
rect -1849 -3894 -1815 3822
rect -1391 -3894 -1357 3822
rect -933 -3894 -899 3822
rect -475 -3894 -441 3822
rect -17 -3894 17 3822
rect 441 -3894 475 3822
rect 899 -3894 933 3822
rect 1357 -3894 1391 3822
rect 1815 -3894 1849 3822
rect 2273 -3894 2307 3822
<< metal1 >>
rect -2165 3915 -1957 3921
rect -2165 3881 -2153 3915
rect -1969 3881 -1957 3915
rect -2165 3875 -1957 3881
rect -1707 3915 -1499 3921
rect -1707 3881 -1695 3915
rect -1511 3881 -1499 3915
rect -1707 3875 -1499 3881
rect -1249 3915 -1041 3921
rect -1249 3881 -1237 3915
rect -1053 3881 -1041 3915
rect -1249 3875 -1041 3881
rect -791 3915 -583 3921
rect -791 3881 -779 3915
rect -595 3881 -583 3915
rect -791 3875 -583 3881
rect -333 3915 -125 3921
rect -333 3881 -321 3915
rect -137 3881 -125 3915
rect -333 3875 -125 3881
rect 125 3915 333 3921
rect 125 3881 137 3915
rect 321 3881 333 3915
rect 125 3875 333 3881
rect 583 3915 791 3921
rect 583 3881 595 3915
rect 779 3881 791 3915
rect 583 3875 791 3881
rect 1041 3915 1249 3921
rect 1041 3881 1053 3915
rect 1237 3881 1249 3915
rect 1041 3875 1249 3881
rect 1499 3915 1707 3921
rect 1499 3881 1511 3915
rect 1695 3881 1707 3915
rect 1499 3875 1707 3881
rect 1957 3915 2165 3921
rect 1957 3881 1969 3915
rect 2153 3881 2165 3915
rect 1957 3875 2165 3881
rect -2313 3822 -2267 3834
rect -2313 -3894 -2307 3822
rect -2273 -3894 -2267 3822
rect -2313 -3906 -2267 -3894
rect -1855 3822 -1809 3834
rect -1855 -3894 -1849 3822
rect -1815 -3894 -1809 3822
rect -1855 -3906 -1809 -3894
rect -1397 3822 -1351 3834
rect -1397 -3894 -1391 3822
rect -1357 -3894 -1351 3822
rect -1397 -3906 -1351 -3894
rect -939 3822 -893 3834
rect -939 -3894 -933 3822
rect -899 -3894 -893 3822
rect -939 -3906 -893 -3894
rect -481 3822 -435 3834
rect -481 -3894 -475 3822
rect -441 -3894 -435 3822
rect -481 -3906 -435 -3894
rect -23 3822 23 3834
rect -23 -3894 -17 3822
rect 17 -3894 23 3822
rect -23 -3906 23 -3894
rect 435 3822 481 3834
rect 435 -3894 441 3822
rect 475 -3894 481 3822
rect 435 -3906 481 -3894
rect 893 3822 939 3834
rect 893 -3894 899 3822
rect 933 -3894 939 3822
rect 893 -3906 939 -3894
rect 1351 3822 1397 3834
rect 1351 -3894 1357 3822
rect 1391 -3894 1397 3822
rect 1351 -3906 1397 -3894
rect 1809 3822 1855 3834
rect 1809 -3894 1815 3822
rect 1849 -3894 1855 3822
rect 1809 -3906 1855 -3894
rect 2267 3822 2313 3834
rect 2267 -3894 2273 3822
rect 2307 -3894 2313 3822
rect 2267 -3906 2313 -3894
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 38.7 l 2 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 50 viadrn 100 viasrc 100
string library sky130
<< end >>
