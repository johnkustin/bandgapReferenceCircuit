magic
tech sky130A
timestamp 1620324069
<< nwell >>
rect -4956 -1381 4956 1381
<< pmoslvt >>
rect -4909 -1350 -4709 1350
rect -4680 -1350 -4480 1350
rect -4451 -1350 -4251 1350
rect -4222 -1350 -4022 1350
rect -3993 -1350 -3793 1350
rect -3764 -1350 -3564 1350
rect -3535 -1350 -3335 1350
rect -3306 -1350 -3106 1350
rect -3077 -1350 -2877 1350
rect -2848 -1350 -2648 1350
rect -2619 -1350 -2419 1350
rect -2390 -1350 -2190 1350
rect -2161 -1350 -1961 1350
rect -1932 -1350 -1732 1350
rect -1703 -1350 -1503 1350
rect -1474 -1350 -1274 1350
rect -1245 -1350 -1045 1350
rect -1016 -1350 -816 1350
rect -787 -1350 -587 1350
rect -558 -1350 -358 1350
rect -329 -1350 -129 1350
rect -100 -1350 100 1350
rect 129 -1350 329 1350
rect 358 -1350 558 1350
rect 587 -1350 787 1350
rect 816 -1350 1016 1350
rect 1045 -1350 1245 1350
rect 1274 -1350 1474 1350
rect 1503 -1350 1703 1350
rect 1732 -1350 1932 1350
rect 1961 -1350 2161 1350
rect 2190 -1350 2390 1350
rect 2419 -1350 2619 1350
rect 2648 -1350 2848 1350
rect 2877 -1350 3077 1350
rect 3106 -1350 3306 1350
rect 3335 -1350 3535 1350
rect 3564 -1350 3764 1350
rect 3793 -1350 3993 1350
rect 4022 -1350 4222 1350
rect 4251 -1350 4451 1350
rect 4480 -1350 4680 1350
rect 4709 -1350 4909 1350
<< pdiff >>
rect -4938 1344 -4909 1350
rect -4938 -1344 -4932 1344
rect -4915 -1344 -4909 1344
rect -4938 -1350 -4909 -1344
rect -4709 1344 -4680 1350
rect -4709 -1344 -4703 1344
rect -4686 -1344 -4680 1344
rect -4709 -1350 -4680 -1344
rect -4480 1344 -4451 1350
rect -4480 -1344 -4474 1344
rect -4457 -1344 -4451 1344
rect -4480 -1350 -4451 -1344
rect -4251 1344 -4222 1350
rect -4251 -1344 -4245 1344
rect -4228 -1344 -4222 1344
rect -4251 -1350 -4222 -1344
rect -4022 1344 -3993 1350
rect -4022 -1344 -4016 1344
rect -3999 -1344 -3993 1344
rect -4022 -1350 -3993 -1344
rect -3793 1344 -3764 1350
rect -3793 -1344 -3787 1344
rect -3770 -1344 -3764 1344
rect -3793 -1350 -3764 -1344
rect -3564 1344 -3535 1350
rect -3564 -1344 -3558 1344
rect -3541 -1344 -3535 1344
rect -3564 -1350 -3535 -1344
rect -3335 1344 -3306 1350
rect -3335 -1344 -3329 1344
rect -3312 -1344 -3306 1344
rect -3335 -1350 -3306 -1344
rect -3106 1344 -3077 1350
rect -3106 -1344 -3100 1344
rect -3083 -1344 -3077 1344
rect -3106 -1350 -3077 -1344
rect -2877 1344 -2848 1350
rect -2877 -1344 -2871 1344
rect -2854 -1344 -2848 1344
rect -2877 -1350 -2848 -1344
rect -2648 1344 -2619 1350
rect -2648 -1344 -2642 1344
rect -2625 -1344 -2619 1344
rect -2648 -1350 -2619 -1344
rect -2419 1344 -2390 1350
rect -2419 -1344 -2413 1344
rect -2396 -1344 -2390 1344
rect -2419 -1350 -2390 -1344
rect -2190 1344 -2161 1350
rect -2190 -1344 -2184 1344
rect -2167 -1344 -2161 1344
rect -2190 -1350 -2161 -1344
rect -1961 1344 -1932 1350
rect -1961 -1344 -1955 1344
rect -1938 -1344 -1932 1344
rect -1961 -1350 -1932 -1344
rect -1732 1344 -1703 1350
rect -1732 -1344 -1726 1344
rect -1709 -1344 -1703 1344
rect -1732 -1350 -1703 -1344
rect -1503 1344 -1474 1350
rect -1503 -1344 -1497 1344
rect -1480 -1344 -1474 1344
rect -1503 -1350 -1474 -1344
rect -1274 1344 -1245 1350
rect -1274 -1344 -1268 1344
rect -1251 -1344 -1245 1344
rect -1274 -1350 -1245 -1344
rect -1045 1344 -1016 1350
rect -1045 -1344 -1039 1344
rect -1022 -1344 -1016 1344
rect -1045 -1350 -1016 -1344
rect -816 1344 -787 1350
rect -816 -1344 -810 1344
rect -793 -1344 -787 1344
rect -816 -1350 -787 -1344
rect -587 1344 -558 1350
rect -587 -1344 -581 1344
rect -564 -1344 -558 1344
rect -587 -1350 -558 -1344
rect -358 1344 -329 1350
rect -358 -1344 -352 1344
rect -335 -1344 -329 1344
rect -358 -1350 -329 -1344
rect -129 1344 -100 1350
rect -129 -1344 -123 1344
rect -106 -1344 -100 1344
rect -129 -1350 -100 -1344
rect 100 1344 129 1350
rect 100 -1344 106 1344
rect 123 -1344 129 1344
rect 100 -1350 129 -1344
rect 329 1344 358 1350
rect 329 -1344 335 1344
rect 352 -1344 358 1344
rect 329 -1350 358 -1344
rect 558 1344 587 1350
rect 558 -1344 564 1344
rect 581 -1344 587 1344
rect 558 -1350 587 -1344
rect 787 1344 816 1350
rect 787 -1344 793 1344
rect 810 -1344 816 1344
rect 787 -1350 816 -1344
rect 1016 1344 1045 1350
rect 1016 -1344 1022 1344
rect 1039 -1344 1045 1344
rect 1016 -1350 1045 -1344
rect 1245 1344 1274 1350
rect 1245 -1344 1251 1344
rect 1268 -1344 1274 1344
rect 1245 -1350 1274 -1344
rect 1474 1344 1503 1350
rect 1474 -1344 1480 1344
rect 1497 -1344 1503 1344
rect 1474 -1350 1503 -1344
rect 1703 1344 1732 1350
rect 1703 -1344 1709 1344
rect 1726 -1344 1732 1344
rect 1703 -1350 1732 -1344
rect 1932 1344 1961 1350
rect 1932 -1344 1938 1344
rect 1955 -1344 1961 1344
rect 1932 -1350 1961 -1344
rect 2161 1344 2190 1350
rect 2161 -1344 2167 1344
rect 2184 -1344 2190 1344
rect 2161 -1350 2190 -1344
rect 2390 1344 2419 1350
rect 2390 -1344 2396 1344
rect 2413 -1344 2419 1344
rect 2390 -1350 2419 -1344
rect 2619 1344 2648 1350
rect 2619 -1344 2625 1344
rect 2642 -1344 2648 1344
rect 2619 -1350 2648 -1344
rect 2848 1344 2877 1350
rect 2848 -1344 2854 1344
rect 2871 -1344 2877 1344
rect 2848 -1350 2877 -1344
rect 3077 1344 3106 1350
rect 3077 -1344 3083 1344
rect 3100 -1344 3106 1344
rect 3077 -1350 3106 -1344
rect 3306 1344 3335 1350
rect 3306 -1344 3312 1344
rect 3329 -1344 3335 1344
rect 3306 -1350 3335 -1344
rect 3535 1344 3564 1350
rect 3535 -1344 3541 1344
rect 3558 -1344 3564 1344
rect 3535 -1350 3564 -1344
rect 3764 1344 3793 1350
rect 3764 -1344 3770 1344
rect 3787 -1344 3793 1344
rect 3764 -1350 3793 -1344
rect 3993 1344 4022 1350
rect 3993 -1344 3999 1344
rect 4016 -1344 4022 1344
rect 3993 -1350 4022 -1344
rect 4222 1344 4251 1350
rect 4222 -1344 4228 1344
rect 4245 -1344 4251 1344
rect 4222 -1350 4251 -1344
rect 4451 1344 4480 1350
rect 4451 -1344 4457 1344
rect 4474 -1344 4480 1344
rect 4451 -1350 4480 -1344
rect 4680 1344 4709 1350
rect 4680 -1344 4686 1344
rect 4703 -1344 4709 1344
rect 4680 -1350 4709 -1344
rect 4909 1344 4938 1350
rect 4909 -1344 4915 1344
rect 4932 -1344 4938 1344
rect 4909 -1350 4938 -1344
<< pdiffc >>
rect -4932 -1344 -4915 1344
rect -4703 -1344 -4686 1344
rect -4474 -1344 -4457 1344
rect -4245 -1344 -4228 1344
rect -4016 -1344 -3999 1344
rect -3787 -1344 -3770 1344
rect -3558 -1344 -3541 1344
rect -3329 -1344 -3312 1344
rect -3100 -1344 -3083 1344
rect -2871 -1344 -2854 1344
rect -2642 -1344 -2625 1344
rect -2413 -1344 -2396 1344
rect -2184 -1344 -2167 1344
rect -1955 -1344 -1938 1344
rect -1726 -1344 -1709 1344
rect -1497 -1344 -1480 1344
rect -1268 -1344 -1251 1344
rect -1039 -1344 -1022 1344
rect -810 -1344 -793 1344
rect -581 -1344 -564 1344
rect -352 -1344 -335 1344
rect -123 -1344 -106 1344
rect 106 -1344 123 1344
rect 335 -1344 352 1344
rect 564 -1344 581 1344
rect 793 -1344 810 1344
rect 1022 -1344 1039 1344
rect 1251 -1344 1268 1344
rect 1480 -1344 1497 1344
rect 1709 -1344 1726 1344
rect 1938 -1344 1955 1344
rect 2167 -1344 2184 1344
rect 2396 -1344 2413 1344
rect 2625 -1344 2642 1344
rect 2854 -1344 2871 1344
rect 3083 -1344 3100 1344
rect 3312 -1344 3329 1344
rect 3541 -1344 3558 1344
rect 3770 -1344 3787 1344
rect 3999 -1344 4016 1344
rect 4228 -1344 4245 1344
rect 4457 -1344 4474 1344
rect 4686 -1344 4703 1344
rect 4915 -1344 4932 1344
<< poly >>
rect -4909 1350 -4709 1363
rect -4680 1350 -4480 1363
rect -4451 1350 -4251 1363
rect -4222 1350 -4022 1363
rect -3993 1350 -3793 1363
rect -3764 1350 -3564 1363
rect -3535 1350 -3335 1363
rect -3306 1350 -3106 1363
rect -3077 1350 -2877 1363
rect -2848 1350 -2648 1363
rect -2619 1350 -2419 1363
rect -2390 1350 -2190 1363
rect -2161 1350 -1961 1363
rect -1932 1350 -1732 1363
rect -1703 1350 -1503 1363
rect -1474 1350 -1274 1363
rect -1245 1350 -1045 1363
rect -1016 1350 -816 1363
rect -787 1350 -587 1363
rect -558 1350 -358 1363
rect -329 1350 -129 1363
rect -100 1350 100 1363
rect 129 1350 329 1363
rect 358 1350 558 1363
rect 587 1350 787 1363
rect 816 1350 1016 1363
rect 1045 1350 1245 1363
rect 1274 1350 1474 1363
rect 1503 1350 1703 1363
rect 1732 1350 1932 1363
rect 1961 1350 2161 1363
rect 2190 1350 2390 1363
rect 2419 1350 2619 1363
rect 2648 1350 2848 1363
rect 2877 1350 3077 1363
rect 3106 1350 3306 1363
rect 3335 1350 3535 1363
rect 3564 1350 3764 1363
rect 3793 1350 3993 1363
rect 4022 1350 4222 1363
rect 4251 1350 4451 1363
rect 4480 1350 4680 1363
rect 4709 1350 4909 1363
rect -4909 -1363 -4709 -1350
rect -4680 -1363 -4480 -1350
rect -4451 -1363 -4251 -1350
rect -4222 -1363 -4022 -1350
rect -3993 -1363 -3793 -1350
rect -3764 -1363 -3564 -1350
rect -3535 -1363 -3335 -1350
rect -3306 -1363 -3106 -1350
rect -3077 -1363 -2877 -1350
rect -2848 -1363 -2648 -1350
rect -2619 -1363 -2419 -1350
rect -2390 -1363 -2190 -1350
rect -2161 -1363 -1961 -1350
rect -1932 -1363 -1732 -1350
rect -1703 -1363 -1503 -1350
rect -1474 -1363 -1274 -1350
rect -1245 -1363 -1045 -1350
rect -1016 -1363 -816 -1350
rect -787 -1363 -587 -1350
rect -558 -1363 -358 -1350
rect -329 -1363 -129 -1350
rect -100 -1363 100 -1350
rect 129 -1363 329 -1350
rect 358 -1363 558 -1350
rect 587 -1363 787 -1350
rect 816 -1363 1016 -1350
rect 1045 -1363 1245 -1350
rect 1274 -1363 1474 -1350
rect 1503 -1363 1703 -1350
rect 1732 -1363 1932 -1350
rect 1961 -1363 2161 -1350
rect 2190 -1363 2390 -1350
rect 2419 -1363 2619 -1350
rect 2648 -1363 2848 -1350
rect 2877 -1363 3077 -1350
rect 3106 -1363 3306 -1350
rect 3335 -1363 3535 -1350
rect 3564 -1363 3764 -1350
rect 3793 -1363 3993 -1350
rect 4022 -1363 4222 -1350
rect 4251 -1363 4451 -1350
rect 4480 -1363 4680 -1350
rect 4709 -1363 4909 -1350
<< locali >>
rect -4932 1344 -4915 1352
rect -4932 -1352 -4915 -1344
rect -4703 1344 -4686 1352
rect -4703 -1352 -4686 -1344
rect -4474 1344 -4457 1352
rect -4474 -1352 -4457 -1344
rect -4245 1344 -4228 1352
rect -4245 -1352 -4228 -1344
rect -4016 1344 -3999 1352
rect -4016 -1352 -3999 -1344
rect -3787 1344 -3770 1352
rect -3787 -1352 -3770 -1344
rect -3558 1344 -3541 1352
rect -3558 -1352 -3541 -1344
rect -3329 1344 -3312 1352
rect -3329 -1352 -3312 -1344
rect -3100 1344 -3083 1352
rect -3100 -1352 -3083 -1344
rect -2871 1344 -2854 1352
rect -2871 -1352 -2854 -1344
rect -2642 1344 -2625 1352
rect -2642 -1352 -2625 -1344
rect -2413 1344 -2396 1352
rect -2413 -1352 -2396 -1344
rect -2184 1344 -2167 1352
rect -2184 -1352 -2167 -1344
rect -1955 1344 -1938 1352
rect -1955 -1352 -1938 -1344
rect -1726 1344 -1709 1352
rect -1726 -1352 -1709 -1344
rect -1497 1344 -1480 1352
rect -1497 -1352 -1480 -1344
rect -1268 1344 -1251 1352
rect -1268 -1352 -1251 -1344
rect -1039 1344 -1022 1352
rect -1039 -1352 -1022 -1344
rect -810 1344 -793 1352
rect -810 -1352 -793 -1344
rect -581 1344 -564 1352
rect -581 -1352 -564 -1344
rect -352 1344 -335 1352
rect -352 -1352 -335 -1344
rect -123 1344 -106 1352
rect -123 -1352 -106 -1344
rect 106 1344 123 1352
rect 106 -1352 123 -1344
rect 335 1344 352 1352
rect 335 -1352 352 -1344
rect 564 1344 581 1352
rect 564 -1352 581 -1344
rect 793 1344 810 1352
rect 793 -1352 810 -1344
rect 1022 1344 1039 1352
rect 1022 -1352 1039 -1344
rect 1251 1344 1268 1352
rect 1251 -1352 1268 -1344
rect 1480 1344 1497 1352
rect 1480 -1352 1497 -1344
rect 1709 1344 1726 1352
rect 1709 -1352 1726 -1344
rect 1938 1344 1955 1352
rect 1938 -1352 1955 -1344
rect 2167 1344 2184 1352
rect 2167 -1352 2184 -1344
rect 2396 1344 2413 1352
rect 2396 -1352 2413 -1344
rect 2625 1344 2642 1352
rect 2625 -1352 2642 -1344
rect 2854 1344 2871 1352
rect 2854 -1352 2871 -1344
rect 3083 1344 3100 1352
rect 3083 -1352 3100 -1344
rect 3312 1344 3329 1352
rect 3312 -1352 3329 -1344
rect 3541 1344 3558 1352
rect 3541 -1352 3558 -1344
rect 3770 1344 3787 1352
rect 3770 -1352 3787 -1344
rect 3999 1344 4016 1352
rect 3999 -1352 4016 -1344
rect 4228 1344 4245 1352
rect 4228 -1352 4245 -1344
rect 4457 1344 4474 1352
rect 4457 -1352 4474 -1344
rect 4686 1344 4703 1352
rect 4686 -1352 4703 -1344
rect 4915 1344 4932 1352
rect 4915 -1352 4932 -1344
<< viali >>
rect -4932 -1344 -4915 1344
rect -4703 -1344 -4686 1344
rect -4474 -1344 -4457 1344
rect -4245 -1344 -4228 1344
rect -4016 -1344 -3999 1344
rect -3787 -1344 -3770 1344
rect -3558 -1344 -3541 1344
rect -3329 -1344 -3312 1344
rect -3100 -1344 -3083 1344
rect -2871 -1344 -2854 1344
rect -2642 -1344 -2625 1344
rect -2413 -1344 -2396 1344
rect -2184 -1344 -2167 1344
rect -1955 -1344 -1938 1344
rect -1726 -1344 -1709 1344
rect -1497 -1344 -1480 1344
rect -1268 -1344 -1251 1344
rect -1039 -1344 -1022 1344
rect -810 -1344 -793 1344
rect -581 -1344 -564 1344
rect -352 -1344 -335 1344
rect -123 -1344 -106 1344
rect 106 -1344 123 1344
rect 335 -1344 352 1344
rect 564 -1344 581 1344
rect 793 -1344 810 1344
rect 1022 -1344 1039 1344
rect 1251 -1344 1268 1344
rect 1480 -1344 1497 1344
rect 1709 -1344 1726 1344
rect 1938 -1344 1955 1344
rect 2167 -1344 2184 1344
rect 2396 -1344 2413 1344
rect 2625 -1344 2642 1344
rect 2854 -1344 2871 1344
rect 3083 -1344 3100 1344
rect 3312 -1344 3329 1344
rect 3541 -1344 3558 1344
rect 3770 -1344 3787 1344
rect 3999 -1344 4016 1344
rect 4228 -1344 4245 1344
rect 4457 -1344 4474 1344
rect 4686 -1344 4703 1344
rect 4915 -1344 4932 1344
<< metal1 >>
rect -4935 1344 -4912 1350
rect -4935 -1344 -4932 1344
rect -4915 -1344 -4912 1344
rect -4935 -1350 -4912 -1344
rect -4706 1344 -4683 1350
rect -4706 -1344 -4703 1344
rect -4686 -1344 -4683 1344
rect -4706 -1350 -4683 -1344
rect -4477 1344 -4454 1350
rect -4477 -1344 -4474 1344
rect -4457 -1344 -4454 1344
rect -4477 -1350 -4454 -1344
rect -4248 1344 -4225 1350
rect -4248 -1344 -4245 1344
rect -4228 -1344 -4225 1344
rect -4248 -1350 -4225 -1344
rect -4019 1344 -3996 1350
rect -4019 -1344 -4016 1344
rect -3999 -1344 -3996 1344
rect -4019 -1350 -3996 -1344
rect -3790 1344 -3767 1350
rect -3790 -1344 -3787 1344
rect -3770 -1344 -3767 1344
rect -3790 -1350 -3767 -1344
rect -3561 1344 -3538 1350
rect -3561 -1344 -3558 1344
rect -3541 -1344 -3538 1344
rect -3561 -1350 -3538 -1344
rect -3332 1344 -3309 1350
rect -3332 -1344 -3329 1344
rect -3312 -1344 -3309 1344
rect -3332 -1350 -3309 -1344
rect -3103 1344 -3080 1350
rect -3103 -1344 -3100 1344
rect -3083 -1344 -3080 1344
rect -3103 -1350 -3080 -1344
rect -2874 1344 -2851 1350
rect -2874 -1344 -2871 1344
rect -2854 -1344 -2851 1344
rect -2874 -1350 -2851 -1344
rect -2645 1344 -2622 1350
rect -2645 -1344 -2642 1344
rect -2625 -1344 -2622 1344
rect -2645 -1350 -2622 -1344
rect -2416 1344 -2393 1350
rect -2416 -1344 -2413 1344
rect -2396 -1344 -2393 1344
rect -2416 -1350 -2393 -1344
rect -2187 1344 -2164 1350
rect -2187 -1344 -2184 1344
rect -2167 -1344 -2164 1344
rect -2187 -1350 -2164 -1344
rect -1958 1344 -1935 1350
rect -1958 -1344 -1955 1344
rect -1938 -1344 -1935 1344
rect -1958 -1350 -1935 -1344
rect -1729 1344 -1706 1350
rect -1729 -1344 -1726 1344
rect -1709 -1344 -1706 1344
rect -1729 -1350 -1706 -1344
rect -1500 1344 -1477 1350
rect -1500 -1344 -1497 1344
rect -1480 -1344 -1477 1344
rect -1500 -1350 -1477 -1344
rect -1271 1344 -1248 1350
rect -1271 -1344 -1268 1344
rect -1251 -1344 -1248 1344
rect -1271 -1350 -1248 -1344
rect -1042 1344 -1019 1350
rect -1042 -1344 -1039 1344
rect -1022 -1344 -1019 1344
rect -1042 -1350 -1019 -1344
rect -813 1344 -790 1350
rect -813 -1344 -810 1344
rect -793 -1344 -790 1344
rect -813 -1350 -790 -1344
rect -584 1344 -561 1350
rect -584 -1344 -581 1344
rect -564 -1344 -561 1344
rect -584 -1350 -561 -1344
rect -355 1344 -332 1350
rect -355 -1344 -352 1344
rect -335 -1344 -332 1344
rect -355 -1350 -332 -1344
rect -126 1344 -103 1350
rect -126 -1344 -123 1344
rect -106 -1344 -103 1344
rect -126 -1350 -103 -1344
rect 103 1344 126 1350
rect 103 -1344 106 1344
rect 123 -1344 126 1344
rect 103 -1350 126 -1344
rect 332 1344 355 1350
rect 332 -1344 335 1344
rect 352 -1344 355 1344
rect 332 -1350 355 -1344
rect 561 1344 584 1350
rect 561 -1344 564 1344
rect 581 -1344 584 1344
rect 561 -1350 584 -1344
rect 790 1344 813 1350
rect 790 -1344 793 1344
rect 810 -1344 813 1344
rect 790 -1350 813 -1344
rect 1019 1344 1042 1350
rect 1019 -1344 1022 1344
rect 1039 -1344 1042 1344
rect 1019 -1350 1042 -1344
rect 1248 1344 1271 1350
rect 1248 -1344 1251 1344
rect 1268 -1344 1271 1344
rect 1248 -1350 1271 -1344
rect 1477 1344 1500 1350
rect 1477 -1344 1480 1344
rect 1497 -1344 1500 1344
rect 1477 -1350 1500 -1344
rect 1706 1344 1729 1350
rect 1706 -1344 1709 1344
rect 1726 -1344 1729 1344
rect 1706 -1350 1729 -1344
rect 1935 1344 1958 1350
rect 1935 -1344 1938 1344
rect 1955 -1344 1958 1344
rect 1935 -1350 1958 -1344
rect 2164 1344 2187 1350
rect 2164 -1344 2167 1344
rect 2184 -1344 2187 1344
rect 2164 -1350 2187 -1344
rect 2393 1344 2416 1350
rect 2393 -1344 2396 1344
rect 2413 -1344 2416 1344
rect 2393 -1350 2416 -1344
rect 2622 1344 2645 1350
rect 2622 -1344 2625 1344
rect 2642 -1344 2645 1344
rect 2622 -1350 2645 -1344
rect 2851 1344 2874 1350
rect 2851 -1344 2854 1344
rect 2871 -1344 2874 1344
rect 2851 -1350 2874 -1344
rect 3080 1344 3103 1350
rect 3080 -1344 3083 1344
rect 3100 -1344 3103 1344
rect 3080 -1350 3103 -1344
rect 3309 1344 3332 1350
rect 3309 -1344 3312 1344
rect 3329 -1344 3332 1344
rect 3309 -1350 3332 -1344
rect 3538 1344 3561 1350
rect 3538 -1344 3541 1344
rect 3558 -1344 3561 1344
rect 3538 -1350 3561 -1344
rect 3767 1344 3790 1350
rect 3767 -1344 3770 1344
rect 3787 -1344 3790 1344
rect 3767 -1350 3790 -1344
rect 3996 1344 4019 1350
rect 3996 -1344 3999 1344
rect 4016 -1344 4019 1344
rect 3996 -1350 4019 -1344
rect 4225 1344 4248 1350
rect 4225 -1344 4228 1344
rect 4245 -1344 4248 1344
rect 4225 -1350 4248 -1344
rect 4454 1344 4477 1350
rect 4454 -1344 4457 1344
rect 4474 -1344 4477 1344
rect 4454 -1350 4477 -1344
rect 4683 1344 4706 1350
rect 4683 -1344 4686 1344
rect 4703 -1344 4706 1344
rect 4683 -1350 4706 -1344
rect 4912 1344 4935 1350
rect 4912 -1344 4915 1344
rect 4932 -1344 4935 1344
rect 4912 -1350 4935 -1344
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 27 l 2 m 1 nf 43 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
