magic
tech sky130A
magscale 1 2
timestamp 1621229569
<< error_p >>
rect 16156 -20900 16162 -20894
rect 16162 -20906 16168 -20900
<< error_s >>
rect 16162 -19966 16168 -19960
rect 16674 -19966 16680 -19960
rect 16156 -19972 16162 -19966
rect 16680 -19972 16686 -19966
<< pwell >>
rect 16590 -17702 16652 -17564
<< psubdiff >>
rect 7278 -16480 13630 -16456
rect 7278 -17050 7302 -16480
rect 13606 -17050 13630 -16480
rect 7278 -17074 13630 -17050
rect 16590 -17702 16652 -17564
rect 7278 -31168 13630 -31144
rect 7278 -31738 7302 -31168
rect 13606 -31738 13630 -31168
rect 7278 -31762 13630 -31738
rect 7278 -36128 13630 -36104
rect 7278 -36698 7302 -36128
rect 13606 -36698 13630 -36128
rect 7278 -36722 13630 -36698
rect 7278 -39372 13630 -39348
rect 7278 -39942 7302 -39372
rect 13606 -39942 13630 -39372
rect 7278 -39966 13630 -39942
<< psubdiffcont >>
rect 7302 -17050 13606 -16480
rect 7302 -31738 13606 -31168
rect 7302 -36698 13606 -36128
rect 7302 -39942 13606 -39372
<< xpolycontact >>
rect 6870 -17850 7302 -17280
rect 13606 -17850 14038 -17280
rect 13612 -18668 14038 -18098
rect 13612 -20304 14038 -19734
rect 13606 -21940 14038 -21370
rect 13606 -24394 14038 -23824
rect 13606 -25212 14038 -24642
rect 13606 -27666 14038 -27096
rect 13606 -28484 14038 -27914
rect 6870 -29302 7302 -28732
rect 13606 -30120 14038 -29550
<< locali >>
rect 16584 -11502 26884 -11302
rect 16584 -12802 26784 -12402
rect 16584 -14102 26784 -13702
rect 16584 -15402 26784 -15002
rect 6870 -16464 7302 -16456
rect 13606 -16464 14038 -16456
rect 6870 -16480 14038 -16464
rect 6870 -17050 7302 -16480
rect 13606 -17050 14038 -16480
rect 16584 -16702 26884 -16202
rect 6870 -17066 14038 -17050
rect 6870 -17280 7302 -17066
rect 13606 -17280 14038 -17066
rect 16584 -17562 26884 -17502
rect 16582 -17564 26884 -17562
rect 16582 -17580 16630 -17564
rect 16652 -17580 26884 -17564
rect 16582 -17702 26884 -17580
rect 16582 -17720 16630 -17702
rect 6870 -31152 7302 -30368
rect 13606 -31152 14038 -30368
rect 6870 -31168 14038 -31152
rect 6870 -31422 7302 -31168
rect 6808 -31738 7302 -31422
rect 13606 -31738 14038 -31168
rect 6808 -31754 14038 -31738
rect 6808 -31762 7302 -31754
rect 6808 -33392 7244 -31762
rect 6808 -36116 7240 -35276
rect 11540 -35846 12070 -31754
rect 13606 -31762 14038 -31754
rect 11544 -36112 12070 -35846
rect 12692 -36112 13200 -36102
rect 7286 -36116 13622 -36112
rect 6808 -36128 13622 -36116
rect 6808 -36698 7302 -36128
rect 13606 -36698 13622 -36128
rect 6808 -36714 13622 -36698
rect 6808 -36720 7798 -36714
rect 8194 -39356 8636 -36714
rect 11950 -37482 12382 -36714
rect 12692 -37742 13200 -36714
rect 12692 -38548 13200 -38290
rect 11950 -39118 13200 -38548
rect 12696 -39356 13200 -39118
rect 7286 -39372 13622 -39356
rect 7286 -39942 7302 -39372
rect 13606 -39942 13622 -39372
rect 7286 -39958 13622 -39942
rect 8194 -39968 8636 -39958
rect 12696 -39962 13200 -39958
<< viali >>
rect 13623 -18652 14020 -18114
rect 13623 -20288 14020 -19750
rect 13624 -21924 14021 -21386
rect 13623 -24378 14020 -23840
rect 13624 -25196 14021 -24658
rect 13624 -27650 14021 -27112
rect 13624 -30104 14021 -29566
<< metal1 >>
rect 16884 -14112 26584 -11602
rect 16884 -14932 20666 -14112
rect 20724 -14176 21428 -14170
rect 20724 -14868 20730 -14176
rect 21422 -14868 21428 -14176
rect 20724 -14874 21428 -14868
rect 21484 -14932 26584 -14112
rect 16884 -15468 26584 -14932
rect 16884 -16150 25886 -15468
rect 26562 -16150 26584 -15468
rect 16884 -16762 26584 -16150
rect 6882 -17296 7291 -17284
rect 6882 -17834 6888 -17296
rect 7285 -17834 7291 -17296
rect 6882 -17846 7291 -17834
rect 13617 -17296 14026 -17284
rect 13617 -17834 13623 -17296
rect 14020 -17834 14026 -17296
rect 16884 -17444 25894 -16762
rect 26570 -17444 26584 -16762
rect 16884 -17446 26584 -17444
rect 13617 -17846 14026 -17834
rect 13606 -18048 14304 -18042
rect 6070 -18104 6640 -18098
rect 6070 -18662 6076 -18104
rect 6634 -18662 6640 -18104
rect 5270 -19740 5840 -19728
rect 5270 -20298 5276 -19740
rect 5834 -20298 5840 -19740
rect 5270 -22194 5840 -20298
rect 6070 -20558 6640 -18662
rect 6870 -18104 7302 -18098
rect 6870 -18662 6876 -18104
rect 7296 -18662 7302 -18104
rect 6870 -18668 7302 -18662
rect 13606 -18740 13612 -18048
rect 13606 -18746 14304 -18740
rect 13606 -18866 21430 -18860
rect 6870 -18922 7302 -18916
rect 6870 -19480 6876 -18922
rect 7296 -19480 7302 -18922
rect 6870 -19486 7302 -19480
rect 7532 -18922 8102 -18916
rect 7532 -19480 7538 -18922
rect 8096 -19480 8102 -18922
rect 6870 -19740 7302 -19734
rect 6870 -20298 6876 -19740
rect 7296 -20298 7302 -19740
rect 6870 -20304 7302 -20298
rect 6070 -21116 6076 -20558
rect 6634 -21116 6640 -20558
rect 6070 -21236 6640 -21116
rect 6870 -20558 7302 -20552
rect 6870 -21116 6876 -20558
rect 7296 -21116 7302 -20558
rect 6870 -21122 7302 -21116
rect 6870 -21376 7302 -21370
rect 6870 -21934 6876 -21376
rect 7296 -21934 7302 -21376
rect 6870 -21940 7302 -21934
rect 7532 -21376 8102 -19480
rect 13606 -19558 13612 -18866
rect 14304 -19558 20730 -18866
rect 21422 -19558 21430 -18866
rect 13606 -19564 21430 -19558
rect 13606 -19684 14310 -19678
rect 13606 -20376 13612 -19684
rect 14304 -20376 14310 -19684
rect 16680 -19966 26582 -19960
rect 13606 -20382 14310 -20376
rect 7532 -21934 7538 -21376
rect 8096 -21934 8102 -21376
rect 7532 -21940 8102 -21934
rect 12006 -20558 12576 -20552
rect 12006 -21116 12012 -20558
rect 12570 -21116 12576 -20558
rect 5270 -22752 5276 -22194
rect 5834 -22752 5840 -22194
rect 5270 -22926 5840 -22752
rect 6870 -22194 7302 -22188
rect 6870 -22752 6876 -22194
rect 7296 -22752 7302 -22194
rect 6870 -22758 7302 -22752
rect 6070 -23012 6640 -23006
rect 6070 -23570 6076 -23012
rect 6634 -23570 6640 -23012
rect 6070 -25466 6640 -23570
rect 6870 -23012 7302 -23006
rect 6870 -23570 6876 -23012
rect 7296 -23570 7302 -23012
rect 12006 -23012 12576 -21116
rect 13606 -20558 14038 -20552
rect 13606 -21116 13612 -20558
rect 14032 -21116 14038 -20558
rect 16680 -20902 25640 -19966
rect 26576 -20902 26582 -19966
rect 16680 -20908 26582 -20902
rect 13606 -21122 14038 -21116
rect 13606 -21376 14038 -21370
rect 13606 -21934 13612 -21376
rect 14032 -21934 14038 -21376
rect 13606 -21940 14038 -21934
rect 14268 -21376 14838 -21370
rect 14268 -21934 14274 -21376
rect 14832 -21934 14838 -21376
rect 12006 -23570 12012 -23012
rect 12570 -23570 12576 -23012
rect 12806 -22194 13376 -22188
rect 12806 -22752 12812 -22194
rect 13370 -22752 13376 -22194
rect 6870 -23576 7302 -23570
rect 6870 -23830 7302 -23824
rect 6870 -24388 6876 -23830
rect 7296 -24388 7302 -23830
rect 6870 -24394 7302 -24388
rect 6870 -24648 7302 -24642
rect 6870 -25206 6876 -24648
rect 7296 -25206 7302 -24648
rect 6870 -25212 7302 -25206
rect 7532 -24648 8102 -24642
rect 7532 -25206 7538 -24648
rect 8096 -25206 8102 -24648
rect 6070 -26024 6076 -25466
rect 6634 -26024 6640 -25466
rect 6070 -26152 6640 -26024
rect 6870 -25466 7302 -25460
rect 6870 -26024 6876 -25466
rect 7296 -26024 7302 -25466
rect 6870 -26030 7302 -26024
rect 5270 -26284 5840 -26278
rect 5270 -26842 5276 -26284
rect 5834 -26842 5840 -26284
rect 5270 -27908 5840 -26842
rect 6870 -26284 7302 -26278
rect 6870 -26842 6876 -26284
rect 7296 -26842 7302 -26284
rect 6870 -26848 7302 -26842
rect 6870 -27102 7302 -27096
rect 6870 -27660 6876 -27102
rect 7296 -27660 7302 -27102
rect 6870 -27666 7302 -27660
rect 7532 -27102 8102 -25206
rect 7532 -27660 7538 -27102
rect 8096 -27660 8102 -27102
rect 7532 -27666 8102 -27660
rect 12006 -25466 12576 -25460
rect 12006 -26024 12012 -25466
rect 12570 -26024 12576 -25466
rect 5270 -28466 5276 -27908
rect 5834 -28466 5840 -27908
rect 5270 -28472 5840 -28466
rect 6870 -27920 7302 -27914
rect 6870 -28478 6876 -27920
rect 7296 -28478 7302 -27920
rect 6870 -28484 7302 -28478
rect 6070 -28738 6640 -28732
rect 6070 -29296 6076 -28738
rect 6634 -29296 6640 -28738
rect 6070 -34336 6640 -29296
rect 6870 -28738 7302 -28732
rect 6870 -29296 6876 -28738
rect 7296 -29296 7302 -28738
rect 6870 -29302 7302 -29296
rect 12006 -28738 12576 -26024
rect 12806 -26284 13376 -22752
rect 13606 -22194 14038 -22188
rect 13606 -22752 13612 -22194
rect 14032 -22752 14038 -22194
rect 13606 -22758 14038 -22752
rect 13606 -23012 14038 -23006
rect 13606 -23570 13612 -23012
rect 14032 -23570 14038 -23012
rect 13606 -23576 14038 -23570
rect 13606 -23774 14162 -23768
rect 13606 -23830 13644 -23774
rect 13606 -24388 13612 -23830
rect 13606 -24466 13644 -24388
rect 13606 -24472 14162 -24466
rect 13606 -24648 14038 -24642
rect 13606 -25206 13612 -24648
rect 14032 -25206 14038 -24648
rect 13606 -25212 14038 -25206
rect 14268 -24648 14838 -21934
rect 14268 -25206 14274 -24648
rect 14832 -25206 14838 -24648
rect 14268 -25212 14838 -25206
rect 13606 -25466 14038 -25460
rect 13606 -26024 13612 -25466
rect 14032 -26024 14038 -25466
rect 13606 -26030 14038 -26024
rect 12806 -26842 12812 -26284
rect 13370 -26842 13376 -26284
rect 12806 -26848 13376 -26842
rect 13606 -26284 14038 -26278
rect 13606 -26842 13612 -26284
rect 14032 -26842 14038 -26284
rect 13606 -26848 14038 -26842
rect 13606 -27102 14038 -27096
rect 13606 -27660 13612 -27102
rect 14032 -27660 14038 -27102
rect 13606 -27666 14038 -27660
rect 14268 -27102 14838 -27096
rect 14268 -27660 14274 -27102
rect 14832 -27660 14838 -27102
rect 12006 -29296 12012 -28738
rect 12570 -29296 12576 -28738
rect 12006 -29302 12576 -29296
rect 12806 -27920 13376 -27914
rect 12806 -28478 12812 -27920
rect 13370 -28478 13376 -27920
rect 6870 -29556 7302 -29550
rect 6870 -30114 6876 -29556
rect 7296 -30114 7302 -29556
rect 6870 -30120 7302 -30114
rect 7532 -29556 8102 -29550
rect 7532 -30114 7538 -29556
rect 8096 -30114 8102 -29556
rect 7532 -33638 8102 -30114
rect 6808 -34210 8102 -33638
rect 6068 -34458 6640 -34336
rect 6068 -35028 7240 -34458
rect 11961 -37742 12370 -37740
rect 12806 -37742 13376 -28478
rect 13606 -27920 14038 -27914
rect 13606 -28478 13612 -27920
rect 14032 -28478 14038 -27920
rect 13606 -28484 14038 -28478
rect 13606 -28738 14038 -28732
rect 13606 -29296 13612 -28738
rect 14032 -29296 14038 -28738
rect 13606 -29302 14038 -29296
rect 13606 -29556 14038 -29550
rect 13606 -30114 13612 -29556
rect 14032 -30114 14038 -29556
rect 13606 -30120 14038 -30114
rect 14268 -29556 14838 -27660
rect 14268 -30114 14274 -29556
rect 14832 -30114 14838 -29556
rect 14268 -30120 14838 -30114
rect 11961 -37746 13376 -37742
rect 11961 -38284 11967 -37746
rect 12364 -38284 13376 -37746
rect 11961 -38290 13376 -38284
<< via1 >>
rect 20730 -14868 21422 -14176
rect 25886 -16150 26562 -15468
rect 25894 -17444 26570 -16762
rect 6076 -18662 6634 -18104
rect 5276 -20298 5834 -19740
rect 6876 -18662 7296 -18104
rect 13612 -18114 14304 -18048
rect 13612 -18652 13623 -18114
rect 13623 -18652 14020 -18114
rect 14020 -18652 14304 -18114
rect 13612 -18740 14304 -18652
rect 6876 -19480 7296 -18922
rect 7538 -19480 8096 -18922
rect 6876 -20298 7296 -19740
rect 6076 -21116 6634 -20558
rect 6876 -21116 7296 -20558
rect 6876 -21934 7296 -21376
rect 13612 -19558 14304 -18866
rect 20730 -19558 21422 -18866
rect 13612 -19750 14304 -19684
rect 13612 -20288 13623 -19750
rect 13623 -20288 14020 -19750
rect 14020 -20288 14304 -19750
rect 13612 -20376 14304 -20288
rect 7538 -21934 8096 -21376
rect 12012 -21116 12570 -20558
rect 5276 -22752 5834 -22194
rect 6876 -22752 7296 -22194
rect 6076 -23570 6634 -23012
rect 6876 -23570 7296 -23012
rect 13612 -21116 14032 -20558
rect 16162 -20900 16680 -19966
rect 25640 -20902 26576 -19966
rect 13612 -21386 14032 -21376
rect 13612 -21924 13624 -21386
rect 13624 -21924 14021 -21386
rect 14021 -21924 14032 -21386
rect 13612 -21934 14032 -21924
rect 14274 -21934 14832 -21376
rect 12012 -23570 12570 -23012
rect 12812 -22752 13370 -22194
rect 6876 -24388 7296 -23830
rect 6876 -25206 7296 -24648
rect 7538 -25206 8096 -24648
rect 6076 -26024 6634 -25466
rect 6876 -26024 7296 -25466
rect 5276 -26842 5834 -26284
rect 6876 -26842 7296 -26284
rect 6876 -27660 7296 -27102
rect 7538 -27660 8096 -27102
rect 12012 -26024 12570 -25466
rect 5276 -28466 5834 -27908
rect 6876 -28478 7296 -27920
rect 6076 -29296 6634 -28738
rect 6876 -29296 7296 -28738
rect 13612 -22752 14032 -22194
rect 13612 -23570 14032 -23012
rect 13644 -23830 14162 -23774
rect 13612 -23840 14162 -23830
rect 13612 -24378 13623 -23840
rect 13623 -24378 14020 -23840
rect 14020 -24378 14162 -23840
rect 13612 -24388 14162 -24378
rect 13644 -24466 14162 -24388
rect 13612 -24658 14032 -24648
rect 13612 -25196 13624 -24658
rect 13624 -25196 14021 -24658
rect 14021 -25196 14032 -24658
rect 13612 -25206 14032 -25196
rect 14274 -25206 14832 -24648
rect 13612 -26024 14032 -25466
rect 12812 -26842 13370 -26284
rect 13612 -26842 14032 -26284
rect 13612 -27112 14032 -27102
rect 13612 -27650 13624 -27112
rect 13624 -27650 14021 -27112
rect 14021 -27650 14032 -27112
rect 13612 -27660 14032 -27650
rect 14274 -27660 14832 -27102
rect 12012 -29296 12570 -28738
rect 12812 -28478 13370 -27920
rect 6876 -30114 7296 -29556
rect 7538 -30114 8096 -29556
rect 13612 -28478 14032 -27920
rect 13612 -29296 14032 -28738
rect 13612 -29566 14032 -29556
rect 13612 -30104 13624 -29566
rect 13624 -30104 14021 -29566
rect 14021 -30104 14032 -29566
rect 13612 -30114 14032 -30104
rect 14274 -30114 14832 -29556
<< metal2 >>
rect 20724 -14176 21428 -14170
rect 20724 -14868 20730 -14176
rect 21422 -14868 21428 -14176
rect 13606 -18048 14310 -18042
rect 6070 -18104 7302 -18098
rect 6070 -18662 6076 -18104
rect 6634 -18662 6876 -18104
rect 7296 -18662 7302 -18104
rect 13606 -18110 13612 -18048
rect 6070 -18668 7302 -18662
rect 9732 -18680 13612 -18110
rect 6870 -18922 8102 -18916
rect 6870 -19480 6876 -18922
rect 7296 -19480 7538 -18922
rect 8096 -19480 8102 -18922
rect 6870 -19486 8102 -19480
rect 5270 -19740 7302 -19734
rect 5270 -20298 5276 -19740
rect 5834 -20298 6876 -19740
rect 7296 -20298 7302 -19740
rect 5840 -20304 7302 -20298
rect 6070 -20558 7302 -20552
rect 6070 -21116 6076 -20558
rect 6634 -21116 6876 -20558
rect 7296 -21116 7302 -20558
rect 6070 -21122 7302 -21116
rect 6870 -21376 8102 -21370
rect 6870 -21934 6876 -21376
rect 7296 -21934 7538 -21376
rect 8096 -21934 8102 -21376
rect 6870 -21940 8102 -21934
rect 5270 -22194 7302 -22188
rect 5270 -22752 5276 -22194
rect 5834 -22752 6876 -22194
rect 7296 -22752 7302 -22194
rect 5270 -22758 7302 -22752
rect 6070 -23012 7302 -23006
rect 6070 -23570 6076 -23012
rect 6634 -23570 6876 -23012
rect 7296 -23570 7302 -23012
rect 6070 -23576 7302 -23570
rect 9732 -23824 10302 -18680
rect 13606 -18740 13612 -18680
rect 14304 -18740 14310 -18048
rect 13606 -18746 14310 -18740
rect 13606 -18866 14304 -18860
rect 13606 -19558 13612 -18866
rect 13606 -19564 14304 -19558
rect 20724 -18866 21428 -14868
rect 20724 -19558 20730 -18866
rect 21422 -19558 21428 -18866
rect 20724 -19564 21428 -19558
rect 25634 -15468 26582 -15418
rect 25634 -16150 25886 -15468
rect 26562 -16150 26582 -15468
rect 25634 -16762 26582 -16150
rect 25634 -17444 25894 -16762
rect 26570 -17444 26582 -16762
rect 13606 -19684 14310 -19678
rect 13606 -20376 13612 -19684
rect 14304 -20376 14310 -19684
rect 25634 -19966 26582 -17444
rect 13606 -20382 14310 -20376
rect 12006 -20558 14038 -20552
rect 12006 -21116 12012 -20558
rect 12570 -21116 13612 -20558
rect 14032 -21116 14038 -20558
rect 12006 -21122 14038 -21116
rect 13606 -21376 14838 -21370
rect 13606 -21934 13612 -21376
rect 14032 -21934 14274 -21376
rect 14832 -21934 14838 -21376
rect 13606 -21940 14838 -21934
rect 12806 -22194 14038 -22188
rect 12806 -22752 12812 -22194
rect 13370 -22752 13612 -22194
rect 14032 -22752 14038 -22194
rect 12806 -22758 14038 -22752
rect 12006 -23012 14038 -23006
rect 12006 -23570 12012 -23012
rect 12570 -23570 13612 -23012
rect 14032 -23570 14038 -23012
rect 12006 -23576 14038 -23570
rect 13644 -23770 14910 -23768
rect 16156 -23770 16686 -20900
rect 25634 -20902 25640 -19966
rect 26576 -20902 26582 -19966
rect 25634 -20908 26582 -20902
rect 13644 -23774 16686 -23770
rect 6870 -23830 10302 -23824
rect 6870 -24388 6876 -23830
rect 7296 -24388 10302 -23830
rect 6870 -24394 10302 -24388
rect 13606 -23830 13644 -23824
rect 13606 -24388 13612 -23830
rect 13606 -24394 13644 -24388
rect 14162 -24466 16686 -23774
rect 13644 -24472 16686 -24466
rect 6870 -24648 8102 -24642
rect 6870 -25206 6876 -24648
rect 7296 -25206 7538 -24648
rect 8096 -25206 8102 -24648
rect 6870 -25212 8102 -25206
rect 13606 -24648 14832 -24642
rect 13606 -25206 13612 -24648
rect 14032 -25206 14274 -24648
rect 14832 -25206 14838 -24648
rect 13606 -25212 14838 -25206
rect 6070 -25466 7302 -25460
rect 6070 -26024 6076 -25466
rect 6634 -26024 6876 -25466
rect 7296 -26024 7302 -25466
rect 6070 -26030 7302 -26024
rect 12006 -25466 14038 -25460
rect 12006 -26024 12012 -25466
rect 12570 -26024 13612 -25466
rect 14032 -26024 14038 -25466
rect 12006 -26030 14038 -26024
rect 5270 -26284 7302 -26278
rect 5270 -26842 5276 -26284
rect 5834 -26842 6876 -26284
rect 7296 -26842 7302 -26284
rect 5270 -26848 7302 -26842
rect 12806 -26284 14038 -26278
rect 12806 -26842 12812 -26284
rect 13370 -26842 13612 -26284
rect 14032 -26842 14038 -26284
rect 12806 -26848 14038 -26842
rect 6870 -27102 8102 -27096
rect 6870 -27660 6876 -27102
rect 7296 -27660 7538 -27102
rect 8096 -27660 8102 -27102
rect 6870 -27666 8102 -27660
rect 13606 -27102 14832 -27096
rect 13606 -27660 13612 -27102
rect 14032 -27660 14274 -27102
rect 14832 -27660 14838 -27102
rect 13606 -27666 14838 -27660
rect 5270 -27908 7284 -27902
rect 5270 -28466 5276 -27908
rect 5834 -27914 7284 -27908
rect 5834 -27920 7302 -27914
rect 5834 -28466 6876 -27920
rect 5270 -28472 6876 -28466
rect 6870 -28478 6876 -28472
rect 7296 -28478 7302 -27920
rect 6870 -28484 7302 -28478
rect 12806 -27920 14038 -27914
rect 12806 -28478 12812 -27920
rect 13370 -28478 13612 -27920
rect 14032 -28478 14038 -27920
rect 12806 -28484 14038 -28478
rect 6070 -28738 7302 -28732
rect 6070 -29296 6076 -28738
rect 6634 -29296 6876 -28738
rect 7296 -29296 7302 -28738
rect 6070 -29302 7302 -29296
rect 12006 -28738 14038 -28732
rect 12006 -29296 12012 -28738
rect 12570 -29296 13612 -28738
rect 14032 -29296 14038 -28738
rect 12006 -29302 14038 -29296
rect 6870 -29556 8102 -29550
rect 6870 -30114 6876 -29556
rect 7296 -30114 7538 -29556
rect 8096 -30114 8102 -29556
rect 6870 -30120 8102 -30114
rect 13606 -29556 14832 -29550
rect 13606 -30114 13612 -29556
rect 14032 -30114 14274 -29556
rect 14832 -30114 14838 -29556
rect 13606 -30120 14838 -30114
use sky130_fd_pr__res_xhigh_po_2p85_EDZVPS  sky130_fd_pr__res_xhigh_po_2p85_EDZVPS_0
timestamp 1621208350
transform 0 1 10454 1 0 -24109
box -6831 -3584 6831 3584
use sky130_fd_pr__res_xhigh_po_2p85_R3CJ3X  sky130_fd_pr__res_xhigh_po_2p85_R3CJ3X_0
timestamp 1621223045
transform 0 -1 10288 -1 0 -38015
box -1105 -2094 1105 2094
use sky130_fd_pr__res_xhigh_po_2p85_W28W8W  sky130_fd_pr__res_xhigh_po_2p85_W28W8W_0
timestamp 1621223045
transform 0 -1 9390 -1 0 -34334
box -1514 -2582 1514 2582
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1288 0 7 1288
timestamp 1620883575
transform 0 1 16542 -1 0 -11276
box 26 26 1314 1314
<< labels >>
flabel metal2 25634 -18580 26582 -17444 5 FreeSans 1600 0 0 0 Vbneg
flabel locali 11698 -34850 11988 -33746 7 FreeSans 800 90 0 0 GND!
port 4 n
flabel metal2 6870 -29302 7302 -28732 7 FreeSans 800 90 0 0 VbEnd
flabel metal2 13606 -28484 14038 -27914 7 FreeSans 800 90 0 0 VbgEnd
flabel metal2 6870 -30120 8102 -29550 7 FreeSans 800 90 0 0 VaEnd
flabel metal2 13612 -20376 14304 -19684 7 FreeSans 1600 90 0 0 Vbg
port 3 n
flabel metal2 13606 -18746 14310 -18042 7 FreeSans 1600 90 0 0 Vb
port 1 n
flabel metal1 14304 -19564 14876 -18860 1 FreeSans 1600 0 0 0 Va
port 5 n
<< end >>
