magic
tech sky130A
magscale 1 2
timestamp 1621617037
<< psubdiff >>
rect -960 670 2860 694
rect -960 594 454 670
rect 1446 594 2860 670
rect -960 570 2860 594
rect -956 516 -508 570
rect -956 -60 -932 516
rect -532 -60 -508 516
rect 2410 516 2858 570
rect -956 -84 -508 -60
rect 2410 -60 2434 516
rect 2834 -60 2858 516
rect 2410 -84 2858 -60
<< psubdiffcont >>
rect 454 594 1446 670
rect -932 -60 -532 516
rect 2434 -60 2834 516
<< poly >>
rect 1438 404 1762 438
<< locali >>
rect 438 670 1462 686
rect 438 594 454 670
rect 1446 594 1462 670
rect 438 554 1462 594
rect -948 516 -516 532
rect -948 -60 -932 516
rect -532 438 -516 516
rect 438 502 466 554
rect 518 502 1382 554
rect 1434 502 1462 554
rect 438 490 1462 502
rect 2418 516 2850 532
rect 2418 438 2434 516
rect -532 404 -378 438
rect 464 404 522 438
rect 922 404 980 438
rect 1380 404 1438 438
rect 2280 404 2434 438
rect -532 -38 -406 404
rect 2308 -38 2434 404
rect -532 -60 -516 -38
rect -948 -76 -516 -60
rect 2418 -60 2434 -38
rect 2834 -60 2850 516
rect 2418 -76 2850 -60
<< viali >>
rect 466 502 518 554
rect 1382 502 1434 554
<< metal1 >>
rect 454 554 530 566
rect 454 502 466 554
rect 518 502 530 554
rect 454 490 530 502
rect 1370 554 1446 566
rect 1370 502 1382 554
rect 1434 502 1446 554
rect 1370 490 1446 502
rect 148 438 380 450
rect 12 404 380 438
rect 12 366 56 404
rect 148 386 380 404
rect 12 -164 58 366
rect 470 -22 516 490
rect 2 -170 66 -164
rect 2 -222 8 -170
rect 60 -222 66 -170
rect 2 -228 66 -222
rect 928 -370 974 366
rect 1386 -22 1432 490
rect 1512 438 1744 450
rect 1512 404 1890 438
rect 1512 386 1744 404
rect 1844 -158 1890 404
rect 1836 -164 1900 -158
rect 1836 -216 1842 -164
rect 1894 -216 1900 -164
rect 1836 -222 1900 -216
rect 920 -376 984 -370
rect 920 -428 926 -376
rect 978 -428 984 -376
rect 920 -434 984 -428
<< via1 >>
rect 8 -222 60 -170
rect 1842 -216 1894 -164
rect 926 -428 978 -376
<< metal2 >>
rect 2 -164 1900 -158
rect 2 -170 1842 -164
rect 2 -222 8 -170
rect 60 -216 1842 -170
rect 1894 -216 1900 -164
rect 60 -222 1900 -216
rect 2 -228 1900 -222
rect 60 -376 1842 -368
rect 60 -428 926 -376
rect 978 -428 1842 -376
rect 60 -438 1842 -428
use sky130_fd_pr__nfet_01v8_lvt_NHDRMS  sky130_fd_pr__nfet_01v8_lvt_NHDRMS_0
timestamp 1621616995
transform 1 0 951 0 1 197
box -1403 -257 1403 257
<< labels >>
flabel metal2 60 -438 1842 -368 1 FreeSans 800 0 0 0 Vq
port 2 n
flabel metal2 60 -228 1842 -158 1 FreeSans 800 0 0 0 Vx
port 1 n
flabel locali 920 532 1002 560 1 FreeSans 800 0 0 0 GND!
port 3 n
<< end >>
