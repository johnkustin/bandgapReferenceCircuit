magic
tech sky130A
magscale 1 2
timestamp 1622139266
<< nwell >>
rect 312604 625006 329982 625008
rect 302804 616506 312332 619848
rect 312604 617108 330870 625006
rect 312604 617106 318524 617108
rect 319314 617106 324024 617108
rect 324814 617106 330870 617108
<< pwell >>
rect 334648 627639 341088 627740
rect 334648 626553 334749 627639
rect 335835 626553 336037 627639
rect 337123 626553 337325 627639
rect 338411 626553 338613 627639
rect 339699 626553 339901 627639
rect 340987 626553 341088 627639
rect 334648 626351 341088 626553
rect 334648 625265 334749 626351
rect 335835 625265 336037 626351
rect 337123 625265 337325 626351
rect 338411 625265 338613 626351
rect 339699 625265 339901 626351
rect 340987 625265 341088 626351
rect 334648 625063 341088 625265
rect 334648 623977 334749 625063
rect 335835 623977 336037 625063
rect 337123 623977 337325 625063
rect 338411 623977 338613 625063
rect 339699 623977 339901 625063
rect 340987 623977 341088 625063
rect 334648 623775 341088 623977
rect 334648 622689 334749 623775
rect 335835 622689 336037 623775
rect 337123 622689 337325 623775
rect 338411 622689 338613 623775
rect 339699 622689 339901 623775
rect 340987 622689 341088 623775
rect 334648 622487 341088 622689
rect 334648 621401 334749 622487
rect 335835 621401 336037 622487
rect 337123 621401 337325 622487
rect 338411 621401 338613 622487
rect 339699 621401 339901 622487
rect 340987 621401 341088 622487
rect 334648 621199 341088 621401
rect 334648 620113 334749 621199
rect 335835 620113 336037 621199
rect 337123 620113 337325 621199
rect 338411 620113 338613 621199
rect 339699 620113 339901 621199
rect 340987 620113 341088 621199
rect 334648 619911 341088 620113
rect 334648 618825 334749 619911
rect 335835 618825 336037 619911
rect 337123 618825 337325 619911
rect 338411 618825 338613 619911
rect 339699 618825 339901 619911
rect 340987 618825 341088 619911
rect 334648 618623 341088 618825
rect 334648 617537 334749 618623
rect 335835 617537 336037 618623
rect 337123 617537 337325 618623
rect 338411 617537 338613 618623
rect 339699 617537 339901 618623
rect 340987 617537 341088 618623
rect 334648 617436 341088 617537
<< nbase >>
rect 334775 626579 335809 627613
rect 336063 626579 337097 627613
rect 337351 626579 338385 627613
rect 338639 626579 339673 627613
rect 339927 626579 340961 627613
rect 334775 625291 335809 626325
rect 336063 625291 337097 626325
rect 337351 625291 338385 626325
rect 338639 625291 339673 626325
rect 339927 625291 340961 626325
rect 334775 624003 335809 625037
rect 336063 624003 337097 625037
rect 337351 624003 338385 625037
rect 338639 624003 339673 625037
rect 339927 624003 340961 625037
rect 334775 622715 335809 623749
rect 336063 622715 337097 623749
rect 337351 622715 338385 623749
rect 338639 622715 339673 623749
rect 339927 622715 340961 623749
rect 334775 621427 335809 622461
rect 336063 621427 337097 622461
rect 337351 621427 338385 622461
rect 338639 621427 339673 622461
rect 339927 621427 340961 622461
rect 334775 620139 335809 621173
rect 336063 620139 337097 621173
rect 337351 620139 338385 621173
rect 338639 620139 339673 621173
rect 339927 620139 340961 621173
rect 334775 618851 335809 619885
rect 336063 618851 337097 619885
rect 337351 618851 338385 619885
rect 338639 618851 339673 619885
rect 339927 618851 340961 619885
rect 334775 617563 335809 618597
rect 336063 617563 337097 618597
rect 337351 617563 338385 618597
rect 338639 617563 339673 618597
rect 339927 617563 340961 618597
<< pmoslvt >>
rect 303642 617168 304042 619748
rect 304214 617168 304614 619748
rect 304786 617168 305186 619748
rect 305358 617168 305758 619748
rect 305930 617168 306330 619748
rect 306502 617168 306902 619748
rect 307074 617168 307474 619748
rect 307646 617168 308046 619748
rect 308218 617168 308618 619748
rect 308790 617168 309190 619748
rect 309362 617168 309762 619748
rect 309934 617168 310334 619748
rect 310506 617168 310906 619748
rect 311078 617168 311478 619748
rect 313450 617206 313850 624946
rect 313908 617206 314308 624946
rect 314366 617206 314766 624946
rect 314824 617206 315224 624946
rect 315282 617206 315682 624946
rect 315740 617206 316140 624946
rect 316198 617206 316598 624946
rect 316656 617206 317056 624946
rect 317114 617206 317514 624946
rect 317572 617206 317972 624946
rect 318030 617206 318430 624946
rect 319408 617206 319808 624946
rect 319866 617206 320266 624946
rect 320324 617206 320724 624946
rect 320782 617206 321182 624946
rect 321240 617206 321640 624946
rect 321698 617206 322098 624946
rect 322156 617206 322556 624946
rect 322614 617206 323014 624946
rect 323072 617206 323472 624946
rect 323530 617206 323930 624946
rect 324908 617206 325308 624946
rect 325366 617206 325766 624946
rect 325824 617206 326224 624946
rect 326282 617206 326682 624946
rect 326740 617206 327140 624946
rect 327198 617206 327598 624946
rect 327656 617206 328056 624946
rect 328114 617206 328514 624946
rect 328572 617206 328972 624946
rect 329030 617206 329430 624946
rect 329488 617206 329888 624946
<< nmoslvt >>
rect 305028 623912 310428 624312
rect 300438 620638 300838 621038
rect 300896 620638 301296 621038
rect 301354 620638 301754 621038
rect 301812 620638 302212 621038
rect 302270 620638 302670 621038
rect 302728 620638 303128 621038
rect 305368 620360 305768 622160
rect 305940 620360 306340 622160
rect 306512 620360 306912 622160
rect 307084 620360 307484 622160
rect 307656 620360 308056 622160
rect 308228 620360 308628 622160
rect 308800 620360 309200 622160
rect 309372 620360 309772 622160
<< ndiff >>
rect 305028 624358 310428 624370
rect 305028 624324 305040 624358
rect 310416 624324 310428 624358
rect 305028 624312 310428 624324
rect 305028 623900 310428 623912
rect 305028 623866 305040 623900
rect 310416 623866 310428 623900
rect 305028 623854 310428 623866
rect 300380 621026 300438 621038
rect 300380 620650 300392 621026
rect 300426 620650 300438 621026
rect 300380 620638 300438 620650
rect 300838 621026 300896 621038
rect 300838 620650 300850 621026
rect 300884 620650 300896 621026
rect 300838 620638 300896 620650
rect 301296 621026 301354 621038
rect 301296 620650 301308 621026
rect 301342 620650 301354 621026
rect 301296 620638 301354 620650
rect 301754 621026 301812 621038
rect 301754 620650 301766 621026
rect 301800 620650 301812 621026
rect 301754 620638 301812 620650
rect 302212 621026 302270 621038
rect 302212 620650 302224 621026
rect 302258 620650 302270 621026
rect 302212 620638 302270 620650
rect 302670 621026 302728 621038
rect 302670 620650 302682 621026
rect 302716 620650 302728 621026
rect 302670 620638 302728 620650
rect 303128 621026 303186 621038
rect 303128 620650 303140 621026
rect 303174 620650 303186 621026
rect 303128 620638 303186 620650
rect 305310 622148 305368 622160
rect 305310 620372 305322 622148
rect 305356 620372 305368 622148
rect 305310 620360 305368 620372
rect 305768 622148 305826 622160
rect 305768 620372 305780 622148
rect 305814 620372 305826 622148
rect 305768 620360 305826 620372
rect 305882 622148 305940 622160
rect 305882 620372 305894 622148
rect 305928 620372 305940 622148
rect 305882 620360 305940 620372
rect 306340 622148 306398 622160
rect 306340 620372 306352 622148
rect 306386 620372 306398 622148
rect 306340 620360 306398 620372
rect 306454 622148 306512 622160
rect 306454 620372 306466 622148
rect 306500 620372 306512 622148
rect 306454 620360 306512 620372
rect 306912 622148 306970 622160
rect 306912 620372 306924 622148
rect 306958 620372 306970 622148
rect 306912 620360 306970 620372
rect 307026 622148 307084 622160
rect 307026 620372 307038 622148
rect 307072 620372 307084 622148
rect 307026 620360 307084 620372
rect 307484 622148 307542 622160
rect 307484 620372 307496 622148
rect 307530 620372 307542 622148
rect 307484 620360 307542 620372
rect 307598 622148 307656 622160
rect 307598 620372 307610 622148
rect 307644 620372 307656 622148
rect 307598 620360 307656 620372
rect 308056 622148 308114 622160
rect 308056 620372 308068 622148
rect 308102 620372 308114 622148
rect 308056 620360 308114 620372
rect 308170 622148 308228 622160
rect 308170 620372 308182 622148
rect 308216 620372 308228 622148
rect 308170 620360 308228 620372
rect 308628 622148 308686 622160
rect 308628 620372 308640 622148
rect 308674 620372 308686 622148
rect 308628 620360 308686 620372
rect 308742 622148 308800 622160
rect 308742 620372 308754 622148
rect 308788 620372 308800 622148
rect 308742 620360 308800 620372
rect 309200 622148 309258 622160
rect 309200 620372 309212 622148
rect 309246 620372 309258 622148
rect 309200 620360 309258 620372
rect 309314 622148 309372 622160
rect 309314 620372 309326 622148
rect 309360 620372 309372 622148
rect 309314 620360 309372 620372
rect 309772 622148 309830 622160
rect 309772 620372 309784 622148
rect 309818 620372 309830 622148
rect 309772 620360 309830 620372
<< pdiff >>
rect 334952 627382 335632 627436
rect 334952 627348 335004 627382
rect 335038 627348 335094 627382
rect 335128 627348 335184 627382
rect 335218 627348 335274 627382
rect 335308 627348 335364 627382
rect 335398 627348 335454 627382
rect 335488 627348 335544 627382
rect 335578 627348 335632 627382
rect 334952 627292 335632 627348
rect 334952 627258 335004 627292
rect 335038 627258 335094 627292
rect 335128 627258 335184 627292
rect 335218 627258 335274 627292
rect 335308 627258 335364 627292
rect 335398 627258 335454 627292
rect 335488 627258 335544 627292
rect 335578 627258 335632 627292
rect 334952 627202 335632 627258
rect 334952 627168 335004 627202
rect 335038 627168 335094 627202
rect 335128 627168 335184 627202
rect 335218 627168 335274 627202
rect 335308 627168 335364 627202
rect 335398 627168 335454 627202
rect 335488 627168 335544 627202
rect 335578 627168 335632 627202
rect 334952 627112 335632 627168
rect 334952 627078 335004 627112
rect 335038 627078 335094 627112
rect 335128 627078 335184 627112
rect 335218 627078 335274 627112
rect 335308 627078 335364 627112
rect 335398 627078 335454 627112
rect 335488 627078 335544 627112
rect 335578 627078 335632 627112
rect 334952 627022 335632 627078
rect 334952 626988 335004 627022
rect 335038 626988 335094 627022
rect 335128 626988 335184 627022
rect 335218 626988 335274 627022
rect 335308 626988 335364 627022
rect 335398 626988 335454 627022
rect 335488 626988 335544 627022
rect 335578 626988 335632 627022
rect 334952 626932 335632 626988
rect 334952 626898 335004 626932
rect 335038 626898 335094 626932
rect 335128 626898 335184 626932
rect 335218 626898 335274 626932
rect 335308 626898 335364 626932
rect 335398 626898 335454 626932
rect 335488 626898 335544 626932
rect 335578 626898 335632 626932
rect 334952 626842 335632 626898
rect 334952 626808 335004 626842
rect 335038 626808 335094 626842
rect 335128 626808 335184 626842
rect 335218 626808 335274 626842
rect 335308 626808 335364 626842
rect 335398 626808 335454 626842
rect 335488 626808 335544 626842
rect 335578 626808 335632 626842
rect 334952 626756 335632 626808
rect 336240 627382 336920 627436
rect 336240 627348 336292 627382
rect 336326 627348 336382 627382
rect 336416 627348 336472 627382
rect 336506 627348 336562 627382
rect 336596 627348 336652 627382
rect 336686 627348 336742 627382
rect 336776 627348 336832 627382
rect 336866 627348 336920 627382
rect 336240 627292 336920 627348
rect 336240 627258 336292 627292
rect 336326 627258 336382 627292
rect 336416 627258 336472 627292
rect 336506 627258 336562 627292
rect 336596 627258 336652 627292
rect 336686 627258 336742 627292
rect 336776 627258 336832 627292
rect 336866 627258 336920 627292
rect 336240 627202 336920 627258
rect 336240 627168 336292 627202
rect 336326 627168 336382 627202
rect 336416 627168 336472 627202
rect 336506 627168 336562 627202
rect 336596 627168 336652 627202
rect 336686 627168 336742 627202
rect 336776 627168 336832 627202
rect 336866 627168 336920 627202
rect 336240 627112 336920 627168
rect 336240 627078 336292 627112
rect 336326 627078 336382 627112
rect 336416 627078 336472 627112
rect 336506 627078 336562 627112
rect 336596 627078 336652 627112
rect 336686 627078 336742 627112
rect 336776 627078 336832 627112
rect 336866 627078 336920 627112
rect 336240 627022 336920 627078
rect 336240 626988 336292 627022
rect 336326 626988 336382 627022
rect 336416 626988 336472 627022
rect 336506 626988 336562 627022
rect 336596 626988 336652 627022
rect 336686 626988 336742 627022
rect 336776 626988 336832 627022
rect 336866 626988 336920 627022
rect 336240 626932 336920 626988
rect 336240 626898 336292 626932
rect 336326 626898 336382 626932
rect 336416 626898 336472 626932
rect 336506 626898 336562 626932
rect 336596 626898 336652 626932
rect 336686 626898 336742 626932
rect 336776 626898 336832 626932
rect 336866 626898 336920 626932
rect 336240 626842 336920 626898
rect 336240 626808 336292 626842
rect 336326 626808 336382 626842
rect 336416 626808 336472 626842
rect 336506 626808 336562 626842
rect 336596 626808 336652 626842
rect 336686 626808 336742 626842
rect 336776 626808 336832 626842
rect 336866 626808 336920 626842
rect 336240 626756 336920 626808
rect 337528 627382 338208 627436
rect 337528 627348 337580 627382
rect 337614 627348 337670 627382
rect 337704 627348 337760 627382
rect 337794 627348 337850 627382
rect 337884 627348 337940 627382
rect 337974 627348 338030 627382
rect 338064 627348 338120 627382
rect 338154 627348 338208 627382
rect 337528 627292 338208 627348
rect 337528 627258 337580 627292
rect 337614 627258 337670 627292
rect 337704 627258 337760 627292
rect 337794 627258 337850 627292
rect 337884 627258 337940 627292
rect 337974 627258 338030 627292
rect 338064 627258 338120 627292
rect 338154 627258 338208 627292
rect 337528 627202 338208 627258
rect 337528 627168 337580 627202
rect 337614 627168 337670 627202
rect 337704 627168 337760 627202
rect 337794 627168 337850 627202
rect 337884 627168 337940 627202
rect 337974 627168 338030 627202
rect 338064 627168 338120 627202
rect 338154 627168 338208 627202
rect 337528 627112 338208 627168
rect 337528 627078 337580 627112
rect 337614 627078 337670 627112
rect 337704 627078 337760 627112
rect 337794 627078 337850 627112
rect 337884 627078 337940 627112
rect 337974 627078 338030 627112
rect 338064 627078 338120 627112
rect 338154 627078 338208 627112
rect 337528 627022 338208 627078
rect 337528 626988 337580 627022
rect 337614 626988 337670 627022
rect 337704 626988 337760 627022
rect 337794 626988 337850 627022
rect 337884 626988 337940 627022
rect 337974 626988 338030 627022
rect 338064 626988 338120 627022
rect 338154 626988 338208 627022
rect 337528 626932 338208 626988
rect 337528 626898 337580 626932
rect 337614 626898 337670 626932
rect 337704 626898 337760 626932
rect 337794 626898 337850 626932
rect 337884 626898 337940 626932
rect 337974 626898 338030 626932
rect 338064 626898 338120 626932
rect 338154 626898 338208 626932
rect 337528 626842 338208 626898
rect 337528 626808 337580 626842
rect 337614 626808 337670 626842
rect 337704 626808 337760 626842
rect 337794 626808 337850 626842
rect 337884 626808 337940 626842
rect 337974 626808 338030 626842
rect 338064 626808 338120 626842
rect 338154 626808 338208 626842
rect 337528 626756 338208 626808
rect 338816 627382 339496 627436
rect 338816 627348 338868 627382
rect 338902 627348 338958 627382
rect 338992 627348 339048 627382
rect 339082 627348 339138 627382
rect 339172 627348 339228 627382
rect 339262 627348 339318 627382
rect 339352 627348 339408 627382
rect 339442 627348 339496 627382
rect 338816 627292 339496 627348
rect 338816 627258 338868 627292
rect 338902 627258 338958 627292
rect 338992 627258 339048 627292
rect 339082 627258 339138 627292
rect 339172 627258 339228 627292
rect 339262 627258 339318 627292
rect 339352 627258 339408 627292
rect 339442 627258 339496 627292
rect 338816 627202 339496 627258
rect 338816 627168 338868 627202
rect 338902 627168 338958 627202
rect 338992 627168 339048 627202
rect 339082 627168 339138 627202
rect 339172 627168 339228 627202
rect 339262 627168 339318 627202
rect 339352 627168 339408 627202
rect 339442 627168 339496 627202
rect 338816 627112 339496 627168
rect 338816 627078 338868 627112
rect 338902 627078 338958 627112
rect 338992 627078 339048 627112
rect 339082 627078 339138 627112
rect 339172 627078 339228 627112
rect 339262 627078 339318 627112
rect 339352 627078 339408 627112
rect 339442 627078 339496 627112
rect 338816 627022 339496 627078
rect 338816 626988 338868 627022
rect 338902 626988 338958 627022
rect 338992 626988 339048 627022
rect 339082 626988 339138 627022
rect 339172 626988 339228 627022
rect 339262 626988 339318 627022
rect 339352 626988 339408 627022
rect 339442 626988 339496 627022
rect 338816 626932 339496 626988
rect 338816 626898 338868 626932
rect 338902 626898 338958 626932
rect 338992 626898 339048 626932
rect 339082 626898 339138 626932
rect 339172 626898 339228 626932
rect 339262 626898 339318 626932
rect 339352 626898 339408 626932
rect 339442 626898 339496 626932
rect 338816 626842 339496 626898
rect 338816 626808 338868 626842
rect 338902 626808 338958 626842
rect 338992 626808 339048 626842
rect 339082 626808 339138 626842
rect 339172 626808 339228 626842
rect 339262 626808 339318 626842
rect 339352 626808 339408 626842
rect 339442 626808 339496 626842
rect 338816 626756 339496 626808
rect 340104 627382 340784 627436
rect 340104 627348 340156 627382
rect 340190 627348 340246 627382
rect 340280 627348 340336 627382
rect 340370 627348 340426 627382
rect 340460 627348 340516 627382
rect 340550 627348 340606 627382
rect 340640 627348 340696 627382
rect 340730 627348 340784 627382
rect 340104 627292 340784 627348
rect 340104 627258 340156 627292
rect 340190 627258 340246 627292
rect 340280 627258 340336 627292
rect 340370 627258 340426 627292
rect 340460 627258 340516 627292
rect 340550 627258 340606 627292
rect 340640 627258 340696 627292
rect 340730 627258 340784 627292
rect 340104 627202 340784 627258
rect 340104 627168 340156 627202
rect 340190 627168 340246 627202
rect 340280 627168 340336 627202
rect 340370 627168 340426 627202
rect 340460 627168 340516 627202
rect 340550 627168 340606 627202
rect 340640 627168 340696 627202
rect 340730 627168 340784 627202
rect 340104 627112 340784 627168
rect 340104 627078 340156 627112
rect 340190 627078 340246 627112
rect 340280 627078 340336 627112
rect 340370 627078 340426 627112
rect 340460 627078 340516 627112
rect 340550 627078 340606 627112
rect 340640 627078 340696 627112
rect 340730 627078 340784 627112
rect 340104 627022 340784 627078
rect 340104 626988 340156 627022
rect 340190 626988 340246 627022
rect 340280 626988 340336 627022
rect 340370 626988 340426 627022
rect 340460 626988 340516 627022
rect 340550 626988 340606 627022
rect 340640 626988 340696 627022
rect 340730 626988 340784 627022
rect 340104 626932 340784 626988
rect 340104 626898 340156 626932
rect 340190 626898 340246 626932
rect 340280 626898 340336 626932
rect 340370 626898 340426 626932
rect 340460 626898 340516 626932
rect 340550 626898 340606 626932
rect 340640 626898 340696 626932
rect 340730 626898 340784 626932
rect 340104 626842 340784 626898
rect 340104 626808 340156 626842
rect 340190 626808 340246 626842
rect 340280 626808 340336 626842
rect 340370 626808 340426 626842
rect 340460 626808 340516 626842
rect 340550 626808 340606 626842
rect 340640 626808 340696 626842
rect 340730 626808 340784 626842
rect 340104 626756 340784 626808
rect 334952 626094 335632 626148
rect 334952 626060 335004 626094
rect 335038 626060 335094 626094
rect 335128 626060 335184 626094
rect 335218 626060 335274 626094
rect 335308 626060 335364 626094
rect 335398 626060 335454 626094
rect 335488 626060 335544 626094
rect 335578 626060 335632 626094
rect 334952 626004 335632 626060
rect 334952 625970 335004 626004
rect 335038 625970 335094 626004
rect 335128 625970 335184 626004
rect 335218 625970 335274 626004
rect 335308 625970 335364 626004
rect 335398 625970 335454 626004
rect 335488 625970 335544 626004
rect 335578 625970 335632 626004
rect 334952 625914 335632 625970
rect 334952 625880 335004 625914
rect 335038 625880 335094 625914
rect 335128 625880 335184 625914
rect 335218 625880 335274 625914
rect 335308 625880 335364 625914
rect 335398 625880 335454 625914
rect 335488 625880 335544 625914
rect 335578 625880 335632 625914
rect 334952 625824 335632 625880
rect 334952 625790 335004 625824
rect 335038 625790 335094 625824
rect 335128 625790 335184 625824
rect 335218 625790 335274 625824
rect 335308 625790 335364 625824
rect 335398 625790 335454 625824
rect 335488 625790 335544 625824
rect 335578 625790 335632 625824
rect 334952 625734 335632 625790
rect 334952 625700 335004 625734
rect 335038 625700 335094 625734
rect 335128 625700 335184 625734
rect 335218 625700 335274 625734
rect 335308 625700 335364 625734
rect 335398 625700 335454 625734
rect 335488 625700 335544 625734
rect 335578 625700 335632 625734
rect 334952 625644 335632 625700
rect 334952 625610 335004 625644
rect 335038 625610 335094 625644
rect 335128 625610 335184 625644
rect 335218 625610 335274 625644
rect 335308 625610 335364 625644
rect 335398 625610 335454 625644
rect 335488 625610 335544 625644
rect 335578 625610 335632 625644
rect 334952 625554 335632 625610
rect 334952 625520 335004 625554
rect 335038 625520 335094 625554
rect 335128 625520 335184 625554
rect 335218 625520 335274 625554
rect 335308 625520 335364 625554
rect 335398 625520 335454 625554
rect 335488 625520 335544 625554
rect 335578 625520 335632 625554
rect 334952 625468 335632 625520
rect 336240 626094 336920 626148
rect 336240 626060 336292 626094
rect 336326 626060 336382 626094
rect 336416 626060 336472 626094
rect 336506 626060 336562 626094
rect 336596 626060 336652 626094
rect 336686 626060 336742 626094
rect 336776 626060 336832 626094
rect 336866 626060 336920 626094
rect 336240 626004 336920 626060
rect 336240 625970 336292 626004
rect 336326 625970 336382 626004
rect 336416 625970 336472 626004
rect 336506 625970 336562 626004
rect 336596 625970 336652 626004
rect 336686 625970 336742 626004
rect 336776 625970 336832 626004
rect 336866 625970 336920 626004
rect 336240 625914 336920 625970
rect 336240 625880 336292 625914
rect 336326 625880 336382 625914
rect 336416 625880 336472 625914
rect 336506 625880 336562 625914
rect 336596 625880 336652 625914
rect 336686 625880 336742 625914
rect 336776 625880 336832 625914
rect 336866 625880 336920 625914
rect 336240 625824 336920 625880
rect 336240 625790 336292 625824
rect 336326 625790 336382 625824
rect 336416 625790 336472 625824
rect 336506 625790 336562 625824
rect 336596 625790 336652 625824
rect 336686 625790 336742 625824
rect 336776 625790 336832 625824
rect 336866 625790 336920 625824
rect 336240 625734 336920 625790
rect 336240 625700 336292 625734
rect 336326 625700 336382 625734
rect 336416 625700 336472 625734
rect 336506 625700 336562 625734
rect 336596 625700 336652 625734
rect 336686 625700 336742 625734
rect 336776 625700 336832 625734
rect 336866 625700 336920 625734
rect 336240 625644 336920 625700
rect 336240 625610 336292 625644
rect 336326 625610 336382 625644
rect 336416 625610 336472 625644
rect 336506 625610 336562 625644
rect 336596 625610 336652 625644
rect 336686 625610 336742 625644
rect 336776 625610 336832 625644
rect 336866 625610 336920 625644
rect 336240 625554 336920 625610
rect 336240 625520 336292 625554
rect 336326 625520 336382 625554
rect 336416 625520 336472 625554
rect 336506 625520 336562 625554
rect 336596 625520 336652 625554
rect 336686 625520 336742 625554
rect 336776 625520 336832 625554
rect 336866 625520 336920 625554
rect 336240 625468 336920 625520
rect 337528 626094 338208 626148
rect 337528 626060 337580 626094
rect 337614 626060 337670 626094
rect 337704 626060 337760 626094
rect 337794 626060 337850 626094
rect 337884 626060 337940 626094
rect 337974 626060 338030 626094
rect 338064 626060 338120 626094
rect 338154 626060 338208 626094
rect 337528 626004 338208 626060
rect 337528 625970 337580 626004
rect 337614 625970 337670 626004
rect 337704 625970 337760 626004
rect 337794 625970 337850 626004
rect 337884 625970 337940 626004
rect 337974 625970 338030 626004
rect 338064 625970 338120 626004
rect 338154 625970 338208 626004
rect 337528 625914 338208 625970
rect 337528 625880 337580 625914
rect 337614 625880 337670 625914
rect 337704 625880 337760 625914
rect 337794 625880 337850 625914
rect 337884 625880 337940 625914
rect 337974 625880 338030 625914
rect 338064 625880 338120 625914
rect 338154 625880 338208 625914
rect 337528 625824 338208 625880
rect 337528 625790 337580 625824
rect 337614 625790 337670 625824
rect 337704 625790 337760 625824
rect 337794 625790 337850 625824
rect 337884 625790 337940 625824
rect 337974 625790 338030 625824
rect 338064 625790 338120 625824
rect 338154 625790 338208 625824
rect 337528 625734 338208 625790
rect 337528 625700 337580 625734
rect 337614 625700 337670 625734
rect 337704 625700 337760 625734
rect 337794 625700 337850 625734
rect 337884 625700 337940 625734
rect 337974 625700 338030 625734
rect 338064 625700 338120 625734
rect 338154 625700 338208 625734
rect 337528 625644 338208 625700
rect 337528 625610 337580 625644
rect 337614 625610 337670 625644
rect 337704 625610 337760 625644
rect 337794 625610 337850 625644
rect 337884 625610 337940 625644
rect 337974 625610 338030 625644
rect 338064 625610 338120 625644
rect 338154 625610 338208 625644
rect 337528 625554 338208 625610
rect 337528 625520 337580 625554
rect 337614 625520 337670 625554
rect 337704 625520 337760 625554
rect 337794 625520 337850 625554
rect 337884 625520 337940 625554
rect 337974 625520 338030 625554
rect 338064 625520 338120 625554
rect 338154 625520 338208 625554
rect 337528 625468 338208 625520
rect 338816 626094 339496 626148
rect 338816 626060 338868 626094
rect 338902 626060 338958 626094
rect 338992 626060 339048 626094
rect 339082 626060 339138 626094
rect 339172 626060 339228 626094
rect 339262 626060 339318 626094
rect 339352 626060 339408 626094
rect 339442 626060 339496 626094
rect 338816 626004 339496 626060
rect 338816 625970 338868 626004
rect 338902 625970 338958 626004
rect 338992 625970 339048 626004
rect 339082 625970 339138 626004
rect 339172 625970 339228 626004
rect 339262 625970 339318 626004
rect 339352 625970 339408 626004
rect 339442 625970 339496 626004
rect 338816 625914 339496 625970
rect 338816 625880 338868 625914
rect 338902 625880 338958 625914
rect 338992 625880 339048 625914
rect 339082 625880 339138 625914
rect 339172 625880 339228 625914
rect 339262 625880 339318 625914
rect 339352 625880 339408 625914
rect 339442 625880 339496 625914
rect 338816 625824 339496 625880
rect 338816 625790 338868 625824
rect 338902 625790 338958 625824
rect 338992 625790 339048 625824
rect 339082 625790 339138 625824
rect 339172 625790 339228 625824
rect 339262 625790 339318 625824
rect 339352 625790 339408 625824
rect 339442 625790 339496 625824
rect 338816 625734 339496 625790
rect 338816 625700 338868 625734
rect 338902 625700 338958 625734
rect 338992 625700 339048 625734
rect 339082 625700 339138 625734
rect 339172 625700 339228 625734
rect 339262 625700 339318 625734
rect 339352 625700 339408 625734
rect 339442 625700 339496 625734
rect 338816 625644 339496 625700
rect 338816 625610 338868 625644
rect 338902 625610 338958 625644
rect 338992 625610 339048 625644
rect 339082 625610 339138 625644
rect 339172 625610 339228 625644
rect 339262 625610 339318 625644
rect 339352 625610 339408 625644
rect 339442 625610 339496 625644
rect 338816 625554 339496 625610
rect 338816 625520 338868 625554
rect 338902 625520 338958 625554
rect 338992 625520 339048 625554
rect 339082 625520 339138 625554
rect 339172 625520 339228 625554
rect 339262 625520 339318 625554
rect 339352 625520 339408 625554
rect 339442 625520 339496 625554
rect 338816 625468 339496 625520
rect 340104 626094 340784 626148
rect 340104 626060 340156 626094
rect 340190 626060 340246 626094
rect 340280 626060 340336 626094
rect 340370 626060 340426 626094
rect 340460 626060 340516 626094
rect 340550 626060 340606 626094
rect 340640 626060 340696 626094
rect 340730 626060 340784 626094
rect 340104 626004 340784 626060
rect 340104 625970 340156 626004
rect 340190 625970 340246 626004
rect 340280 625970 340336 626004
rect 340370 625970 340426 626004
rect 340460 625970 340516 626004
rect 340550 625970 340606 626004
rect 340640 625970 340696 626004
rect 340730 625970 340784 626004
rect 340104 625914 340784 625970
rect 340104 625880 340156 625914
rect 340190 625880 340246 625914
rect 340280 625880 340336 625914
rect 340370 625880 340426 625914
rect 340460 625880 340516 625914
rect 340550 625880 340606 625914
rect 340640 625880 340696 625914
rect 340730 625880 340784 625914
rect 340104 625824 340784 625880
rect 340104 625790 340156 625824
rect 340190 625790 340246 625824
rect 340280 625790 340336 625824
rect 340370 625790 340426 625824
rect 340460 625790 340516 625824
rect 340550 625790 340606 625824
rect 340640 625790 340696 625824
rect 340730 625790 340784 625824
rect 340104 625734 340784 625790
rect 340104 625700 340156 625734
rect 340190 625700 340246 625734
rect 340280 625700 340336 625734
rect 340370 625700 340426 625734
rect 340460 625700 340516 625734
rect 340550 625700 340606 625734
rect 340640 625700 340696 625734
rect 340730 625700 340784 625734
rect 340104 625644 340784 625700
rect 340104 625610 340156 625644
rect 340190 625610 340246 625644
rect 340280 625610 340336 625644
rect 340370 625610 340426 625644
rect 340460 625610 340516 625644
rect 340550 625610 340606 625644
rect 340640 625610 340696 625644
rect 340730 625610 340784 625644
rect 340104 625554 340784 625610
rect 340104 625520 340156 625554
rect 340190 625520 340246 625554
rect 340280 625520 340336 625554
rect 340370 625520 340426 625554
rect 340460 625520 340516 625554
rect 340550 625520 340606 625554
rect 340640 625520 340696 625554
rect 340730 625520 340784 625554
rect 340104 625468 340784 625520
rect 313392 624934 313450 624946
rect 303584 619736 303642 619748
rect 303584 617180 303596 619736
rect 303630 617180 303642 619736
rect 303584 617168 303642 617180
rect 304042 619736 304100 619748
rect 304042 617180 304054 619736
rect 304088 617180 304100 619736
rect 304042 617168 304100 617180
rect 304156 619736 304214 619748
rect 304156 617180 304168 619736
rect 304202 617180 304214 619736
rect 304156 617168 304214 617180
rect 304614 619736 304672 619748
rect 304614 617180 304626 619736
rect 304660 617180 304672 619736
rect 304614 617168 304672 617180
rect 304728 619736 304786 619748
rect 304728 617180 304740 619736
rect 304774 617180 304786 619736
rect 304728 617168 304786 617180
rect 305186 619736 305244 619748
rect 305186 617180 305198 619736
rect 305232 617180 305244 619736
rect 305186 617168 305244 617180
rect 305300 619736 305358 619748
rect 305300 617180 305312 619736
rect 305346 617180 305358 619736
rect 305300 617168 305358 617180
rect 305758 619736 305816 619748
rect 305758 617180 305770 619736
rect 305804 617180 305816 619736
rect 305758 617168 305816 617180
rect 305872 619736 305930 619748
rect 305872 617180 305884 619736
rect 305918 617180 305930 619736
rect 305872 617168 305930 617180
rect 306330 619736 306388 619748
rect 306330 617180 306342 619736
rect 306376 617180 306388 619736
rect 306330 617168 306388 617180
rect 306444 619736 306502 619748
rect 306444 617180 306456 619736
rect 306490 617180 306502 619736
rect 306444 617168 306502 617180
rect 306902 619736 306960 619748
rect 306902 617180 306914 619736
rect 306948 617180 306960 619736
rect 306902 617168 306960 617180
rect 307016 619736 307074 619748
rect 307016 617180 307028 619736
rect 307062 617180 307074 619736
rect 307016 617168 307074 617180
rect 307474 619736 307532 619748
rect 307474 617180 307486 619736
rect 307520 617180 307532 619736
rect 307474 617168 307532 617180
rect 307588 619736 307646 619748
rect 307588 617180 307600 619736
rect 307634 617180 307646 619736
rect 307588 617168 307646 617180
rect 308046 619736 308104 619748
rect 308046 617180 308058 619736
rect 308092 617180 308104 619736
rect 308046 617168 308104 617180
rect 308160 619736 308218 619748
rect 308160 617180 308172 619736
rect 308206 617180 308218 619736
rect 308160 617168 308218 617180
rect 308618 619736 308676 619748
rect 308618 617180 308630 619736
rect 308664 617180 308676 619736
rect 308618 617168 308676 617180
rect 308732 619736 308790 619748
rect 308732 617180 308744 619736
rect 308778 617180 308790 619736
rect 308732 617168 308790 617180
rect 309190 619736 309248 619748
rect 309190 617180 309202 619736
rect 309236 617180 309248 619736
rect 309190 617168 309248 617180
rect 309304 619736 309362 619748
rect 309304 617180 309316 619736
rect 309350 617180 309362 619736
rect 309304 617168 309362 617180
rect 309762 619736 309820 619748
rect 309762 617180 309774 619736
rect 309808 617180 309820 619736
rect 309762 617168 309820 617180
rect 309876 619736 309934 619748
rect 309876 617180 309888 619736
rect 309922 617180 309934 619736
rect 309876 617168 309934 617180
rect 310334 619736 310392 619748
rect 310334 617180 310346 619736
rect 310380 617180 310392 619736
rect 310334 617168 310392 617180
rect 310448 619736 310506 619748
rect 310448 617180 310460 619736
rect 310494 617180 310506 619736
rect 310448 617168 310506 617180
rect 310906 619736 310964 619748
rect 310906 617180 310918 619736
rect 310952 617180 310964 619736
rect 310906 617168 310964 617180
rect 311020 619736 311078 619748
rect 311020 617180 311032 619736
rect 311066 617180 311078 619736
rect 311020 617168 311078 617180
rect 311478 619736 311536 619748
rect 311478 617180 311490 619736
rect 311524 617180 311536 619736
rect 313392 617218 313404 624934
rect 313438 617218 313450 624934
rect 313392 617206 313450 617218
rect 313850 624934 313908 624946
rect 313850 617218 313862 624934
rect 313896 617218 313908 624934
rect 313850 617206 313908 617218
rect 314308 624934 314366 624946
rect 314308 617218 314320 624934
rect 314354 617218 314366 624934
rect 314308 617206 314366 617218
rect 314766 624934 314824 624946
rect 314766 617218 314778 624934
rect 314812 617218 314824 624934
rect 314766 617206 314824 617218
rect 315224 624934 315282 624946
rect 315224 617218 315236 624934
rect 315270 617218 315282 624934
rect 315224 617206 315282 617218
rect 315682 624934 315740 624946
rect 315682 617218 315694 624934
rect 315728 617218 315740 624934
rect 315682 617206 315740 617218
rect 316140 624934 316198 624946
rect 316140 617218 316152 624934
rect 316186 617218 316198 624934
rect 316140 617206 316198 617218
rect 316598 624934 316656 624946
rect 316598 617218 316610 624934
rect 316644 617218 316656 624934
rect 316598 617206 316656 617218
rect 317056 624934 317114 624946
rect 317056 617218 317068 624934
rect 317102 617218 317114 624934
rect 317056 617206 317114 617218
rect 317514 624934 317572 624946
rect 317514 617218 317526 624934
rect 317560 617218 317572 624934
rect 317514 617206 317572 617218
rect 317972 624934 318030 624946
rect 317972 617218 317984 624934
rect 318018 617218 318030 624934
rect 317972 617206 318030 617218
rect 318430 624934 318488 624946
rect 318430 617218 318442 624934
rect 318476 617218 318488 624934
rect 319350 624934 319408 624946
rect 318430 617206 318488 617218
rect 319350 617218 319362 624934
rect 319396 617218 319408 624934
rect 319350 617206 319408 617218
rect 319808 624934 319866 624946
rect 319808 617218 319820 624934
rect 319854 617218 319866 624934
rect 319808 617206 319866 617218
rect 320266 624934 320324 624946
rect 320266 617218 320278 624934
rect 320312 617218 320324 624934
rect 320266 617206 320324 617218
rect 320724 624934 320782 624946
rect 320724 617218 320736 624934
rect 320770 617218 320782 624934
rect 320724 617206 320782 617218
rect 321182 624934 321240 624946
rect 321182 617218 321194 624934
rect 321228 617218 321240 624934
rect 321182 617206 321240 617218
rect 321640 624934 321698 624946
rect 321640 617218 321652 624934
rect 321686 617218 321698 624934
rect 321640 617206 321698 617218
rect 322098 624934 322156 624946
rect 322098 617218 322110 624934
rect 322144 617218 322156 624934
rect 322098 617206 322156 617218
rect 322556 624934 322614 624946
rect 322556 617218 322568 624934
rect 322602 617218 322614 624934
rect 322556 617206 322614 617218
rect 323014 624934 323072 624946
rect 323014 617218 323026 624934
rect 323060 617218 323072 624934
rect 323014 617206 323072 617218
rect 323472 624934 323530 624946
rect 323472 617218 323484 624934
rect 323518 617218 323530 624934
rect 323472 617206 323530 617218
rect 323930 624934 323988 624946
rect 323930 617218 323942 624934
rect 323976 617218 323988 624934
rect 324850 624934 324908 624946
rect 323930 617206 323988 617218
rect 324850 617218 324862 624934
rect 324896 617218 324908 624934
rect 324850 617206 324908 617218
rect 325308 624934 325366 624946
rect 325308 617218 325320 624934
rect 325354 617218 325366 624934
rect 325308 617206 325366 617218
rect 325766 624934 325824 624946
rect 325766 617218 325778 624934
rect 325812 617218 325824 624934
rect 325766 617206 325824 617218
rect 326224 624934 326282 624946
rect 326224 617218 326236 624934
rect 326270 617218 326282 624934
rect 326224 617206 326282 617218
rect 326682 624934 326740 624946
rect 326682 617218 326694 624934
rect 326728 617218 326740 624934
rect 326682 617206 326740 617218
rect 327140 624934 327198 624946
rect 327140 617218 327152 624934
rect 327186 617218 327198 624934
rect 327140 617206 327198 617218
rect 327598 624934 327656 624946
rect 327598 617218 327610 624934
rect 327644 617218 327656 624934
rect 327598 617206 327656 617218
rect 328056 624934 328114 624946
rect 328056 617218 328068 624934
rect 328102 617218 328114 624934
rect 328056 617206 328114 617218
rect 328514 624934 328572 624946
rect 328514 617218 328526 624934
rect 328560 617218 328572 624934
rect 328514 617206 328572 617218
rect 328972 624934 329030 624946
rect 328972 617218 328984 624934
rect 329018 617218 329030 624934
rect 328972 617206 329030 617218
rect 329430 624934 329488 624946
rect 329430 617218 329442 624934
rect 329476 617218 329488 624934
rect 329430 617206 329488 617218
rect 329888 624934 329946 624946
rect 329888 617218 329900 624934
rect 329934 617218 329946 624934
rect 334952 624806 335632 624860
rect 334952 624772 335004 624806
rect 335038 624772 335094 624806
rect 335128 624772 335184 624806
rect 335218 624772 335274 624806
rect 335308 624772 335364 624806
rect 335398 624772 335454 624806
rect 335488 624772 335544 624806
rect 335578 624772 335632 624806
rect 334952 624716 335632 624772
rect 334952 624682 335004 624716
rect 335038 624682 335094 624716
rect 335128 624682 335184 624716
rect 335218 624682 335274 624716
rect 335308 624682 335364 624716
rect 335398 624682 335454 624716
rect 335488 624682 335544 624716
rect 335578 624682 335632 624716
rect 334952 624626 335632 624682
rect 334952 624592 335004 624626
rect 335038 624592 335094 624626
rect 335128 624592 335184 624626
rect 335218 624592 335274 624626
rect 335308 624592 335364 624626
rect 335398 624592 335454 624626
rect 335488 624592 335544 624626
rect 335578 624592 335632 624626
rect 334952 624536 335632 624592
rect 334952 624502 335004 624536
rect 335038 624502 335094 624536
rect 335128 624502 335184 624536
rect 335218 624502 335274 624536
rect 335308 624502 335364 624536
rect 335398 624502 335454 624536
rect 335488 624502 335544 624536
rect 335578 624502 335632 624536
rect 334952 624446 335632 624502
rect 334952 624412 335004 624446
rect 335038 624412 335094 624446
rect 335128 624412 335184 624446
rect 335218 624412 335274 624446
rect 335308 624412 335364 624446
rect 335398 624412 335454 624446
rect 335488 624412 335544 624446
rect 335578 624412 335632 624446
rect 334952 624356 335632 624412
rect 334952 624322 335004 624356
rect 335038 624322 335094 624356
rect 335128 624322 335184 624356
rect 335218 624322 335274 624356
rect 335308 624322 335364 624356
rect 335398 624322 335454 624356
rect 335488 624322 335544 624356
rect 335578 624322 335632 624356
rect 334952 624266 335632 624322
rect 334952 624232 335004 624266
rect 335038 624232 335094 624266
rect 335128 624232 335184 624266
rect 335218 624232 335274 624266
rect 335308 624232 335364 624266
rect 335398 624232 335454 624266
rect 335488 624232 335544 624266
rect 335578 624232 335632 624266
rect 334952 624180 335632 624232
rect 336240 624806 336920 624860
rect 336240 624772 336292 624806
rect 336326 624772 336382 624806
rect 336416 624772 336472 624806
rect 336506 624772 336562 624806
rect 336596 624772 336652 624806
rect 336686 624772 336742 624806
rect 336776 624772 336832 624806
rect 336866 624772 336920 624806
rect 336240 624716 336920 624772
rect 336240 624682 336292 624716
rect 336326 624682 336382 624716
rect 336416 624682 336472 624716
rect 336506 624682 336562 624716
rect 336596 624682 336652 624716
rect 336686 624682 336742 624716
rect 336776 624682 336832 624716
rect 336866 624682 336920 624716
rect 336240 624626 336920 624682
rect 336240 624592 336292 624626
rect 336326 624592 336382 624626
rect 336416 624592 336472 624626
rect 336506 624592 336562 624626
rect 336596 624592 336652 624626
rect 336686 624592 336742 624626
rect 336776 624592 336832 624626
rect 336866 624592 336920 624626
rect 336240 624536 336920 624592
rect 336240 624502 336292 624536
rect 336326 624502 336382 624536
rect 336416 624502 336472 624536
rect 336506 624502 336562 624536
rect 336596 624502 336652 624536
rect 336686 624502 336742 624536
rect 336776 624502 336832 624536
rect 336866 624502 336920 624536
rect 336240 624446 336920 624502
rect 336240 624412 336292 624446
rect 336326 624412 336382 624446
rect 336416 624412 336472 624446
rect 336506 624412 336562 624446
rect 336596 624412 336652 624446
rect 336686 624412 336742 624446
rect 336776 624412 336832 624446
rect 336866 624412 336920 624446
rect 336240 624356 336920 624412
rect 336240 624322 336292 624356
rect 336326 624322 336382 624356
rect 336416 624322 336472 624356
rect 336506 624322 336562 624356
rect 336596 624322 336652 624356
rect 336686 624322 336742 624356
rect 336776 624322 336832 624356
rect 336866 624322 336920 624356
rect 336240 624266 336920 624322
rect 336240 624232 336292 624266
rect 336326 624232 336382 624266
rect 336416 624232 336472 624266
rect 336506 624232 336562 624266
rect 336596 624232 336652 624266
rect 336686 624232 336742 624266
rect 336776 624232 336832 624266
rect 336866 624232 336920 624266
rect 336240 624180 336920 624232
rect 337528 624806 338208 624860
rect 337528 624772 337580 624806
rect 337614 624772 337670 624806
rect 337704 624772 337760 624806
rect 337794 624772 337850 624806
rect 337884 624772 337940 624806
rect 337974 624772 338030 624806
rect 338064 624772 338120 624806
rect 338154 624772 338208 624806
rect 337528 624716 338208 624772
rect 337528 624682 337580 624716
rect 337614 624682 337670 624716
rect 337704 624682 337760 624716
rect 337794 624682 337850 624716
rect 337884 624682 337940 624716
rect 337974 624682 338030 624716
rect 338064 624682 338120 624716
rect 338154 624682 338208 624716
rect 337528 624626 338208 624682
rect 337528 624592 337580 624626
rect 337614 624592 337670 624626
rect 337704 624592 337760 624626
rect 337794 624592 337850 624626
rect 337884 624592 337940 624626
rect 337974 624592 338030 624626
rect 338064 624592 338120 624626
rect 338154 624592 338208 624626
rect 337528 624536 338208 624592
rect 337528 624502 337580 624536
rect 337614 624502 337670 624536
rect 337704 624502 337760 624536
rect 337794 624502 337850 624536
rect 337884 624502 337940 624536
rect 337974 624502 338030 624536
rect 338064 624502 338120 624536
rect 338154 624502 338208 624536
rect 337528 624446 338208 624502
rect 337528 624412 337580 624446
rect 337614 624412 337670 624446
rect 337704 624412 337760 624446
rect 337794 624412 337850 624446
rect 337884 624412 337940 624446
rect 337974 624412 338030 624446
rect 338064 624412 338120 624446
rect 338154 624412 338208 624446
rect 337528 624356 338208 624412
rect 337528 624322 337580 624356
rect 337614 624322 337670 624356
rect 337704 624322 337760 624356
rect 337794 624322 337850 624356
rect 337884 624322 337940 624356
rect 337974 624322 338030 624356
rect 338064 624322 338120 624356
rect 338154 624322 338208 624356
rect 337528 624266 338208 624322
rect 337528 624232 337580 624266
rect 337614 624232 337670 624266
rect 337704 624232 337760 624266
rect 337794 624232 337850 624266
rect 337884 624232 337940 624266
rect 337974 624232 338030 624266
rect 338064 624232 338120 624266
rect 338154 624232 338208 624266
rect 337528 624180 338208 624232
rect 338816 624806 339496 624860
rect 338816 624772 338868 624806
rect 338902 624772 338958 624806
rect 338992 624772 339048 624806
rect 339082 624772 339138 624806
rect 339172 624772 339228 624806
rect 339262 624772 339318 624806
rect 339352 624772 339408 624806
rect 339442 624772 339496 624806
rect 338816 624716 339496 624772
rect 338816 624682 338868 624716
rect 338902 624682 338958 624716
rect 338992 624682 339048 624716
rect 339082 624682 339138 624716
rect 339172 624682 339228 624716
rect 339262 624682 339318 624716
rect 339352 624682 339408 624716
rect 339442 624682 339496 624716
rect 338816 624626 339496 624682
rect 338816 624592 338868 624626
rect 338902 624592 338958 624626
rect 338992 624592 339048 624626
rect 339082 624592 339138 624626
rect 339172 624592 339228 624626
rect 339262 624592 339318 624626
rect 339352 624592 339408 624626
rect 339442 624592 339496 624626
rect 338816 624536 339496 624592
rect 338816 624502 338868 624536
rect 338902 624502 338958 624536
rect 338992 624502 339048 624536
rect 339082 624502 339138 624536
rect 339172 624502 339228 624536
rect 339262 624502 339318 624536
rect 339352 624502 339408 624536
rect 339442 624502 339496 624536
rect 338816 624446 339496 624502
rect 338816 624412 338868 624446
rect 338902 624412 338958 624446
rect 338992 624412 339048 624446
rect 339082 624412 339138 624446
rect 339172 624412 339228 624446
rect 339262 624412 339318 624446
rect 339352 624412 339408 624446
rect 339442 624412 339496 624446
rect 338816 624356 339496 624412
rect 338816 624322 338868 624356
rect 338902 624322 338958 624356
rect 338992 624322 339048 624356
rect 339082 624322 339138 624356
rect 339172 624322 339228 624356
rect 339262 624322 339318 624356
rect 339352 624322 339408 624356
rect 339442 624322 339496 624356
rect 338816 624266 339496 624322
rect 338816 624232 338868 624266
rect 338902 624232 338958 624266
rect 338992 624232 339048 624266
rect 339082 624232 339138 624266
rect 339172 624232 339228 624266
rect 339262 624232 339318 624266
rect 339352 624232 339408 624266
rect 339442 624232 339496 624266
rect 338816 624180 339496 624232
rect 340104 624806 340784 624860
rect 340104 624772 340156 624806
rect 340190 624772 340246 624806
rect 340280 624772 340336 624806
rect 340370 624772 340426 624806
rect 340460 624772 340516 624806
rect 340550 624772 340606 624806
rect 340640 624772 340696 624806
rect 340730 624772 340784 624806
rect 340104 624716 340784 624772
rect 340104 624682 340156 624716
rect 340190 624682 340246 624716
rect 340280 624682 340336 624716
rect 340370 624682 340426 624716
rect 340460 624682 340516 624716
rect 340550 624682 340606 624716
rect 340640 624682 340696 624716
rect 340730 624682 340784 624716
rect 340104 624626 340784 624682
rect 340104 624592 340156 624626
rect 340190 624592 340246 624626
rect 340280 624592 340336 624626
rect 340370 624592 340426 624626
rect 340460 624592 340516 624626
rect 340550 624592 340606 624626
rect 340640 624592 340696 624626
rect 340730 624592 340784 624626
rect 340104 624536 340784 624592
rect 340104 624502 340156 624536
rect 340190 624502 340246 624536
rect 340280 624502 340336 624536
rect 340370 624502 340426 624536
rect 340460 624502 340516 624536
rect 340550 624502 340606 624536
rect 340640 624502 340696 624536
rect 340730 624502 340784 624536
rect 340104 624446 340784 624502
rect 340104 624412 340156 624446
rect 340190 624412 340246 624446
rect 340280 624412 340336 624446
rect 340370 624412 340426 624446
rect 340460 624412 340516 624446
rect 340550 624412 340606 624446
rect 340640 624412 340696 624446
rect 340730 624412 340784 624446
rect 340104 624356 340784 624412
rect 340104 624322 340156 624356
rect 340190 624322 340246 624356
rect 340280 624322 340336 624356
rect 340370 624322 340426 624356
rect 340460 624322 340516 624356
rect 340550 624322 340606 624356
rect 340640 624322 340696 624356
rect 340730 624322 340784 624356
rect 340104 624266 340784 624322
rect 340104 624232 340156 624266
rect 340190 624232 340246 624266
rect 340280 624232 340336 624266
rect 340370 624232 340426 624266
rect 340460 624232 340516 624266
rect 340550 624232 340606 624266
rect 340640 624232 340696 624266
rect 340730 624232 340784 624266
rect 340104 624180 340784 624232
rect 334952 623518 335632 623572
rect 334952 623484 335004 623518
rect 335038 623484 335094 623518
rect 335128 623484 335184 623518
rect 335218 623484 335274 623518
rect 335308 623484 335364 623518
rect 335398 623484 335454 623518
rect 335488 623484 335544 623518
rect 335578 623484 335632 623518
rect 334952 623428 335632 623484
rect 334952 623394 335004 623428
rect 335038 623394 335094 623428
rect 335128 623394 335184 623428
rect 335218 623394 335274 623428
rect 335308 623394 335364 623428
rect 335398 623394 335454 623428
rect 335488 623394 335544 623428
rect 335578 623394 335632 623428
rect 334952 623338 335632 623394
rect 334952 623304 335004 623338
rect 335038 623304 335094 623338
rect 335128 623304 335184 623338
rect 335218 623304 335274 623338
rect 335308 623304 335364 623338
rect 335398 623304 335454 623338
rect 335488 623304 335544 623338
rect 335578 623304 335632 623338
rect 334952 623248 335632 623304
rect 334952 623214 335004 623248
rect 335038 623214 335094 623248
rect 335128 623214 335184 623248
rect 335218 623214 335274 623248
rect 335308 623214 335364 623248
rect 335398 623214 335454 623248
rect 335488 623214 335544 623248
rect 335578 623214 335632 623248
rect 334952 623158 335632 623214
rect 334952 623124 335004 623158
rect 335038 623124 335094 623158
rect 335128 623124 335184 623158
rect 335218 623124 335274 623158
rect 335308 623124 335364 623158
rect 335398 623124 335454 623158
rect 335488 623124 335544 623158
rect 335578 623124 335632 623158
rect 334952 623068 335632 623124
rect 334952 623034 335004 623068
rect 335038 623034 335094 623068
rect 335128 623034 335184 623068
rect 335218 623034 335274 623068
rect 335308 623034 335364 623068
rect 335398 623034 335454 623068
rect 335488 623034 335544 623068
rect 335578 623034 335632 623068
rect 334952 622978 335632 623034
rect 334952 622944 335004 622978
rect 335038 622944 335094 622978
rect 335128 622944 335184 622978
rect 335218 622944 335274 622978
rect 335308 622944 335364 622978
rect 335398 622944 335454 622978
rect 335488 622944 335544 622978
rect 335578 622944 335632 622978
rect 334952 622892 335632 622944
rect 336240 623518 336920 623572
rect 336240 623484 336292 623518
rect 336326 623484 336382 623518
rect 336416 623484 336472 623518
rect 336506 623484 336562 623518
rect 336596 623484 336652 623518
rect 336686 623484 336742 623518
rect 336776 623484 336832 623518
rect 336866 623484 336920 623518
rect 336240 623428 336920 623484
rect 336240 623394 336292 623428
rect 336326 623394 336382 623428
rect 336416 623394 336472 623428
rect 336506 623394 336562 623428
rect 336596 623394 336652 623428
rect 336686 623394 336742 623428
rect 336776 623394 336832 623428
rect 336866 623394 336920 623428
rect 336240 623338 336920 623394
rect 336240 623304 336292 623338
rect 336326 623304 336382 623338
rect 336416 623304 336472 623338
rect 336506 623304 336562 623338
rect 336596 623304 336652 623338
rect 336686 623304 336742 623338
rect 336776 623304 336832 623338
rect 336866 623304 336920 623338
rect 336240 623248 336920 623304
rect 336240 623214 336292 623248
rect 336326 623214 336382 623248
rect 336416 623214 336472 623248
rect 336506 623214 336562 623248
rect 336596 623214 336652 623248
rect 336686 623214 336742 623248
rect 336776 623214 336832 623248
rect 336866 623214 336920 623248
rect 336240 623158 336920 623214
rect 336240 623124 336292 623158
rect 336326 623124 336382 623158
rect 336416 623124 336472 623158
rect 336506 623124 336562 623158
rect 336596 623124 336652 623158
rect 336686 623124 336742 623158
rect 336776 623124 336832 623158
rect 336866 623124 336920 623158
rect 336240 623068 336920 623124
rect 336240 623034 336292 623068
rect 336326 623034 336382 623068
rect 336416 623034 336472 623068
rect 336506 623034 336562 623068
rect 336596 623034 336652 623068
rect 336686 623034 336742 623068
rect 336776 623034 336832 623068
rect 336866 623034 336920 623068
rect 336240 622978 336920 623034
rect 336240 622944 336292 622978
rect 336326 622944 336382 622978
rect 336416 622944 336472 622978
rect 336506 622944 336562 622978
rect 336596 622944 336652 622978
rect 336686 622944 336742 622978
rect 336776 622944 336832 622978
rect 336866 622944 336920 622978
rect 336240 622892 336920 622944
rect 337528 623518 338208 623572
rect 337528 623484 337580 623518
rect 337614 623484 337670 623518
rect 337704 623484 337760 623518
rect 337794 623484 337850 623518
rect 337884 623484 337940 623518
rect 337974 623484 338030 623518
rect 338064 623484 338120 623518
rect 338154 623484 338208 623518
rect 337528 623428 338208 623484
rect 337528 623394 337580 623428
rect 337614 623394 337670 623428
rect 337704 623394 337760 623428
rect 337794 623394 337850 623428
rect 337884 623394 337940 623428
rect 337974 623394 338030 623428
rect 338064 623394 338120 623428
rect 338154 623394 338208 623428
rect 337528 623338 338208 623394
rect 337528 623304 337580 623338
rect 337614 623304 337670 623338
rect 337704 623304 337760 623338
rect 337794 623304 337850 623338
rect 337884 623304 337940 623338
rect 337974 623304 338030 623338
rect 338064 623304 338120 623338
rect 338154 623304 338208 623338
rect 337528 623248 338208 623304
rect 337528 623214 337580 623248
rect 337614 623214 337670 623248
rect 337704 623214 337760 623248
rect 337794 623214 337850 623248
rect 337884 623214 337940 623248
rect 337974 623214 338030 623248
rect 338064 623214 338120 623248
rect 338154 623214 338208 623248
rect 337528 623158 338208 623214
rect 337528 623124 337580 623158
rect 337614 623124 337670 623158
rect 337704 623124 337760 623158
rect 337794 623124 337850 623158
rect 337884 623124 337940 623158
rect 337974 623124 338030 623158
rect 338064 623124 338120 623158
rect 338154 623124 338208 623158
rect 337528 623068 338208 623124
rect 337528 623034 337580 623068
rect 337614 623034 337670 623068
rect 337704 623034 337760 623068
rect 337794 623034 337850 623068
rect 337884 623034 337940 623068
rect 337974 623034 338030 623068
rect 338064 623034 338120 623068
rect 338154 623034 338208 623068
rect 337528 622978 338208 623034
rect 337528 622944 337580 622978
rect 337614 622944 337670 622978
rect 337704 622944 337760 622978
rect 337794 622944 337850 622978
rect 337884 622944 337940 622978
rect 337974 622944 338030 622978
rect 338064 622944 338120 622978
rect 338154 622944 338208 622978
rect 337528 622892 338208 622944
rect 338816 623518 339496 623572
rect 338816 623484 338868 623518
rect 338902 623484 338958 623518
rect 338992 623484 339048 623518
rect 339082 623484 339138 623518
rect 339172 623484 339228 623518
rect 339262 623484 339318 623518
rect 339352 623484 339408 623518
rect 339442 623484 339496 623518
rect 338816 623428 339496 623484
rect 338816 623394 338868 623428
rect 338902 623394 338958 623428
rect 338992 623394 339048 623428
rect 339082 623394 339138 623428
rect 339172 623394 339228 623428
rect 339262 623394 339318 623428
rect 339352 623394 339408 623428
rect 339442 623394 339496 623428
rect 338816 623338 339496 623394
rect 338816 623304 338868 623338
rect 338902 623304 338958 623338
rect 338992 623304 339048 623338
rect 339082 623304 339138 623338
rect 339172 623304 339228 623338
rect 339262 623304 339318 623338
rect 339352 623304 339408 623338
rect 339442 623304 339496 623338
rect 338816 623248 339496 623304
rect 338816 623214 338868 623248
rect 338902 623214 338958 623248
rect 338992 623214 339048 623248
rect 339082 623214 339138 623248
rect 339172 623214 339228 623248
rect 339262 623214 339318 623248
rect 339352 623214 339408 623248
rect 339442 623214 339496 623248
rect 338816 623158 339496 623214
rect 338816 623124 338868 623158
rect 338902 623124 338958 623158
rect 338992 623124 339048 623158
rect 339082 623124 339138 623158
rect 339172 623124 339228 623158
rect 339262 623124 339318 623158
rect 339352 623124 339408 623158
rect 339442 623124 339496 623158
rect 338816 623068 339496 623124
rect 338816 623034 338868 623068
rect 338902 623034 338958 623068
rect 338992 623034 339048 623068
rect 339082 623034 339138 623068
rect 339172 623034 339228 623068
rect 339262 623034 339318 623068
rect 339352 623034 339408 623068
rect 339442 623034 339496 623068
rect 338816 622978 339496 623034
rect 338816 622944 338868 622978
rect 338902 622944 338958 622978
rect 338992 622944 339048 622978
rect 339082 622944 339138 622978
rect 339172 622944 339228 622978
rect 339262 622944 339318 622978
rect 339352 622944 339408 622978
rect 339442 622944 339496 622978
rect 338816 622892 339496 622944
rect 340104 623518 340784 623572
rect 340104 623484 340156 623518
rect 340190 623484 340246 623518
rect 340280 623484 340336 623518
rect 340370 623484 340426 623518
rect 340460 623484 340516 623518
rect 340550 623484 340606 623518
rect 340640 623484 340696 623518
rect 340730 623484 340784 623518
rect 340104 623428 340784 623484
rect 340104 623394 340156 623428
rect 340190 623394 340246 623428
rect 340280 623394 340336 623428
rect 340370 623394 340426 623428
rect 340460 623394 340516 623428
rect 340550 623394 340606 623428
rect 340640 623394 340696 623428
rect 340730 623394 340784 623428
rect 340104 623338 340784 623394
rect 340104 623304 340156 623338
rect 340190 623304 340246 623338
rect 340280 623304 340336 623338
rect 340370 623304 340426 623338
rect 340460 623304 340516 623338
rect 340550 623304 340606 623338
rect 340640 623304 340696 623338
rect 340730 623304 340784 623338
rect 340104 623248 340784 623304
rect 340104 623214 340156 623248
rect 340190 623214 340246 623248
rect 340280 623214 340336 623248
rect 340370 623214 340426 623248
rect 340460 623214 340516 623248
rect 340550 623214 340606 623248
rect 340640 623214 340696 623248
rect 340730 623214 340784 623248
rect 340104 623158 340784 623214
rect 340104 623124 340156 623158
rect 340190 623124 340246 623158
rect 340280 623124 340336 623158
rect 340370 623124 340426 623158
rect 340460 623124 340516 623158
rect 340550 623124 340606 623158
rect 340640 623124 340696 623158
rect 340730 623124 340784 623158
rect 340104 623068 340784 623124
rect 340104 623034 340156 623068
rect 340190 623034 340246 623068
rect 340280 623034 340336 623068
rect 340370 623034 340426 623068
rect 340460 623034 340516 623068
rect 340550 623034 340606 623068
rect 340640 623034 340696 623068
rect 340730 623034 340784 623068
rect 340104 622978 340784 623034
rect 340104 622944 340156 622978
rect 340190 622944 340246 622978
rect 340280 622944 340336 622978
rect 340370 622944 340426 622978
rect 340460 622944 340516 622978
rect 340550 622944 340606 622978
rect 340640 622944 340696 622978
rect 340730 622944 340784 622978
rect 340104 622892 340784 622944
rect 334952 622230 335632 622284
rect 334952 622196 335004 622230
rect 335038 622196 335094 622230
rect 335128 622196 335184 622230
rect 335218 622196 335274 622230
rect 335308 622196 335364 622230
rect 335398 622196 335454 622230
rect 335488 622196 335544 622230
rect 335578 622196 335632 622230
rect 334952 622140 335632 622196
rect 334952 622106 335004 622140
rect 335038 622106 335094 622140
rect 335128 622106 335184 622140
rect 335218 622106 335274 622140
rect 335308 622106 335364 622140
rect 335398 622106 335454 622140
rect 335488 622106 335544 622140
rect 335578 622106 335632 622140
rect 334952 622050 335632 622106
rect 334952 622016 335004 622050
rect 335038 622016 335094 622050
rect 335128 622016 335184 622050
rect 335218 622016 335274 622050
rect 335308 622016 335364 622050
rect 335398 622016 335454 622050
rect 335488 622016 335544 622050
rect 335578 622016 335632 622050
rect 334952 621960 335632 622016
rect 334952 621926 335004 621960
rect 335038 621926 335094 621960
rect 335128 621926 335184 621960
rect 335218 621926 335274 621960
rect 335308 621926 335364 621960
rect 335398 621926 335454 621960
rect 335488 621926 335544 621960
rect 335578 621926 335632 621960
rect 334952 621870 335632 621926
rect 334952 621836 335004 621870
rect 335038 621836 335094 621870
rect 335128 621836 335184 621870
rect 335218 621836 335274 621870
rect 335308 621836 335364 621870
rect 335398 621836 335454 621870
rect 335488 621836 335544 621870
rect 335578 621836 335632 621870
rect 334952 621780 335632 621836
rect 334952 621746 335004 621780
rect 335038 621746 335094 621780
rect 335128 621746 335184 621780
rect 335218 621746 335274 621780
rect 335308 621746 335364 621780
rect 335398 621746 335454 621780
rect 335488 621746 335544 621780
rect 335578 621746 335632 621780
rect 334952 621690 335632 621746
rect 334952 621656 335004 621690
rect 335038 621656 335094 621690
rect 335128 621656 335184 621690
rect 335218 621656 335274 621690
rect 335308 621656 335364 621690
rect 335398 621656 335454 621690
rect 335488 621656 335544 621690
rect 335578 621656 335632 621690
rect 334952 621604 335632 621656
rect 336240 622230 336920 622284
rect 336240 622196 336292 622230
rect 336326 622196 336382 622230
rect 336416 622196 336472 622230
rect 336506 622196 336562 622230
rect 336596 622196 336652 622230
rect 336686 622196 336742 622230
rect 336776 622196 336832 622230
rect 336866 622196 336920 622230
rect 336240 622140 336920 622196
rect 336240 622106 336292 622140
rect 336326 622106 336382 622140
rect 336416 622106 336472 622140
rect 336506 622106 336562 622140
rect 336596 622106 336652 622140
rect 336686 622106 336742 622140
rect 336776 622106 336832 622140
rect 336866 622106 336920 622140
rect 336240 622050 336920 622106
rect 336240 622016 336292 622050
rect 336326 622016 336382 622050
rect 336416 622016 336472 622050
rect 336506 622016 336562 622050
rect 336596 622016 336652 622050
rect 336686 622016 336742 622050
rect 336776 622016 336832 622050
rect 336866 622016 336920 622050
rect 336240 621960 336920 622016
rect 336240 621926 336292 621960
rect 336326 621926 336382 621960
rect 336416 621926 336472 621960
rect 336506 621926 336562 621960
rect 336596 621926 336652 621960
rect 336686 621926 336742 621960
rect 336776 621926 336832 621960
rect 336866 621926 336920 621960
rect 336240 621870 336920 621926
rect 336240 621836 336292 621870
rect 336326 621836 336382 621870
rect 336416 621836 336472 621870
rect 336506 621836 336562 621870
rect 336596 621836 336652 621870
rect 336686 621836 336742 621870
rect 336776 621836 336832 621870
rect 336866 621836 336920 621870
rect 336240 621780 336920 621836
rect 336240 621746 336292 621780
rect 336326 621746 336382 621780
rect 336416 621746 336472 621780
rect 336506 621746 336562 621780
rect 336596 621746 336652 621780
rect 336686 621746 336742 621780
rect 336776 621746 336832 621780
rect 336866 621746 336920 621780
rect 336240 621690 336920 621746
rect 336240 621656 336292 621690
rect 336326 621656 336382 621690
rect 336416 621656 336472 621690
rect 336506 621656 336562 621690
rect 336596 621656 336652 621690
rect 336686 621656 336742 621690
rect 336776 621656 336832 621690
rect 336866 621656 336920 621690
rect 336240 621604 336920 621656
rect 337528 622230 338208 622284
rect 337528 622196 337580 622230
rect 337614 622196 337670 622230
rect 337704 622196 337760 622230
rect 337794 622196 337850 622230
rect 337884 622196 337940 622230
rect 337974 622196 338030 622230
rect 338064 622196 338120 622230
rect 338154 622196 338208 622230
rect 337528 622140 338208 622196
rect 337528 622106 337580 622140
rect 337614 622106 337670 622140
rect 337704 622106 337760 622140
rect 337794 622106 337850 622140
rect 337884 622106 337940 622140
rect 337974 622106 338030 622140
rect 338064 622106 338120 622140
rect 338154 622106 338208 622140
rect 337528 622050 338208 622106
rect 337528 622016 337580 622050
rect 337614 622016 337670 622050
rect 337704 622016 337760 622050
rect 337794 622016 337850 622050
rect 337884 622016 337940 622050
rect 337974 622016 338030 622050
rect 338064 622016 338120 622050
rect 338154 622016 338208 622050
rect 337528 621960 338208 622016
rect 337528 621926 337580 621960
rect 337614 621926 337670 621960
rect 337704 621926 337760 621960
rect 337794 621926 337850 621960
rect 337884 621926 337940 621960
rect 337974 621926 338030 621960
rect 338064 621926 338120 621960
rect 338154 621926 338208 621960
rect 337528 621870 338208 621926
rect 337528 621836 337580 621870
rect 337614 621836 337670 621870
rect 337704 621836 337760 621870
rect 337794 621836 337850 621870
rect 337884 621836 337940 621870
rect 337974 621836 338030 621870
rect 338064 621836 338120 621870
rect 338154 621836 338208 621870
rect 337528 621780 338208 621836
rect 337528 621746 337580 621780
rect 337614 621746 337670 621780
rect 337704 621746 337760 621780
rect 337794 621746 337850 621780
rect 337884 621746 337940 621780
rect 337974 621746 338030 621780
rect 338064 621746 338120 621780
rect 338154 621746 338208 621780
rect 337528 621690 338208 621746
rect 337528 621656 337580 621690
rect 337614 621656 337670 621690
rect 337704 621656 337760 621690
rect 337794 621656 337850 621690
rect 337884 621656 337940 621690
rect 337974 621656 338030 621690
rect 338064 621656 338120 621690
rect 338154 621656 338208 621690
rect 337528 621604 338208 621656
rect 338816 622230 339496 622284
rect 338816 622196 338868 622230
rect 338902 622196 338958 622230
rect 338992 622196 339048 622230
rect 339082 622196 339138 622230
rect 339172 622196 339228 622230
rect 339262 622196 339318 622230
rect 339352 622196 339408 622230
rect 339442 622196 339496 622230
rect 338816 622140 339496 622196
rect 338816 622106 338868 622140
rect 338902 622106 338958 622140
rect 338992 622106 339048 622140
rect 339082 622106 339138 622140
rect 339172 622106 339228 622140
rect 339262 622106 339318 622140
rect 339352 622106 339408 622140
rect 339442 622106 339496 622140
rect 338816 622050 339496 622106
rect 338816 622016 338868 622050
rect 338902 622016 338958 622050
rect 338992 622016 339048 622050
rect 339082 622016 339138 622050
rect 339172 622016 339228 622050
rect 339262 622016 339318 622050
rect 339352 622016 339408 622050
rect 339442 622016 339496 622050
rect 338816 621960 339496 622016
rect 338816 621926 338868 621960
rect 338902 621926 338958 621960
rect 338992 621926 339048 621960
rect 339082 621926 339138 621960
rect 339172 621926 339228 621960
rect 339262 621926 339318 621960
rect 339352 621926 339408 621960
rect 339442 621926 339496 621960
rect 338816 621870 339496 621926
rect 338816 621836 338868 621870
rect 338902 621836 338958 621870
rect 338992 621836 339048 621870
rect 339082 621836 339138 621870
rect 339172 621836 339228 621870
rect 339262 621836 339318 621870
rect 339352 621836 339408 621870
rect 339442 621836 339496 621870
rect 338816 621780 339496 621836
rect 338816 621746 338868 621780
rect 338902 621746 338958 621780
rect 338992 621746 339048 621780
rect 339082 621746 339138 621780
rect 339172 621746 339228 621780
rect 339262 621746 339318 621780
rect 339352 621746 339408 621780
rect 339442 621746 339496 621780
rect 338816 621690 339496 621746
rect 338816 621656 338868 621690
rect 338902 621656 338958 621690
rect 338992 621656 339048 621690
rect 339082 621656 339138 621690
rect 339172 621656 339228 621690
rect 339262 621656 339318 621690
rect 339352 621656 339408 621690
rect 339442 621656 339496 621690
rect 338816 621604 339496 621656
rect 340104 622230 340784 622284
rect 340104 622196 340156 622230
rect 340190 622196 340246 622230
rect 340280 622196 340336 622230
rect 340370 622196 340426 622230
rect 340460 622196 340516 622230
rect 340550 622196 340606 622230
rect 340640 622196 340696 622230
rect 340730 622196 340784 622230
rect 340104 622140 340784 622196
rect 340104 622106 340156 622140
rect 340190 622106 340246 622140
rect 340280 622106 340336 622140
rect 340370 622106 340426 622140
rect 340460 622106 340516 622140
rect 340550 622106 340606 622140
rect 340640 622106 340696 622140
rect 340730 622106 340784 622140
rect 340104 622050 340784 622106
rect 340104 622016 340156 622050
rect 340190 622016 340246 622050
rect 340280 622016 340336 622050
rect 340370 622016 340426 622050
rect 340460 622016 340516 622050
rect 340550 622016 340606 622050
rect 340640 622016 340696 622050
rect 340730 622016 340784 622050
rect 340104 621960 340784 622016
rect 340104 621926 340156 621960
rect 340190 621926 340246 621960
rect 340280 621926 340336 621960
rect 340370 621926 340426 621960
rect 340460 621926 340516 621960
rect 340550 621926 340606 621960
rect 340640 621926 340696 621960
rect 340730 621926 340784 621960
rect 340104 621870 340784 621926
rect 340104 621836 340156 621870
rect 340190 621836 340246 621870
rect 340280 621836 340336 621870
rect 340370 621836 340426 621870
rect 340460 621836 340516 621870
rect 340550 621836 340606 621870
rect 340640 621836 340696 621870
rect 340730 621836 340784 621870
rect 340104 621780 340784 621836
rect 340104 621746 340156 621780
rect 340190 621746 340246 621780
rect 340280 621746 340336 621780
rect 340370 621746 340426 621780
rect 340460 621746 340516 621780
rect 340550 621746 340606 621780
rect 340640 621746 340696 621780
rect 340730 621746 340784 621780
rect 340104 621690 340784 621746
rect 340104 621656 340156 621690
rect 340190 621656 340246 621690
rect 340280 621656 340336 621690
rect 340370 621656 340426 621690
rect 340460 621656 340516 621690
rect 340550 621656 340606 621690
rect 340640 621656 340696 621690
rect 340730 621656 340784 621690
rect 340104 621604 340784 621656
rect 334952 620942 335632 620996
rect 334952 620908 335004 620942
rect 335038 620908 335094 620942
rect 335128 620908 335184 620942
rect 335218 620908 335274 620942
rect 335308 620908 335364 620942
rect 335398 620908 335454 620942
rect 335488 620908 335544 620942
rect 335578 620908 335632 620942
rect 334952 620852 335632 620908
rect 334952 620818 335004 620852
rect 335038 620818 335094 620852
rect 335128 620818 335184 620852
rect 335218 620818 335274 620852
rect 335308 620818 335364 620852
rect 335398 620818 335454 620852
rect 335488 620818 335544 620852
rect 335578 620818 335632 620852
rect 334952 620762 335632 620818
rect 334952 620728 335004 620762
rect 335038 620728 335094 620762
rect 335128 620728 335184 620762
rect 335218 620728 335274 620762
rect 335308 620728 335364 620762
rect 335398 620728 335454 620762
rect 335488 620728 335544 620762
rect 335578 620728 335632 620762
rect 334952 620672 335632 620728
rect 334952 620638 335004 620672
rect 335038 620638 335094 620672
rect 335128 620638 335184 620672
rect 335218 620638 335274 620672
rect 335308 620638 335364 620672
rect 335398 620638 335454 620672
rect 335488 620638 335544 620672
rect 335578 620638 335632 620672
rect 334952 620582 335632 620638
rect 334952 620548 335004 620582
rect 335038 620548 335094 620582
rect 335128 620548 335184 620582
rect 335218 620548 335274 620582
rect 335308 620548 335364 620582
rect 335398 620548 335454 620582
rect 335488 620548 335544 620582
rect 335578 620548 335632 620582
rect 334952 620492 335632 620548
rect 334952 620458 335004 620492
rect 335038 620458 335094 620492
rect 335128 620458 335184 620492
rect 335218 620458 335274 620492
rect 335308 620458 335364 620492
rect 335398 620458 335454 620492
rect 335488 620458 335544 620492
rect 335578 620458 335632 620492
rect 334952 620402 335632 620458
rect 334952 620368 335004 620402
rect 335038 620368 335094 620402
rect 335128 620368 335184 620402
rect 335218 620368 335274 620402
rect 335308 620368 335364 620402
rect 335398 620368 335454 620402
rect 335488 620368 335544 620402
rect 335578 620368 335632 620402
rect 334952 620316 335632 620368
rect 336240 620942 336920 620996
rect 336240 620908 336292 620942
rect 336326 620908 336382 620942
rect 336416 620908 336472 620942
rect 336506 620908 336562 620942
rect 336596 620908 336652 620942
rect 336686 620908 336742 620942
rect 336776 620908 336832 620942
rect 336866 620908 336920 620942
rect 336240 620852 336920 620908
rect 336240 620818 336292 620852
rect 336326 620818 336382 620852
rect 336416 620818 336472 620852
rect 336506 620818 336562 620852
rect 336596 620818 336652 620852
rect 336686 620818 336742 620852
rect 336776 620818 336832 620852
rect 336866 620818 336920 620852
rect 336240 620762 336920 620818
rect 336240 620728 336292 620762
rect 336326 620728 336382 620762
rect 336416 620728 336472 620762
rect 336506 620728 336562 620762
rect 336596 620728 336652 620762
rect 336686 620728 336742 620762
rect 336776 620728 336832 620762
rect 336866 620728 336920 620762
rect 336240 620672 336920 620728
rect 336240 620638 336292 620672
rect 336326 620638 336382 620672
rect 336416 620638 336472 620672
rect 336506 620638 336562 620672
rect 336596 620638 336652 620672
rect 336686 620638 336742 620672
rect 336776 620638 336832 620672
rect 336866 620638 336920 620672
rect 336240 620582 336920 620638
rect 336240 620548 336292 620582
rect 336326 620548 336382 620582
rect 336416 620548 336472 620582
rect 336506 620548 336562 620582
rect 336596 620548 336652 620582
rect 336686 620548 336742 620582
rect 336776 620548 336832 620582
rect 336866 620548 336920 620582
rect 336240 620492 336920 620548
rect 336240 620458 336292 620492
rect 336326 620458 336382 620492
rect 336416 620458 336472 620492
rect 336506 620458 336562 620492
rect 336596 620458 336652 620492
rect 336686 620458 336742 620492
rect 336776 620458 336832 620492
rect 336866 620458 336920 620492
rect 336240 620402 336920 620458
rect 336240 620368 336292 620402
rect 336326 620368 336382 620402
rect 336416 620368 336472 620402
rect 336506 620368 336562 620402
rect 336596 620368 336652 620402
rect 336686 620368 336742 620402
rect 336776 620368 336832 620402
rect 336866 620368 336920 620402
rect 336240 620316 336920 620368
rect 337528 620942 338208 620996
rect 337528 620908 337580 620942
rect 337614 620908 337670 620942
rect 337704 620908 337760 620942
rect 337794 620908 337850 620942
rect 337884 620908 337940 620942
rect 337974 620908 338030 620942
rect 338064 620908 338120 620942
rect 338154 620908 338208 620942
rect 337528 620852 338208 620908
rect 337528 620818 337580 620852
rect 337614 620818 337670 620852
rect 337704 620818 337760 620852
rect 337794 620818 337850 620852
rect 337884 620818 337940 620852
rect 337974 620818 338030 620852
rect 338064 620818 338120 620852
rect 338154 620818 338208 620852
rect 337528 620762 338208 620818
rect 337528 620728 337580 620762
rect 337614 620728 337670 620762
rect 337704 620728 337760 620762
rect 337794 620728 337850 620762
rect 337884 620728 337940 620762
rect 337974 620728 338030 620762
rect 338064 620728 338120 620762
rect 338154 620728 338208 620762
rect 337528 620672 338208 620728
rect 337528 620638 337580 620672
rect 337614 620638 337670 620672
rect 337704 620638 337760 620672
rect 337794 620638 337850 620672
rect 337884 620638 337940 620672
rect 337974 620638 338030 620672
rect 338064 620638 338120 620672
rect 338154 620638 338208 620672
rect 337528 620582 338208 620638
rect 337528 620548 337580 620582
rect 337614 620548 337670 620582
rect 337704 620548 337760 620582
rect 337794 620548 337850 620582
rect 337884 620548 337940 620582
rect 337974 620548 338030 620582
rect 338064 620548 338120 620582
rect 338154 620548 338208 620582
rect 337528 620492 338208 620548
rect 337528 620458 337580 620492
rect 337614 620458 337670 620492
rect 337704 620458 337760 620492
rect 337794 620458 337850 620492
rect 337884 620458 337940 620492
rect 337974 620458 338030 620492
rect 338064 620458 338120 620492
rect 338154 620458 338208 620492
rect 337528 620402 338208 620458
rect 337528 620368 337580 620402
rect 337614 620368 337670 620402
rect 337704 620368 337760 620402
rect 337794 620368 337850 620402
rect 337884 620368 337940 620402
rect 337974 620368 338030 620402
rect 338064 620368 338120 620402
rect 338154 620368 338208 620402
rect 337528 620316 338208 620368
rect 338816 620942 339496 620996
rect 338816 620908 338868 620942
rect 338902 620908 338958 620942
rect 338992 620908 339048 620942
rect 339082 620908 339138 620942
rect 339172 620908 339228 620942
rect 339262 620908 339318 620942
rect 339352 620908 339408 620942
rect 339442 620908 339496 620942
rect 338816 620852 339496 620908
rect 338816 620818 338868 620852
rect 338902 620818 338958 620852
rect 338992 620818 339048 620852
rect 339082 620818 339138 620852
rect 339172 620818 339228 620852
rect 339262 620818 339318 620852
rect 339352 620818 339408 620852
rect 339442 620818 339496 620852
rect 338816 620762 339496 620818
rect 338816 620728 338868 620762
rect 338902 620728 338958 620762
rect 338992 620728 339048 620762
rect 339082 620728 339138 620762
rect 339172 620728 339228 620762
rect 339262 620728 339318 620762
rect 339352 620728 339408 620762
rect 339442 620728 339496 620762
rect 338816 620672 339496 620728
rect 338816 620638 338868 620672
rect 338902 620638 338958 620672
rect 338992 620638 339048 620672
rect 339082 620638 339138 620672
rect 339172 620638 339228 620672
rect 339262 620638 339318 620672
rect 339352 620638 339408 620672
rect 339442 620638 339496 620672
rect 338816 620582 339496 620638
rect 338816 620548 338868 620582
rect 338902 620548 338958 620582
rect 338992 620548 339048 620582
rect 339082 620548 339138 620582
rect 339172 620548 339228 620582
rect 339262 620548 339318 620582
rect 339352 620548 339408 620582
rect 339442 620548 339496 620582
rect 338816 620492 339496 620548
rect 338816 620458 338868 620492
rect 338902 620458 338958 620492
rect 338992 620458 339048 620492
rect 339082 620458 339138 620492
rect 339172 620458 339228 620492
rect 339262 620458 339318 620492
rect 339352 620458 339408 620492
rect 339442 620458 339496 620492
rect 338816 620402 339496 620458
rect 338816 620368 338868 620402
rect 338902 620368 338958 620402
rect 338992 620368 339048 620402
rect 339082 620368 339138 620402
rect 339172 620368 339228 620402
rect 339262 620368 339318 620402
rect 339352 620368 339408 620402
rect 339442 620368 339496 620402
rect 338816 620316 339496 620368
rect 340104 620942 340784 620996
rect 340104 620908 340156 620942
rect 340190 620908 340246 620942
rect 340280 620908 340336 620942
rect 340370 620908 340426 620942
rect 340460 620908 340516 620942
rect 340550 620908 340606 620942
rect 340640 620908 340696 620942
rect 340730 620908 340784 620942
rect 340104 620852 340784 620908
rect 340104 620818 340156 620852
rect 340190 620818 340246 620852
rect 340280 620818 340336 620852
rect 340370 620818 340426 620852
rect 340460 620818 340516 620852
rect 340550 620818 340606 620852
rect 340640 620818 340696 620852
rect 340730 620818 340784 620852
rect 340104 620762 340784 620818
rect 340104 620728 340156 620762
rect 340190 620728 340246 620762
rect 340280 620728 340336 620762
rect 340370 620728 340426 620762
rect 340460 620728 340516 620762
rect 340550 620728 340606 620762
rect 340640 620728 340696 620762
rect 340730 620728 340784 620762
rect 340104 620672 340784 620728
rect 340104 620638 340156 620672
rect 340190 620638 340246 620672
rect 340280 620638 340336 620672
rect 340370 620638 340426 620672
rect 340460 620638 340516 620672
rect 340550 620638 340606 620672
rect 340640 620638 340696 620672
rect 340730 620638 340784 620672
rect 340104 620582 340784 620638
rect 340104 620548 340156 620582
rect 340190 620548 340246 620582
rect 340280 620548 340336 620582
rect 340370 620548 340426 620582
rect 340460 620548 340516 620582
rect 340550 620548 340606 620582
rect 340640 620548 340696 620582
rect 340730 620548 340784 620582
rect 340104 620492 340784 620548
rect 340104 620458 340156 620492
rect 340190 620458 340246 620492
rect 340280 620458 340336 620492
rect 340370 620458 340426 620492
rect 340460 620458 340516 620492
rect 340550 620458 340606 620492
rect 340640 620458 340696 620492
rect 340730 620458 340784 620492
rect 340104 620402 340784 620458
rect 340104 620368 340156 620402
rect 340190 620368 340246 620402
rect 340280 620368 340336 620402
rect 340370 620368 340426 620402
rect 340460 620368 340516 620402
rect 340550 620368 340606 620402
rect 340640 620368 340696 620402
rect 340730 620368 340784 620402
rect 340104 620316 340784 620368
rect 334952 619654 335632 619708
rect 334952 619620 335004 619654
rect 335038 619620 335094 619654
rect 335128 619620 335184 619654
rect 335218 619620 335274 619654
rect 335308 619620 335364 619654
rect 335398 619620 335454 619654
rect 335488 619620 335544 619654
rect 335578 619620 335632 619654
rect 334952 619564 335632 619620
rect 334952 619530 335004 619564
rect 335038 619530 335094 619564
rect 335128 619530 335184 619564
rect 335218 619530 335274 619564
rect 335308 619530 335364 619564
rect 335398 619530 335454 619564
rect 335488 619530 335544 619564
rect 335578 619530 335632 619564
rect 334952 619474 335632 619530
rect 334952 619440 335004 619474
rect 335038 619440 335094 619474
rect 335128 619440 335184 619474
rect 335218 619440 335274 619474
rect 335308 619440 335364 619474
rect 335398 619440 335454 619474
rect 335488 619440 335544 619474
rect 335578 619440 335632 619474
rect 334952 619384 335632 619440
rect 334952 619350 335004 619384
rect 335038 619350 335094 619384
rect 335128 619350 335184 619384
rect 335218 619350 335274 619384
rect 335308 619350 335364 619384
rect 335398 619350 335454 619384
rect 335488 619350 335544 619384
rect 335578 619350 335632 619384
rect 334952 619294 335632 619350
rect 334952 619260 335004 619294
rect 335038 619260 335094 619294
rect 335128 619260 335184 619294
rect 335218 619260 335274 619294
rect 335308 619260 335364 619294
rect 335398 619260 335454 619294
rect 335488 619260 335544 619294
rect 335578 619260 335632 619294
rect 334952 619204 335632 619260
rect 334952 619170 335004 619204
rect 335038 619170 335094 619204
rect 335128 619170 335184 619204
rect 335218 619170 335274 619204
rect 335308 619170 335364 619204
rect 335398 619170 335454 619204
rect 335488 619170 335544 619204
rect 335578 619170 335632 619204
rect 334952 619114 335632 619170
rect 334952 619080 335004 619114
rect 335038 619080 335094 619114
rect 335128 619080 335184 619114
rect 335218 619080 335274 619114
rect 335308 619080 335364 619114
rect 335398 619080 335454 619114
rect 335488 619080 335544 619114
rect 335578 619080 335632 619114
rect 334952 619028 335632 619080
rect 336240 619654 336920 619708
rect 336240 619620 336292 619654
rect 336326 619620 336382 619654
rect 336416 619620 336472 619654
rect 336506 619620 336562 619654
rect 336596 619620 336652 619654
rect 336686 619620 336742 619654
rect 336776 619620 336832 619654
rect 336866 619620 336920 619654
rect 336240 619564 336920 619620
rect 336240 619530 336292 619564
rect 336326 619530 336382 619564
rect 336416 619530 336472 619564
rect 336506 619530 336562 619564
rect 336596 619530 336652 619564
rect 336686 619530 336742 619564
rect 336776 619530 336832 619564
rect 336866 619530 336920 619564
rect 336240 619474 336920 619530
rect 336240 619440 336292 619474
rect 336326 619440 336382 619474
rect 336416 619440 336472 619474
rect 336506 619440 336562 619474
rect 336596 619440 336652 619474
rect 336686 619440 336742 619474
rect 336776 619440 336832 619474
rect 336866 619440 336920 619474
rect 336240 619384 336920 619440
rect 336240 619350 336292 619384
rect 336326 619350 336382 619384
rect 336416 619350 336472 619384
rect 336506 619350 336562 619384
rect 336596 619350 336652 619384
rect 336686 619350 336742 619384
rect 336776 619350 336832 619384
rect 336866 619350 336920 619384
rect 336240 619294 336920 619350
rect 336240 619260 336292 619294
rect 336326 619260 336382 619294
rect 336416 619260 336472 619294
rect 336506 619260 336562 619294
rect 336596 619260 336652 619294
rect 336686 619260 336742 619294
rect 336776 619260 336832 619294
rect 336866 619260 336920 619294
rect 336240 619204 336920 619260
rect 336240 619170 336292 619204
rect 336326 619170 336382 619204
rect 336416 619170 336472 619204
rect 336506 619170 336562 619204
rect 336596 619170 336652 619204
rect 336686 619170 336742 619204
rect 336776 619170 336832 619204
rect 336866 619170 336920 619204
rect 336240 619114 336920 619170
rect 336240 619080 336292 619114
rect 336326 619080 336382 619114
rect 336416 619080 336472 619114
rect 336506 619080 336562 619114
rect 336596 619080 336652 619114
rect 336686 619080 336742 619114
rect 336776 619080 336832 619114
rect 336866 619080 336920 619114
rect 336240 619028 336920 619080
rect 337528 619654 338208 619708
rect 337528 619620 337580 619654
rect 337614 619620 337670 619654
rect 337704 619620 337760 619654
rect 337794 619620 337850 619654
rect 337884 619620 337940 619654
rect 337974 619620 338030 619654
rect 338064 619620 338120 619654
rect 338154 619620 338208 619654
rect 337528 619564 338208 619620
rect 337528 619530 337580 619564
rect 337614 619530 337670 619564
rect 337704 619530 337760 619564
rect 337794 619530 337850 619564
rect 337884 619530 337940 619564
rect 337974 619530 338030 619564
rect 338064 619530 338120 619564
rect 338154 619530 338208 619564
rect 337528 619474 338208 619530
rect 337528 619440 337580 619474
rect 337614 619440 337670 619474
rect 337704 619440 337760 619474
rect 337794 619440 337850 619474
rect 337884 619440 337940 619474
rect 337974 619440 338030 619474
rect 338064 619440 338120 619474
rect 338154 619440 338208 619474
rect 337528 619384 338208 619440
rect 337528 619350 337580 619384
rect 337614 619350 337670 619384
rect 337704 619350 337760 619384
rect 337794 619350 337850 619384
rect 337884 619350 337940 619384
rect 337974 619350 338030 619384
rect 338064 619350 338120 619384
rect 338154 619350 338208 619384
rect 337528 619294 338208 619350
rect 337528 619260 337580 619294
rect 337614 619260 337670 619294
rect 337704 619260 337760 619294
rect 337794 619260 337850 619294
rect 337884 619260 337940 619294
rect 337974 619260 338030 619294
rect 338064 619260 338120 619294
rect 338154 619260 338208 619294
rect 337528 619204 338208 619260
rect 337528 619170 337580 619204
rect 337614 619170 337670 619204
rect 337704 619170 337760 619204
rect 337794 619170 337850 619204
rect 337884 619170 337940 619204
rect 337974 619170 338030 619204
rect 338064 619170 338120 619204
rect 338154 619170 338208 619204
rect 337528 619114 338208 619170
rect 337528 619080 337580 619114
rect 337614 619080 337670 619114
rect 337704 619080 337760 619114
rect 337794 619080 337850 619114
rect 337884 619080 337940 619114
rect 337974 619080 338030 619114
rect 338064 619080 338120 619114
rect 338154 619080 338208 619114
rect 337528 619028 338208 619080
rect 338816 619654 339496 619708
rect 338816 619620 338868 619654
rect 338902 619620 338958 619654
rect 338992 619620 339048 619654
rect 339082 619620 339138 619654
rect 339172 619620 339228 619654
rect 339262 619620 339318 619654
rect 339352 619620 339408 619654
rect 339442 619620 339496 619654
rect 338816 619564 339496 619620
rect 338816 619530 338868 619564
rect 338902 619530 338958 619564
rect 338992 619530 339048 619564
rect 339082 619530 339138 619564
rect 339172 619530 339228 619564
rect 339262 619530 339318 619564
rect 339352 619530 339408 619564
rect 339442 619530 339496 619564
rect 338816 619474 339496 619530
rect 338816 619440 338868 619474
rect 338902 619440 338958 619474
rect 338992 619440 339048 619474
rect 339082 619440 339138 619474
rect 339172 619440 339228 619474
rect 339262 619440 339318 619474
rect 339352 619440 339408 619474
rect 339442 619440 339496 619474
rect 338816 619384 339496 619440
rect 338816 619350 338868 619384
rect 338902 619350 338958 619384
rect 338992 619350 339048 619384
rect 339082 619350 339138 619384
rect 339172 619350 339228 619384
rect 339262 619350 339318 619384
rect 339352 619350 339408 619384
rect 339442 619350 339496 619384
rect 338816 619294 339496 619350
rect 338816 619260 338868 619294
rect 338902 619260 338958 619294
rect 338992 619260 339048 619294
rect 339082 619260 339138 619294
rect 339172 619260 339228 619294
rect 339262 619260 339318 619294
rect 339352 619260 339408 619294
rect 339442 619260 339496 619294
rect 338816 619204 339496 619260
rect 338816 619170 338868 619204
rect 338902 619170 338958 619204
rect 338992 619170 339048 619204
rect 339082 619170 339138 619204
rect 339172 619170 339228 619204
rect 339262 619170 339318 619204
rect 339352 619170 339408 619204
rect 339442 619170 339496 619204
rect 338816 619114 339496 619170
rect 338816 619080 338868 619114
rect 338902 619080 338958 619114
rect 338992 619080 339048 619114
rect 339082 619080 339138 619114
rect 339172 619080 339228 619114
rect 339262 619080 339318 619114
rect 339352 619080 339408 619114
rect 339442 619080 339496 619114
rect 338816 619028 339496 619080
rect 340104 619654 340784 619708
rect 340104 619620 340156 619654
rect 340190 619620 340246 619654
rect 340280 619620 340336 619654
rect 340370 619620 340426 619654
rect 340460 619620 340516 619654
rect 340550 619620 340606 619654
rect 340640 619620 340696 619654
rect 340730 619620 340784 619654
rect 340104 619564 340784 619620
rect 340104 619530 340156 619564
rect 340190 619530 340246 619564
rect 340280 619530 340336 619564
rect 340370 619530 340426 619564
rect 340460 619530 340516 619564
rect 340550 619530 340606 619564
rect 340640 619530 340696 619564
rect 340730 619530 340784 619564
rect 340104 619474 340784 619530
rect 340104 619440 340156 619474
rect 340190 619440 340246 619474
rect 340280 619440 340336 619474
rect 340370 619440 340426 619474
rect 340460 619440 340516 619474
rect 340550 619440 340606 619474
rect 340640 619440 340696 619474
rect 340730 619440 340784 619474
rect 340104 619384 340784 619440
rect 340104 619350 340156 619384
rect 340190 619350 340246 619384
rect 340280 619350 340336 619384
rect 340370 619350 340426 619384
rect 340460 619350 340516 619384
rect 340550 619350 340606 619384
rect 340640 619350 340696 619384
rect 340730 619350 340784 619384
rect 340104 619294 340784 619350
rect 340104 619260 340156 619294
rect 340190 619260 340246 619294
rect 340280 619260 340336 619294
rect 340370 619260 340426 619294
rect 340460 619260 340516 619294
rect 340550 619260 340606 619294
rect 340640 619260 340696 619294
rect 340730 619260 340784 619294
rect 340104 619204 340784 619260
rect 340104 619170 340156 619204
rect 340190 619170 340246 619204
rect 340280 619170 340336 619204
rect 340370 619170 340426 619204
rect 340460 619170 340516 619204
rect 340550 619170 340606 619204
rect 340640 619170 340696 619204
rect 340730 619170 340784 619204
rect 340104 619114 340784 619170
rect 340104 619080 340156 619114
rect 340190 619080 340246 619114
rect 340280 619080 340336 619114
rect 340370 619080 340426 619114
rect 340460 619080 340516 619114
rect 340550 619080 340606 619114
rect 340640 619080 340696 619114
rect 340730 619080 340784 619114
rect 340104 619028 340784 619080
rect 334952 618366 335632 618420
rect 334952 618332 335004 618366
rect 335038 618332 335094 618366
rect 335128 618332 335184 618366
rect 335218 618332 335274 618366
rect 335308 618332 335364 618366
rect 335398 618332 335454 618366
rect 335488 618332 335544 618366
rect 335578 618332 335632 618366
rect 334952 618276 335632 618332
rect 334952 618242 335004 618276
rect 335038 618242 335094 618276
rect 335128 618242 335184 618276
rect 335218 618242 335274 618276
rect 335308 618242 335364 618276
rect 335398 618242 335454 618276
rect 335488 618242 335544 618276
rect 335578 618242 335632 618276
rect 334952 618186 335632 618242
rect 334952 618152 335004 618186
rect 335038 618152 335094 618186
rect 335128 618152 335184 618186
rect 335218 618152 335274 618186
rect 335308 618152 335364 618186
rect 335398 618152 335454 618186
rect 335488 618152 335544 618186
rect 335578 618152 335632 618186
rect 334952 618096 335632 618152
rect 334952 618062 335004 618096
rect 335038 618062 335094 618096
rect 335128 618062 335184 618096
rect 335218 618062 335274 618096
rect 335308 618062 335364 618096
rect 335398 618062 335454 618096
rect 335488 618062 335544 618096
rect 335578 618062 335632 618096
rect 334952 618006 335632 618062
rect 334952 617972 335004 618006
rect 335038 617972 335094 618006
rect 335128 617972 335184 618006
rect 335218 617972 335274 618006
rect 335308 617972 335364 618006
rect 335398 617972 335454 618006
rect 335488 617972 335544 618006
rect 335578 617972 335632 618006
rect 334952 617916 335632 617972
rect 334952 617882 335004 617916
rect 335038 617882 335094 617916
rect 335128 617882 335184 617916
rect 335218 617882 335274 617916
rect 335308 617882 335364 617916
rect 335398 617882 335454 617916
rect 335488 617882 335544 617916
rect 335578 617882 335632 617916
rect 334952 617826 335632 617882
rect 334952 617792 335004 617826
rect 335038 617792 335094 617826
rect 335128 617792 335184 617826
rect 335218 617792 335274 617826
rect 335308 617792 335364 617826
rect 335398 617792 335454 617826
rect 335488 617792 335544 617826
rect 335578 617792 335632 617826
rect 334952 617740 335632 617792
rect 336240 618366 336920 618420
rect 336240 618332 336292 618366
rect 336326 618332 336382 618366
rect 336416 618332 336472 618366
rect 336506 618332 336562 618366
rect 336596 618332 336652 618366
rect 336686 618332 336742 618366
rect 336776 618332 336832 618366
rect 336866 618332 336920 618366
rect 336240 618276 336920 618332
rect 336240 618242 336292 618276
rect 336326 618242 336382 618276
rect 336416 618242 336472 618276
rect 336506 618242 336562 618276
rect 336596 618242 336652 618276
rect 336686 618242 336742 618276
rect 336776 618242 336832 618276
rect 336866 618242 336920 618276
rect 336240 618186 336920 618242
rect 336240 618152 336292 618186
rect 336326 618152 336382 618186
rect 336416 618152 336472 618186
rect 336506 618152 336562 618186
rect 336596 618152 336652 618186
rect 336686 618152 336742 618186
rect 336776 618152 336832 618186
rect 336866 618152 336920 618186
rect 336240 618096 336920 618152
rect 336240 618062 336292 618096
rect 336326 618062 336382 618096
rect 336416 618062 336472 618096
rect 336506 618062 336562 618096
rect 336596 618062 336652 618096
rect 336686 618062 336742 618096
rect 336776 618062 336832 618096
rect 336866 618062 336920 618096
rect 336240 618006 336920 618062
rect 336240 617972 336292 618006
rect 336326 617972 336382 618006
rect 336416 617972 336472 618006
rect 336506 617972 336562 618006
rect 336596 617972 336652 618006
rect 336686 617972 336742 618006
rect 336776 617972 336832 618006
rect 336866 617972 336920 618006
rect 336240 617916 336920 617972
rect 336240 617882 336292 617916
rect 336326 617882 336382 617916
rect 336416 617882 336472 617916
rect 336506 617882 336562 617916
rect 336596 617882 336652 617916
rect 336686 617882 336742 617916
rect 336776 617882 336832 617916
rect 336866 617882 336920 617916
rect 336240 617826 336920 617882
rect 336240 617792 336292 617826
rect 336326 617792 336382 617826
rect 336416 617792 336472 617826
rect 336506 617792 336562 617826
rect 336596 617792 336652 617826
rect 336686 617792 336742 617826
rect 336776 617792 336832 617826
rect 336866 617792 336920 617826
rect 336240 617740 336920 617792
rect 337528 618366 338208 618420
rect 337528 618332 337580 618366
rect 337614 618332 337670 618366
rect 337704 618332 337760 618366
rect 337794 618332 337850 618366
rect 337884 618332 337940 618366
rect 337974 618332 338030 618366
rect 338064 618332 338120 618366
rect 338154 618332 338208 618366
rect 337528 618276 338208 618332
rect 337528 618242 337580 618276
rect 337614 618242 337670 618276
rect 337704 618242 337760 618276
rect 337794 618242 337850 618276
rect 337884 618242 337940 618276
rect 337974 618242 338030 618276
rect 338064 618242 338120 618276
rect 338154 618242 338208 618276
rect 337528 618186 338208 618242
rect 337528 618152 337580 618186
rect 337614 618152 337670 618186
rect 337704 618152 337760 618186
rect 337794 618152 337850 618186
rect 337884 618152 337940 618186
rect 337974 618152 338030 618186
rect 338064 618152 338120 618186
rect 338154 618152 338208 618186
rect 337528 618096 338208 618152
rect 337528 618062 337580 618096
rect 337614 618062 337670 618096
rect 337704 618062 337760 618096
rect 337794 618062 337850 618096
rect 337884 618062 337940 618096
rect 337974 618062 338030 618096
rect 338064 618062 338120 618096
rect 338154 618062 338208 618096
rect 337528 618006 338208 618062
rect 337528 617972 337580 618006
rect 337614 617972 337670 618006
rect 337704 617972 337760 618006
rect 337794 617972 337850 618006
rect 337884 617972 337940 618006
rect 337974 617972 338030 618006
rect 338064 617972 338120 618006
rect 338154 617972 338208 618006
rect 337528 617916 338208 617972
rect 337528 617882 337580 617916
rect 337614 617882 337670 617916
rect 337704 617882 337760 617916
rect 337794 617882 337850 617916
rect 337884 617882 337940 617916
rect 337974 617882 338030 617916
rect 338064 617882 338120 617916
rect 338154 617882 338208 617916
rect 337528 617826 338208 617882
rect 337528 617792 337580 617826
rect 337614 617792 337670 617826
rect 337704 617792 337760 617826
rect 337794 617792 337850 617826
rect 337884 617792 337940 617826
rect 337974 617792 338030 617826
rect 338064 617792 338120 617826
rect 338154 617792 338208 617826
rect 337528 617740 338208 617792
rect 338816 618366 339496 618420
rect 338816 618332 338868 618366
rect 338902 618332 338958 618366
rect 338992 618332 339048 618366
rect 339082 618332 339138 618366
rect 339172 618332 339228 618366
rect 339262 618332 339318 618366
rect 339352 618332 339408 618366
rect 339442 618332 339496 618366
rect 338816 618276 339496 618332
rect 338816 618242 338868 618276
rect 338902 618242 338958 618276
rect 338992 618242 339048 618276
rect 339082 618242 339138 618276
rect 339172 618242 339228 618276
rect 339262 618242 339318 618276
rect 339352 618242 339408 618276
rect 339442 618242 339496 618276
rect 338816 618186 339496 618242
rect 338816 618152 338868 618186
rect 338902 618152 338958 618186
rect 338992 618152 339048 618186
rect 339082 618152 339138 618186
rect 339172 618152 339228 618186
rect 339262 618152 339318 618186
rect 339352 618152 339408 618186
rect 339442 618152 339496 618186
rect 338816 618096 339496 618152
rect 338816 618062 338868 618096
rect 338902 618062 338958 618096
rect 338992 618062 339048 618096
rect 339082 618062 339138 618096
rect 339172 618062 339228 618096
rect 339262 618062 339318 618096
rect 339352 618062 339408 618096
rect 339442 618062 339496 618096
rect 338816 618006 339496 618062
rect 338816 617972 338868 618006
rect 338902 617972 338958 618006
rect 338992 617972 339048 618006
rect 339082 617972 339138 618006
rect 339172 617972 339228 618006
rect 339262 617972 339318 618006
rect 339352 617972 339408 618006
rect 339442 617972 339496 618006
rect 338816 617916 339496 617972
rect 338816 617882 338868 617916
rect 338902 617882 338958 617916
rect 338992 617882 339048 617916
rect 339082 617882 339138 617916
rect 339172 617882 339228 617916
rect 339262 617882 339318 617916
rect 339352 617882 339408 617916
rect 339442 617882 339496 617916
rect 338816 617826 339496 617882
rect 338816 617792 338868 617826
rect 338902 617792 338958 617826
rect 338992 617792 339048 617826
rect 339082 617792 339138 617826
rect 339172 617792 339228 617826
rect 339262 617792 339318 617826
rect 339352 617792 339408 617826
rect 339442 617792 339496 617826
rect 338816 617740 339496 617792
rect 340104 618366 340784 618420
rect 340104 618332 340156 618366
rect 340190 618332 340246 618366
rect 340280 618332 340336 618366
rect 340370 618332 340426 618366
rect 340460 618332 340516 618366
rect 340550 618332 340606 618366
rect 340640 618332 340696 618366
rect 340730 618332 340784 618366
rect 340104 618276 340784 618332
rect 340104 618242 340156 618276
rect 340190 618242 340246 618276
rect 340280 618242 340336 618276
rect 340370 618242 340426 618276
rect 340460 618242 340516 618276
rect 340550 618242 340606 618276
rect 340640 618242 340696 618276
rect 340730 618242 340784 618276
rect 340104 618186 340784 618242
rect 340104 618152 340156 618186
rect 340190 618152 340246 618186
rect 340280 618152 340336 618186
rect 340370 618152 340426 618186
rect 340460 618152 340516 618186
rect 340550 618152 340606 618186
rect 340640 618152 340696 618186
rect 340730 618152 340784 618186
rect 340104 618096 340784 618152
rect 340104 618062 340156 618096
rect 340190 618062 340246 618096
rect 340280 618062 340336 618096
rect 340370 618062 340426 618096
rect 340460 618062 340516 618096
rect 340550 618062 340606 618096
rect 340640 618062 340696 618096
rect 340730 618062 340784 618096
rect 340104 618006 340784 618062
rect 340104 617972 340156 618006
rect 340190 617972 340246 618006
rect 340280 617972 340336 618006
rect 340370 617972 340426 618006
rect 340460 617972 340516 618006
rect 340550 617972 340606 618006
rect 340640 617972 340696 618006
rect 340730 617972 340784 618006
rect 340104 617916 340784 617972
rect 340104 617882 340156 617916
rect 340190 617882 340246 617916
rect 340280 617882 340336 617916
rect 340370 617882 340426 617916
rect 340460 617882 340516 617916
rect 340550 617882 340606 617916
rect 340640 617882 340696 617916
rect 340730 617882 340784 617916
rect 340104 617826 340784 617882
rect 340104 617792 340156 617826
rect 340190 617792 340246 617826
rect 340280 617792 340336 617826
rect 340370 617792 340426 617826
rect 340460 617792 340516 617826
rect 340550 617792 340606 617826
rect 340640 617792 340696 617826
rect 340730 617792 340784 617826
rect 340104 617740 340784 617792
rect 329888 617206 329946 617218
rect 311478 617168 311536 617180
<< ndiffc >>
rect 305040 624324 310416 624358
rect 305040 623866 310416 623900
rect 300392 620650 300426 621026
rect 300850 620650 300884 621026
rect 301308 620650 301342 621026
rect 301766 620650 301800 621026
rect 302224 620650 302258 621026
rect 302682 620650 302716 621026
rect 303140 620650 303174 621026
rect 305322 620372 305356 622148
rect 305780 620372 305814 622148
rect 305894 620372 305928 622148
rect 306352 620372 306386 622148
rect 306466 620372 306500 622148
rect 306924 620372 306958 622148
rect 307038 620372 307072 622148
rect 307496 620372 307530 622148
rect 307610 620372 307644 622148
rect 308068 620372 308102 622148
rect 308182 620372 308216 622148
rect 308640 620372 308674 622148
rect 308754 620372 308788 622148
rect 309212 620372 309246 622148
rect 309326 620372 309360 622148
rect 309784 620372 309818 622148
<< pdiffc >>
rect 335004 627348 335038 627382
rect 335094 627348 335128 627382
rect 335184 627348 335218 627382
rect 335274 627348 335308 627382
rect 335364 627348 335398 627382
rect 335454 627348 335488 627382
rect 335544 627348 335578 627382
rect 335004 627258 335038 627292
rect 335094 627258 335128 627292
rect 335184 627258 335218 627292
rect 335274 627258 335308 627292
rect 335364 627258 335398 627292
rect 335454 627258 335488 627292
rect 335544 627258 335578 627292
rect 335004 627168 335038 627202
rect 335094 627168 335128 627202
rect 335184 627168 335218 627202
rect 335274 627168 335308 627202
rect 335364 627168 335398 627202
rect 335454 627168 335488 627202
rect 335544 627168 335578 627202
rect 335004 627078 335038 627112
rect 335094 627078 335128 627112
rect 335184 627078 335218 627112
rect 335274 627078 335308 627112
rect 335364 627078 335398 627112
rect 335454 627078 335488 627112
rect 335544 627078 335578 627112
rect 335004 626988 335038 627022
rect 335094 626988 335128 627022
rect 335184 626988 335218 627022
rect 335274 626988 335308 627022
rect 335364 626988 335398 627022
rect 335454 626988 335488 627022
rect 335544 626988 335578 627022
rect 335004 626898 335038 626932
rect 335094 626898 335128 626932
rect 335184 626898 335218 626932
rect 335274 626898 335308 626932
rect 335364 626898 335398 626932
rect 335454 626898 335488 626932
rect 335544 626898 335578 626932
rect 335004 626808 335038 626842
rect 335094 626808 335128 626842
rect 335184 626808 335218 626842
rect 335274 626808 335308 626842
rect 335364 626808 335398 626842
rect 335454 626808 335488 626842
rect 335544 626808 335578 626842
rect 336292 627348 336326 627382
rect 336382 627348 336416 627382
rect 336472 627348 336506 627382
rect 336562 627348 336596 627382
rect 336652 627348 336686 627382
rect 336742 627348 336776 627382
rect 336832 627348 336866 627382
rect 336292 627258 336326 627292
rect 336382 627258 336416 627292
rect 336472 627258 336506 627292
rect 336562 627258 336596 627292
rect 336652 627258 336686 627292
rect 336742 627258 336776 627292
rect 336832 627258 336866 627292
rect 336292 627168 336326 627202
rect 336382 627168 336416 627202
rect 336472 627168 336506 627202
rect 336562 627168 336596 627202
rect 336652 627168 336686 627202
rect 336742 627168 336776 627202
rect 336832 627168 336866 627202
rect 336292 627078 336326 627112
rect 336382 627078 336416 627112
rect 336472 627078 336506 627112
rect 336562 627078 336596 627112
rect 336652 627078 336686 627112
rect 336742 627078 336776 627112
rect 336832 627078 336866 627112
rect 336292 626988 336326 627022
rect 336382 626988 336416 627022
rect 336472 626988 336506 627022
rect 336562 626988 336596 627022
rect 336652 626988 336686 627022
rect 336742 626988 336776 627022
rect 336832 626988 336866 627022
rect 336292 626898 336326 626932
rect 336382 626898 336416 626932
rect 336472 626898 336506 626932
rect 336562 626898 336596 626932
rect 336652 626898 336686 626932
rect 336742 626898 336776 626932
rect 336832 626898 336866 626932
rect 336292 626808 336326 626842
rect 336382 626808 336416 626842
rect 336472 626808 336506 626842
rect 336562 626808 336596 626842
rect 336652 626808 336686 626842
rect 336742 626808 336776 626842
rect 336832 626808 336866 626842
rect 337580 627348 337614 627382
rect 337670 627348 337704 627382
rect 337760 627348 337794 627382
rect 337850 627348 337884 627382
rect 337940 627348 337974 627382
rect 338030 627348 338064 627382
rect 338120 627348 338154 627382
rect 337580 627258 337614 627292
rect 337670 627258 337704 627292
rect 337760 627258 337794 627292
rect 337850 627258 337884 627292
rect 337940 627258 337974 627292
rect 338030 627258 338064 627292
rect 338120 627258 338154 627292
rect 337580 627168 337614 627202
rect 337670 627168 337704 627202
rect 337760 627168 337794 627202
rect 337850 627168 337884 627202
rect 337940 627168 337974 627202
rect 338030 627168 338064 627202
rect 338120 627168 338154 627202
rect 337580 627078 337614 627112
rect 337670 627078 337704 627112
rect 337760 627078 337794 627112
rect 337850 627078 337884 627112
rect 337940 627078 337974 627112
rect 338030 627078 338064 627112
rect 338120 627078 338154 627112
rect 337580 626988 337614 627022
rect 337670 626988 337704 627022
rect 337760 626988 337794 627022
rect 337850 626988 337884 627022
rect 337940 626988 337974 627022
rect 338030 626988 338064 627022
rect 338120 626988 338154 627022
rect 337580 626898 337614 626932
rect 337670 626898 337704 626932
rect 337760 626898 337794 626932
rect 337850 626898 337884 626932
rect 337940 626898 337974 626932
rect 338030 626898 338064 626932
rect 338120 626898 338154 626932
rect 337580 626808 337614 626842
rect 337670 626808 337704 626842
rect 337760 626808 337794 626842
rect 337850 626808 337884 626842
rect 337940 626808 337974 626842
rect 338030 626808 338064 626842
rect 338120 626808 338154 626842
rect 338868 627348 338902 627382
rect 338958 627348 338992 627382
rect 339048 627348 339082 627382
rect 339138 627348 339172 627382
rect 339228 627348 339262 627382
rect 339318 627348 339352 627382
rect 339408 627348 339442 627382
rect 338868 627258 338902 627292
rect 338958 627258 338992 627292
rect 339048 627258 339082 627292
rect 339138 627258 339172 627292
rect 339228 627258 339262 627292
rect 339318 627258 339352 627292
rect 339408 627258 339442 627292
rect 338868 627168 338902 627202
rect 338958 627168 338992 627202
rect 339048 627168 339082 627202
rect 339138 627168 339172 627202
rect 339228 627168 339262 627202
rect 339318 627168 339352 627202
rect 339408 627168 339442 627202
rect 338868 627078 338902 627112
rect 338958 627078 338992 627112
rect 339048 627078 339082 627112
rect 339138 627078 339172 627112
rect 339228 627078 339262 627112
rect 339318 627078 339352 627112
rect 339408 627078 339442 627112
rect 338868 626988 338902 627022
rect 338958 626988 338992 627022
rect 339048 626988 339082 627022
rect 339138 626988 339172 627022
rect 339228 626988 339262 627022
rect 339318 626988 339352 627022
rect 339408 626988 339442 627022
rect 338868 626898 338902 626932
rect 338958 626898 338992 626932
rect 339048 626898 339082 626932
rect 339138 626898 339172 626932
rect 339228 626898 339262 626932
rect 339318 626898 339352 626932
rect 339408 626898 339442 626932
rect 338868 626808 338902 626842
rect 338958 626808 338992 626842
rect 339048 626808 339082 626842
rect 339138 626808 339172 626842
rect 339228 626808 339262 626842
rect 339318 626808 339352 626842
rect 339408 626808 339442 626842
rect 340156 627348 340190 627382
rect 340246 627348 340280 627382
rect 340336 627348 340370 627382
rect 340426 627348 340460 627382
rect 340516 627348 340550 627382
rect 340606 627348 340640 627382
rect 340696 627348 340730 627382
rect 340156 627258 340190 627292
rect 340246 627258 340280 627292
rect 340336 627258 340370 627292
rect 340426 627258 340460 627292
rect 340516 627258 340550 627292
rect 340606 627258 340640 627292
rect 340696 627258 340730 627292
rect 340156 627168 340190 627202
rect 340246 627168 340280 627202
rect 340336 627168 340370 627202
rect 340426 627168 340460 627202
rect 340516 627168 340550 627202
rect 340606 627168 340640 627202
rect 340696 627168 340730 627202
rect 340156 627078 340190 627112
rect 340246 627078 340280 627112
rect 340336 627078 340370 627112
rect 340426 627078 340460 627112
rect 340516 627078 340550 627112
rect 340606 627078 340640 627112
rect 340696 627078 340730 627112
rect 340156 626988 340190 627022
rect 340246 626988 340280 627022
rect 340336 626988 340370 627022
rect 340426 626988 340460 627022
rect 340516 626988 340550 627022
rect 340606 626988 340640 627022
rect 340696 626988 340730 627022
rect 340156 626898 340190 626932
rect 340246 626898 340280 626932
rect 340336 626898 340370 626932
rect 340426 626898 340460 626932
rect 340516 626898 340550 626932
rect 340606 626898 340640 626932
rect 340696 626898 340730 626932
rect 340156 626808 340190 626842
rect 340246 626808 340280 626842
rect 340336 626808 340370 626842
rect 340426 626808 340460 626842
rect 340516 626808 340550 626842
rect 340606 626808 340640 626842
rect 340696 626808 340730 626842
rect 335004 626060 335038 626094
rect 335094 626060 335128 626094
rect 335184 626060 335218 626094
rect 335274 626060 335308 626094
rect 335364 626060 335398 626094
rect 335454 626060 335488 626094
rect 335544 626060 335578 626094
rect 335004 625970 335038 626004
rect 335094 625970 335128 626004
rect 335184 625970 335218 626004
rect 335274 625970 335308 626004
rect 335364 625970 335398 626004
rect 335454 625970 335488 626004
rect 335544 625970 335578 626004
rect 335004 625880 335038 625914
rect 335094 625880 335128 625914
rect 335184 625880 335218 625914
rect 335274 625880 335308 625914
rect 335364 625880 335398 625914
rect 335454 625880 335488 625914
rect 335544 625880 335578 625914
rect 335004 625790 335038 625824
rect 335094 625790 335128 625824
rect 335184 625790 335218 625824
rect 335274 625790 335308 625824
rect 335364 625790 335398 625824
rect 335454 625790 335488 625824
rect 335544 625790 335578 625824
rect 335004 625700 335038 625734
rect 335094 625700 335128 625734
rect 335184 625700 335218 625734
rect 335274 625700 335308 625734
rect 335364 625700 335398 625734
rect 335454 625700 335488 625734
rect 335544 625700 335578 625734
rect 335004 625610 335038 625644
rect 335094 625610 335128 625644
rect 335184 625610 335218 625644
rect 335274 625610 335308 625644
rect 335364 625610 335398 625644
rect 335454 625610 335488 625644
rect 335544 625610 335578 625644
rect 335004 625520 335038 625554
rect 335094 625520 335128 625554
rect 335184 625520 335218 625554
rect 335274 625520 335308 625554
rect 335364 625520 335398 625554
rect 335454 625520 335488 625554
rect 335544 625520 335578 625554
rect 336292 626060 336326 626094
rect 336382 626060 336416 626094
rect 336472 626060 336506 626094
rect 336562 626060 336596 626094
rect 336652 626060 336686 626094
rect 336742 626060 336776 626094
rect 336832 626060 336866 626094
rect 336292 625970 336326 626004
rect 336382 625970 336416 626004
rect 336472 625970 336506 626004
rect 336562 625970 336596 626004
rect 336652 625970 336686 626004
rect 336742 625970 336776 626004
rect 336832 625970 336866 626004
rect 336292 625880 336326 625914
rect 336382 625880 336416 625914
rect 336472 625880 336506 625914
rect 336562 625880 336596 625914
rect 336652 625880 336686 625914
rect 336742 625880 336776 625914
rect 336832 625880 336866 625914
rect 336292 625790 336326 625824
rect 336382 625790 336416 625824
rect 336472 625790 336506 625824
rect 336562 625790 336596 625824
rect 336652 625790 336686 625824
rect 336742 625790 336776 625824
rect 336832 625790 336866 625824
rect 336292 625700 336326 625734
rect 336382 625700 336416 625734
rect 336472 625700 336506 625734
rect 336562 625700 336596 625734
rect 336652 625700 336686 625734
rect 336742 625700 336776 625734
rect 336832 625700 336866 625734
rect 336292 625610 336326 625644
rect 336382 625610 336416 625644
rect 336472 625610 336506 625644
rect 336562 625610 336596 625644
rect 336652 625610 336686 625644
rect 336742 625610 336776 625644
rect 336832 625610 336866 625644
rect 336292 625520 336326 625554
rect 336382 625520 336416 625554
rect 336472 625520 336506 625554
rect 336562 625520 336596 625554
rect 336652 625520 336686 625554
rect 336742 625520 336776 625554
rect 336832 625520 336866 625554
rect 337580 626060 337614 626094
rect 337670 626060 337704 626094
rect 337760 626060 337794 626094
rect 337850 626060 337884 626094
rect 337940 626060 337974 626094
rect 338030 626060 338064 626094
rect 338120 626060 338154 626094
rect 337580 625970 337614 626004
rect 337670 625970 337704 626004
rect 337760 625970 337794 626004
rect 337850 625970 337884 626004
rect 337940 625970 337974 626004
rect 338030 625970 338064 626004
rect 338120 625970 338154 626004
rect 337580 625880 337614 625914
rect 337670 625880 337704 625914
rect 337760 625880 337794 625914
rect 337850 625880 337884 625914
rect 337940 625880 337974 625914
rect 338030 625880 338064 625914
rect 338120 625880 338154 625914
rect 337580 625790 337614 625824
rect 337670 625790 337704 625824
rect 337760 625790 337794 625824
rect 337850 625790 337884 625824
rect 337940 625790 337974 625824
rect 338030 625790 338064 625824
rect 338120 625790 338154 625824
rect 337580 625700 337614 625734
rect 337670 625700 337704 625734
rect 337760 625700 337794 625734
rect 337850 625700 337884 625734
rect 337940 625700 337974 625734
rect 338030 625700 338064 625734
rect 338120 625700 338154 625734
rect 337580 625610 337614 625644
rect 337670 625610 337704 625644
rect 337760 625610 337794 625644
rect 337850 625610 337884 625644
rect 337940 625610 337974 625644
rect 338030 625610 338064 625644
rect 338120 625610 338154 625644
rect 337580 625520 337614 625554
rect 337670 625520 337704 625554
rect 337760 625520 337794 625554
rect 337850 625520 337884 625554
rect 337940 625520 337974 625554
rect 338030 625520 338064 625554
rect 338120 625520 338154 625554
rect 338868 626060 338902 626094
rect 338958 626060 338992 626094
rect 339048 626060 339082 626094
rect 339138 626060 339172 626094
rect 339228 626060 339262 626094
rect 339318 626060 339352 626094
rect 339408 626060 339442 626094
rect 338868 625970 338902 626004
rect 338958 625970 338992 626004
rect 339048 625970 339082 626004
rect 339138 625970 339172 626004
rect 339228 625970 339262 626004
rect 339318 625970 339352 626004
rect 339408 625970 339442 626004
rect 338868 625880 338902 625914
rect 338958 625880 338992 625914
rect 339048 625880 339082 625914
rect 339138 625880 339172 625914
rect 339228 625880 339262 625914
rect 339318 625880 339352 625914
rect 339408 625880 339442 625914
rect 338868 625790 338902 625824
rect 338958 625790 338992 625824
rect 339048 625790 339082 625824
rect 339138 625790 339172 625824
rect 339228 625790 339262 625824
rect 339318 625790 339352 625824
rect 339408 625790 339442 625824
rect 338868 625700 338902 625734
rect 338958 625700 338992 625734
rect 339048 625700 339082 625734
rect 339138 625700 339172 625734
rect 339228 625700 339262 625734
rect 339318 625700 339352 625734
rect 339408 625700 339442 625734
rect 338868 625610 338902 625644
rect 338958 625610 338992 625644
rect 339048 625610 339082 625644
rect 339138 625610 339172 625644
rect 339228 625610 339262 625644
rect 339318 625610 339352 625644
rect 339408 625610 339442 625644
rect 338868 625520 338902 625554
rect 338958 625520 338992 625554
rect 339048 625520 339082 625554
rect 339138 625520 339172 625554
rect 339228 625520 339262 625554
rect 339318 625520 339352 625554
rect 339408 625520 339442 625554
rect 340156 626060 340190 626094
rect 340246 626060 340280 626094
rect 340336 626060 340370 626094
rect 340426 626060 340460 626094
rect 340516 626060 340550 626094
rect 340606 626060 340640 626094
rect 340696 626060 340730 626094
rect 340156 625970 340190 626004
rect 340246 625970 340280 626004
rect 340336 625970 340370 626004
rect 340426 625970 340460 626004
rect 340516 625970 340550 626004
rect 340606 625970 340640 626004
rect 340696 625970 340730 626004
rect 340156 625880 340190 625914
rect 340246 625880 340280 625914
rect 340336 625880 340370 625914
rect 340426 625880 340460 625914
rect 340516 625880 340550 625914
rect 340606 625880 340640 625914
rect 340696 625880 340730 625914
rect 340156 625790 340190 625824
rect 340246 625790 340280 625824
rect 340336 625790 340370 625824
rect 340426 625790 340460 625824
rect 340516 625790 340550 625824
rect 340606 625790 340640 625824
rect 340696 625790 340730 625824
rect 340156 625700 340190 625734
rect 340246 625700 340280 625734
rect 340336 625700 340370 625734
rect 340426 625700 340460 625734
rect 340516 625700 340550 625734
rect 340606 625700 340640 625734
rect 340696 625700 340730 625734
rect 340156 625610 340190 625644
rect 340246 625610 340280 625644
rect 340336 625610 340370 625644
rect 340426 625610 340460 625644
rect 340516 625610 340550 625644
rect 340606 625610 340640 625644
rect 340696 625610 340730 625644
rect 340156 625520 340190 625554
rect 340246 625520 340280 625554
rect 340336 625520 340370 625554
rect 340426 625520 340460 625554
rect 340516 625520 340550 625554
rect 340606 625520 340640 625554
rect 340696 625520 340730 625554
rect 303596 617180 303630 619736
rect 304054 617180 304088 619736
rect 304168 617180 304202 619736
rect 304626 617180 304660 619736
rect 304740 617180 304774 619736
rect 305198 617180 305232 619736
rect 305312 617180 305346 619736
rect 305770 617180 305804 619736
rect 305884 617180 305918 619736
rect 306342 617180 306376 619736
rect 306456 617180 306490 619736
rect 306914 617180 306948 619736
rect 307028 617180 307062 619736
rect 307486 617180 307520 619736
rect 307600 617180 307634 619736
rect 308058 617180 308092 619736
rect 308172 617180 308206 619736
rect 308630 617180 308664 619736
rect 308744 617180 308778 619736
rect 309202 617180 309236 619736
rect 309316 617180 309350 619736
rect 309774 617180 309808 619736
rect 309888 617180 309922 619736
rect 310346 617180 310380 619736
rect 310460 617180 310494 619736
rect 310918 617180 310952 619736
rect 311032 617180 311066 619736
rect 311490 617180 311524 619736
rect 313404 617218 313438 624934
rect 313862 617218 313896 624934
rect 314320 617218 314354 624934
rect 314778 617218 314812 624934
rect 315236 617218 315270 624934
rect 315694 617218 315728 624934
rect 316152 617218 316186 624934
rect 316610 617218 316644 624934
rect 317068 617218 317102 624934
rect 317526 617218 317560 624934
rect 317984 617218 318018 624934
rect 318442 617218 318476 624934
rect 319362 617218 319396 624934
rect 319820 617218 319854 624934
rect 320278 617218 320312 624934
rect 320736 617218 320770 624934
rect 321194 617218 321228 624934
rect 321652 617218 321686 624934
rect 322110 617218 322144 624934
rect 322568 617218 322602 624934
rect 323026 617218 323060 624934
rect 323484 617218 323518 624934
rect 323942 617218 323976 624934
rect 324862 617218 324896 624934
rect 325320 617218 325354 624934
rect 325778 617218 325812 624934
rect 326236 617218 326270 624934
rect 326694 617218 326728 624934
rect 327152 617218 327186 624934
rect 327610 617218 327644 624934
rect 328068 617218 328102 624934
rect 328526 617218 328560 624934
rect 328984 617218 329018 624934
rect 329442 617218 329476 624934
rect 329900 617218 329934 624934
rect 335004 624772 335038 624806
rect 335094 624772 335128 624806
rect 335184 624772 335218 624806
rect 335274 624772 335308 624806
rect 335364 624772 335398 624806
rect 335454 624772 335488 624806
rect 335544 624772 335578 624806
rect 335004 624682 335038 624716
rect 335094 624682 335128 624716
rect 335184 624682 335218 624716
rect 335274 624682 335308 624716
rect 335364 624682 335398 624716
rect 335454 624682 335488 624716
rect 335544 624682 335578 624716
rect 335004 624592 335038 624626
rect 335094 624592 335128 624626
rect 335184 624592 335218 624626
rect 335274 624592 335308 624626
rect 335364 624592 335398 624626
rect 335454 624592 335488 624626
rect 335544 624592 335578 624626
rect 335004 624502 335038 624536
rect 335094 624502 335128 624536
rect 335184 624502 335218 624536
rect 335274 624502 335308 624536
rect 335364 624502 335398 624536
rect 335454 624502 335488 624536
rect 335544 624502 335578 624536
rect 335004 624412 335038 624446
rect 335094 624412 335128 624446
rect 335184 624412 335218 624446
rect 335274 624412 335308 624446
rect 335364 624412 335398 624446
rect 335454 624412 335488 624446
rect 335544 624412 335578 624446
rect 335004 624322 335038 624356
rect 335094 624322 335128 624356
rect 335184 624322 335218 624356
rect 335274 624322 335308 624356
rect 335364 624322 335398 624356
rect 335454 624322 335488 624356
rect 335544 624322 335578 624356
rect 335004 624232 335038 624266
rect 335094 624232 335128 624266
rect 335184 624232 335218 624266
rect 335274 624232 335308 624266
rect 335364 624232 335398 624266
rect 335454 624232 335488 624266
rect 335544 624232 335578 624266
rect 336292 624772 336326 624806
rect 336382 624772 336416 624806
rect 336472 624772 336506 624806
rect 336562 624772 336596 624806
rect 336652 624772 336686 624806
rect 336742 624772 336776 624806
rect 336832 624772 336866 624806
rect 336292 624682 336326 624716
rect 336382 624682 336416 624716
rect 336472 624682 336506 624716
rect 336562 624682 336596 624716
rect 336652 624682 336686 624716
rect 336742 624682 336776 624716
rect 336832 624682 336866 624716
rect 336292 624592 336326 624626
rect 336382 624592 336416 624626
rect 336472 624592 336506 624626
rect 336562 624592 336596 624626
rect 336652 624592 336686 624626
rect 336742 624592 336776 624626
rect 336832 624592 336866 624626
rect 336292 624502 336326 624536
rect 336382 624502 336416 624536
rect 336472 624502 336506 624536
rect 336562 624502 336596 624536
rect 336652 624502 336686 624536
rect 336742 624502 336776 624536
rect 336832 624502 336866 624536
rect 336292 624412 336326 624446
rect 336382 624412 336416 624446
rect 336472 624412 336506 624446
rect 336562 624412 336596 624446
rect 336652 624412 336686 624446
rect 336742 624412 336776 624446
rect 336832 624412 336866 624446
rect 336292 624322 336326 624356
rect 336382 624322 336416 624356
rect 336472 624322 336506 624356
rect 336562 624322 336596 624356
rect 336652 624322 336686 624356
rect 336742 624322 336776 624356
rect 336832 624322 336866 624356
rect 336292 624232 336326 624266
rect 336382 624232 336416 624266
rect 336472 624232 336506 624266
rect 336562 624232 336596 624266
rect 336652 624232 336686 624266
rect 336742 624232 336776 624266
rect 336832 624232 336866 624266
rect 337580 624772 337614 624806
rect 337670 624772 337704 624806
rect 337760 624772 337794 624806
rect 337850 624772 337884 624806
rect 337940 624772 337974 624806
rect 338030 624772 338064 624806
rect 338120 624772 338154 624806
rect 337580 624682 337614 624716
rect 337670 624682 337704 624716
rect 337760 624682 337794 624716
rect 337850 624682 337884 624716
rect 337940 624682 337974 624716
rect 338030 624682 338064 624716
rect 338120 624682 338154 624716
rect 337580 624592 337614 624626
rect 337670 624592 337704 624626
rect 337760 624592 337794 624626
rect 337850 624592 337884 624626
rect 337940 624592 337974 624626
rect 338030 624592 338064 624626
rect 338120 624592 338154 624626
rect 337580 624502 337614 624536
rect 337670 624502 337704 624536
rect 337760 624502 337794 624536
rect 337850 624502 337884 624536
rect 337940 624502 337974 624536
rect 338030 624502 338064 624536
rect 338120 624502 338154 624536
rect 337580 624412 337614 624446
rect 337670 624412 337704 624446
rect 337760 624412 337794 624446
rect 337850 624412 337884 624446
rect 337940 624412 337974 624446
rect 338030 624412 338064 624446
rect 338120 624412 338154 624446
rect 337580 624322 337614 624356
rect 337670 624322 337704 624356
rect 337760 624322 337794 624356
rect 337850 624322 337884 624356
rect 337940 624322 337974 624356
rect 338030 624322 338064 624356
rect 338120 624322 338154 624356
rect 337580 624232 337614 624266
rect 337670 624232 337704 624266
rect 337760 624232 337794 624266
rect 337850 624232 337884 624266
rect 337940 624232 337974 624266
rect 338030 624232 338064 624266
rect 338120 624232 338154 624266
rect 338868 624772 338902 624806
rect 338958 624772 338992 624806
rect 339048 624772 339082 624806
rect 339138 624772 339172 624806
rect 339228 624772 339262 624806
rect 339318 624772 339352 624806
rect 339408 624772 339442 624806
rect 338868 624682 338902 624716
rect 338958 624682 338992 624716
rect 339048 624682 339082 624716
rect 339138 624682 339172 624716
rect 339228 624682 339262 624716
rect 339318 624682 339352 624716
rect 339408 624682 339442 624716
rect 338868 624592 338902 624626
rect 338958 624592 338992 624626
rect 339048 624592 339082 624626
rect 339138 624592 339172 624626
rect 339228 624592 339262 624626
rect 339318 624592 339352 624626
rect 339408 624592 339442 624626
rect 338868 624502 338902 624536
rect 338958 624502 338992 624536
rect 339048 624502 339082 624536
rect 339138 624502 339172 624536
rect 339228 624502 339262 624536
rect 339318 624502 339352 624536
rect 339408 624502 339442 624536
rect 338868 624412 338902 624446
rect 338958 624412 338992 624446
rect 339048 624412 339082 624446
rect 339138 624412 339172 624446
rect 339228 624412 339262 624446
rect 339318 624412 339352 624446
rect 339408 624412 339442 624446
rect 338868 624322 338902 624356
rect 338958 624322 338992 624356
rect 339048 624322 339082 624356
rect 339138 624322 339172 624356
rect 339228 624322 339262 624356
rect 339318 624322 339352 624356
rect 339408 624322 339442 624356
rect 338868 624232 338902 624266
rect 338958 624232 338992 624266
rect 339048 624232 339082 624266
rect 339138 624232 339172 624266
rect 339228 624232 339262 624266
rect 339318 624232 339352 624266
rect 339408 624232 339442 624266
rect 340156 624772 340190 624806
rect 340246 624772 340280 624806
rect 340336 624772 340370 624806
rect 340426 624772 340460 624806
rect 340516 624772 340550 624806
rect 340606 624772 340640 624806
rect 340696 624772 340730 624806
rect 340156 624682 340190 624716
rect 340246 624682 340280 624716
rect 340336 624682 340370 624716
rect 340426 624682 340460 624716
rect 340516 624682 340550 624716
rect 340606 624682 340640 624716
rect 340696 624682 340730 624716
rect 340156 624592 340190 624626
rect 340246 624592 340280 624626
rect 340336 624592 340370 624626
rect 340426 624592 340460 624626
rect 340516 624592 340550 624626
rect 340606 624592 340640 624626
rect 340696 624592 340730 624626
rect 340156 624502 340190 624536
rect 340246 624502 340280 624536
rect 340336 624502 340370 624536
rect 340426 624502 340460 624536
rect 340516 624502 340550 624536
rect 340606 624502 340640 624536
rect 340696 624502 340730 624536
rect 340156 624412 340190 624446
rect 340246 624412 340280 624446
rect 340336 624412 340370 624446
rect 340426 624412 340460 624446
rect 340516 624412 340550 624446
rect 340606 624412 340640 624446
rect 340696 624412 340730 624446
rect 340156 624322 340190 624356
rect 340246 624322 340280 624356
rect 340336 624322 340370 624356
rect 340426 624322 340460 624356
rect 340516 624322 340550 624356
rect 340606 624322 340640 624356
rect 340696 624322 340730 624356
rect 340156 624232 340190 624266
rect 340246 624232 340280 624266
rect 340336 624232 340370 624266
rect 340426 624232 340460 624266
rect 340516 624232 340550 624266
rect 340606 624232 340640 624266
rect 340696 624232 340730 624266
rect 335004 623484 335038 623518
rect 335094 623484 335128 623518
rect 335184 623484 335218 623518
rect 335274 623484 335308 623518
rect 335364 623484 335398 623518
rect 335454 623484 335488 623518
rect 335544 623484 335578 623518
rect 335004 623394 335038 623428
rect 335094 623394 335128 623428
rect 335184 623394 335218 623428
rect 335274 623394 335308 623428
rect 335364 623394 335398 623428
rect 335454 623394 335488 623428
rect 335544 623394 335578 623428
rect 335004 623304 335038 623338
rect 335094 623304 335128 623338
rect 335184 623304 335218 623338
rect 335274 623304 335308 623338
rect 335364 623304 335398 623338
rect 335454 623304 335488 623338
rect 335544 623304 335578 623338
rect 335004 623214 335038 623248
rect 335094 623214 335128 623248
rect 335184 623214 335218 623248
rect 335274 623214 335308 623248
rect 335364 623214 335398 623248
rect 335454 623214 335488 623248
rect 335544 623214 335578 623248
rect 335004 623124 335038 623158
rect 335094 623124 335128 623158
rect 335184 623124 335218 623158
rect 335274 623124 335308 623158
rect 335364 623124 335398 623158
rect 335454 623124 335488 623158
rect 335544 623124 335578 623158
rect 335004 623034 335038 623068
rect 335094 623034 335128 623068
rect 335184 623034 335218 623068
rect 335274 623034 335308 623068
rect 335364 623034 335398 623068
rect 335454 623034 335488 623068
rect 335544 623034 335578 623068
rect 335004 622944 335038 622978
rect 335094 622944 335128 622978
rect 335184 622944 335218 622978
rect 335274 622944 335308 622978
rect 335364 622944 335398 622978
rect 335454 622944 335488 622978
rect 335544 622944 335578 622978
rect 336292 623484 336326 623518
rect 336382 623484 336416 623518
rect 336472 623484 336506 623518
rect 336562 623484 336596 623518
rect 336652 623484 336686 623518
rect 336742 623484 336776 623518
rect 336832 623484 336866 623518
rect 336292 623394 336326 623428
rect 336382 623394 336416 623428
rect 336472 623394 336506 623428
rect 336562 623394 336596 623428
rect 336652 623394 336686 623428
rect 336742 623394 336776 623428
rect 336832 623394 336866 623428
rect 336292 623304 336326 623338
rect 336382 623304 336416 623338
rect 336472 623304 336506 623338
rect 336562 623304 336596 623338
rect 336652 623304 336686 623338
rect 336742 623304 336776 623338
rect 336832 623304 336866 623338
rect 336292 623214 336326 623248
rect 336382 623214 336416 623248
rect 336472 623214 336506 623248
rect 336562 623214 336596 623248
rect 336652 623214 336686 623248
rect 336742 623214 336776 623248
rect 336832 623214 336866 623248
rect 336292 623124 336326 623158
rect 336382 623124 336416 623158
rect 336472 623124 336506 623158
rect 336562 623124 336596 623158
rect 336652 623124 336686 623158
rect 336742 623124 336776 623158
rect 336832 623124 336866 623158
rect 336292 623034 336326 623068
rect 336382 623034 336416 623068
rect 336472 623034 336506 623068
rect 336562 623034 336596 623068
rect 336652 623034 336686 623068
rect 336742 623034 336776 623068
rect 336832 623034 336866 623068
rect 336292 622944 336326 622978
rect 336382 622944 336416 622978
rect 336472 622944 336506 622978
rect 336562 622944 336596 622978
rect 336652 622944 336686 622978
rect 336742 622944 336776 622978
rect 336832 622944 336866 622978
rect 337580 623484 337614 623518
rect 337670 623484 337704 623518
rect 337760 623484 337794 623518
rect 337850 623484 337884 623518
rect 337940 623484 337974 623518
rect 338030 623484 338064 623518
rect 338120 623484 338154 623518
rect 337580 623394 337614 623428
rect 337670 623394 337704 623428
rect 337760 623394 337794 623428
rect 337850 623394 337884 623428
rect 337940 623394 337974 623428
rect 338030 623394 338064 623428
rect 338120 623394 338154 623428
rect 337580 623304 337614 623338
rect 337670 623304 337704 623338
rect 337760 623304 337794 623338
rect 337850 623304 337884 623338
rect 337940 623304 337974 623338
rect 338030 623304 338064 623338
rect 338120 623304 338154 623338
rect 337580 623214 337614 623248
rect 337670 623214 337704 623248
rect 337760 623214 337794 623248
rect 337850 623214 337884 623248
rect 337940 623214 337974 623248
rect 338030 623214 338064 623248
rect 338120 623214 338154 623248
rect 337580 623124 337614 623158
rect 337670 623124 337704 623158
rect 337760 623124 337794 623158
rect 337850 623124 337884 623158
rect 337940 623124 337974 623158
rect 338030 623124 338064 623158
rect 338120 623124 338154 623158
rect 337580 623034 337614 623068
rect 337670 623034 337704 623068
rect 337760 623034 337794 623068
rect 337850 623034 337884 623068
rect 337940 623034 337974 623068
rect 338030 623034 338064 623068
rect 338120 623034 338154 623068
rect 337580 622944 337614 622978
rect 337670 622944 337704 622978
rect 337760 622944 337794 622978
rect 337850 622944 337884 622978
rect 337940 622944 337974 622978
rect 338030 622944 338064 622978
rect 338120 622944 338154 622978
rect 338868 623484 338902 623518
rect 338958 623484 338992 623518
rect 339048 623484 339082 623518
rect 339138 623484 339172 623518
rect 339228 623484 339262 623518
rect 339318 623484 339352 623518
rect 339408 623484 339442 623518
rect 338868 623394 338902 623428
rect 338958 623394 338992 623428
rect 339048 623394 339082 623428
rect 339138 623394 339172 623428
rect 339228 623394 339262 623428
rect 339318 623394 339352 623428
rect 339408 623394 339442 623428
rect 338868 623304 338902 623338
rect 338958 623304 338992 623338
rect 339048 623304 339082 623338
rect 339138 623304 339172 623338
rect 339228 623304 339262 623338
rect 339318 623304 339352 623338
rect 339408 623304 339442 623338
rect 338868 623214 338902 623248
rect 338958 623214 338992 623248
rect 339048 623214 339082 623248
rect 339138 623214 339172 623248
rect 339228 623214 339262 623248
rect 339318 623214 339352 623248
rect 339408 623214 339442 623248
rect 338868 623124 338902 623158
rect 338958 623124 338992 623158
rect 339048 623124 339082 623158
rect 339138 623124 339172 623158
rect 339228 623124 339262 623158
rect 339318 623124 339352 623158
rect 339408 623124 339442 623158
rect 338868 623034 338902 623068
rect 338958 623034 338992 623068
rect 339048 623034 339082 623068
rect 339138 623034 339172 623068
rect 339228 623034 339262 623068
rect 339318 623034 339352 623068
rect 339408 623034 339442 623068
rect 338868 622944 338902 622978
rect 338958 622944 338992 622978
rect 339048 622944 339082 622978
rect 339138 622944 339172 622978
rect 339228 622944 339262 622978
rect 339318 622944 339352 622978
rect 339408 622944 339442 622978
rect 340156 623484 340190 623518
rect 340246 623484 340280 623518
rect 340336 623484 340370 623518
rect 340426 623484 340460 623518
rect 340516 623484 340550 623518
rect 340606 623484 340640 623518
rect 340696 623484 340730 623518
rect 340156 623394 340190 623428
rect 340246 623394 340280 623428
rect 340336 623394 340370 623428
rect 340426 623394 340460 623428
rect 340516 623394 340550 623428
rect 340606 623394 340640 623428
rect 340696 623394 340730 623428
rect 340156 623304 340190 623338
rect 340246 623304 340280 623338
rect 340336 623304 340370 623338
rect 340426 623304 340460 623338
rect 340516 623304 340550 623338
rect 340606 623304 340640 623338
rect 340696 623304 340730 623338
rect 340156 623214 340190 623248
rect 340246 623214 340280 623248
rect 340336 623214 340370 623248
rect 340426 623214 340460 623248
rect 340516 623214 340550 623248
rect 340606 623214 340640 623248
rect 340696 623214 340730 623248
rect 340156 623124 340190 623158
rect 340246 623124 340280 623158
rect 340336 623124 340370 623158
rect 340426 623124 340460 623158
rect 340516 623124 340550 623158
rect 340606 623124 340640 623158
rect 340696 623124 340730 623158
rect 340156 623034 340190 623068
rect 340246 623034 340280 623068
rect 340336 623034 340370 623068
rect 340426 623034 340460 623068
rect 340516 623034 340550 623068
rect 340606 623034 340640 623068
rect 340696 623034 340730 623068
rect 340156 622944 340190 622978
rect 340246 622944 340280 622978
rect 340336 622944 340370 622978
rect 340426 622944 340460 622978
rect 340516 622944 340550 622978
rect 340606 622944 340640 622978
rect 340696 622944 340730 622978
rect 335004 622196 335038 622230
rect 335094 622196 335128 622230
rect 335184 622196 335218 622230
rect 335274 622196 335308 622230
rect 335364 622196 335398 622230
rect 335454 622196 335488 622230
rect 335544 622196 335578 622230
rect 335004 622106 335038 622140
rect 335094 622106 335128 622140
rect 335184 622106 335218 622140
rect 335274 622106 335308 622140
rect 335364 622106 335398 622140
rect 335454 622106 335488 622140
rect 335544 622106 335578 622140
rect 335004 622016 335038 622050
rect 335094 622016 335128 622050
rect 335184 622016 335218 622050
rect 335274 622016 335308 622050
rect 335364 622016 335398 622050
rect 335454 622016 335488 622050
rect 335544 622016 335578 622050
rect 335004 621926 335038 621960
rect 335094 621926 335128 621960
rect 335184 621926 335218 621960
rect 335274 621926 335308 621960
rect 335364 621926 335398 621960
rect 335454 621926 335488 621960
rect 335544 621926 335578 621960
rect 335004 621836 335038 621870
rect 335094 621836 335128 621870
rect 335184 621836 335218 621870
rect 335274 621836 335308 621870
rect 335364 621836 335398 621870
rect 335454 621836 335488 621870
rect 335544 621836 335578 621870
rect 335004 621746 335038 621780
rect 335094 621746 335128 621780
rect 335184 621746 335218 621780
rect 335274 621746 335308 621780
rect 335364 621746 335398 621780
rect 335454 621746 335488 621780
rect 335544 621746 335578 621780
rect 335004 621656 335038 621690
rect 335094 621656 335128 621690
rect 335184 621656 335218 621690
rect 335274 621656 335308 621690
rect 335364 621656 335398 621690
rect 335454 621656 335488 621690
rect 335544 621656 335578 621690
rect 336292 622196 336326 622230
rect 336382 622196 336416 622230
rect 336472 622196 336506 622230
rect 336562 622196 336596 622230
rect 336652 622196 336686 622230
rect 336742 622196 336776 622230
rect 336832 622196 336866 622230
rect 336292 622106 336326 622140
rect 336382 622106 336416 622140
rect 336472 622106 336506 622140
rect 336562 622106 336596 622140
rect 336652 622106 336686 622140
rect 336742 622106 336776 622140
rect 336832 622106 336866 622140
rect 336292 622016 336326 622050
rect 336382 622016 336416 622050
rect 336472 622016 336506 622050
rect 336562 622016 336596 622050
rect 336652 622016 336686 622050
rect 336742 622016 336776 622050
rect 336832 622016 336866 622050
rect 336292 621926 336326 621960
rect 336382 621926 336416 621960
rect 336472 621926 336506 621960
rect 336562 621926 336596 621960
rect 336652 621926 336686 621960
rect 336742 621926 336776 621960
rect 336832 621926 336866 621960
rect 336292 621836 336326 621870
rect 336382 621836 336416 621870
rect 336472 621836 336506 621870
rect 336562 621836 336596 621870
rect 336652 621836 336686 621870
rect 336742 621836 336776 621870
rect 336832 621836 336866 621870
rect 336292 621746 336326 621780
rect 336382 621746 336416 621780
rect 336472 621746 336506 621780
rect 336562 621746 336596 621780
rect 336652 621746 336686 621780
rect 336742 621746 336776 621780
rect 336832 621746 336866 621780
rect 336292 621656 336326 621690
rect 336382 621656 336416 621690
rect 336472 621656 336506 621690
rect 336562 621656 336596 621690
rect 336652 621656 336686 621690
rect 336742 621656 336776 621690
rect 336832 621656 336866 621690
rect 337580 622196 337614 622230
rect 337670 622196 337704 622230
rect 337760 622196 337794 622230
rect 337850 622196 337884 622230
rect 337940 622196 337974 622230
rect 338030 622196 338064 622230
rect 338120 622196 338154 622230
rect 337580 622106 337614 622140
rect 337670 622106 337704 622140
rect 337760 622106 337794 622140
rect 337850 622106 337884 622140
rect 337940 622106 337974 622140
rect 338030 622106 338064 622140
rect 338120 622106 338154 622140
rect 337580 622016 337614 622050
rect 337670 622016 337704 622050
rect 337760 622016 337794 622050
rect 337850 622016 337884 622050
rect 337940 622016 337974 622050
rect 338030 622016 338064 622050
rect 338120 622016 338154 622050
rect 337580 621926 337614 621960
rect 337670 621926 337704 621960
rect 337760 621926 337794 621960
rect 337850 621926 337884 621960
rect 337940 621926 337974 621960
rect 338030 621926 338064 621960
rect 338120 621926 338154 621960
rect 337580 621836 337614 621870
rect 337670 621836 337704 621870
rect 337760 621836 337794 621870
rect 337850 621836 337884 621870
rect 337940 621836 337974 621870
rect 338030 621836 338064 621870
rect 338120 621836 338154 621870
rect 337580 621746 337614 621780
rect 337670 621746 337704 621780
rect 337760 621746 337794 621780
rect 337850 621746 337884 621780
rect 337940 621746 337974 621780
rect 338030 621746 338064 621780
rect 338120 621746 338154 621780
rect 337580 621656 337614 621690
rect 337670 621656 337704 621690
rect 337760 621656 337794 621690
rect 337850 621656 337884 621690
rect 337940 621656 337974 621690
rect 338030 621656 338064 621690
rect 338120 621656 338154 621690
rect 338868 622196 338902 622230
rect 338958 622196 338992 622230
rect 339048 622196 339082 622230
rect 339138 622196 339172 622230
rect 339228 622196 339262 622230
rect 339318 622196 339352 622230
rect 339408 622196 339442 622230
rect 338868 622106 338902 622140
rect 338958 622106 338992 622140
rect 339048 622106 339082 622140
rect 339138 622106 339172 622140
rect 339228 622106 339262 622140
rect 339318 622106 339352 622140
rect 339408 622106 339442 622140
rect 338868 622016 338902 622050
rect 338958 622016 338992 622050
rect 339048 622016 339082 622050
rect 339138 622016 339172 622050
rect 339228 622016 339262 622050
rect 339318 622016 339352 622050
rect 339408 622016 339442 622050
rect 338868 621926 338902 621960
rect 338958 621926 338992 621960
rect 339048 621926 339082 621960
rect 339138 621926 339172 621960
rect 339228 621926 339262 621960
rect 339318 621926 339352 621960
rect 339408 621926 339442 621960
rect 338868 621836 338902 621870
rect 338958 621836 338992 621870
rect 339048 621836 339082 621870
rect 339138 621836 339172 621870
rect 339228 621836 339262 621870
rect 339318 621836 339352 621870
rect 339408 621836 339442 621870
rect 338868 621746 338902 621780
rect 338958 621746 338992 621780
rect 339048 621746 339082 621780
rect 339138 621746 339172 621780
rect 339228 621746 339262 621780
rect 339318 621746 339352 621780
rect 339408 621746 339442 621780
rect 338868 621656 338902 621690
rect 338958 621656 338992 621690
rect 339048 621656 339082 621690
rect 339138 621656 339172 621690
rect 339228 621656 339262 621690
rect 339318 621656 339352 621690
rect 339408 621656 339442 621690
rect 340156 622196 340190 622230
rect 340246 622196 340280 622230
rect 340336 622196 340370 622230
rect 340426 622196 340460 622230
rect 340516 622196 340550 622230
rect 340606 622196 340640 622230
rect 340696 622196 340730 622230
rect 340156 622106 340190 622140
rect 340246 622106 340280 622140
rect 340336 622106 340370 622140
rect 340426 622106 340460 622140
rect 340516 622106 340550 622140
rect 340606 622106 340640 622140
rect 340696 622106 340730 622140
rect 340156 622016 340190 622050
rect 340246 622016 340280 622050
rect 340336 622016 340370 622050
rect 340426 622016 340460 622050
rect 340516 622016 340550 622050
rect 340606 622016 340640 622050
rect 340696 622016 340730 622050
rect 340156 621926 340190 621960
rect 340246 621926 340280 621960
rect 340336 621926 340370 621960
rect 340426 621926 340460 621960
rect 340516 621926 340550 621960
rect 340606 621926 340640 621960
rect 340696 621926 340730 621960
rect 340156 621836 340190 621870
rect 340246 621836 340280 621870
rect 340336 621836 340370 621870
rect 340426 621836 340460 621870
rect 340516 621836 340550 621870
rect 340606 621836 340640 621870
rect 340696 621836 340730 621870
rect 340156 621746 340190 621780
rect 340246 621746 340280 621780
rect 340336 621746 340370 621780
rect 340426 621746 340460 621780
rect 340516 621746 340550 621780
rect 340606 621746 340640 621780
rect 340696 621746 340730 621780
rect 340156 621656 340190 621690
rect 340246 621656 340280 621690
rect 340336 621656 340370 621690
rect 340426 621656 340460 621690
rect 340516 621656 340550 621690
rect 340606 621656 340640 621690
rect 340696 621656 340730 621690
rect 335004 620908 335038 620942
rect 335094 620908 335128 620942
rect 335184 620908 335218 620942
rect 335274 620908 335308 620942
rect 335364 620908 335398 620942
rect 335454 620908 335488 620942
rect 335544 620908 335578 620942
rect 335004 620818 335038 620852
rect 335094 620818 335128 620852
rect 335184 620818 335218 620852
rect 335274 620818 335308 620852
rect 335364 620818 335398 620852
rect 335454 620818 335488 620852
rect 335544 620818 335578 620852
rect 335004 620728 335038 620762
rect 335094 620728 335128 620762
rect 335184 620728 335218 620762
rect 335274 620728 335308 620762
rect 335364 620728 335398 620762
rect 335454 620728 335488 620762
rect 335544 620728 335578 620762
rect 335004 620638 335038 620672
rect 335094 620638 335128 620672
rect 335184 620638 335218 620672
rect 335274 620638 335308 620672
rect 335364 620638 335398 620672
rect 335454 620638 335488 620672
rect 335544 620638 335578 620672
rect 335004 620548 335038 620582
rect 335094 620548 335128 620582
rect 335184 620548 335218 620582
rect 335274 620548 335308 620582
rect 335364 620548 335398 620582
rect 335454 620548 335488 620582
rect 335544 620548 335578 620582
rect 335004 620458 335038 620492
rect 335094 620458 335128 620492
rect 335184 620458 335218 620492
rect 335274 620458 335308 620492
rect 335364 620458 335398 620492
rect 335454 620458 335488 620492
rect 335544 620458 335578 620492
rect 335004 620368 335038 620402
rect 335094 620368 335128 620402
rect 335184 620368 335218 620402
rect 335274 620368 335308 620402
rect 335364 620368 335398 620402
rect 335454 620368 335488 620402
rect 335544 620368 335578 620402
rect 336292 620908 336326 620942
rect 336382 620908 336416 620942
rect 336472 620908 336506 620942
rect 336562 620908 336596 620942
rect 336652 620908 336686 620942
rect 336742 620908 336776 620942
rect 336832 620908 336866 620942
rect 336292 620818 336326 620852
rect 336382 620818 336416 620852
rect 336472 620818 336506 620852
rect 336562 620818 336596 620852
rect 336652 620818 336686 620852
rect 336742 620818 336776 620852
rect 336832 620818 336866 620852
rect 336292 620728 336326 620762
rect 336382 620728 336416 620762
rect 336472 620728 336506 620762
rect 336562 620728 336596 620762
rect 336652 620728 336686 620762
rect 336742 620728 336776 620762
rect 336832 620728 336866 620762
rect 336292 620638 336326 620672
rect 336382 620638 336416 620672
rect 336472 620638 336506 620672
rect 336562 620638 336596 620672
rect 336652 620638 336686 620672
rect 336742 620638 336776 620672
rect 336832 620638 336866 620672
rect 336292 620548 336326 620582
rect 336382 620548 336416 620582
rect 336472 620548 336506 620582
rect 336562 620548 336596 620582
rect 336652 620548 336686 620582
rect 336742 620548 336776 620582
rect 336832 620548 336866 620582
rect 336292 620458 336326 620492
rect 336382 620458 336416 620492
rect 336472 620458 336506 620492
rect 336562 620458 336596 620492
rect 336652 620458 336686 620492
rect 336742 620458 336776 620492
rect 336832 620458 336866 620492
rect 336292 620368 336326 620402
rect 336382 620368 336416 620402
rect 336472 620368 336506 620402
rect 336562 620368 336596 620402
rect 336652 620368 336686 620402
rect 336742 620368 336776 620402
rect 336832 620368 336866 620402
rect 337580 620908 337614 620942
rect 337670 620908 337704 620942
rect 337760 620908 337794 620942
rect 337850 620908 337884 620942
rect 337940 620908 337974 620942
rect 338030 620908 338064 620942
rect 338120 620908 338154 620942
rect 337580 620818 337614 620852
rect 337670 620818 337704 620852
rect 337760 620818 337794 620852
rect 337850 620818 337884 620852
rect 337940 620818 337974 620852
rect 338030 620818 338064 620852
rect 338120 620818 338154 620852
rect 337580 620728 337614 620762
rect 337670 620728 337704 620762
rect 337760 620728 337794 620762
rect 337850 620728 337884 620762
rect 337940 620728 337974 620762
rect 338030 620728 338064 620762
rect 338120 620728 338154 620762
rect 337580 620638 337614 620672
rect 337670 620638 337704 620672
rect 337760 620638 337794 620672
rect 337850 620638 337884 620672
rect 337940 620638 337974 620672
rect 338030 620638 338064 620672
rect 338120 620638 338154 620672
rect 337580 620548 337614 620582
rect 337670 620548 337704 620582
rect 337760 620548 337794 620582
rect 337850 620548 337884 620582
rect 337940 620548 337974 620582
rect 338030 620548 338064 620582
rect 338120 620548 338154 620582
rect 337580 620458 337614 620492
rect 337670 620458 337704 620492
rect 337760 620458 337794 620492
rect 337850 620458 337884 620492
rect 337940 620458 337974 620492
rect 338030 620458 338064 620492
rect 338120 620458 338154 620492
rect 337580 620368 337614 620402
rect 337670 620368 337704 620402
rect 337760 620368 337794 620402
rect 337850 620368 337884 620402
rect 337940 620368 337974 620402
rect 338030 620368 338064 620402
rect 338120 620368 338154 620402
rect 338868 620908 338902 620942
rect 338958 620908 338992 620942
rect 339048 620908 339082 620942
rect 339138 620908 339172 620942
rect 339228 620908 339262 620942
rect 339318 620908 339352 620942
rect 339408 620908 339442 620942
rect 338868 620818 338902 620852
rect 338958 620818 338992 620852
rect 339048 620818 339082 620852
rect 339138 620818 339172 620852
rect 339228 620818 339262 620852
rect 339318 620818 339352 620852
rect 339408 620818 339442 620852
rect 338868 620728 338902 620762
rect 338958 620728 338992 620762
rect 339048 620728 339082 620762
rect 339138 620728 339172 620762
rect 339228 620728 339262 620762
rect 339318 620728 339352 620762
rect 339408 620728 339442 620762
rect 338868 620638 338902 620672
rect 338958 620638 338992 620672
rect 339048 620638 339082 620672
rect 339138 620638 339172 620672
rect 339228 620638 339262 620672
rect 339318 620638 339352 620672
rect 339408 620638 339442 620672
rect 338868 620548 338902 620582
rect 338958 620548 338992 620582
rect 339048 620548 339082 620582
rect 339138 620548 339172 620582
rect 339228 620548 339262 620582
rect 339318 620548 339352 620582
rect 339408 620548 339442 620582
rect 338868 620458 338902 620492
rect 338958 620458 338992 620492
rect 339048 620458 339082 620492
rect 339138 620458 339172 620492
rect 339228 620458 339262 620492
rect 339318 620458 339352 620492
rect 339408 620458 339442 620492
rect 338868 620368 338902 620402
rect 338958 620368 338992 620402
rect 339048 620368 339082 620402
rect 339138 620368 339172 620402
rect 339228 620368 339262 620402
rect 339318 620368 339352 620402
rect 339408 620368 339442 620402
rect 340156 620908 340190 620942
rect 340246 620908 340280 620942
rect 340336 620908 340370 620942
rect 340426 620908 340460 620942
rect 340516 620908 340550 620942
rect 340606 620908 340640 620942
rect 340696 620908 340730 620942
rect 340156 620818 340190 620852
rect 340246 620818 340280 620852
rect 340336 620818 340370 620852
rect 340426 620818 340460 620852
rect 340516 620818 340550 620852
rect 340606 620818 340640 620852
rect 340696 620818 340730 620852
rect 340156 620728 340190 620762
rect 340246 620728 340280 620762
rect 340336 620728 340370 620762
rect 340426 620728 340460 620762
rect 340516 620728 340550 620762
rect 340606 620728 340640 620762
rect 340696 620728 340730 620762
rect 340156 620638 340190 620672
rect 340246 620638 340280 620672
rect 340336 620638 340370 620672
rect 340426 620638 340460 620672
rect 340516 620638 340550 620672
rect 340606 620638 340640 620672
rect 340696 620638 340730 620672
rect 340156 620548 340190 620582
rect 340246 620548 340280 620582
rect 340336 620548 340370 620582
rect 340426 620548 340460 620582
rect 340516 620548 340550 620582
rect 340606 620548 340640 620582
rect 340696 620548 340730 620582
rect 340156 620458 340190 620492
rect 340246 620458 340280 620492
rect 340336 620458 340370 620492
rect 340426 620458 340460 620492
rect 340516 620458 340550 620492
rect 340606 620458 340640 620492
rect 340696 620458 340730 620492
rect 340156 620368 340190 620402
rect 340246 620368 340280 620402
rect 340336 620368 340370 620402
rect 340426 620368 340460 620402
rect 340516 620368 340550 620402
rect 340606 620368 340640 620402
rect 340696 620368 340730 620402
rect 335004 619620 335038 619654
rect 335094 619620 335128 619654
rect 335184 619620 335218 619654
rect 335274 619620 335308 619654
rect 335364 619620 335398 619654
rect 335454 619620 335488 619654
rect 335544 619620 335578 619654
rect 335004 619530 335038 619564
rect 335094 619530 335128 619564
rect 335184 619530 335218 619564
rect 335274 619530 335308 619564
rect 335364 619530 335398 619564
rect 335454 619530 335488 619564
rect 335544 619530 335578 619564
rect 335004 619440 335038 619474
rect 335094 619440 335128 619474
rect 335184 619440 335218 619474
rect 335274 619440 335308 619474
rect 335364 619440 335398 619474
rect 335454 619440 335488 619474
rect 335544 619440 335578 619474
rect 335004 619350 335038 619384
rect 335094 619350 335128 619384
rect 335184 619350 335218 619384
rect 335274 619350 335308 619384
rect 335364 619350 335398 619384
rect 335454 619350 335488 619384
rect 335544 619350 335578 619384
rect 335004 619260 335038 619294
rect 335094 619260 335128 619294
rect 335184 619260 335218 619294
rect 335274 619260 335308 619294
rect 335364 619260 335398 619294
rect 335454 619260 335488 619294
rect 335544 619260 335578 619294
rect 335004 619170 335038 619204
rect 335094 619170 335128 619204
rect 335184 619170 335218 619204
rect 335274 619170 335308 619204
rect 335364 619170 335398 619204
rect 335454 619170 335488 619204
rect 335544 619170 335578 619204
rect 335004 619080 335038 619114
rect 335094 619080 335128 619114
rect 335184 619080 335218 619114
rect 335274 619080 335308 619114
rect 335364 619080 335398 619114
rect 335454 619080 335488 619114
rect 335544 619080 335578 619114
rect 336292 619620 336326 619654
rect 336382 619620 336416 619654
rect 336472 619620 336506 619654
rect 336562 619620 336596 619654
rect 336652 619620 336686 619654
rect 336742 619620 336776 619654
rect 336832 619620 336866 619654
rect 336292 619530 336326 619564
rect 336382 619530 336416 619564
rect 336472 619530 336506 619564
rect 336562 619530 336596 619564
rect 336652 619530 336686 619564
rect 336742 619530 336776 619564
rect 336832 619530 336866 619564
rect 336292 619440 336326 619474
rect 336382 619440 336416 619474
rect 336472 619440 336506 619474
rect 336562 619440 336596 619474
rect 336652 619440 336686 619474
rect 336742 619440 336776 619474
rect 336832 619440 336866 619474
rect 336292 619350 336326 619384
rect 336382 619350 336416 619384
rect 336472 619350 336506 619384
rect 336562 619350 336596 619384
rect 336652 619350 336686 619384
rect 336742 619350 336776 619384
rect 336832 619350 336866 619384
rect 336292 619260 336326 619294
rect 336382 619260 336416 619294
rect 336472 619260 336506 619294
rect 336562 619260 336596 619294
rect 336652 619260 336686 619294
rect 336742 619260 336776 619294
rect 336832 619260 336866 619294
rect 336292 619170 336326 619204
rect 336382 619170 336416 619204
rect 336472 619170 336506 619204
rect 336562 619170 336596 619204
rect 336652 619170 336686 619204
rect 336742 619170 336776 619204
rect 336832 619170 336866 619204
rect 336292 619080 336326 619114
rect 336382 619080 336416 619114
rect 336472 619080 336506 619114
rect 336562 619080 336596 619114
rect 336652 619080 336686 619114
rect 336742 619080 336776 619114
rect 336832 619080 336866 619114
rect 337580 619620 337614 619654
rect 337670 619620 337704 619654
rect 337760 619620 337794 619654
rect 337850 619620 337884 619654
rect 337940 619620 337974 619654
rect 338030 619620 338064 619654
rect 338120 619620 338154 619654
rect 337580 619530 337614 619564
rect 337670 619530 337704 619564
rect 337760 619530 337794 619564
rect 337850 619530 337884 619564
rect 337940 619530 337974 619564
rect 338030 619530 338064 619564
rect 338120 619530 338154 619564
rect 337580 619440 337614 619474
rect 337670 619440 337704 619474
rect 337760 619440 337794 619474
rect 337850 619440 337884 619474
rect 337940 619440 337974 619474
rect 338030 619440 338064 619474
rect 338120 619440 338154 619474
rect 337580 619350 337614 619384
rect 337670 619350 337704 619384
rect 337760 619350 337794 619384
rect 337850 619350 337884 619384
rect 337940 619350 337974 619384
rect 338030 619350 338064 619384
rect 338120 619350 338154 619384
rect 337580 619260 337614 619294
rect 337670 619260 337704 619294
rect 337760 619260 337794 619294
rect 337850 619260 337884 619294
rect 337940 619260 337974 619294
rect 338030 619260 338064 619294
rect 338120 619260 338154 619294
rect 337580 619170 337614 619204
rect 337670 619170 337704 619204
rect 337760 619170 337794 619204
rect 337850 619170 337884 619204
rect 337940 619170 337974 619204
rect 338030 619170 338064 619204
rect 338120 619170 338154 619204
rect 337580 619080 337614 619114
rect 337670 619080 337704 619114
rect 337760 619080 337794 619114
rect 337850 619080 337884 619114
rect 337940 619080 337974 619114
rect 338030 619080 338064 619114
rect 338120 619080 338154 619114
rect 338868 619620 338902 619654
rect 338958 619620 338992 619654
rect 339048 619620 339082 619654
rect 339138 619620 339172 619654
rect 339228 619620 339262 619654
rect 339318 619620 339352 619654
rect 339408 619620 339442 619654
rect 338868 619530 338902 619564
rect 338958 619530 338992 619564
rect 339048 619530 339082 619564
rect 339138 619530 339172 619564
rect 339228 619530 339262 619564
rect 339318 619530 339352 619564
rect 339408 619530 339442 619564
rect 338868 619440 338902 619474
rect 338958 619440 338992 619474
rect 339048 619440 339082 619474
rect 339138 619440 339172 619474
rect 339228 619440 339262 619474
rect 339318 619440 339352 619474
rect 339408 619440 339442 619474
rect 338868 619350 338902 619384
rect 338958 619350 338992 619384
rect 339048 619350 339082 619384
rect 339138 619350 339172 619384
rect 339228 619350 339262 619384
rect 339318 619350 339352 619384
rect 339408 619350 339442 619384
rect 338868 619260 338902 619294
rect 338958 619260 338992 619294
rect 339048 619260 339082 619294
rect 339138 619260 339172 619294
rect 339228 619260 339262 619294
rect 339318 619260 339352 619294
rect 339408 619260 339442 619294
rect 338868 619170 338902 619204
rect 338958 619170 338992 619204
rect 339048 619170 339082 619204
rect 339138 619170 339172 619204
rect 339228 619170 339262 619204
rect 339318 619170 339352 619204
rect 339408 619170 339442 619204
rect 338868 619080 338902 619114
rect 338958 619080 338992 619114
rect 339048 619080 339082 619114
rect 339138 619080 339172 619114
rect 339228 619080 339262 619114
rect 339318 619080 339352 619114
rect 339408 619080 339442 619114
rect 340156 619620 340190 619654
rect 340246 619620 340280 619654
rect 340336 619620 340370 619654
rect 340426 619620 340460 619654
rect 340516 619620 340550 619654
rect 340606 619620 340640 619654
rect 340696 619620 340730 619654
rect 340156 619530 340190 619564
rect 340246 619530 340280 619564
rect 340336 619530 340370 619564
rect 340426 619530 340460 619564
rect 340516 619530 340550 619564
rect 340606 619530 340640 619564
rect 340696 619530 340730 619564
rect 340156 619440 340190 619474
rect 340246 619440 340280 619474
rect 340336 619440 340370 619474
rect 340426 619440 340460 619474
rect 340516 619440 340550 619474
rect 340606 619440 340640 619474
rect 340696 619440 340730 619474
rect 340156 619350 340190 619384
rect 340246 619350 340280 619384
rect 340336 619350 340370 619384
rect 340426 619350 340460 619384
rect 340516 619350 340550 619384
rect 340606 619350 340640 619384
rect 340696 619350 340730 619384
rect 340156 619260 340190 619294
rect 340246 619260 340280 619294
rect 340336 619260 340370 619294
rect 340426 619260 340460 619294
rect 340516 619260 340550 619294
rect 340606 619260 340640 619294
rect 340696 619260 340730 619294
rect 340156 619170 340190 619204
rect 340246 619170 340280 619204
rect 340336 619170 340370 619204
rect 340426 619170 340460 619204
rect 340516 619170 340550 619204
rect 340606 619170 340640 619204
rect 340696 619170 340730 619204
rect 340156 619080 340190 619114
rect 340246 619080 340280 619114
rect 340336 619080 340370 619114
rect 340426 619080 340460 619114
rect 340516 619080 340550 619114
rect 340606 619080 340640 619114
rect 340696 619080 340730 619114
rect 335004 618332 335038 618366
rect 335094 618332 335128 618366
rect 335184 618332 335218 618366
rect 335274 618332 335308 618366
rect 335364 618332 335398 618366
rect 335454 618332 335488 618366
rect 335544 618332 335578 618366
rect 335004 618242 335038 618276
rect 335094 618242 335128 618276
rect 335184 618242 335218 618276
rect 335274 618242 335308 618276
rect 335364 618242 335398 618276
rect 335454 618242 335488 618276
rect 335544 618242 335578 618276
rect 335004 618152 335038 618186
rect 335094 618152 335128 618186
rect 335184 618152 335218 618186
rect 335274 618152 335308 618186
rect 335364 618152 335398 618186
rect 335454 618152 335488 618186
rect 335544 618152 335578 618186
rect 335004 618062 335038 618096
rect 335094 618062 335128 618096
rect 335184 618062 335218 618096
rect 335274 618062 335308 618096
rect 335364 618062 335398 618096
rect 335454 618062 335488 618096
rect 335544 618062 335578 618096
rect 335004 617972 335038 618006
rect 335094 617972 335128 618006
rect 335184 617972 335218 618006
rect 335274 617972 335308 618006
rect 335364 617972 335398 618006
rect 335454 617972 335488 618006
rect 335544 617972 335578 618006
rect 335004 617882 335038 617916
rect 335094 617882 335128 617916
rect 335184 617882 335218 617916
rect 335274 617882 335308 617916
rect 335364 617882 335398 617916
rect 335454 617882 335488 617916
rect 335544 617882 335578 617916
rect 335004 617792 335038 617826
rect 335094 617792 335128 617826
rect 335184 617792 335218 617826
rect 335274 617792 335308 617826
rect 335364 617792 335398 617826
rect 335454 617792 335488 617826
rect 335544 617792 335578 617826
rect 336292 618332 336326 618366
rect 336382 618332 336416 618366
rect 336472 618332 336506 618366
rect 336562 618332 336596 618366
rect 336652 618332 336686 618366
rect 336742 618332 336776 618366
rect 336832 618332 336866 618366
rect 336292 618242 336326 618276
rect 336382 618242 336416 618276
rect 336472 618242 336506 618276
rect 336562 618242 336596 618276
rect 336652 618242 336686 618276
rect 336742 618242 336776 618276
rect 336832 618242 336866 618276
rect 336292 618152 336326 618186
rect 336382 618152 336416 618186
rect 336472 618152 336506 618186
rect 336562 618152 336596 618186
rect 336652 618152 336686 618186
rect 336742 618152 336776 618186
rect 336832 618152 336866 618186
rect 336292 618062 336326 618096
rect 336382 618062 336416 618096
rect 336472 618062 336506 618096
rect 336562 618062 336596 618096
rect 336652 618062 336686 618096
rect 336742 618062 336776 618096
rect 336832 618062 336866 618096
rect 336292 617972 336326 618006
rect 336382 617972 336416 618006
rect 336472 617972 336506 618006
rect 336562 617972 336596 618006
rect 336652 617972 336686 618006
rect 336742 617972 336776 618006
rect 336832 617972 336866 618006
rect 336292 617882 336326 617916
rect 336382 617882 336416 617916
rect 336472 617882 336506 617916
rect 336562 617882 336596 617916
rect 336652 617882 336686 617916
rect 336742 617882 336776 617916
rect 336832 617882 336866 617916
rect 336292 617792 336326 617826
rect 336382 617792 336416 617826
rect 336472 617792 336506 617826
rect 336562 617792 336596 617826
rect 336652 617792 336686 617826
rect 336742 617792 336776 617826
rect 336832 617792 336866 617826
rect 337580 618332 337614 618366
rect 337670 618332 337704 618366
rect 337760 618332 337794 618366
rect 337850 618332 337884 618366
rect 337940 618332 337974 618366
rect 338030 618332 338064 618366
rect 338120 618332 338154 618366
rect 337580 618242 337614 618276
rect 337670 618242 337704 618276
rect 337760 618242 337794 618276
rect 337850 618242 337884 618276
rect 337940 618242 337974 618276
rect 338030 618242 338064 618276
rect 338120 618242 338154 618276
rect 337580 618152 337614 618186
rect 337670 618152 337704 618186
rect 337760 618152 337794 618186
rect 337850 618152 337884 618186
rect 337940 618152 337974 618186
rect 338030 618152 338064 618186
rect 338120 618152 338154 618186
rect 337580 618062 337614 618096
rect 337670 618062 337704 618096
rect 337760 618062 337794 618096
rect 337850 618062 337884 618096
rect 337940 618062 337974 618096
rect 338030 618062 338064 618096
rect 338120 618062 338154 618096
rect 337580 617972 337614 618006
rect 337670 617972 337704 618006
rect 337760 617972 337794 618006
rect 337850 617972 337884 618006
rect 337940 617972 337974 618006
rect 338030 617972 338064 618006
rect 338120 617972 338154 618006
rect 337580 617882 337614 617916
rect 337670 617882 337704 617916
rect 337760 617882 337794 617916
rect 337850 617882 337884 617916
rect 337940 617882 337974 617916
rect 338030 617882 338064 617916
rect 338120 617882 338154 617916
rect 337580 617792 337614 617826
rect 337670 617792 337704 617826
rect 337760 617792 337794 617826
rect 337850 617792 337884 617826
rect 337940 617792 337974 617826
rect 338030 617792 338064 617826
rect 338120 617792 338154 617826
rect 338868 618332 338902 618366
rect 338958 618332 338992 618366
rect 339048 618332 339082 618366
rect 339138 618332 339172 618366
rect 339228 618332 339262 618366
rect 339318 618332 339352 618366
rect 339408 618332 339442 618366
rect 338868 618242 338902 618276
rect 338958 618242 338992 618276
rect 339048 618242 339082 618276
rect 339138 618242 339172 618276
rect 339228 618242 339262 618276
rect 339318 618242 339352 618276
rect 339408 618242 339442 618276
rect 338868 618152 338902 618186
rect 338958 618152 338992 618186
rect 339048 618152 339082 618186
rect 339138 618152 339172 618186
rect 339228 618152 339262 618186
rect 339318 618152 339352 618186
rect 339408 618152 339442 618186
rect 338868 618062 338902 618096
rect 338958 618062 338992 618096
rect 339048 618062 339082 618096
rect 339138 618062 339172 618096
rect 339228 618062 339262 618096
rect 339318 618062 339352 618096
rect 339408 618062 339442 618096
rect 338868 617972 338902 618006
rect 338958 617972 338992 618006
rect 339048 617972 339082 618006
rect 339138 617972 339172 618006
rect 339228 617972 339262 618006
rect 339318 617972 339352 618006
rect 339408 617972 339442 618006
rect 338868 617882 338902 617916
rect 338958 617882 338992 617916
rect 339048 617882 339082 617916
rect 339138 617882 339172 617916
rect 339228 617882 339262 617916
rect 339318 617882 339352 617916
rect 339408 617882 339442 617916
rect 338868 617792 338902 617826
rect 338958 617792 338992 617826
rect 339048 617792 339082 617826
rect 339138 617792 339172 617826
rect 339228 617792 339262 617826
rect 339318 617792 339352 617826
rect 339408 617792 339442 617826
rect 340156 618332 340190 618366
rect 340246 618332 340280 618366
rect 340336 618332 340370 618366
rect 340426 618332 340460 618366
rect 340516 618332 340550 618366
rect 340606 618332 340640 618366
rect 340696 618332 340730 618366
rect 340156 618242 340190 618276
rect 340246 618242 340280 618276
rect 340336 618242 340370 618276
rect 340426 618242 340460 618276
rect 340516 618242 340550 618276
rect 340606 618242 340640 618276
rect 340696 618242 340730 618276
rect 340156 618152 340190 618186
rect 340246 618152 340280 618186
rect 340336 618152 340370 618186
rect 340426 618152 340460 618186
rect 340516 618152 340550 618186
rect 340606 618152 340640 618186
rect 340696 618152 340730 618186
rect 340156 618062 340190 618096
rect 340246 618062 340280 618096
rect 340336 618062 340370 618096
rect 340426 618062 340460 618096
rect 340516 618062 340550 618096
rect 340606 618062 340640 618096
rect 340696 618062 340730 618096
rect 340156 617972 340190 618006
rect 340246 617972 340280 618006
rect 340336 617972 340370 618006
rect 340426 617972 340460 618006
rect 340516 617972 340550 618006
rect 340606 617972 340640 618006
rect 340696 617972 340730 618006
rect 340156 617882 340190 617916
rect 340246 617882 340280 617916
rect 340336 617882 340370 617916
rect 340426 617882 340460 617916
rect 340516 617882 340550 617916
rect 340606 617882 340640 617916
rect 340696 617882 340730 617916
rect 340156 617792 340190 617826
rect 340246 617792 340280 617826
rect 340336 617792 340370 617826
rect 340426 617792 340460 617826
rect 340516 617792 340550 617826
rect 340606 617792 340640 617826
rect 340696 617792 340730 617826
<< psubdiff >>
rect 297800 642672 343160 642696
rect 297800 641672 297824 642672
rect 343136 641672 343160 642672
rect 297800 641648 343160 641672
rect 342088 640648 343136 640672
rect 297848 640624 298896 640648
rect 297848 616472 297872 640624
rect 298872 616472 298896 640624
rect 300664 640542 311896 640566
rect 300664 639776 300688 640542
rect 311872 639776 311896 640542
rect 300664 639752 311896 639776
rect 312424 637006 313042 637030
rect 312424 630702 312448 637006
rect 313018 630702 313042 637006
rect 315668 637006 316286 637030
rect 312424 630678 313042 630702
rect 315668 630702 315692 637006
rect 316262 630702 316286 637006
rect 320628 637006 321246 637030
rect 315668 630678 316286 630702
rect 320628 630702 320652 637006
rect 321222 630702 321246 637006
rect 320628 630678 321246 630702
rect 335316 637006 335934 637030
rect 335316 630702 335340 637006
rect 335910 630702 335934 637006
rect 335316 630678 335934 630702
rect 334648 627708 341088 627740
rect 334648 627674 334782 627708
rect 334816 627674 334872 627708
rect 334906 627674 334962 627708
rect 334996 627674 335052 627708
rect 335086 627674 335142 627708
rect 335176 627674 335232 627708
rect 335266 627674 335322 627708
rect 335356 627674 335412 627708
rect 335446 627674 335502 627708
rect 335536 627674 335592 627708
rect 335626 627674 335682 627708
rect 335716 627674 335772 627708
rect 335806 627674 336070 627708
rect 336104 627674 336160 627708
rect 336194 627674 336250 627708
rect 336284 627674 336340 627708
rect 336374 627674 336430 627708
rect 336464 627674 336520 627708
rect 336554 627674 336610 627708
rect 336644 627674 336700 627708
rect 336734 627674 336790 627708
rect 336824 627674 336880 627708
rect 336914 627674 336970 627708
rect 337004 627674 337060 627708
rect 337094 627674 337358 627708
rect 337392 627674 337448 627708
rect 337482 627674 337538 627708
rect 337572 627674 337628 627708
rect 337662 627674 337718 627708
rect 337752 627674 337808 627708
rect 337842 627674 337898 627708
rect 337932 627674 337988 627708
rect 338022 627674 338078 627708
rect 338112 627674 338168 627708
rect 338202 627674 338258 627708
rect 338292 627674 338348 627708
rect 338382 627674 338646 627708
rect 338680 627674 338736 627708
rect 338770 627674 338826 627708
rect 338860 627674 338916 627708
rect 338950 627674 339006 627708
rect 339040 627674 339096 627708
rect 339130 627674 339186 627708
rect 339220 627674 339276 627708
rect 339310 627674 339366 627708
rect 339400 627674 339456 627708
rect 339490 627674 339546 627708
rect 339580 627674 339636 627708
rect 339670 627674 339934 627708
rect 339968 627674 340024 627708
rect 340058 627674 340114 627708
rect 340148 627674 340204 627708
rect 340238 627674 340294 627708
rect 340328 627674 340384 627708
rect 340418 627674 340474 627708
rect 340508 627674 340564 627708
rect 340598 627674 340654 627708
rect 340688 627674 340744 627708
rect 340778 627674 340834 627708
rect 340868 627674 340924 627708
rect 340958 627674 341088 627708
rect 334648 627639 341088 627674
rect 334648 627624 334749 627639
rect 334648 627590 334681 627624
rect 334715 627590 334749 627624
rect 334648 627534 334749 627590
rect 335835 627624 336037 627639
rect 335835 627590 335868 627624
rect 335902 627590 335969 627624
rect 336003 627590 336037 627624
rect 334648 627500 334681 627534
rect 334715 627500 334749 627534
rect 334648 627444 334749 627500
rect 334648 627410 334681 627444
rect 334715 627410 334749 627444
rect 334648 627354 334749 627410
rect 334648 627320 334681 627354
rect 334715 627320 334749 627354
rect 334648 627264 334749 627320
rect 334648 627230 334681 627264
rect 334715 627230 334749 627264
rect 334648 627174 334749 627230
rect 334648 627140 334681 627174
rect 334715 627140 334749 627174
rect 334648 627084 334749 627140
rect 334648 627050 334681 627084
rect 334715 627050 334749 627084
rect 334648 626994 334749 627050
rect 334648 626960 334681 626994
rect 334715 626960 334749 626994
rect 334648 626904 334749 626960
rect 334648 626870 334681 626904
rect 334715 626870 334749 626904
rect 334648 626814 334749 626870
rect 334648 626780 334681 626814
rect 334715 626780 334749 626814
rect 334648 626724 334749 626780
rect 334648 626690 334681 626724
rect 334715 626690 334749 626724
rect 334648 626634 334749 626690
rect 334648 626600 334681 626634
rect 334715 626600 334749 626634
rect 335835 627534 336037 627590
rect 337123 627624 337325 627639
rect 337123 627590 337156 627624
rect 337190 627590 337257 627624
rect 337291 627590 337325 627624
rect 335835 627500 335868 627534
rect 335902 627500 335969 627534
rect 336003 627500 336037 627534
rect 335835 627444 336037 627500
rect 335835 627410 335868 627444
rect 335902 627410 335969 627444
rect 336003 627410 336037 627444
rect 335835 627354 336037 627410
rect 335835 627320 335868 627354
rect 335902 627320 335969 627354
rect 336003 627320 336037 627354
rect 335835 627264 336037 627320
rect 335835 627230 335868 627264
rect 335902 627230 335969 627264
rect 336003 627230 336037 627264
rect 335835 627174 336037 627230
rect 335835 627140 335868 627174
rect 335902 627140 335969 627174
rect 336003 627140 336037 627174
rect 335835 627084 336037 627140
rect 335835 627050 335868 627084
rect 335902 627050 335969 627084
rect 336003 627050 336037 627084
rect 335835 626994 336037 627050
rect 335835 626960 335868 626994
rect 335902 626960 335969 626994
rect 336003 626960 336037 626994
rect 335835 626904 336037 626960
rect 335835 626870 335868 626904
rect 335902 626870 335969 626904
rect 336003 626870 336037 626904
rect 335835 626814 336037 626870
rect 335835 626780 335868 626814
rect 335902 626780 335969 626814
rect 336003 626780 336037 626814
rect 335835 626724 336037 626780
rect 335835 626690 335868 626724
rect 335902 626690 335969 626724
rect 336003 626690 336037 626724
rect 335835 626634 336037 626690
rect 334648 626553 334749 626600
rect 335835 626600 335868 626634
rect 335902 626600 335969 626634
rect 336003 626600 336037 626634
rect 337123 627534 337325 627590
rect 338411 627624 338613 627639
rect 338411 627590 338444 627624
rect 338478 627590 338545 627624
rect 338579 627590 338613 627624
rect 337123 627500 337156 627534
rect 337190 627500 337257 627534
rect 337291 627500 337325 627534
rect 337123 627444 337325 627500
rect 337123 627410 337156 627444
rect 337190 627410 337257 627444
rect 337291 627410 337325 627444
rect 337123 627354 337325 627410
rect 337123 627320 337156 627354
rect 337190 627320 337257 627354
rect 337291 627320 337325 627354
rect 337123 627264 337325 627320
rect 337123 627230 337156 627264
rect 337190 627230 337257 627264
rect 337291 627230 337325 627264
rect 337123 627174 337325 627230
rect 337123 627140 337156 627174
rect 337190 627140 337257 627174
rect 337291 627140 337325 627174
rect 337123 627084 337325 627140
rect 337123 627050 337156 627084
rect 337190 627050 337257 627084
rect 337291 627050 337325 627084
rect 337123 626994 337325 627050
rect 337123 626960 337156 626994
rect 337190 626960 337257 626994
rect 337291 626960 337325 626994
rect 337123 626904 337325 626960
rect 337123 626870 337156 626904
rect 337190 626870 337257 626904
rect 337291 626870 337325 626904
rect 337123 626814 337325 626870
rect 337123 626780 337156 626814
rect 337190 626780 337257 626814
rect 337291 626780 337325 626814
rect 337123 626724 337325 626780
rect 337123 626690 337156 626724
rect 337190 626690 337257 626724
rect 337291 626690 337325 626724
rect 337123 626634 337325 626690
rect 335835 626553 336037 626600
rect 337123 626600 337156 626634
rect 337190 626600 337257 626634
rect 337291 626600 337325 626634
rect 338411 627534 338613 627590
rect 339699 627624 339901 627639
rect 339699 627590 339732 627624
rect 339766 627590 339833 627624
rect 339867 627590 339901 627624
rect 338411 627500 338444 627534
rect 338478 627500 338545 627534
rect 338579 627500 338613 627534
rect 338411 627444 338613 627500
rect 338411 627410 338444 627444
rect 338478 627410 338545 627444
rect 338579 627410 338613 627444
rect 338411 627354 338613 627410
rect 338411 627320 338444 627354
rect 338478 627320 338545 627354
rect 338579 627320 338613 627354
rect 338411 627264 338613 627320
rect 338411 627230 338444 627264
rect 338478 627230 338545 627264
rect 338579 627230 338613 627264
rect 338411 627174 338613 627230
rect 338411 627140 338444 627174
rect 338478 627140 338545 627174
rect 338579 627140 338613 627174
rect 338411 627084 338613 627140
rect 338411 627050 338444 627084
rect 338478 627050 338545 627084
rect 338579 627050 338613 627084
rect 338411 626994 338613 627050
rect 338411 626960 338444 626994
rect 338478 626960 338545 626994
rect 338579 626960 338613 626994
rect 338411 626904 338613 626960
rect 338411 626870 338444 626904
rect 338478 626870 338545 626904
rect 338579 626870 338613 626904
rect 338411 626814 338613 626870
rect 338411 626780 338444 626814
rect 338478 626780 338545 626814
rect 338579 626780 338613 626814
rect 338411 626724 338613 626780
rect 338411 626690 338444 626724
rect 338478 626690 338545 626724
rect 338579 626690 338613 626724
rect 338411 626634 338613 626690
rect 337123 626553 337325 626600
rect 338411 626600 338444 626634
rect 338478 626600 338545 626634
rect 338579 626600 338613 626634
rect 339699 627534 339901 627590
rect 340987 627624 341088 627639
rect 340987 627590 341020 627624
rect 341054 627590 341088 627624
rect 339699 627500 339732 627534
rect 339766 627500 339833 627534
rect 339867 627500 339901 627534
rect 339699 627444 339901 627500
rect 339699 627410 339732 627444
rect 339766 627410 339833 627444
rect 339867 627410 339901 627444
rect 339699 627354 339901 627410
rect 339699 627320 339732 627354
rect 339766 627320 339833 627354
rect 339867 627320 339901 627354
rect 339699 627264 339901 627320
rect 339699 627230 339732 627264
rect 339766 627230 339833 627264
rect 339867 627230 339901 627264
rect 339699 627174 339901 627230
rect 339699 627140 339732 627174
rect 339766 627140 339833 627174
rect 339867 627140 339901 627174
rect 339699 627084 339901 627140
rect 339699 627050 339732 627084
rect 339766 627050 339833 627084
rect 339867 627050 339901 627084
rect 339699 626994 339901 627050
rect 339699 626960 339732 626994
rect 339766 626960 339833 626994
rect 339867 626960 339901 626994
rect 339699 626904 339901 626960
rect 339699 626870 339732 626904
rect 339766 626870 339833 626904
rect 339867 626870 339901 626904
rect 339699 626814 339901 626870
rect 339699 626780 339732 626814
rect 339766 626780 339833 626814
rect 339867 626780 339901 626814
rect 339699 626724 339901 626780
rect 339699 626690 339732 626724
rect 339766 626690 339833 626724
rect 339867 626690 339901 626724
rect 339699 626634 339901 626690
rect 338411 626553 338613 626600
rect 339699 626600 339732 626634
rect 339766 626600 339833 626634
rect 339867 626600 339901 626634
rect 340987 627534 341088 627590
rect 340987 627500 341020 627534
rect 341054 627500 341088 627534
rect 340987 627444 341088 627500
rect 340987 627410 341020 627444
rect 341054 627410 341088 627444
rect 340987 627354 341088 627410
rect 340987 627320 341020 627354
rect 341054 627320 341088 627354
rect 340987 627264 341088 627320
rect 340987 627230 341020 627264
rect 341054 627230 341088 627264
rect 340987 627174 341088 627230
rect 340987 627140 341020 627174
rect 341054 627140 341088 627174
rect 340987 627084 341088 627140
rect 340987 627050 341020 627084
rect 341054 627050 341088 627084
rect 340987 626994 341088 627050
rect 340987 626960 341020 626994
rect 341054 626960 341088 626994
rect 340987 626904 341088 626960
rect 340987 626870 341020 626904
rect 341054 626870 341088 626904
rect 340987 626814 341088 626870
rect 340987 626780 341020 626814
rect 341054 626780 341088 626814
rect 340987 626724 341088 626780
rect 340987 626690 341020 626724
rect 341054 626690 341088 626724
rect 340987 626634 341088 626690
rect 339699 626553 339901 626600
rect 340987 626600 341020 626634
rect 341054 626600 341088 626634
rect 340987 626553 341088 626600
rect 334648 626544 341088 626553
rect 334648 626510 334681 626544
rect 334715 626521 335868 626544
rect 334715 626510 334782 626521
rect 334648 626487 334782 626510
rect 334816 626487 334872 626521
rect 334906 626487 334962 626521
rect 334996 626487 335052 626521
rect 335086 626487 335142 626521
rect 335176 626487 335232 626521
rect 335266 626487 335322 626521
rect 335356 626487 335412 626521
rect 335446 626487 335502 626521
rect 335536 626487 335592 626521
rect 335626 626487 335682 626521
rect 335716 626487 335772 626521
rect 335806 626510 335868 626521
rect 335902 626510 335969 626544
rect 336003 626521 337156 626544
rect 336003 626510 336070 626521
rect 335806 626487 336070 626510
rect 336104 626487 336160 626521
rect 336194 626487 336250 626521
rect 336284 626487 336340 626521
rect 336374 626487 336430 626521
rect 336464 626487 336520 626521
rect 336554 626487 336610 626521
rect 336644 626487 336700 626521
rect 336734 626487 336790 626521
rect 336824 626487 336880 626521
rect 336914 626487 336970 626521
rect 337004 626487 337060 626521
rect 337094 626510 337156 626521
rect 337190 626510 337257 626544
rect 337291 626521 338444 626544
rect 337291 626510 337358 626521
rect 337094 626487 337358 626510
rect 337392 626487 337448 626521
rect 337482 626487 337538 626521
rect 337572 626487 337628 626521
rect 337662 626487 337718 626521
rect 337752 626487 337808 626521
rect 337842 626487 337898 626521
rect 337932 626487 337988 626521
rect 338022 626487 338078 626521
rect 338112 626487 338168 626521
rect 338202 626487 338258 626521
rect 338292 626487 338348 626521
rect 338382 626510 338444 626521
rect 338478 626510 338545 626544
rect 338579 626521 339732 626544
rect 338579 626510 338646 626521
rect 338382 626487 338646 626510
rect 338680 626487 338736 626521
rect 338770 626487 338826 626521
rect 338860 626487 338916 626521
rect 338950 626487 339006 626521
rect 339040 626487 339096 626521
rect 339130 626487 339186 626521
rect 339220 626487 339276 626521
rect 339310 626487 339366 626521
rect 339400 626487 339456 626521
rect 339490 626487 339546 626521
rect 339580 626487 339636 626521
rect 339670 626510 339732 626521
rect 339766 626510 339833 626544
rect 339867 626521 341020 626544
rect 339867 626510 339934 626521
rect 339670 626487 339934 626510
rect 339968 626487 340024 626521
rect 340058 626487 340114 626521
rect 340148 626487 340204 626521
rect 340238 626487 340294 626521
rect 340328 626487 340384 626521
rect 340418 626487 340474 626521
rect 340508 626487 340564 626521
rect 340598 626487 340654 626521
rect 340688 626487 340744 626521
rect 340778 626487 340834 626521
rect 340868 626487 340924 626521
rect 340958 626510 341020 626521
rect 341054 626510 341088 626544
rect 340958 626487 341088 626510
rect 334648 626420 341088 626487
rect 334648 626386 334782 626420
rect 334816 626386 334872 626420
rect 334906 626386 334962 626420
rect 334996 626386 335052 626420
rect 335086 626386 335142 626420
rect 335176 626386 335232 626420
rect 335266 626386 335322 626420
rect 335356 626386 335412 626420
rect 335446 626386 335502 626420
rect 335536 626386 335592 626420
rect 335626 626386 335682 626420
rect 335716 626386 335772 626420
rect 335806 626386 336070 626420
rect 336104 626386 336160 626420
rect 336194 626386 336250 626420
rect 336284 626386 336340 626420
rect 336374 626386 336430 626420
rect 336464 626386 336520 626420
rect 336554 626386 336610 626420
rect 336644 626386 336700 626420
rect 336734 626386 336790 626420
rect 336824 626386 336880 626420
rect 336914 626386 336970 626420
rect 337004 626386 337060 626420
rect 337094 626386 337358 626420
rect 337392 626386 337448 626420
rect 337482 626386 337538 626420
rect 337572 626386 337628 626420
rect 337662 626386 337718 626420
rect 337752 626386 337808 626420
rect 337842 626386 337898 626420
rect 337932 626386 337988 626420
rect 338022 626386 338078 626420
rect 338112 626386 338168 626420
rect 338202 626386 338258 626420
rect 338292 626386 338348 626420
rect 338382 626386 338646 626420
rect 338680 626386 338736 626420
rect 338770 626386 338826 626420
rect 338860 626386 338916 626420
rect 338950 626386 339006 626420
rect 339040 626386 339096 626420
rect 339130 626386 339186 626420
rect 339220 626386 339276 626420
rect 339310 626386 339366 626420
rect 339400 626386 339456 626420
rect 339490 626386 339546 626420
rect 339580 626386 339636 626420
rect 339670 626386 339934 626420
rect 339968 626386 340024 626420
rect 340058 626386 340114 626420
rect 340148 626386 340204 626420
rect 340238 626386 340294 626420
rect 340328 626386 340384 626420
rect 340418 626386 340474 626420
rect 340508 626386 340564 626420
rect 340598 626386 340654 626420
rect 340688 626386 340744 626420
rect 340778 626386 340834 626420
rect 340868 626386 340924 626420
rect 340958 626386 341088 626420
rect 334648 626351 341088 626386
rect 334648 626336 334749 626351
rect 334648 626302 334681 626336
rect 334715 626302 334749 626336
rect 334648 626246 334749 626302
rect 335835 626336 336037 626351
rect 335835 626302 335868 626336
rect 335902 626302 335969 626336
rect 336003 626302 336037 626336
rect 334648 626212 334681 626246
rect 334715 626212 334749 626246
rect 334648 626156 334749 626212
rect 334648 626122 334681 626156
rect 334715 626122 334749 626156
rect 334648 626066 334749 626122
rect 334648 626032 334681 626066
rect 334715 626032 334749 626066
rect 334648 625976 334749 626032
rect 334648 625942 334681 625976
rect 334715 625942 334749 625976
rect 334648 625886 334749 625942
rect 334648 625852 334681 625886
rect 334715 625852 334749 625886
rect 334648 625796 334749 625852
rect 334648 625762 334681 625796
rect 334715 625762 334749 625796
rect 334648 625706 334749 625762
rect 334648 625672 334681 625706
rect 334715 625672 334749 625706
rect 334648 625616 334749 625672
rect 334648 625582 334681 625616
rect 334715 625582 334749 625616
rect 334648 625526 334749 625582
rect 334648 625492 334681 625526
rect 334715 625492 334749 625526
rect 334648 625436 334749 625492
rect 334648 625402 334681 625436
rect 334715 625402 334749 625436
rect 334648 625346 334749 625402
rect 334648 625312 334681 625346
rect 334715 625312 334749 625346
rect 335835 626246 336037 626302
rect 337123 626336 337325 626351
rect 337123 626302 337156 626336
rect 337190 626302 337257 626336
rect 337291 626302 337325 626336
rect 335835 626212 335868 626246
rect 335902 626212 335969 626246
rect 336003 626212 336037 626246
rect 335835 626156 336037 626212
rect 335835 626122 335868 626156
rect 335902 626122 335969 626156
rect 336003 626122 336037 626156
rect 335835 626066 336037 626122
rect 335835 626032 335868 626066
rect 335902 626032 335969 626066
rect 336003 626032 336037 626066
rect 335835 625976 336037 626032
rect 335835 625942 335868 625976
rect 335902 625942 335969 625976
rect 336003 625942 336037 625976
rect 335835 625886 336037 625942
rect 335835 625852 335868 625886
rect 335902 625852 335969 625886
rect 336003 625852 336037 625886
rect 335835 625796 336037 625852
rect 335835 625762 335868 625796
rect 335902 625762 335969 625796
rect 336003 625762 336037 625796
rect 335835 625706 336037 625762
rect 335835 625672 335868 625706
rect 335902 625672 335969 625706
rect 336003 625672 336037 625706
rect 335835 625616 336037 625672
rect 335835 625582 335868 625616
rect 335902 625582 335969 625616
rect 336003 625582 336037 625616
rect 335835 625526 336037 625582
rect 335835 625492 335868 625526
rect 335902 625492 335969 625526
rect 336003 625492 336037 625526
rect 335835 625436 336037 625492
rect 335835 625402 335868 625436
rect 335902 625402 335969 625436
rect 336003 625402 336037 625436
rect 335835 625346 336037 625402
rect 334648 625265 334749 625312
rect 335835 625312 335868 625346
rect 335902 625312 335969 625346
rect 336003 625312 336037 625346
rect 337123 626246 337325 626302
rect 338411 626336 338613 626351
rect 338411 626302 338444 626336
rect 338478 626302 338545 626336
rect 338579 626302 338613 626336
rect 337123 626212 337156 626246
rect 337190 626212 337257 626246
rect 337291 626212 337325 626246
rect 337123 626156 337325 626212
rect 337123 626122 337156 626156
rect 337190 626122 337257 626156
rect 337291 626122 337325 626156
rect 337123 626066 337325 626122
rect 337123 626032 337156 626066
rect 337190 626032 337257 626066
rect 337291 626032 337325 626066
rect 337123 625976 337325 626032
rect 337123 625942 337156 625976
rect 337190 625942 337257 625976
rect 337291 625942 337325 625976
rect 337123 625886 337325 625942
rect 337123 625852 337156 625886
rect 337190 625852 337257 625886
rect 337291 625852 337325 625886
rect 337123 625796 337325 625852
rect 337123 625762 337156 625796
rect 337190 625762 337257 625796
rect 337291 625762 337325 625796
rect 337123 625706 337325 625762
rect 337123 625672 337156 625706
rect 337190 625672 337257 625706
rect 337291 625672 337325 625706
rect 337123 625616 337325 625672
rect 337123 625582 337156 625616
rect 337190 625582 337257 625616
rect 337291 625582 337325 625616
rect 337123 625526 337325 625582
rect 337123 625492 337156 625526
rect 337190 625492 337257 625526
rect 337291 625492 337325 625526
rect 337123 625436 337325 625492
rect 337123 625402 337156 625436
rect 337190 625402 337257 625436
rect 337291 625402 337325 625436
rect 337123 625346 337325 625402
rect 335835 625265 336037 625312
rect 337123 625312 337156 625346
rect 337190 625312 337257 625346
rect 337291 625312 337325 625346
rect 338411 626246 338613 626302
rect 339699 626336 339901 626351
rect 339699 626302 339732 626336
rect 339766 626302 339833 626336
rect 339867 626302 339901 626336
rect 338411 626212 338444 626246
rect 338478 626212 338545 626246
rect 338579 626212 338613 626246
rect 338411 626156 338613 626212
rect 338411 626122 338444 626156
rect 338478 626122 338545 626156
rect 338579 626122 338613 626156
rect 338411 626066 338613 626122
rect 338411 626032 338444 626066
rect 338478 626032 338545 626066
rect 338579 626032 338613 626066
rect 338411 625976 338613 626032
rect 338411 625942 338444 625976
rect 338478 625942 338545 625976
rect 338579 625942 338613 625976
rect 338411 625886 338613 625942
rect 338411 625852 338444 625886
rect 338478 625852 338545 625886
rect 338579 625852 338613 625886
rect 338411 625796 338613 625852
rect 338411 625762 338444 625796
rect 338478 625762 338545 625796
rect 338579 625762 338613 625796
rect 338411 625706 338613 625762
rect 338411 625672 338444 625706
rect 338478 625672 338545 625706
rect 338579 625672 338613 625706
rect 338411 625616 338613 625672
rect 338411 625582 338444 625616
rect 338478 625582 338545 625616
rect 338579 625582 338613 625616
rect 338411 625526 338613 625582
rect 338411 625492 338444 625526
rect 338478 625492 338545 625526
rect 338579 625492 338613 625526
rect 338411 625436 338613 625492
rect 338411 625402 338444 625436
rect 338478 625402 338545 625436
rect 338579 625402 338613 625436
rect 338411 625346 338613 625402
rect 337123 625265 337325 625312
rect 338411 625312 338444 625346
rect 338478 625312 338545 625346
rect 338579 625312 338613 625346
rect 339699 626246 339901 626302
rect 340987 626336 341088 626351
rect 340987 626302 341020 626336
rect 341054 626302 341088 626336
rect 339699 626212 339732 626246
rect 339766 626212 339833 626246
rect 339867 626212 339901 626246
rect 339699 626156 339901 626212
rect 339699 626122 339732 626156
rect 339766 626122 339833 626156
rect 339867 626122 339901 626156
rect 339699 626066 339901 626122
rect 339699 626032 339732 626066
rect 339766 626032 339833 626066
rect 339867 626032 339901 626066
rect 339699 625976 339901 626032
rect 339699 625942 339732 625976
rect 339766 625942 339833 625976
rect 339867 625942 339901 625976
rect 339699 625886 339901 625942
rect 339699 625852 339732 625886
rect 339766 625852 339833 625886
rect 339867 625852 339901 625886
rect 339699 625796 339901 625852
rect 339699 625762 339732 625796
rect 339766 625762 339833 625796
rect 339867 625762 339901 625796
rect 339699 625706 339901 625762
rect 339699 625672 339732 625706
rect 339766 625672 339833 625706
rect 339867 625672 339901 625706
rect 339699 625616 339901 625672
rect 339699 625582 339732 625616
rect 339766 625582 339833 625616
rect 339867 625582 339901 625616
rect 339699 625526 339901 625582
rect 339699 625492 339732 625526
rect 339766 625492 339833 625526
rect 339867 625492 339901 625526
rect 339699 625436 339901 625492
rect 339699 625402 339732 625436
rect 339766 625402 339833 625436
rect 339867 625402 339901 625436
rect 339699 625346 339901 625402
rect 338411 625265 338613 625312
rect 339699 625312 339732 625346
rect 339766 625312 339833 625346
rect 339867 625312 339901 625346
rect 340987 626246 341088 626302
rect 340987 626212 341020 626246
rect 341054 626212 341088 626246
rect 340987 626156 341088 626212
rect 340987 626122 341020 626156
rect 341054 626122 341088 626156
rect 340987 626066 341088 626122
rect 340987 626032 341020 626066
rect 341054 626032 341088 626066
rect 340987 625976 341088 626032
rect 340987 625942 341020 625976
rect 341054 625942 341088 625976
rect 340987 625886 341088 625942
rect 340987 625852 341020 625886
rect 341054 625852 341088 625886
rect 340987 625796 341088 625852
rect 340987 625762 341020 625796
rect 341054 625762 341088 625796
rect 340987 625706 341088 625762
rect 340987 625672 341020 625706
rect 341054 625672 341088 625706
rect 340987 625616 341088 625672
rect 340987 625582 341020 625616
rect 341054 625582 341088 625616
rect 340987 625526 341088 625582
rect 340987 625492 341020 625526
rect 341054 625492 341088 625526
rect 340987 625436 341088 625492
rect 340987 625402 341020 625436
rect 341054 625402 341088 625436
rect 340987 625346 341088 625402
rect 339699 625265 339901 625312
rect 340987 625312 341020 625346
rect 341054 625312 341088 625346
rect 340987 625265 341088 625312
rect 334648 625256 341088 625265
rect 334648 625222 334681 625256
rect 334715 625233 335868 625256
rect 334715 625222 334782 625233
rect 334648 625199 334782 625222
rect 334816 625199 334872 625233
rect 334906 625199 334962 625233
rect 334996 625199 335052 625233
rect 335086 625199 335142 625233
rect 335176 625199 335232 625233
rect 335266 625199 335322 625233
rect 335356 625199 335412 625233
rect 335446 625199 335502 625233
rect 335536 625199 335592 625233
rect 335626 625199 335682 625233
rect 335716 625199 335772 625233
rect 335806 625222 335868 625233
rect 335902 625222 335969 625256
rect 336003 625233 337156 625256
rect 336003 625222 336070 625233
rect 335806 625199 336070 625222
rect 336104 625199 336160 625233
rect 336194 625199 336250 625233
rect 336284 625199 336340 625233
rect 336374 625199 336430 625233
rect 336464 625199 336520 625233
rect 336554 625199 336610 625233
rect 336644 625199 336700 625233
rect 336734 625199 336790 625233
rect 336824 625199 336880 625233
rect 336914 625199 336970 625233
rect 337004 625199 337060 625233
rect 337094 625222 337156 625233
rect 337190 625222 337257 625256
rect 337291 625233 338444 625256
rect 337291 625222 337358 625233
rect 337094 625199 337358 625222
rect 337392 625199 337448 625233
rect 337482 625199 337538 625233
rect 337572 625199 337628 625233
rect 337662 625199 337718 625233
rect 337752 625199 337808 625233
rect 337842 625199 337898 625233
rect 337932 625199 337988 625233
rect 338022 625199 338078 625233
rect 338112 625199 338168 625233
rect 338202 625199 338258 625233
rect 338292 625199 338348 625233
rect 338382 625222 338444 625233
rect 338478 625222 338545 625256
rect 338579 625233 339732 625256
rect 338579 625222 338646 625233
rect 338382 625199 338646 625222
rect 338680 625199 338736 625233
rect 338770 625199 338826 625233
rect 338860 625199 338916 625233
rect 338950 625199 339006 625233
rect 339040 625199 339096 625233
rect 339130 625199 339186 625233
rect 339220 625199 339276 625233
rect 339310 625199 339366 625233
rect 339400 625199 339456 625233
rect 339490 625199 339546 625233
rect 339580 625199 339636 625233
rect 339670 625222 339732 625233
rect 339766 625222 339833 625256
rect 339867 625233 341020 625256
rect 339867 625222 339934 625233
rect 339670 625199 339934 625222
rect 339968 625199 340024 625233
rect 340058 625199 340114 625233
rect 340148 625199 340204 625233
rect 340238 625199 340294 625233
rect 340328 625199 340384 625233
rect 340418 625199 340474 625233
rect 340508 625199 340564 625233
rect 340598 625199 340654 625233
rect 340688 625199 340744 625233
rect 340778 625199 340834 625233
rect 340868 625199 340924 625233
rect 340958 625222 341020 625233
rect 341054 625222 341088 625256
rect 340958 625199 341088 625222
rect 334648 625132 341088 625199
rect 334648 625098 334782 625132
rect 334816 625098 334872 625132
rect 334906 625098 334962 625132
rect 334996 625098 335052 625132
rect 335086 625098 335142 625132
rect 335176 625098 335232 625132
rect 335266 625098 335322 625132
rect 335356 625098 335412 625132
rect 335446 625098 335502 625132
rect 335536 625098 335592 625132
rect 335626 625098 335682 625132
rect 335716 625098 335772 625132
rect 335806 625098 336070 625132
rect 336104 625098 336160 625132
rect 336194 625098 336250 625132
rect 336284 625098 336340 625132
rect 336374 625098 336430 625132
rect 336464 625098 336520 625132
rect 336554 625098 336610 625132
rect 336644 625098 336700 625132
rect 336734 625098 336790 625132
rect 336824 625098 336880 625132
rect 336914 625098 336970 625132
rect 337004 625098 337060 625132
rect 337094 625098 337358 625132
rect 337392 625098 337448 625132
rect 337482 625098 337538 625132
rect 337572 625098 337628 625132
rect 337662 625098 337718 625132
rect 337752 625098 337808 625132
rect 337842 625098 337898 625132
rect 337932 625098 337988 625132
rect 338022 625098 338078 625132
rect 338112 625098 338168 625132
rect 338202 625098 338258 625132
rect 338292 625098 338348 625132
rect 338382 625098 338646 625132
rect 338680 625098 338736 625132
rect 338770 625098 338826 625132
rect 338860 625098 338916 625132
rect 338950 625098 339006 625132
rect 339040 625098 339096 625132
rect 339130 625098 339186 625132
rect 339220 625098 339276 625132
rect 339310 625098 339366 625132
rect 339400 625098 339456 625132
rect 339490 625098 339546 625132
rect 339580 625098 339636 625132
rect 339670 625098 339934 625132
rect 339968 625098 340024 625132
rect 340058 625098 340114 625132
rect 340148 625098 340204 625132
rect 340238 625098 340294 625132
rect 340328 625098 340384 625132
rect 340418 625098 340474 625132
rect 340508 625098 340564 625132
rect 340598 625098 340654 625132
rect 340688 625098 340744 625132
rect 340778 625098 340834 625132
rect 340868 625098 340924 625132
rect 340958 625098 341088 625132
rect 334648 625063 341088 625098
rect 334648 625048 334749 625063
rect 334648 625014 334681 625048
rect 334715 625014 334749 625048
rect 334648 624958 334749 625014
rect 335835 625048 336037 625063
rect 335835 625014 335868 625048
rect 335902 625014 335969 625048
rect 336003 625014 336037 625048
rect 304298 624888 310798 624912
rect 304298 624556 304322 624888
rect 310774 624556 310798 624888
rect 304298 624532 310798 624556
rect 304720 622148 304920 622248
rect 299872 621342 303692 621366
rect 299872 621266 301286 621342
rect 302278 621266 303692 621342
rect 299872 621242 303692 621266
rect 299876 621188 300324 621242
rect 299876 620612 299900 621188
rect 300300 620612 300324 621188
rect 303242 621188 303690 621242
rect 303242 620612 303266 621188
rect 303666 620612 303690 621188
rect 299876 620588 300324 620612
rect 303242 620588 303690 620612
rect 304720 620548 304770 622148
rect 304870 620548 304920 622148
rect 304720 620448 304920 620548
rect 310220 622148 310420 622248
rect 310220 620548 310270 622148
rect 310370 620548 310420 622148
rect 310220 620448 310420 620548
rect 334648 624924 334681 624958
rect 334715 624924 334749 624958
rect 334648 624868 334749 624924
rect 334648 624834 334681 624868
rect 334715 624834 334749 624868
rect 334648 624778 334749 624834
rect 334648 624744 334681 624778
rect 334715 624744 334749 624778
rect 334648 624688 334749 624744
rect 334648 624654 334681 624688
rect 334715 624654 334749 624688
rect 334648 624598 334749 624654
rect 334648 624564 334681 624598
rect 334715 624564 334749 624598
rect 334648 624508 334749 624564
rect 334648 624474 334681 624508
rect 334715 624474 334749 624508
rect 334648 624418 334749 624474
rect 334648 624384 334681 624418
rect 334715 624384 334749 624418
rect 334648 624328 334749 624384
rect 334648 624294 334681 624328
rect 334715 624294 334749 624328
rect 334648 624238 334749 624294
rect 334648 624204 334681 624238
rect 334715 624204 334749 624238
rect 334648 624148 334749 624204
rect 334648 624114 334681 624148
rect 334715 624114 334749 624148
rect 334648 624058 334749 624114
rect 334648 624024 334681 624058
rect 334715 624024 334749 624058
rect 335835 624958 336037 625014
rect 337123 625048 337325 625063
rect 337123 625014 337156 625048
rect 337190 625014 337257 625048
rect 337291 625014 337325 625048
rect 335835 624924 335868 624958
rect 335902 624924 335969 624958
rect 336003 624924 336037 624958
rect 335835 624868 336037 624924
rect 335835 624834 335868 624868
rect 335902 624834 335969 624868
rect 336003 624834 336037 624868
rect 335835 624778 336037 624834
rect 335835 624744 335868 624778
rect 335902 624744 335969 624778
rect 336003 624744 336037 624778
rect 335835 624688 336037 624744
rect 335835 624654 335868 624688
rect 335902 624654 335969 624688
rect 336003 624654 336037 624688
rect 335835 624598 336037 624654
rect 335835 624564 335868 624598
rect 335902 624564 335969 624598
rect 336003 624564 336037 624598
rect 335835 624508 336037 624564
rect 335835 624474 335868 624508
rect 335902 624474 335969 624508
rect 336003 624474 336037 624508
rect 335835 624418 336037 624474
rect 335835 624384 335868 624418
rect 335902 624384 335969 624418
rect 336003 624384 336037 624418
rect 335835 624328 336037 624384
rect 335835 624294 335868 624328
rect 335902 624294 335969 624328
rect 336003 624294 336037 624328
rect 335835 624238 336037 624294
rect 335835 624204 335868 624238
rect 335902 624204 335969 624238
rect 336003 624204 336037 624238
rect 335835 624148 336037 624204
rect 335835 624114 335868 624148
rect 335902 624114 335969 624148
rect 336003 624114 336037 624148
rect 335835 624058 336037 624114
rect 334648 623977 334749 624024
rect 335835 624024 335868 624058
rect 335902 624024 335969 624058
rect 336003 624024 336037 624058
rect 337123 624958 337325 625014
rect 338411 625048 338613 625063
rect 338411 625014 338444 625048
rect 338478 625014 338545 625048
rect 338579 625014 338613 625048
rect 337123 624924 337156 624958
rect 337190 624924 337257 624958
rect 337291 624924 337325 624958
rect 337123 624868 337325 624924
rect 337123 624834 337156 624868
rect 337190 624834 337257 624868
rect 337291 624834 337325 624868
rect 337123 624778 337325 624834
rect 337123 624744 337156 624778
rect 337190 624744 337257 624778
rect 337291 624744 337325 624778
rect 337123 624688 337325 624744
rect 337123 624654 337156 624688
rect 337190 624654 337257 624688
rect 337291 624654 337325 624688
rect 337123 624598 337325 624654
rect 337123 624564 337156 624598
rect 337190 624564 337257 624598
rect 337291 624564 337325 624598
rect 337123 624508 337325 624564
rect 337123 624474 337156 624508
rect 337190 624474 337257 624508
rect 337291 624474 337325 624508
rect 337123 624418 337325 624474
rect 337123 624384 337156 624418
rect 337190 624384 337257 624418
rect 337291 624384 337325 624418
rect 337123 624328 337325 624384
rect 337123 624294 337156 624328
rect 337190 624294 337257 624328
rect 337291 624294 337325 624328
rect 337123 624238 337325 624294
rect 337123 624204 337156 624238
rect 337190 624204 337257 624238
rect 337291 624204 337325 624238
rect 337123 624148 337325 624204
rect 337123 624114 337156 624148
rect 337190 624114 337257 624148
rect 337291 624114 337325 624148
rect 337123 624058 337325 624114
rect 335835 623977 336037 624024
rect 337123 624024 337156 624058
rect 337190 624024 337257 624058
rect 337291 624024 337325 624058
rect 338411 624958 338613 625014
rect 339699 625048 339901 625063
rect 339699 625014 339732 625048
rect 339766 625014 339833 625048
rect 339867 625014 339901 625048
rect 338411 624924 338444 624958
rect 338478 624924 338545 624958
rect 338579 624924 338613 624958
rect 338411 624868 338613 624924
rect 338411 624834 338444 624868
rect 338478 624834 338545 624868
rect 338579 624834 338613 624868
rect 338411 624778 338613 624834
rect 338411 624744 338444 624778
rect 338478 624744 338545 624778
rect 338579 624744 338613 624778
rect 338411 624688 338613 624744
rect 338411 624654 338444 624688
rect 338478 624654 338545 624688
rect 338579 624654 338613 624688
rect 338411 624598 338613 624654
rect 338411 624564 338444 624598
rect 338478 624564 338545 624598
rect 338579 624564 338613 624598
rect 338411 624508 338613 624564
rect 338411 624474 338444 624508
rect 338478 624474 338545 624508
rect 338579 624474 338613 624508
rect 338411 624418 338613 624474
rect 338411 624384 338444 624418
rect 338478 624384 338545 624418
rect 338579 624384 338613 624418
rect 338411 624328 338613 624384
rect 338411 624294 338444 624328
rect 338478 624294 338545 624328
rect 338579 624294 338613 624328
rect 338411 624238 338613 624294
rect 338411 624204 338444 624238
rect 338478 624204 338545 624238
rect 338579 624204 338613 624238
rect 338411 624148 338613 624204
rect 338411 624114 338444 624148
rect 338478 624114 338545 624148
rect 338579 624114 338613 624148
rect 338411 624058 338613 624114
rect 337123 623977 337325 624024
rect 338411 624024 338444 624058
rect 338478 624024 338545 624058
rect 338579 624024 338613 624058
rect 339699 624958 339901 625014
rect 340987 625048 341088 625063
rect 340987 625014 341020 625048
rect 341054 625014 341088 625048
rect 339699 624924 339732 624958
rect 339766 624924 339833 624958
rect 339867 624924 339901 624958
rect 339699 624868 339901 624924
rect 339699 624834 339732 624868
rect 339766 624834 339833 624868
rect 339867 624834 339901 624868
rect 339699 624778 339901 624834
rect 339699 624744 339732 624778
rect 339766 624744 339833 624778
rect 339867 624744 339901 624778
rect 339699 624688 339901 624744
rect 339699 624654 339732 624688
rect 339766 624654 339833 624688
rect 339867 624654 339901 624688
rect 339699 624598 339901 624654
rect 339699 624564 339732 624598
rect 339766 624564 339833 624598
rect 339867 624564 339901 624598
rect 339699 624508 339901 624564
rect 339699 624474 339732 624508
rect 339766 624474 339833 624508
rect 339867 624474 339901 624508
rect 339699 624418 339901 624474
rect 339699 624384 339732 624418
rect 339766 624384 339833 624418
rect 339867 624384 339901 624418
rect 339699 624328 339901 624384
rect 339699 624294 339732 624328
rect 339766 624294 339833 624328
rect 339867 624294 339901 624328
rect 339699 624238 339901 624294
rect 339699 624204 339732 624238
rect 339766 624204 339833 624238
rect 339867 624204 339901 624238
rect 339699 624148 339901 624204
rect 339699 624114 339732 624148
rect 339766 624114 339833 624148
rect 339867 624114 339901 624148
rect 339699 624058 339901 624114
rect 338411 623977 338613 624024
rect 339699 624024 339732 624058
rect 339766 624024 339833 624058
rect 339867 624024 339901 624058
rect 340987 624958 341088 625014
rect 340987 624924 341020 624958
rect 341054 624924 341088 624958
rect 340987 624868 341088 624924
rect 340987 624834 341020 624868
rect 341054 624834 341088 624868
rect 340987 624778 341088 624834
rect 340987 624744 341020 624778
rect 341054 624744 341088 624778
rect 340987 624688 341088 624744
rect 340987 624654 341020 624688
rect 341054 624654 341088 624688
rect 340987 624598 341088 624654
rect 340987 624564 341020 624598
rect 341054 624564 341088 624598
rect 340987 624508 341088 624564
rect 340987 624474 341020 624508
rect 341054 624474 341088 624508
rect 340987 624418 341088 624474
rect 340987 624384 341020 624418
rect 341054 624384 341088 624418
rect 340987 624328 341088 624384
rect 340987 624294 341020 624328
rect 341054 624294 341088 624328
rect 340987 624238 341088 624294
rect 340987 624204 341020 624238
rect 341054 624204 341088 624238
rect 340987 624148 341088 624204
rect 340987 624114 341020 624148
rect 341054 624114 341088 624148
rect 340987 624058 341088 624114
rect 339699 623977 339901 624024
rect 340987 624024 341020 624058
rect 341054 624024 341088 624058
rect 340987 623977 341088 624024
rect 334648 623968 341088 623977
rect 334648 623934 334681 623968
rect 334715 623945 335868 623968
rect 334715 623934 334782 623945
rect 334648 623911 334782 623934
rect 334816 623911 334872 623945
rect 334906 623911 334962 623945
rect 334996 623911 335052 623945
rect 335086 623911 335142 623945
rect 335176 623911 335232 623945
rect 335266 623911 335322 623945
rect 335356 623911 335412 623945
rect 335446 623911 335502 623945
rect 335536 623911 335592 623945
rect 335626 623911 335682 623945
rect 335716 623911 335772 623945
rect 335806 623934 335868 623945
rect 335902 623934 335969 623968
rect 336003 623945 337156 623968
rect 336003 623934 336070 623945
rect 335806 623911 336070 623934
rect 336104 623911 336160 623945
rect 336194 623911 336250 623945
rect 336284 623911 336340 623945
rect 336374 623911 336430 623945
rect 336464 623911 336520 623945
rect 336554 623911 336610 623945
rect 336644 623911 336700 623945
rect 336734 623911 336790 623945
rect 336824 623911 336880 623945
rect 336914 623911 336970 623945
rect 337004 623911 337060 623945
rect 337094 623934 337156 623945
rect 337190 623934 337257 623968
rect 337291 623945 338444 623968
rect 337291 623934 337358 623945
rect 337094 623911 337358 623934
rect 337392 623911 337448 623945
rect 337482 623911 337538 623945
rect 337572 623911 337628 623945
rect 337662 623911 337718 623945
rect 337752 623911 337808 623945
rect 337842 623911 337898 623945
rect 337932 623911 337988 623945
rect 338022 623911 338078 623945
rect 338112 623911 338168 623945
rect 338202 623911 338258 623945
rect 338292 623911 338348 623945
rect 338382 623934 338444 623945
rect 338478 623934 338545 623968
rect 338579 623945 339732 623968
rect 338579 623934 338646 623945
rect 338382 623911 338646 623934
rect 338680 623911 338736 623945
rect 338770 623911 338826 623945
rect 338860 623911 338916 623945
rect 338950 623911 339006 623945
rect 339040 623911 339096 623945
rect 339130 623911 339186 623945
rect 339220 623911 339276 623945
rect 339310 623911 339366 623945
rect 339400 623911 339456 623945
rect 339490 623911 339546 623945
rect 339580 623911 339636 623945
rect 339670 623934 339732 623945
rect 339766 623934 339833 623968
rect 339867 623945 341020 623968
rect 339867 623934 339934 623945
rect 339670 623911 339934 623934
rect 339968 623911 340024 623945
rect 340058 623911 340114 623945
rect 340148 623911 340204 623945
rect 340238 623911 340294 623945
rect 340328 623911 340384 623945
rect 340418 623911 340474 623945
rect 340508 623911 340564 623945
rect 340598 623911 340654 623945
rect 340688 623911 340744 623945
rect 340778 623911 340834 623945
rect 340868 623911 340924 623945
rect 340958 623934 341020 623945
rect 341054 623934 341088 623968
rect 340958 623911 341088 623934
rect 334648 623844 341088 623911
rect 334648 623810 334782 623844
rect 334816 623810 334872 623844
rect 334906 623810 334962 623844
rect 334996 623810 335052 623844
rect 335086 623810 335142 623844
rect 335176 623810 335232 623844
rect 335266 623810 335322 623844
rect 335356 623810 335412 623844
rect 335446 623810 335502 623844
rect 335536 623810 335592 623844
rect 335626 623810 335682 623844
rect 335716 623810 335772 623844
rect 335806 623810 336070 623844
rect 336104 623810 336160 623844
rect 336194 623810 336250 623844
rect 336284 623810 336340 623844
rect 336374 623810 336430 623844
rect 336464 623810 336520 623844
rect 336554 623810 336610 623844
rect 336644 623810 336700 623844
rect 336734 623810 336790 623844
rect 336824 623810 336880 623844
rect 336914 623810 336970 623844
rect 337004 623810 337060 623844
rect 337094 623810 337358 623844
rect 337392 623810 337448 623844
rect 337482 623810 337538 623844
rect 337572 623810 337628 623844
rect 337662 623810 337718 623844
rect 337752 623810 337808 623844
rect 337842 623810 337898 623844
rect 337932 623810 337988 623844
rect 338022 623810 338078 623844
rect 338112 623810 338168 623844
rect 338202 623810 338258 623844
rect 338292 623810 338348 623844
rect 338382 623810 338646 623844
rect 338680 623810 338736 623844
rect 338770 623810 338826 623844
rect 338860 623810 338916 623844
rect 338950 623810 339006 623844
rect 339040 623810 339096 623844
rect 339130 623810 339186 623844
rect 339220 623810 339276 623844
rect 339310 623810 339366 623844
rect 339400 623810 339456 623844
rect 339490 623810 339546 623844
rect 339580 623810 339636 623844
rect 339670 623810 339934 623844
rect 339968 623810 340024 623844
rect 340058 623810 340114 623844
rect 340148 623810 340204 623844
rect 340238 623810 340294 623844
rect 340328 623810 340384 623844
rect 340418 623810 340474 623844
rect 340508 623810 340564 623844
rect 340598 623810 340654 623844
rect 340688 623810 340744 623844
rect 340778 623810 340834 623844
rect 340868 623810 340924 623844
rect 340958 623810 341088 623844
rect 334648 623775 341088 623810
rect 334648 623760 334749 623775
rect 334648 623726 334681 623760
rect 334715 623726 334749 623760
rect 334648 623670 334749 623726
rect 335835 623760 336037 623775
rect 335835 623726 335868 623760
rect 335902 623726 335969 623760
rect 336003 623726 336037 623760
rect 334648 623636 334681 623670
rect 334715 623636 334749 623670
rect 334648 623580 334749 623636
rect 334648 623546 334681 623580
rect 334715 623546 334749 623580
rect 334648 623490 334749 623546
rect 334648 623456 334681 623490
rect 334715 623456 334749 623490
rect 334648 623400 334749 623456
rect 334648 623366 334681 623400
rect 334715 623366 334749 623400
rect 334648 623310 334749 623366
rect 334648 623276 334681 623310
rect 334715 623276 334749 623310
rect 334648 623220 334749 623276
rect 334648 623186 334681 623220
rect 334715 623186 334749 623220
rect 334648 623130 334749 623186
rect 334648 623096 334681 623130
rect 334715 623096 334749 623130
rect 334648 623040 334749 623096
rect 334648 623006 334681 623040
rect 334715 623006 334749 623040
rect 334648 622950 334749 623006
rect 334648 622916 334681 622950
rect 334715 622916 334749 622950
rect 334648 622860 334749 622916
rect 334648 622826 334681 622860
rect 334715 622826 334749 622860
rect 334648 622770 334749 622826
rect 334648 622736 334681 622770
rect 334715 622736 334749 622770
rect 335835 623670 336037 623726
rect 337123 623760 337325 623775
rect 337123 623726 337156 623760
rect 337190 623726 337257 623760
rect 337291 623726 337325 623760
rect 335835 623636 335868 623670
rect 335902 623636 335969 623670
rect 336003 623636 336037 623670
rect 335835 623580 336037 623636
rect 335835 623546 335868 623580
rect 335902 623546 335969 623580
rect 336003 623546 336037 623580
rect 335835 623490 336037 623546
rect 335835 623456 335868 623490
rect 335902 623456 335969 623490
rect 336003 623456 336037 623490
rect 335835 623400 336037 623456
rect 335835 623366 335868 623400
rect 335902 623366 335969 623400
rect 336003 623366 336037 623400
rect 335835 623310 336037 623366
rect 335835 623276 335868 623310
rect 335902 623276 335969 623310
rect 336003 623276 336037 623310
rect 335835 623220 336037 623276
rect 335835 623186 335868 623220
rect 335902 623186 335969 623220
rect 336003 623186 336037 623220
rect 335835 623130 336037 623186
rect 335835 623096 335868 623130
rect 335902 623096 335969 623130
rect 336003 623096 336037 623130
rect 335835 623040 336037 623096
rect 335835 623006 335868 623040
rect 335902 623006 335969 623040
rect 336003 623006 336037 623040
rect 335835 622950 336037 623006
rect 335835 622916 335868 622950
rect 335902 622916 335969 622950
rect 336003 622916 336037 622950
rect 335835 622860 336037 622916
rect 335835 622826 335868 622860
rect 335902 622826 335969 622860
rect 336003 622826 336037 622860
rect 335835 622770 336037 622826
rect 334648 622689 334749 622736
rect 335835 622736 335868 622770
rect 335902 622736 335969 622770
rect 336003 622736 336037 622770
rect 337123 623670 337325 623726
rect 338411 623760 338613 623775
rect 338411 623726 338444 623760
rect 338478 623726 338545 623760
rect 338579 623726 338613 623760
rect 337123 623636 337156 623670
rect 337190 623636 337257 623670
rect 337291 623636 337325 623670
rect 337123 623580 337325 623636
rect 337123 623546 337156 623580
rect 337190 623546 337257 623580
rect 337291 623546 337325 623580
rect 337123 623490 337325 623546
rect 337123 623456 337156 623490
rect 337190 623456 337257 623490
rect 337291 623456 337325 623490
rect 337123 623400 337325 623456
rect 337123 623366 337156 623400
rect 337190 623366 337257 623400
rect 337291 623366 337325 623400
rect 337123 623310 337325 623366
rect 337123 623276 337156 623310
rect 337190 623276 337257 623310
rect 337291 623276 337325 623310
rect 337123 623220 337325 623276
rect 337123 623186 337156 623220
rect 337190 623186 337257 623220
rect 337291 623186 337325 623220
rect 337123 623130 337325 623186
rect 337123 623096 337156 623130
rect 337190 623096 337257 623130
rect 337291 623096 337325 623130
rect 337123 623040 337325 623096
rect 337123 623006 337156 623040
rect 337190 623006 337257 623040
rect 337291 623006 337325 623040
rect 337123 622950 337325 623006
rect 337123 622916 337156 622950
rect 337190 622916 337257 622950
rect 337291 622916 337325 622950
rect 337123 622860 337325 622916
rect 337123 622826 337156 622860
rect 337190 622826 337257 622860
rect 337291 622826 337325 622860
rect 337123 622770 337325 622826
rect 335835 622689 336037 622736
rect 337123 622736 337156 622770
rect 337190 622736 337257 622770
rect 337291 622736 337325 622770
rect 338411 623670 338613 623726
rect 339699 623760 339901 623775
rect 339699 623726 339732 623760
rect 339766 623726 339833 623760
rect 339867 623726 339901 623760
rect 338411 623636 338444 623670
rect 338478 623636 338545 623670
rect 338579 623636 338613 623670
rect 338411 623580 338613 623636
rect 338411 623546 338444 623580
rect 338478 623546 338545 623580
rect 338579 623546 338613 623580
rect 338411 623490 338613 623546
rect 338411 623456 338444 623490
rect 338478 623456 338545 623490
rect 338579 623456 338613 623490
rect 338411 623400 338613 623456
rect 338411 623366 338444 623400
rect 338478 623366 338545 623400
rect 338579 623366 338613 623400
rect 338411 623310 338613 623366
rect 338411 623276 338444 623310
rect 338478 623276 338545 623310
rect 338579 623276 338613 623310
rect 338411 623220 338613 623276
rect 338411 623186 338444 623220
rect 338478 623186 338545 623220
rect 338579 623186 338613 623220
rect 338411 623130 338613 623186
rect 338411 623096 338444 623130
rect 338478 623096 338545 623130
rect 338579 623096 338613 623130
rect 338411 623040 338613 623096
rect 338411 623006 338444 623040
rect 338478 623006 338545 623040
rect 338579 623006 338613 623040
rect 338411 622950 338613 623006
rect 338411 622916 338444 622950
rect 338478 622916 338545 622950
rect 338579 622916 338613 622950
rect 338411 622860 338613 622916
rect 338411 622826 338444 622860
rect 338478 622826 338545 622860
rect 338579 622826 338613 622860
rect 338411 622770 338613 622826
rect 337123 622689 337325 622736
rect 338411 622736 338444 622770
rect 338478 622736 338545 622770
rect 338579 622736 338613 622770
rect 339699 623670 339901 623726
rect 340987 623760 341088 623775
rect 340987 623726 341020 623760
rect 341054 623726 341088 623760
rect 339699 623636 339732 623670
rect 339766 623636 339833 623670
rect 339867 623636 339901 623670
rect 339699 623580 339901 623636
rect 339699 623546 339732 623580
rect 339766 623546 339833 623580
rect 339867 623546 339901 623580
rect 339699 623490 339901 623546
rect 339699 623456 339732 623490
rect 339766 623456 339833 623490
rect 339867 623456 339901 623490
rect 339699 623400 339901 623456
rect 339699 623366 339732 623400
rect 339766 623366 339833 623400
rect 339867 623366 339901 623400
rect 339699 623310 339901 623366
rect 339699 623276 339732 623310
rect 339766 623276 339833 623310
rect 339867 623276 339901 623310
rect 339699 623220 339901 623276
rect 339699 623186 339732 623220
rect 339766 623186 339833 623220
rect 339867 623186 339901 623220
rect 339699 623130 339901 623186
rect 339699 623096 339732 623130
rect 339766 623096 339833 623130
rect 339867 623096 339901 623130
rect 339699 623040 339901 623096
rect 339699 623006 339732 623040
rect 339766 623006 339833 623040
rect 339867 623006 339901 623040
rect 339699 622950 339901 623006
rect 339699 622916 339732 622950
rect 339766 622916 339833 622950
rect 339867 622916 339901 622950
rect 339699 622860 339901 622916
rect 339699 622826 339732 622860
rect 339766 622826 339833 622860
rect 339867 622826 339901 622860
rect 339699 622770 339901 622826
rect 338411 622689 338613 622736
rect 339699 622736 339732 622770
rect 339766 622736 339833 622770
rect 339867 622736 339901 622770
rect 340987 623670 341088 623726
rect 340987 623636 341020 623670
rect 341054 623636 341088 623670
rect 340987 623580 341088 623636
rect 340987 623546 341020 623580
rect 341054 623546 341088 623580
rect 340987 623490 341088 623546
rect 340987 623456 341020 623490
rect 341054 623456 341088 623490
rect 340987 623400 341088 623456
rect 340987 623366 341020 623400
rect 341054 623366 341088 623400
rect 340987 623310 341088 623366
rect 340987 623276 341020 623310
rect 341054 623276 341088 623310
rect 340987 623220 341088 623276
rect 340987 623186 341020 623220
rect 341054 623186 341088 623220
rect 340987 623130 341088 623186
rect 340987 623096 341020 623130
rect 341054 623096 341088 623130
rect 340987 623040 341088 623096
rect 340987 623006 341020 623040
rect 341054 623006 341088 623040
rect 340987 622950 341088 623006
rect 340987 622916 341020 622950
rect 341054 622916 341088 622950
rect 340987 622860 341088 622916
rect 340987 622826 341020 622860
rect 341054 622826 341088 622860
rect 340987 622770 341088 622826
rect 339699 622689 339901 622736
rect 340987 622736 341020 622770
rect 341054 622736 341088 622770
rect 340987 622689 341088 622736
rect 334648 622680 341088 622689
rect 334648 622646 334681 622680
rect 334715 622657 335868 622680
rect 334715 622646 334782 622657
rect 334648 622623 334782 622646
rect 334816 622623 334872 622657
rect 334906 622623 334962 622657
rect 334996 622623 335052 622657
rect 335086 622623 335142 622657
rect 335176 622623 335232 622657
rect 335266 622623 335322 622657
rect 335356 622623 335412 622657
rect 335446 622623 335502 622657
rect 335536 622623 335592 622657
rect 335626 622623 335682 622657
rect 335716 622623 335772 622657
rect 335806 622646 335868 622657
rect 335902 622646 335969 622680
rect 336003 622657 337156 622680
rect 336003 622646 336070 622657
rect 335806 622623 336070 622646
rect 336104 622623 336160 622657
rect 336194 622623 336250 622657
rect 336284 622623 336340 622657
rect 336374 622623 336430 622657
rect 336464 622623 336520 622657
rect 336554 622623 336610 622657
rect 336644 622623 336700 622657
rect 336734 622623 336790 622657
rect 336824 622623 336880 622657
rect 336914 622623 336970 622657
rect 337004 622623 337060 622657
rect 337094 622646 337156 622657
rect 337190 622646 337257 622680
rect 337291 622657 338444 622680
rect 337291 622646 337358 622657
rect 337094 622623 337358 622646
rect 337392 622623 337448 622657
rect 337482 622623 337538 622657
rect 337572 622623 337628 622657
rect 337662 622623 337718 622657
rect 337752 622623 337808 622657
rect 337842 622623 337898 622657
rect 337932 622623 337988 622657
rect 338022 622623 338078 622657
rect 338112 622623 338168 622657
rect 338202 622623 338258 622657
rect 338292 622623 338348 622657
rect 338382 622646 338444 622657
rect 338478 622646 338545 622680
rect 338579 622657 339732 622680
rect 338579 622646 338646 622657
rect 338382 622623 338646 622646
rect 338680 622623 338736 622657
rect 338770 622623 338826 622657
rect 338860 622623 338916 622657
rect 338950 622623 339006 622657
rect 339040 622623 339096 622657
rect 339130 622623 339186 622657
rect 339220 622623 339276 622657
rect 339310 622623 339366 622657
rect 339400 622623 339456 622657
rect 339490 622623 339546 622657
rect 339580 622623 339636 622657
rect 339670 622646 339732 622657
rect 339766 622646 339833 622680
rect 339867 622657 341020 622680
rect 339867 622646 339934 622657
rect 339670 622623 339934 622646
rect 339968 622623 340024 622657
rect 340058 622623 340114 622657
rect 340148 622623 340204 622657
rect 340238 622623 340294 622657
rect 340328 622623 340384 622657
rect 340418 622623 340474 622657
rect 340508 622623 340564 622657
rect 340598 622623 340654 622657
rect 340688 622623 340744 622657
rect 340778 622623 340834 622657
rect 340868 622623 340924 622657
rect 340958 622646 341020 622657
rect 341054 622646 341088 622680
rect 340958 622623 341088 622646
rect 334648 622556 341088 622623
rect 334648 622522 334782 622556
rect 334816 622522 334872 622556
rect 334906 622522 334962 622556
rect 334996 622522 335052 622556
rect 335086 622522 335142 622556
rect 335176 622522 335232 622556
rect 335266 622522 335322 622556
rect 335356 622522 335412 622556
rect 335446 622522 335502 622556
rect 335536 622522 335592 622556
rect 335626 622522 335682 622556
rect 335716 622522 335772 622556
rect 335806 622522 336070 622556
rect 336104 622522 336160 622556
rect 336194 622522 336250 622556
rect 336284 622522 336340 622556
rect 336374 622522 336430 622556
rect 336464 622522 336520 622556
rect 336554 622522 336610 622556
rect 336644 622522 336700 622556
rect 336734 622522 336790 622556
rect 336824 622522 336880 622556
rect 336914 622522 336970 622556
rect 337004 622522 337060 622556
rect 337094 622522 337358 622556
rect 337392 622522 337448 622556
rect 337482 622522 337538 622556
rect 337572 622522 337628 622556
rect 337662 622522 337718 622556
rect 337752 622522 337808 622556
rect 337842 622522 337898 622556
rect 337932 622522 337988 622556
rect 338022 622522 338078 622556
rect 338112 622522 338168 622556
rect 338202 622522 338258 622556
rect 338292 622522 338348 622556
rect 338382 622522 338646 622556
rect 338680 622522 338736 622556
rect 338770 622522 338826 622556
rect 338860 622522 338916 622556
rect 338950 622522 339006 622556
rect 339040 622522 339096 622556
rect 339130 622522 339186 622556
rect 339220 622522 339276 622556
rect 339310 622522 339366 622556
rect 339400 622522 339456 622556
rect 339490 622522 339546 622556
rect 339580 622522 339636 622556
rect 339670 622522 339934 622556
rect 339968 622522 340024 622556
rect 340058 622522 340114 622556
rect 340148 622522 340204 622556
rect 340238 622522 340294 622556
rect 340328 622522 340384 622556
rect 340418 622522 340474 622556
rect 340508 622522 340564 622556
rect 340598 622522 340654 622556
rect 340688 622522 340744 622556
rect 340778 622522 340834 622556
rect 340868 622522 340924 622556
rect 340958 622522 341088 622556
rect 334648 622487 341088 622522
rect 334648 622472 334749 622487
rect 334648 622438 334681 622472
rect 334715 622438 334749 622472
rect 334648 622382 334749 622438
rect 335835 622472 336037 622487
rect 335835 622438 335868 622472
rect 335902 622438 335969 622472
rect 336003 622438 336037 622472
rect 334648 622348 334681 622382
rect 334715 622348 334749 622382
rect 334648 622292 334749 622348
rect 334648 622258 334681 622292
rect 334715 622258 334749 622292
rect 334648 622202 334749 622258
rect 334648 622168 334681 622202
rect 334715 622168 334749 622202
rect 334648 622112 334749 622168
rect 334648 622078 334681 622112
rect 334715 622078 334749 622112
rect 334648 622022 334749 622078
rect 334648 621988 334681 622022
rect 334715 621988 334749 622022
rect 334648 621932 334749 621988
rect 334648 621898 334681 621932
rect 334715 621898 334749 621932
rect 334648 621842 334749 621898
rect 334648 621808 334681 621842
rect 334715 621808 334749 621842
rect 334648 621752 334749 621808
rect 334648 621718 334681 621752
rect 334715 621718 334749 621752
rect 334648 621662 334749 621718
rect 334648 621628 334681 621662
rect 334715 621628 334749 621662
rect 334648 621572 334749 621628
rect 334648 621538 334681 621572
rect 334715 621538 334749 621572
rect 334648 621482 334749 621538
rect 334648 621448 334681 621482
rect 334715 621448 334749 621482
rect 335835 622382 336037 622438
rect 337123 622472 337325 622487
rect 337123 622438 337156 622472
rect 337190 622438 337257 622472
rect 337291 622438 337325 622472
rect 335835 622348 335868 622382
rect 335902 622348 335969 622382
rect 336003 622348 336037 622382
rect 335835 622292 336037 622348
rect 335835 622258 335868 622292
rect 335902 622258 335969 622292
rect 336003 622258 336037 622292
rect 335835 622202 336037 622258
rect 335835 622168 335868 622202
rect 335902 622168 335969 622202
rect 336003 622168 336037 622202
rect 335835 622112 336037 622168
rect 335835 622078 335868 622112
rect 335902 622078 335969 622112
rect 336003 622078 336037 622112
rect 335835 622022 336037 622078
rect 335835 621988 335868 622022
rect 335902 621988 335969 622022
rect 336003 621988 336037 622022
rect 335835 621932 336037 621988
rect 335835 621898 335868 621932
rect 335902 621898 335969 621932
rect 336003 621898 336037 621932
rect 335835 621842 336037 621898
rect 335835 621808 335868 621842
rect 335902 621808 335969 621842
rect 336003 621808 336037 621842
rect 335835 621752 336037 621808
rect 335835 621718 335868 621752
rect 335902 621718 335969 621752
rect 336003 621718 336037 621752
rect 335835 621662 336037 621718
rect 335835 621628 335868 621662
rect 335902 621628 335969 621662
rect 336003 621628 336037 621662
rect 335835 621572 336037 621628
rect 335835 621538 335868 621572
rect 335902 621538 335969 621572
rect 336003 621538 336037 621572
rect 335835 621482 336037 621538
rect 334648 621401 334749 621448
rect 335835 621448 335868 621482
rect 335902 621448 335969 621482
rect 336003 621448 336037 621482
rect 337123 622382 337325 622438
rect 338411 622472 338613 622487
rect 338411 622438 338444 622472
rect 338478 622438 338545 622472
rect 338579 622438 338613 622472
rect 337123 622348 337156 622382
rect 337190 622348 337257 622382
rect 337291 622348 337325 622382
rect 337123 622292 337325 622348
rect 337123 622258 337156 622292
rect 337190 622258 337257 622292
rect 337291 622258 337325 622292
rect 337123 622202 337325 622258
rect 337123 622168 337156 622202
rect 337190 622168 337257 622202
rect 337291 622168 337325 622202
rect 337123 622112 337325 622168
rect 337123 622078 337156 622112
rect 337190 622078 337257 622112
rect 337291 622078 337325 622112
rect 337123 622022 337325 622078
rect 337123 621988 337156 622022
rect 337190 621988 337257 622022
rect 337291 621988 337325 622022
rect 337123 621932 337325 621988
rect 337123 621898 337156 621932
rect 337190 621898 337257 621932
rect 337291 621898 337325 621932
rect 337123 621842 337325 621898
rect 337123 621808 337156 621842
rect 337190 621808 337257 621842
rect 337291 621808 337325 621842
rect 337123 621752 337325 621808
rect 337123 621718 337156 621752
rect 337190 621718 337257 621752
rect 337291 621718 337325 621752
rect 337123 621662 337325 621718
rect 337123 621628 337156 621662
rect 337190 621628 337257 621662
rect 337291 621628 337325 621662
rect 337123 621572 337325 621628
rect 337123 621538 337156 621572
rect 337190 621538 337257 621572
rect 337291 621538 337325 621572
rect 337123 621482 337325 621538
rect 335835 621401 336037 621448
rect 337123 621448 337156 621482
rect 337190 621448 337257 621482
rect 337291 621448 337325 621482
rect 338411 622382 338613 622438
rect 339699 622472 339901 622487
rect 339699 622438 339732 622472
rect 339766 622438 339833 622472
rect 339867 622438 339901 622472
rect 338411 622348 338444 622382
rect 338478 622348 338545 622382
rect 338579 622348 338613 622382
rect 338411 622292 338613 622348
rect 338411 622258 338444 622292
rect 338478 622258 338545 622292
rect 338579 622258 338613 622292
rect 338411 622202 338613 622258
rect 338411 622168 338444 622202
rect 338478 622168 338545 622202
rect 338579 622168 338613 622202
rect 338411 622112 338613 622168
rect 338411 622078 338444 622112
rect 338478 622078 338545 622112
rect 338579 622078 338613 622112
rect 338411 622022 338613 622078
rect 338411 621988 338444 622022
rect 338478 621988 338545 622022
rect 338579 621988 338613 622022
rect 338411 621932 338613 621988
rect 338411 621898 338444 621932
rect 338478 621898 338545 621932
rect 338579 621898 338613 621932
rect 338411 621842 338613 621898
rect 338411 621808 338444 621842
rect 338478 621808 338545 621842
rect 338579 621808 338613 621842
rect 338411 621752 338613 621808
rect 338411 621718 338444 621752
rect 338478 621718 338545 621752
rect 338579 621718 338613 621752
rect 338411 621662 338613 621718
rect 338411 621628 338444 621662
rect 338478 621628 338545 621662
rect 338579 621628 338613 621662
rect 338411 621572 338613 621628
rect 338411 621538 338444 621572
rect 338478 621538 338545 621572
rect 338579 621538 338613 621572
rect 338411 621482 338613 621538
rect 337123 621401 337325 621448
rect 338411 621448 338444 621482
rect 338478 621448 338545 621482
rect 338579 621448 338613 621482
rect 339699 622382 339901 622438
rect 340987 622472 341088 622487
rect 340987 622438 341020 622472
rect 341054 622438 341088 622472
rect 339699 622348 339732 622382
rect 339766 622348 339833 622382
rect 339867 622348 339901 622382
rect 339699 622292 339901 622348
rect 339699 622258 339732 622292
rect 339766 622258 339833 622292
rect 339867 622258 339901 622292
rect 339699 622202 339901 622258
rect 339699 622168 339732 622202
rect 339766 622168 339833 622202
rect 339867 622168 339901 622202
rect 339699 622112 339901 622168
rect 339699 622078 339732 622112
rect 339766 622078 339833 622112
rect 339867 622078 339901 622112
rect 339699 622022 339901 622078
rect 339699 621988 339732 622022
rect 339766 621988 339833 622022
rect 339867 621988 339901 622022
rect 339699 621932 339901 621988
rect 339699 621898 339732 621932
rect 339766 621898 339833 621932
rect 339867 621898 339901 621932
rect 339699 621842 339901 621898
rect 339699 621808 339732 621842
rect 339766 621808 339833 621842
rect 339867 621808 339901 621842
rect 339699 621752 339901 621808
rect 339699 621718 339732 621752
rect 339766 621718 339833 621752
rect 339867 621718 339901 621752
rect 339699 621662 339901 621718
rect 339699 621628 339732 621662
rect 339766 621628 339833 621662
rect 339867 621628 339901 621662
rect 339699 621572 339901 621628
rect 339699 621538 339732 621572
rect 339766 621538 339833 621572
rect 339867 621538 339901 621572
rect 339699 621482 339901 621538
rect 338411 621401 338613 621448
rect 339699 621448 339732 621482
rect 339766 621448 339833 621482
rect 339867 621448 339901 621482
rect 340987 622382 341088 622438
rect 340987 622348 341020 622382
rect 341054 622348 341088 622382
rect 340987 622292 341088 622348
rect 340987 622258 341020 622292
rect 341054 622258 341088 622292
rect 340987 622202 341088 622258
rect 340987 622168 341020 622202
rect 341054 622168 341088 622202
rect 340987 622112 341088 622168
rect 340987 622078 341020 622112
rect 341054 622078 341088 622112
rect 340987 622022 341088 622078
rect 340987 621988 341020 622022
rect 341054 621988 341088 622022
rect 340987 621932 341088 621988
rect 340987 621898 341020 621932
rect 341054 621898 341088 621932
rect 340987 621842 341088 621898
rect 340987 621808 341020 621842
rect 341054 621808 341088 621842
rect 340987 621752 341088 621808
rect 340987 621718 341020 621752
rect 341054 621718 341088 621752
rect 340987 621662 341088 621718
rect 340987 621628 341020 621662
rect 341054 621628 341088 621662
rect 340987 621572 341088 621628
rect 340987 621538 341020 621572
rect 341054 621538 341088 621572
rect 340987 621482 341088 621538
rect 339699 621401 339901 621448
rect 340987 621448 341020 621482
rect 341054 621448 341088 621482
rect 340987 621401 341088 621448
rect 334648 621392 341088 621401
rect 334648 621358 334681 621392
rect 334715 621369 335868 621392
rect 334715 621358 334782 621369
rect 334648 621335 334782 621358
rect 334816 621335 334872 621369
rect 334906 621335 334962 621369
rect 334996 621335 335052 621369
rect 335086 621335 335142 621369
rect 335176 621335 335232 621369
rect 335266 621335 335322 621369
rect 335356 621335 335412 621369
rect 335446 621335 335502 621369
rect 335536 621335 335592 621369
rect 335626 621335 335682 621369
rect 335716 621335 335772 621369
rect 335806 621358 335868 621369
rect 335902 621358 335969 621392
rect 336003 621369 337156 621392
rect 336003 621358 336070 621369
rect 335806 621335 336070 621358
rect 336104 621335 336160 621369
rect 336194 621335 336250 621369
rect 336284 621335 336340 621369
rect 336374 621335 336430 621369
rect 336464 621335 336520 621369
rect 336554 621335 336610 621369
rect 336644 621335 336700 621369
rect 336734 621335 336790 621369
rect 336824 621335 336880 621369
rect 336914 621335 336970 621369
rect 337004 621335 337060 621369
rect 337094 621358 337156 621369
rect 337190 621358 337257 621392
rect 337291 621369 338444 621392
rect 337291 621358 337358 621369
rect 337094 621335 337358 621358
rect 337392 621335 337448 621369
rect 337482 621335 337538 621369
rect 337572 621335 337628 621369
rect 337662 621335 337718 621369
rect 337752 621335 337808 621369
rect 337842 621335 337898 621369
rect 337932 621335 337988 621369
rect 338022 621335 338078 621369
rect 338112 621335 338168 621369
rect 338202 621335 338258 621369
rect 338292 621335 338348 621369
rect 338382 621358 338444 621369
rect 338478 621358 338545 621392
rect 338579 621369 339732 621392
rect 338579 621358 338646 621369
rect 338382 621335 338646 621358
rect 338680 621335 338736 621369
rect 338770 621335 338826 621369
rect 338860 621335 338916 621369
rect 338950 621335 339006 621369
rect 339040 621335 339096 621369
rect 339130 621335 339186 621369
rect 339220 621335 339276 621369
rect 339310 621335 339366 621369
rect 339400 621335 339456 621369
rect 339490 621335 339546 621369
rect 339580 621335 339636 621369
rect 339670 621358 339732 621369
rect 339766 621358 339833 621392
rect 339867 621369 341020 621392
rect 339867 621358 339934 621369
rect 339670 621335 339934 621358
rect 339968 621335 340024 621369
rect 340058 621335 340114 621369
rect 340148 621335 340204 621369
rect 340238 621335 340294 621369
rect 340328 621335 340384 621369
rect 340418 621335 340474 621369
rect 340508 621335 340564 621369
rect 340598 621335 340654 621369
rect 340688 621335 340744 621369
rect 340778 621335 340834 621369
rect 340868 621335 340924 621369
rect 340958 621358 341020 621369
rect 341054 621358 341088 621392
rect 340958 621335 341088 621358
rect 334648 621268 341088 621335
rect 334648 621234 334782 621268
rect 334816 621234 334872 621268
rect 334906 621234 334962 621268
rect 334996 621234 335052 621268
rect 335086 621234 335142 621268
rect 335176 621234 335232 621268
rect 335266 621234 335322 621268
rect 335356 621234 335412 621268
rect 335446 621234 335502 621268
rect 335536 621234 335592 621268
rect 335626 621234 335682 621268
rect 335716 621234 335772 621268
rect 335806 621234 336070 621268
rect 336104 621234 336160 621268
rect 336194 621234 336250 621268
rect 336284 621234 336340 621268
rect 336374 621234 336430 621268
rect 336464 621234 336520 621268
rect 336554 621234 336610 621268
rect 336644 621234 336700 621268
rect 336734 621234 336790 621268
rect 336824 621234 336880 621268
rect 336914 621234 336970 621268
rect 337004 621234 337060 621268
rect 337094 621234 337358 621268
rect 337392 621234 337448 621268
rect 337482 621234 337538 621268
rect 337572 621234 337628 621268
rect 337662 621234 337718 621268
rect 337752 621234 337808 621268
rect 337842 621234 337898 621268
rect 337932 621234 337988 621268
rect 338022 621234 338078 621268
rect 338112 621234 338168 621268
rect 338202 621234 338258 621268
rect 338292 621234 338348 621268
rect 338382 621234 338646 621268
rect 338680 621234 338736 621268
rect 338770 621234 338826 621268
rect 338860 621234 338916 621268
rect 338950 621234 339006 621268
rect 339040 621234 339096 621268
rect 339130 621234 339186 621268
rect 339220 621234 339276 621268
rect 339310 621234 339366 621268
rect 339400 621234 339456 621268
rect 339490 621234 339546 621268
rect 339580 621234 339636 621268
rect 339670 621234 339934 621268
rect 339968 621234 340024 621268
rect 340058 621234 340114 621268
rect 340148 621234 340204 621268
rect 340238 621234 340294 621268
rect 340328 621234 340384 621268
rect 340418 621234 340474 621268
rect 340508 621234 340564 621268
rect 340598 621234 340654 621268
rect 340688 621234 340744 621268
rect 340778 621234 340834 621268
rect 340868 621234 340924 621268
rect 340958 621234 341088 621268
rect 334648 621199 341088 621234
rect 334648 621184 334749 621199
rect 334648 621150 334681 621184
rect 334715 621150 334749 621184
rect 334648 621094 334749 621150
rect 335835 621184 336037 621199
rect 335835 621150 335868 621184
rect 335902 621150 335969 621184
rect 336003 621150 336037 621184
rect 334648 621060 334681 621094
rect 334715 621060 334749 621094
rect 334648 621004 334749 621060
rect 334648 620970 334681 621004
rect 334715 620970 334749 621004
rect 334648 620914 334749 620970
rect 334648 620880 334681 620914
rect 334715 620880 334749 620914
rect 334648 620824 334749 620880
rect 334648 620790 334681 620824
rect 334715 620790 334749 620824
rect 334648 620734 334749 620790
rect 334648 620700 334681 620734
rect 334715 620700 334749 620734
rect 334648 620644 334749 620700
rect 334648 620610 334681 620644
rect 334715 620610 334749 620644
rect 334648 620554 334749 620610
rect 334648 620520 334681 620554
rect 334715 620520 334749 620554
rect 334648 620464 334749 620520
rect 334648 620430 334681 620464
rect 334715 620430 334749 620464
rect 334648 620374 334749 620430
rect 334648 620340 334681 620374
rect 334715 620340 334749 620374
rect 334648 620284 334749 620340
rect 334648 620250 334681 620284
rect 334715 620250 334749 620284
rect 334648 620194 334749 620250
rect 334648 620160 334681 620194
rect 334715 620160 334749 620194
rect 335835 621094 336037 621150
rect 337123 621184 337325 621199
rect 337123 621150 337156 621184
rect 337190 621150 337257 621184
rect 337291 621150 337325 621184
rect 335835 621060 335868 621094
rect 335902 621060 335969 621094
rect 336003 621060 336037 621094
rect 335835 621004 336037 621060
rect 335835 620970 335868 621004
rect 335902 620970 335969 621004
rect 336003 620970 336037 621004
rect 335835 620914 336037 620970
rect 335835 620880 335868 620914
rect 335902 620880 335969 620914
rect 336003 620880 336037 620914
rect 335835 620824 336037 620880
rect 335835 620790 335868 620824
rect 335902 620790 335969 620824
rect 336003 620790 336037 620824
rect 335835 620734 336037 620790
rect 335835 620700 335868 620734
rect 335902 620700 335969 620734
rect 336003 620700 336037 620734
rect 335835 620644 336037 620700
rect 335835 620610 335868 620644
rect 335902 620610 335969 620644
rect 336003 620610 336037 620644
rect 335835 620554 336037 620610
rect 335835 620520 335868 620554
rect 335902 620520 335969 620554
rect 336003 620520 336037 620554
rect 335835 620464 336037 620520
rect 335835 620430 335868 620464
rect 335902 620430 335969 620464
rect 336003 620430 336037 620464
rect 335835 620374 336037 620430
rect 335835 620340 335868 620374
rect 335902 620340 335969 620374
rect 336003 620340 336037 620374
rect 335835 620284 336037 620340
rect 335835 620250 335868 620284
rect 335902 620250 335969 620284
rect 336003 620250 336037 620284
rect 335835 620194 336037 620250
rect 334648 620113 334749 620160
rect 335835 620160 335868 620194
rect 335902 620160 335969 620194
rect 336003 620160 336037 620194
rect 337123 621094 337325 621150
rect 338411 621184 338613 621199
rect 338411 621150 338444 621184
rect 338478 621150 338545 621184
rect 338579 621150 338613 621184
rect 337123 621060 337156 621094
rect 337190 621060 337257 621094
rect 337291 621060 337325 621094
rect 337123 621004 337325 621060
rect 337123 620970 337156 621004
rect 337190 620970 337257 621004
rect 337291 620970 337325 621004
rect 337123 620914 337325 620970
rect 337123 620880 337156 620914
rect 337190 620880 337257 620914
rect 337291 620880 337325 620914
rect 337123 620824 337325 620880
rect 337123 620790 337156 620824
rect 337190 620790 337257 620824
rect 337291 620790 337325 620824
rect 337123 620734 337325 620790
rect 337123 620700 337156 620734
rect 337190 620700 337257 620734
rect 337291 620700 337325 620734
rect 337123 620644 337325 620700
rect 337123 620610 337156 620644
rect 337190 620610 337257 620644
rect 337291 620610 337325 620644
rect 337123 620554 337325 620610
rect 337123 620520 337156 620554
rect 337190 620520 337257 620554
rect 337291 620520 337325 620554
rect 337123 620464 337325 620520
rect 337123 620430 337156 620464
rect 337190 620430 337257 620464
rect 337291 620430 337325 620464
rect 337123 620374 337325 620430
rect 337123 620340 337156 620374
rect 337190 620340 337257 620374
rect 337291 620340 337325 620374
rect 337123 620284 337325 620340
rect 337123 620250 337156 620284
rect 337190 620250 337257 620284
rect 337291 620250 337325 620284
rect 337123 620194 337325 620250
rect 335835 620113 336037 620160
rect 337123 620160 337156 620194
rect 337190 620160 337257 620194
rect 337291 620160 337325 620194
rect 338411 621094 338613 621150
rect 339699 621184 339901 621199
rect 339699 621150 339732 621184
rect 339766 621150 339833 621184
rect 339867 621150 339901 621184
rect 338411 621060 338444 621094
rect 338478 621060 338545 621094
rect 338579 621060 338613 621094
rect 338411 621004 338613 621060
rect 338411 620970 338444 621004
rect 338478 620970 338545 621004
rect 338579 620970 338613 621004
rect 338411 620914 338613 620970
rect 338411 620880 338444 620914
rect 338478 620880 338545 620914
rect 338579 620880 338613 620914
rect 338411 620824 338613 620880
rect 338411 620790 338444 620824
rect 338478 620790 338545 620824
rect 338579 620790 338613 620824
rect 338411 620734 338613 620790
rect 338411 620700 338444 620734
rect 338478 620700 338545 620734
rect 338579 620700 338613 620734
rect 338411 620644 338613 620700
rect 338411 620610 338444 620644
rect 338478 620610 338545 620644
rect 338579 620610 338613 620644
rect 338411 620554 338613 620610
rect 338411 620520 338444 620554
rect 338478 620520 338545 620554
rect 338579 620520 338613 620554
rect 338411 620464 338613 620520
rect 338411 620430 338444 620464
rect 338478 620430 338545 620464
rect 338579 620430 338613 620464
rect 338411 620374 338613 620430
rect 338411 620340 338444 620374
rect 338478 620340 338545 620374
rect 338579 620340 338613 620374
rect 338411 620284 338613 620340
rect 338411 620250 338444 620284
rect 338478 620250 338545 620284
rect 338579 620250 338613 620284
rect 338411 620194 338613 620250
rect 337123 620113 337325 620160
rect 338411 620160 338444 620194
rect 338478 620160 338545 620194
rect 338579 620160 338613 620194
rect 339699 621094 339901 621150
rect 340987 621184 341088 621199
rect 340987 621150 341020 621184
rect 341054 621150 341088 621184
rect 339699 621060 339732 621094
rect 339766 621060 339833 621094
rect 339867 621060 339901 621094
rect 339699 621004 339901 621060
rect 339699 620970 339732 621004
rect 339766 620970 339833 621004
rect 339867 620970 339901 621004
rect 339699 620914 339901 620970
rect 339699 620880 339732 620914
rect 339766 620880 339833 620914
rect 339867 620880 339901 620914
rect 339699 620824 339901 620880
rect 339699 620790 339732 620824
rect 339766 620790 339833 620824
rect 339867 620790 339901 620824
rect 339699 620734 339901 620790
rect 339699 620700 339732 620734
rect 339766 620700 339833 620734
rect 339867 620700 339901 620734
rect 339699 620644 339901 620700
rect 339699 620610 339732 620644
rect 339766 620610 339833 620644
rect 339867 620610 339901 620644
rect 339699 620554 339901 620610
rect 339699 620520 339732 620554
rect 339766 620520 339833 620554
rect 339867 620520 339901 620554
rect 339699 620464 339901 620520
rect 339699 620430 339732 620464
rect 339766 620430 339833 620464
rect 339867 620430 339901 620464
rect 339699 620374 339901 620430
rect 339699 620340 339732 620374
rect 339766 620340 339833 620374
rect 339867 620340 339901 620374
rect 339699 620284 339901 620340
rect 339699 620250 339732 620284
rect 339766 620250 339833 620284
rect 339867 620250 339901 620284
rect 339699 620194 339901 620250
rect 338411 620113 338613 620160
rect 339699 620160 339732 620194
rect 339766 620160 339833 620194
rect 339867 620160 339901 620194
rect 340987 621094 341088 621150
rect 340987 621060 341020 621094
rect 341054 621060 341088 621094
rect 340987 621004 341088 621060
rect 340987 620970 341020 621004
rect 341054 620970 341088 621004
rect 340987 620914 341088 620970
rect 340987 620880 341020 620914
rect 341054 620880 341088 620914
rect 340987 620824 341088 620880
rect 340987 620790 341020 620824
rect 341054 620790 341088 620824
rect 340987 620734 341088 620790
rect 340987 620700 341020 620734
rect 341054 620700 341088 620734
rect 340987 620644 341088 620700
rect 340987 620610 341020 620644
rect 341054 620610 341088 620644
rect 340987 620554 341088 620610
rect 340987 620520 341020 620554
rect 341054 620520 341088 620554
rect 340987 620464 341088 620520
rect 340987 620430 341020 620464
rect 341054 620430 341088 620464
rect 340987 620374 341088 620430
rect 340987 620340 341020 620374
rect 341054 620340 341088 620374
rect 340987 620284 341088 620340
rect 340987 620250 341020 620284
rect 341054 620250 341088 620284
rect 340987 620194 341088 620250
rect 339699 620113 339901 620160
rect 340987 620160 341020 620194
rect 341054 620160 341088 620194
rect 340987 620113 341088 620160
rect 334648 620104 341088 620113
rect 334648 620070 334681 620104
rect 334715 620081 335868 620104
rect 334715 620070 334782 620081
rect 334648 620047 334782 620070
rect 334816 620047 334872 620081
rect 334906 620047 334962 620081
rect 334996 620047 335052 620081
rect 335086 620047 335142 620081
rect 335176 620047 335232 620081
rect 335266 620047 335322 620081
rect 335356 620047 335412 620081
rect 335446 620047 335502 620081
rect 335536 620047 335592 620081
rect 335626 620047 335682 620081
rect 335716 620047 335772 620081
rect 335806 620070 335868 620081
rect 335902 620070 335969 620104
rect 336003 620081 337156 620104
rect 336003 620070 336070 620081
rect 335806 620047 336070 620070
rect 336104 620047 336160 620081
rect 336194 620047 336250 620081
rect 336284 620047 336340 620081
rect 336374 620047 336430 620081
rect 336464 620047 336520 620081
rect 336554 620047 336610 620081
rect 336644 620047 336700 620081
rect 336734 620047 336790 620081
rect 336824 620047 336880 620081
rect 336914 620047 336970 620081
rect 337004 620047 337060 620081
rect 337094 620070 337156 620081
rect 337190 620070 337257 620104
rect 337291 620081 338444 620104
rect 337291 620070 337358 620081
rect 337094 620047 337358 620070
rect 337392 620047 337448 620081
rect 337482 620047 337538 620081
rect 337572 620047 337628 620081
rect 337662 620047 337718 620081
rect 337752 620047 337808 620081
rect 337842 620047 337898 620081
rect 337932 620047 337988 620081
rect 338022 620047 338078 620081
rect 338112 620047 338168 620081
rect 338202 620047 338258 620081
rect 338292 620047 338348 620081
rect 338382 620070 338444 620081
rect 338478 620070 338545 620104
rect 338579 620081 339732 620104
rect 338579 620070 338646 620081
rect 338382 620047 338646 620070
rect 338680 620047 338736 620081
rect 338770 620047 338826 620081
rect 338860 620047 338916 620081
rect 338950 620047 339006 620081
rect 339040 620047 339096 620081
rect 339130 620047 339186 620081
rect 339220 620047 339276 620081
rect 339310 620047 339366 620081
rect 339400 620047 339456 620081
rect 339490 620047 339546 620081
rect 339580 620047 339636 620081
rect 339670 620070 339732 620081
rect 339766 620070 339833 620104
rect 339867 620081 341020 620104
rect 339867 620070 339934 620081
rect 339670 620047 339934 620070
rect 339968 620047 340024 620081
rect 340058 620047 340114 620081
rect 340148 620047 340204 620081
rect 340238 620047 340294 620081
rect 340328 620047 340384 620081
rect 340418 620047 340474 620081
rect 340508 620047 340564 620081
rect 340598 620047 340654 620081
rect 340688 620047 340744 620081
rect 340778 620047 340834 620081
rect 340868 620047 340924 620081
rect 340958 620070 341020 620081
rect 341054 620070 341088 620104
rect 340958 620047 341088 620070
rect 334648 619980 341088 620047
rect 334648 619946 334782 619980
rect 334816 619946 334872 619980
rect 334906 619946 334962 619980
rect 334996 619946 335052 619980
rect 335086 619946 335142 619980
rect 335176 619946 335232 619980
rect 335266 619946 335322 619980
rect 335356 619946 335412 619980
rect 335446 619946 335502 619980
rect 335536 619946 335592 619980
rect 335626 619946 335682 619980
rect 335716 619946 335772 619980
rect 335806 619946 336070 619980
rect 336104 619946 336160 619980
rect 336194 619946 336250 619980
rect 336284 619946 336340 619980
rect 336374 619946 336430 619980
rect 336464 619946 336520 619980
rect 336554 619946 336610 619980
rect 336644 619946 336700 619980
rect 336734 619946 336790 619980
rect 336824 619946 336880 619980
rect 336914 619946 336970 619980
rect 337004 619946 337060 619980
rect 337094 619946 337358 619980
rect 337392 619946 337448 619980
rect 337482 619946 337538 619980
rect 337572 619946 337628 619980
rect 337662 619946 337718 619980
rect 337752 619946 337808 619980
rect 337842 619946 337898 619980
rect 337932 619946 337988 619980
rect 338022 619946 338078 619980
rect 338112 619946 338168 619980
rect 338202 619946 338258 619980
rect 338292 619946 338348 619980
rect 338382 619946 338646 619980
rect 338680 619946 338736 619980
rect 338770 619946 338826 619980
rect 338860 619946 338916 619980
rect 338950 619946 339006 619980
rect 339040 619946 339096 619980
rect 339130 619946 339186 619980
rect 339220 619946 339276 619980
rect 339310 619946 339366 619980
rect 339400 619946 339456 619980
rect 339490 619946 339546 619980
rect 339580 619946 339636 619980
rect 339670 619946 339934 619980
rect 339968 619946 340024 619980
rect 340058 619946 340114 619980
rect 340148 619946 340204 619980
rect 340238 619946 340294 619980
rect 340328 619946 340384 619980
rect 340418 619946 340474 619980
rect 340508 619946 340564 619980
rect 340598 619946 340654 619980
rect 340688 619946 340744 619980
rect 340778 619946 340834 619980
rect 340868 619946 340924 619980
rect 340958 619946 341088 619980
rect 334648 619911 341088 619946
rect 334648 619896 334749 619911
rect 334648 619862 334681 619896
rect 334715 619862 334749 619896
rect 334648 619806 334749 619862
rect 335835 619896 336037 619911
rect 335835 619862 335868 619896
rect 335902 619862 335969 619896
rect 336003 619862 336037 619896
rect 334648 619772 334681 619806
rect 334715 619772 334749 619806
rect 334648 619716 334749 619772
rect 334648 619682 334681 619716
rect 334715 619682 334749 619716
rect 334648 619626 334749 619682
rect 334648 619592 334681 619626
rect 334715 619592 334749 619626
rect 334648 619536 334749 619592
rect 334648 619502 334681 619536
rect 334715 619502 334749 619536
rect 334648 619446 334749 619502
rect 334648 619412 334681 619446
rect 334715 619412 334749 619446
rect 334648 619356 334749 619412
rect 334648 619322 334681 619356
rect 334715 619322 334749 619356
rect 334648 619266 334749 619322
rect 334648 619232 334681 619266
rect 334715 619232 334749 619266
rect 334648 619176 334749 619232
rect 334648 619142 334681 619176
rect 334715 619142 334749 619176
rect 334648 619086 334749 619142
rect 334648 619052 334681 619086
rect 334715 619052 334749 619086
rect 334648 618996 334749 619052
rect 334648 618962 334681 618996
rect 334715 618962 334749 618996
rect 334648 618906 334749 618962
rect 334648 618872 334681 618906
rect 334715 618872 334749 618906
rect 335835 619806 336037 619862
rect 337123 619896 337325 619911
rect 337123 619862 337156 619896
rect 337190 619862 337257 619896
rect 337291 619862 337325 619896
rect 335835 619772 335868 619806
rect 335902 619772 335969 619806
rect 336003 619772 336037 619806
rect 335835 619716 336037 619772
rect 335835 619682 335868 619716
rect 335902 619682 335969 619716
rect 336003 619682 336037 619716
rect 335835 619626 336037 619682
rect 335835 619592 335868 619626
rect 335902 619592 335969 619626
rect 336003 619592 336037 619626
rect 335835 619536 336037 619592
rect 335835 619502 335868 619536
rect 335902 619502 335969 619536
rect 336003 619502 336037 619536
rect 335835 619446 336037 619502
rect 335835 619412 335868 619446
rect 335902 619412 335969 619446
rect 336003 619412 336037 619446
rect 335835 619356 336037 619412
rect 335835 619322 335868 619356
rect 335902 619322 335969 619356
rect 336003 619322 336037 619356
rect 335835 619266 336037 619322
rect 335835 619232 335868 619266
rect 335902 619232 335969 619266
rect 336003 619232 336037 619266
rect 335835 619176 336037 619232
rect 335835 619142 335868 619176
rect 335902 619142 335969 619176
rect 336003 619142 336037 619176
rect 335835 619086 336037 619142
rect 335835 619052 335868 619086
rect 335902 619052 335969 619086
rect 336003 619052 336037 619086
rect 335835 618996 336037 619052
rect 335835 618962 335868 618996
rect 335902 618962 335969 618996
rect 336003 618962 336037 618996
rect 335835 618906 336037 618962
rect 334648 618825 334749 618872
rect 335835 618872 335868 618906
rect 335902 618872 335969 618906
rect 336003 618872 336037 618906
rect 337123 619806 337325 619862
rect 338411 619896 338613 619911
rect 338411 619862 338444 619896
rect 338478 619862 338545 619896
rect 338579 619862 338613 619896
rect 337123 619772 337156 619806
rect 337190 619772 337257 619806
rect 337291 619772 337325 619806
rect 337123 619716 337325 619772
rect 337123 619682 337156 619716
rect 337190 619682 337257 619716
rect 337291 619682 337325 619716
rect 337123 619626 337325 619682
rect 337123 619592 337156 619626
rect 337190 619592 337257 619626
rect 337291 619592 337325 619626
rect 337123 619536 337325 619592
rect 337123 619502 337156 619536
rect 337190 619502 337257 619536
rect 337291 619502 337325 619536
rect 337123 619446 337325 619502
rect 337123 619412 337156 619446
rect 337190 619412 337257 619446
rect 337291 619412 337325 619446
rect 337123 619356 337325 619412
rect 337123 619322 337156 619356
rect 337190 619322 337257 619356
rect 337291 619322 337325 619356
rect 337123 619266 337325 619322
rect 337123 619232 337156 619266
rect 337190 619232 337257 619266
rect 337291 619232 337325 619266
rect 337123 619176 337325 619232
rect 337123 619142 337156 619176
rect 337190 619142 337257 619176
rect 337291 619142 337325 619176
rect 337123 619086 337325 619142
rect 337123 619052 337156 619086
rect 337190 619052 337257 619086
rect 337291 619052 337325 619086
rect 337123 618996 337325 619052
rect 337123 618962 337156 618996
rect 337190 618962 337257 618996
rect 337291 618962 337325 618996
rect 337123 618906 337325 618962
rect 335835 618825 336037 618872
rect 337123 618872 337156 618906
rect 337190 618872 337257 618906
rect 337291 618872 337325 618906
rect 338411 619806 338613 619862
rect 339699 619896 339901 619911
rect 339699 619862 339732 619896
rect 339766 619862 339833 619896
rect 339867 619862 339901 619896
rect 338411 619772 338444 619806
rect 338478 619772 338545 619806
rect 338579 619772 338613 619806
rect 338411 619716 338613 619772
rect 338411 619682 338444 619716
rect 338478 619682 338545 619716
rect 338579 619682 338613 619716
rect 338411 619626 338613 619682
rect 338411 619592 338444 619626
rect 338478 619592 338545 619626
rect 338579 619592 338613 619626
rect 338411 619536 338613 619592
rect 338411 619502 338444 619536
rect 338478 619502 338545 619536
rect 338579 619502 338613 619536
rect 338411 619446 338613 619502
rect 338411 619412 338444 619446
rect 338478 619412 338545 619446
rect 338579 619412 338613 619446
rect 338411 619356 338613 619412
rect 338411 619322 338444 619356
rect 338478 619322 338545 619356
rect 338579 619322 338613 619356
rect 338411 619266 338613 619322
rect 338411 619232 338444 619266
rect 338478 619232 338545 619266
rect 338579 619232 338613 619266
rect 338411 619176 338613 619232
rect 338411 619142 338444 619176
rect 338478 619142 338545 619176
rect 338579 619142 338613 619176
rect 338411 619086 338613 619142
rect 338411 619052 338444 619086
rect 338478 619052 338545 619086
rect 338579 619052 338613 619086
rect 338411 618996 338613 619052
rect 338411 618962 338444 618996
rect 338478 618962 338545 618996
rect 338579 618962 338613 618996
rect 338411 618906 338613 618962
rect 337123 618825 337325 618872
rect 338411 618872 338444 618906
rect 338478 618872 338545 618906
rect 338579 618872 338613 618906
rect 339699 619806 339901 619862
rect 340987 619896 341088 619911
rect 340987 619862 341020 619896
rect 341054 619862 341088 619896
rect 339699 619772 339732 619806
rect 339766 619772 339833 619806
rect 339867 619772 339901 619806
rect 339699 619716 339901 619772
rect 339699 619682 339732 619716
rect 339766 619682 339833 619716
rect 339867 619682 339901 619716
rect 339699 619626 339901 619682
rect 339699 619592 339732 619626
rect 339766 619592 339833 619626
rect 339867 619592 339901 619626
rect 339699 619536 339901 619592
rect 339699 619502 339732 619536
rect 339766 619502 339833 619536
rect 339867 619502 339901 619536
rect 339699 619446 339901 619502
rect 339699 619412 339732 619446
rect 339766 619412 339833 619446
rect 339867 619412 339901 619446
rect 339699 619356 339901 619412
rect 339699 619322 339732 619356
rect 339766 619322 339833 619356
rect 339867 619322 339901 619356
rect 339699 619266 339901 619322
rect 339699 619232 339732 619266
rect 339766 619232 339833 619266
rect 339867 619232 339901 619266
rect 339699 619176 339901 619232
rect 339699 619142 339732 619176
rect 339766 619142 339833 619176
rect 339867 619142 339901 619176
rect 339699 619086 339901 619142
rect 339699 619052 339732 619086
rect 339766 619052 339833 619086
rect 339867 619052 339901 619086
rect 339699 618996 339901 619052
rect 339699 618962 339732 618996
rect 339766 618962 339833 618996
rect 339867 618962 339901 618996
rect 339699 618906 339901 618962
rect 338411 618825 338613 618872
rect 339699 618872 339732 618906
rect 339766 618872 339833 618906
rect 339867 618872 339901 618906
rect 340987 619806 341088 619862
rect 340987 619772 341020 619806
rect 341054 619772 341088 619806
rect 340987 619716 341088 619772
rect 340987 619682 341020 619716
rect 341054 619682 341088 619716
rect 340987 619626 341088 619682
rect 340987 619592 341020 619626
rect 341054 619592 341088 619626
rect 340987 619536 341088 619592
rect 340987 619502 341020 619536
rect 341054 619502 341088 619536
rect 340987 619446 341088 619502
rect 340987 619412 341020 619446
rect 341054 619412 341088 619446
rect 340987 619356 341088 619412
rect 340987 619322 341020 619356
rect 341054 619322 341088 619356
rect 340987 619266 341088 619322
rect 340987 619232 341020 619266
rect 341054 619232 341088 619266
rect 340987 619176 341088 619232
rect 340987 619142 341020 619176
rect 341054 619142 341088 619176
rect 340987 619086 341088 619142
rect 340987 619052 341020 619086
rect 341054 619052 341088 619086
rect 340987 618996 341088 619052
rect 340987 618962 341020 618996
rect 341054 618962 341088 618996
rect 340987 618906 341088 618962
rect 339699 618825 339901 618872
rect 340987 618872 341020 618906
rect 341054 618872 341088 618906
rect 340987 618825 341088 618872
rect 334648 618816 341088 618825
rect 334648 618782 334681 618816
rect 334715 618793 335868 618816
rect 334715 618782 334782 618793
rect 334648 618759 334782 618782
rect 334816 618759 334872 618793
rect 334906 618759 334962 618793
rect 334996 618759 335052 618793
rect 335086 618759 335142 618793
rect 335176 618759 335232 618793
rect 335266 618759 335322 618793
rect 335356 618759 335412 618793
rect 335446 618759 335502 618793
rect 335536 618759 335592 618793
rect 335626 618759 335682 618793
rect 335716 618759 335772 618793
rect 335806 618782 335868 618793
rect 335902 618782 335969 618816
rect 336003 618793 337156 618816
rect 336003 618782 336070 618793
rect 335806 618759 336070 618782
rect 336104 618759 336160 618793
rect 336194 618759 336250 618793
rect 336284 618759 336340 618793
rect 336374 618759 336430 618793
rect 336464 618759 336520 618793
rect 336554 618759 336610 618793
rect 336644 618759 336700 618793
rect 336734 618759 336790 618793
rect 336824 618759 336880 618793
rect 336914 618759 336970 618793
rect 337004 618759 337060 618793
rect 337094 618782 337156 618793
rect 337190 618782 337257 618816
rect 337291 618793 338444 618816
rect 337291 618782 337358 618793
rect 337094 618759 337358 618782
rect 337392 618759 337448 618793
rect 337482 618759 337538 618793
rect 337572 618759 337628 618793
rect 337662 618759 337718 618793
rect 337752 618759 337808 618793
rect 337842 618759 337898 618793
rect 337932 618759 337988 618793
rect 338022 618759 338078 618793
rect 338112 618759 338168 618793
rect 338202 618759 338258 618793
rect 338292 618759 338348 618793
rect 338382 618782 338444 618793
rect 338478 618782 338545 618816
rect 338579 618793 339732 618816
rect 338579 618782 338646 618793
rect 338382 618759 338646 618782
rect 338680 618759 338736 618793
rect 338770 618759 338826 618793
rect 338860 618759 338916 618793
rect 338950 618759 339006 618793
rect 339040 618759 339096 618793
rect 339130 618759 339186 618793
rect 339220 618759 339276 618793
rect 339310 618759 339366 618793
rect 339400 618759 339456 618793
rect 339490 618759 339546 618793
rect 339580 618759 339636 618793
rect 339670 618782 339732 618793
rect 339766 618782 339833 618816
rect 339867 618793 341020 618816
rect 339867 618782 339934 618793
rect 339670 618759 339934 618782
rect 339968 618759 340024 618793
rect 340058 618759 340114 618793
rect 340148 618759 340204 618793
rect 340238 618759 340294 618793
rect 340328 618759 340384 618793
rect 340418 618759 340474 618793
rect 340508 618759 340564 618793
rect 340598 618759 340654 618793
rect 340688 618759 340744 618793
rect 340778 618759 340834 618793
rect 340868 618759 340924 618793
rect 340958 618782 341020 618793
rect 341054 618782 341088 618816
rect 340958 618759 341088 618782
rect 334648 618692 341088 618759
rect 334648 618658 334782 618692
rect 334816 618658 334872 618692
rect 334906 618658 334962 618692
rect 334996 618658 335052 618692
rect 335086 618658 335142 618692
rect 335176 618658 335232 618692
rect 335266 618658 335322 618692
rect 335356 618658 335412 618692
rect 335446 618658 335502 618692
rect 335536 618658 335592 618692
rect 335626 618658 335682 618692
rect 335716 618658 335772 618692
rect 335806 618658 336070 618692
rect 336104 618658 336160 618692
rect 336194 618658 336250 618692
rect 336284 618658 336340 618692
rect 336374 618658 336430 618692
rect 336464 618658 336520 618692
rect 336554 618658 336610 618692
rect 336644 618658 336700 618692
rect 336734 618658 336790 618692
rect 336824 618658 336880 618692
rect 336914 618658 336970 618692
rect 337004 618658 337060 618692
rect 337094 618658 337358 618692
rect 337392 618658 337448 618692
rect 337482 618658 337538 618692
rect 337572 618658 337628 618692
rect 337662 618658 337718 618692
rect 337752 618658 337808 618692
rect 337842 618658 337898 618692
rect 337932 618658 337988 618692
rect 338022 618658 338078 618692
rect 338112 618658 338168 618692
rect 338202 618658 338258 618692
rect 338292 618658 338348 618692
rect 338382 618658 338646 618692
rect 338680 618658 338736 618692
rect 338770 618658 338826 618692
rect 338860 618658 338916 618692
rect 338950 618658 339006 618692
rect 339040 618658 339096 618692
rect 339130 618658 339186 618692
rect 339220 618658 339276 618692
rect 339310 618658 339366 618692
rect 339400 618658 339456 618692
rect 339490 618658 339546 618692
rect 339580 618658 339636 618692
rect 339670 618658 339934 618692
rect 339968 618658 340024 618692
rect 340058 618658 340114 618692
rect 340148 618658 340204 618692
rect 340238 618658 340294 618692
rect 340328 618658 340384 618692
rect 340418 618658 340474 618692
rect 340508 618658 340564 618692
rect 340598 618658 340654 618692
rect 340688 618658 340744 618692
rect 340778 618658 340834 618692
rect 340868 618658 340924 618692
rect 340958 618658 341088 618692
rect 334648 618623 341088 618658
rect 334648 618608 334749 618623
rect 334648 618574 334681 618608
rect 334715 618574 334749 618608
rect 334648 618518 334749 618574
rect 335835 618608 336037 618623
rect 335835 618574 335868 618608
rect 335902 618574 335969 618608
rect 336003 618574 336037 618608
rect 334648 618484 334681 618518
rect 334715 618484 334749 618518
rect 334648 618428 334749 618484
rect 334648 618394 334681 618428
rect 334715 618394 334749 618428
rect 334648 618338 334749 618394
rect 334648 618304 334681 618338
rect 334715 618304 334749 618338
rect 334648 618248 334749 618304
rect 334648 618214 334681 618248
rect 334715 618214 334749 618248
rect 334648 618158 334749 618214
rect 334648 618124 334681 618158
rect 334715 618124 334749 618158
rect 334648 618068 334749 618124
rect 334648 618034 334681 618068
rect 334715 618034 334749 618068
rect 334648 617978 334749 618034
rect 334648 617944 334681 617978
rect 334715 617944 334749 617978
rect 334648 617888 334749 617944
rect 334648 617854 334681 617888
rect 334715 617854 334749 617888
rect 334648 617798 334749 617854
rect 334648 617764 334681 617798
rect 334715 617764 334749 617798
rect 334648 617708 334749 617764
rect 334648 617674 334681 617708
rect 334715 617674 334749 617708
rect 334648 617618 334749 617674
rect 334648 617584 334681 617618
rect 334715 617584 334749 617618
rect 335835 618518 336037 618574
rect 337123 618608 337325 618623
rect 337123 618574 337156 618608
rect 337190 618574 337257 618608
rect 337291 618574 337325 618608
rect 335835 618484 335868 618518
rect 335902 618484 335969 618518
rect 336003 618484 336037 618518
rect 335835 618428 336037 618484
rect 335835 618394 335868 618428
rect 335902 618394 335969 618428
rect 336003 618394 336037 618428
rect 335835 618338 336037 618394
rect 335835 618304 335868 618338
rect 335902 618304 335969 618338
rect 336003 618304 336037 618338
rect 335835 618248 336037 618304
rect 335835 618214 335868 618248
rect 335902 618214 335969 618248
rect 336003 618214 336037 618248
rect 335835 618158 336037 618214
rect 335835 618124 335868 618158
rect 335902 618124 335969 618158
rect 336003 618124 336037 618158
rect 335835 618068 336037 618124
rect 335835 618034 335868 618068
rect 335902 618034 335969 618068
rect 336003 618034 336037 618068
rect 335835 617978 336037 618034
rect 335835 617944 335868 617978
rect 335902 617944 335969 617978
rect 336003 617944 336037 617978
rect 335835 617888 336037 617944
rect 335835 617854 335868 617888
rect 335902 617854 335969 617888
rect 336003 617854 336037 617888
rect 335835 617798 336037 617854
rect 335835 617764 335868 617798
rect 335902 617764 335969 617798
rect 336003 617764 336037 617798
rect 335835 617708 336037 617764
rect 335835 617674 335868 617708
rect 335902 617674 335969 617708
rect 336003 617674 336037 617708
rect 335835 617618 336037 617674
rect 334648 617537 334749 617584
rect 335835 617584 335868 617618
rect 335902 617584 335969 617618
rect 336003 617584 336037 617618
rect 337123 618518 337325 618574
rect 338411 618608 338613 618623
rect 338411 618574 338444 618608
rect 338478 618574 338545 618608
rect 338579 618574 338613 618608
rect 337123 618484 337156 618518
rect 337190 618484 337257 618518
rect 337291 618484 337325 618518
rect 337123 618428 337325 618484
rect 337123 618394 337156 618428
rect 337190 618394 337257 618428
rect 337291 618394 337325 618428
rect 337123 618338 337325 618394
rect 337123 618304 337156 618338
rect 337190 618304 337257 618338
rect 337291 618304 337325 618338
rect 337123 618248 337325 618304
rect 337123 618214 337156 618248
rect 337190 618214 337257 618248
rect 337291 618214 337325 618248
rect 337123 618158 337325 618214
rect 337123 618124 337156 618158
rect 337190 618124 337257 618158
rect 337291 618124 337325 618158
rect 337123 618068 337325 618124
rect 337123 618034 337156 618068
rect 337190 618034 337257 618068
rect 337291 618034 337325 618068
rect 337123 617978 337325 618034
rect 337123 617944 337156 617978
rect 337190 617944 337257 617978
rect 337291 617944 337325 617978
rect 337123 617888 337325 617944
rect 337123 617854 337156 617888
rect 337190 617854 337257 617888
rect 337291 617854 337325 617888
rect 337123 617798 337325 617854
rect 337123 617764 337156 617798
rect 337190 617764 337257 617798
rect 337291 617764 337325 617798
rect 337123 617708 337325 617764
rect 337123 617674 337156 617708
rect 337190 617674 337257 617708
rect 337291 617674 337325 617708
rect 337123 617618 337325 617674
rect 335835 617537 336037 617584
rect 337123 617584 337156 617618
rect 337190 617584 337257 617618
rect 337291 617584 337325 617618
rect 338411 618518 338613 618574
rect 339699 618608 339901 618623
rect 339699 618574 339732 618608
rect 339766 618574 339833 618608
rect 339867 618574 339901 618608
rect 338411 618484 338444 618518
rect 338478 618484 338545 618518
rect 338579 618484 338613 618518
rect 338411 618428 338613 618484
rect 338411 618394 338444 618428
rect 338478 618394 338545 618428
rect 338579 618394 338613 618428
rect 338411 618338 338613 618394
rect 338411 618304 338444 618338
rect 338478 618304 338545 618338
rect 338579 618304 338613 618338
rect 338411 618248 338613 618304
rect 338411 618214 338444 618248
rect 338478 618214 338545 618248
rect 338579 618214 338613 618248
rect 338411 618158 338613 618214
rect 338411 618124 338444 618158
rect 338478 618124 338545 618158
rect 338579 618124 338613 618158
rect 338411 618068 338613 618124
rect 338411 618034 338444 618068
rect 338478 618034 338545 618068
rect 338579 618034 338613 618068
rect 338411 617978 338613 618034
rect 338411 617944 338444 617978
rect 338478 617944 338545 617978
rect 338579 617944 338613 617978
rect 338411 617888 338613 617944
rect 338411 617854 338444 617888
rect 338478 617854 338545 617888
rect 338579 617854 338613 617888
rect 338411 617798 338613 617854
rect 338411 617764 338444 617798
rect 338478 617764 338545 617798
rect 338579 617764 338613 617798
rect 338411 617708 338613 617764
rect 338411 617674 338444 617708
rect 338478 617674 338545 617708
rect 338579 617674 338613 617708
rect 338411 617618 338613 617674
rect 337123 617537 337325 617584
rect 338411 617584 338444 617618
rect 338478 617584 338545 617618
rect 338579 617584 338613 617618
rect 339699 618518 339901 618574
rect 340987 618608 341088 618623
rect 340987 618574 341020 618608
rect 341054 618574 341088 618608
rect 339699 618484 339732 618518
rect 339766 618484 339833 618518
rect 339867 618484 339901 618518
rect 339699 618428 339901 618484
rect 339699 618394 339732 618428
rect 339766 618394 339833 618428
rect 339867 618394 339901 618428
rect 339699 618338 339901 618394
rect 339699 618304 339732 618338
rect 339766 618304 339833 618338
rect 339867 618304 339901 618338
rect 339699 618248 339901 618304
rect 339699 618214 339732 618248
rect 339766 618214 339833 618248
rect 339867 618214 339901 618248
rect 339699 618158 339901 618214
rect 339699 618124 339732 618158
rect 339766 618124 339833 618158
rect 339867 618124 339901 618158
rect 339699 618068 339901 618124
rect 339699 618034 339732 618068
rect 339766 618034 339833 618068
rect 339867 618034 339901 618068
rect 339699 617978 339901 618034
rect 339699 617944 339732 617978
rect 339766 617944 339833 617978
rect 339867 617944 339901 617978
rect 339699 617888 339901 617944
rect 339699 617854 339732 617888
rect 339766 617854 339833 617888
rect 339867 617854 339901 617888
rect 339699 617798 339901 617854
rect 339699 617764 339732 617798
rect 339766 617764 339833 617798
rect 339867 617764 339901 617798
rect 339699 617708 339901 617764
rect 339699 617674 339732 617708
rect 339766 617674 339833 617708
rect 339867 617674 339901 617708
rect 339699 617618 339901 617674
rect 338411 617537 338613 617584
rect 339699 617584 339732 617618
rect 339766 617584 339833 617618
rect 339867 617584 339901 617618
rect 340987 618518 341088 618574
rect 340987 618484 341020 618518
rect 341054 618484 341088 618518
rect 340987 618428 341088 618484
rect 340987 618394 341020 618428
rect 341054 618394 341088 618428
rect 340987 618338 341088 618394
rect 340987 618304 341020 618338
rect 341054 618304 341088 618338
rect 340987 618248 341088 618304
rect 340987 618214 341020 618248
rect 341054 618214 341088 618248
rect 340987 618158 341088 618214
rect 340987 618124 341020 618158
rect 341054 618124 341088 618158
rect 340987 618068 341088 618124
rect 340987 618034 341020 618068
rect 341054 618034 341088 618068
rect 340987 617978 341088 618034
rect 340987 617944 341020 617978
rect 341054 617944 341088 617978
rect 340987 617888 341088 617944
rect 340987 617854 341020 617888
rect 341054 617854 341088 617888
rect 340987 617798 341088 617854
rect 340987 617764 341020 617798
rect 341054 617764 341088 617798
rect 340987 617708 341088 617764
rect 340987 617674 341020 617708
rect 341054 617674 341088 617708
rect 340987 617618 341088 617674
rect 339699 617537 339901 617584
rect 340987 617584 341020 617618
rect 341054 617584 341088 617618
rect 340987 617537 341088 617584
rect 334648 617528 341088 617537
rect 334648 617494 334681 617528
rect 334715 617505 335868 617528
rect 334715 617494 334782 617505
rect 334648 617471 334782 617494
rect 334816 617471 334872 617505
rect 334906 617471 334962 617505
rect 334996 617471 335052 617505
rect 335086 617471 335142 617505
rect 335176 617471 335232 617505
rect 335266 617471 335322 617505
rect 335356 617471 335412 617505
rect 335446 617471 335502 617505
rect 335536 617471 335592 617505
rect 335626 617471 335682 617505
rect 335716 617471 335772 617505
rect 335806 617494 335868 617505
rect 335902 617494 335969 617528
rect 336003 617505 337156 617528
rect 336003 617494 336070 617505
rect 335806 617471 336070 617494
rect 336104 617471 336160 617505
rect 336194 617471 336250 617505
rect 336284 617471 336340 617505
rect 336374 617471 336430 617505
rect 336464 617471 336520 617505
rect 336554 617471 336610 617505
rect 336644 617471 336700 617505
rect 336734 617471 336790 617505
rect 336824 617471 336880 617505
rect 336914 617471 336970 617505
rect 337004 617471 337060 617505
rect 337094 617494 337156 617505
rect 337190 617494 337257 617528
rect 337291 617505 338444 617528
rect 337291 617494 337358 617505
rect 337094 617471 337358 617494
rect 337392 617471 337448 617505
rect 337482 617471 337538 617505
rect 337572 617471 337628 617505
rect 337662 617471 337718 617505
rect 337752 617471 337808 617505
rect 337842 617471 337898 617505
rect 337932 617471 337988 617505
rect 338022 617471 338078 617505
rect 338112 617471 338168 617505
rect 338202 617471 338258 617505
rect 338292 617471 338348 617505
rect 338382 617494 338444 617505
rect 338478 617494 338545 617528
rect 338579 617505 339732 617528
rect 338579 617494 338646 617505
rect 338382 617471 338646 617494
rect 338680 617471 338736 617505
rect 338770 617471 338826 617505
rect 338860 617471 338916 617505
rect 338950 617471 339006 617505
rect 339040 617471 339096 617505
rect 339130 617471 339186 617505
rect 339220 617471 339276 617505
rect 339310 617471 339366 617505
rect 339400 617471 339456 617505
rect 339490 617471 339546 617505
rect 339580 617471 339636 617505
rect 339670 617494 339732 617505
rect 339766 617494 339833 617528
rect 339867 617505 341020 617528
rect 339867 617494 339934 617505
rect 339670 617471 339934 617494
rect 339968 617471 340024 617505
rect 340058 617471 340114 617505
rect 340148 617471 340204 617505
rect 340238 617471 340294 617505
rect 340328 617471 340384 617505
rect 340418 617471 340474 617505
rect 340508 617471 340564 617505
rect 340598 617471 340654 617505
rect 340688 617471 340744 617505
rect 340778 617471 340834 617505
rect 340868 617471 340924 617505
rect 340958 617494 341020 617505
rect 341054 617494 341088 617528
rect 340958 617471 341088 617494
rect 334648 617436 341088 617471
rect 297848 616448 298896 616472
rect 297824 615448 341112 615472
rect 297824 614448 297848 615448
rect 341088 614448 341112 615448
rect 297824 614424 341112 614448
rect 342088 614424 342112 640648
rect 343112 614424 343136 640648
rect 342088 614400 343136 614424
<< nsubdiff >>
rect 334811 627558 335773 627577
rect 334811 627524 334922 627558
rect 334956 627524 335012 627558
rect 335046 627524 335102 627558
rect 335136 627524 335192 627558
rect 335226 627524 335282 627558
rect 335316 627524 335372 627558
rect 335406 627524 335462 627558
rect 335496 627524 335552 627558
rect 335586 627524 335642 627558
rect 335676 627524 335773 627558
rect 334811 627505 335773 627524
rect 334811 627464 334883 627505
rect 334811 627430 334830 627464
rect 334864 627430 334883 627464
rect 335701 627445 335773 627505
rect 334811 627374 334883 627430
rect 334811 627340 334830 627374
rect 334864 627340 334883 627374
rect 334811 627284 334883 627340
rect 334811 627250 334830 627284
rect 334864 627250 334883 627284
rect 334811 627194 334883 627250
rect 334811 627160 334830 627194
rect 334864 627160 334883 627194
rect 334811 627104 334883 627160
rect 334811 627070 334830 627104
rect 334864 627070 334883 627104
rect 334811 627014 334883 627070
rect 334811 626980 334830 627014
rect 334864 626980 334883 627014
rect 334811 626924 334883 626980
rect 334811 626890 334830 626924
rect 334864 626890 334883 626924
rect 334811 626834 334883 626890
rect 334811 626800 334830 626834
rect 334864 626800 334883 626834
rect 334811 626744 334883 626800
rect 335701 627411 335720 627445
rect 335754 627411 335773 627445
rect 335701 627355 335773 627411
rect 335701 627321 335720 627355
rect 335754 627321 335773 627355
rect 335701 627265 335773 627321
rect 335701 627231 335720 627265
rect 335754 627231 335773 627265
rect 335701 627175 335773 627231
rect 335701 627141 335720 627175
rect 335754 627141 335773 627175
rect 335701 627085 335773 627141
rect 335701 627051 335720 627085
rect 335754 627051 335773 627085
rect 335701 626995 335773 627051
rect 335701 626961 335720 626995
rect 335754 626961 335773 626995
rect 335701 626905 335773 626961
rect 335701 626871 335720 626905
rect 335754 626871 335773 626905
rect 335701 626815 335773 626871
rect 335701 626781 335720 626815
rect 335754 626781 335773 626815
rect 334811 626710 334830 626744
rect 334864 626710 334883 626744
rect 334811 626687 334883 626710
rect 335701 626725 335773 626781
rect 335701 626691 335720 626725
rect 335754 626691 335773 626725
rect 335701 626687 335773 626691
rect 334811 626668 335773 626687
rect 334811 626634 334888 626668
rect 334922 626634 334978 626668
rect 335012 626634 335068 626668
rect 335102 626634 335158 626668
rect 335192 626634 335248 626668
rect 335282 626634 335338 626668
rect 335372 626634 335428 626668
rect 335462 626634 335518 626668
rect 335552 626634 335608 626668
rect 335642 626634 335773 626668
rect 334811 626615 335773 626634
rect 336099 627558 337061 627577
rect 336099 627524 336210 627558
rect 336244 627524 336300 627558
rect 336334 627524 336390 627558
rect 336424 627524 336480 627558
rect 336514 627524 336570 627558
rect 336604 627524 336660 627558
rect 336694 627524 336750 627558
rect 336784 627524 336840 627558
rect 336874 627524 336930 627558
rect 336964 627524 337061 627558
rect 336099 627505 337061 627524
rect 336099 627464 336171 627505
rect 336099 627430 336118 627464
rect 336152 627430 336171 627464
rect 336989 627445 337061 627505
rect 336099 627374 336171 627430
rect 336099 627340 336118 627374
rect 336152 627340 336171 627374
rect 336099 627284 336171 627340
rect 336099 627250 336118 627284
rect 336152 627250 336171 627284
rect 336099 627194 336171 627250
rect 336099 627160 336118 627194
rect 336152 627160 336171 627194
rect 336099 627104 336171 627160
rect 336099 627070 336118 627104
rect 336152 627070 336171 627104
rect 336099 627014 336171 627070
rect 336099 626980 336118 627014
rect 336152 626980 336171 627014
rect 336099 626924 336171 626980
rect 336099 626890 336118 626924
rect 336152 626890 336171 626924
rect 336099 626834 336171 626890
rect 336099 626800 336118 626834
rect 336152 626800 336171 626834
rect 336099 626744 336171 626800
rect 336989 627411 337008 627445
rect 337042 627411 337061 627445
rect 336989 627355 337061 627411
rect 336989 627321 337008 627355
rect 337042 627321 337061 627355
rect 336989 627265 337061 627321
rect 336989 627231 337008 627265
rect 337042 627231 337061 627265
rect 336989 627175 337061 627231
rect 336989 627141 337008 627175
rect 337042 627141 337061 627175
rect 336989 627085 337061 627141
rect 336989 627051 337008 627085
rect 337042 627051 337061 627085
rect 336989 626995 337061 627051
rect 336989 626961 337008 626995
rect 337042 626961 337061 626995
rect 336989 626905 337061 626961
rect 336989 626871 337008 626905
rect 337042 626871 337061 626905
rect 336989 626815 337061 626871
rect 336989 626781 337008 626815
rect 337042 626781 337061 626815
rect 336099 626710 336118 626744
rect 336152 626710 336171 626744
rect 336099 626687 336171 626710
rect 336989 626725 337061 626781
rect 336989 626691 337008 626725
rect 337042 626691 337061 626725
rect 336989 626687 337061 626691
rect 336099 626668 337061 626687
rect 336099 626634 336176 626668
rect 336210 626634 336266 626668
rect 336300 626634 336356 626668
rect 336390 626634 336446 626668
rect 336480 626634 336536 626668
rect 336570 626634 336626 626668
rect 336660 626634 336716 626668
rect 336750 626634 336806 626668
rect 336840 626634 336896 626668
rect 336930 626634 337061 626668
rect 336099 626615 337061 626634
rect 337387 627558 338349 627577
rect 337387 627524 337498 627558
rect 337532 627524 337588 627558
rect 337622 627524 337678 627558
rect 337712 627524 337768 627558
rect 337802 627524 337858 627558
rect 337892 627524 337948 627558
rect 337982 627524 338038 627558
rect 338072 627524 338128 627558
rect 338162 627524 338218 627558
rect 338252 627524 338349 627558
rect 337387 627505 338349 627524
rect 337387 627464 337459 627505
rect 337387 627430 337406 627464
rect 337440 627430 337459 627464
rect 338277 627445 338349 627505
rect 337387 627374 337459 627430
rect 337387 627340 337406 627374
rect 337440 627340 337459 627374
rect 337387 627284 337459 627340
rect 337387 627250 337406 627284
rect 337440 627250 337459 627284
rect 337387 627194 337459 627250
rect 337387 627160 337406 627194
rect 337440 627160 337459 627194
rect 337387 627104 337459 627160
rect 337387 627070 337406 627104
rect 337440 627070 337459 627104
rect 337387 627014 337459 627070
rect 337387 626980 337406 627014
rect 337440 626980 337459 627014
rect 337387 626924 337459 626980
rect 337387 626890 337406 626924
rect 337440 626890 337459 626924
rect 337387 626834 337459 626890
rect 337387 626800 337406 626834
rect 337440 626800 337459 626834
rect 337387 626744 337459 626800
rect 338277 627411 338296 627445
rect 338330 627411 338349 627445
rect 338277 627355 338349 627411
rect 338277 627321 338296 627355
rect 338330 627321 338349 627355
rect 338277 627265 338349 627321
rect 338277 627231 338296 627265
rect 338330 627231 338349 627265
rect 338277 627175 338349 627231
rect 338277 627141 338296 627175
rect 338330 627141 338349 627175
rect 338277 627085 338349 627141
rect 338277 627051 338296 627085
rect 338330 627051 338349 627085
rect 338277 626995 338349 627051
rect 338277 626961 338296 626995
rect 338330 626961 338349 626995
rect 338277 626905 338349 626961
rect 338277 626871 338296 626905
rect 338330 626871 338349 626905
rect 338277 626815 338349 626871
rect 338277 626781 338296 626815
rect 338330 626781 338349 626815
rect 337387 626710 337406 626744
rect 337440 626710 337459 626744
rect 337387 626687 337459 626710
rect 338277 626725 338349 626781
rect 338277 626691 338296 626725
rect 338330 626691 338349 626725
rect 338277 626687 338349 626691
rect 337387 626668 338349 626687
rect 337387 626634 337464 626668
rect 337498 626634 337554 626668
rect 337588 626634 337644 626668
rect 337678 626634 337734 626668
rect 337768 626634 337824 626668
rect 337858 626634 337914 626668
rect 337948 626634 338004 626668
rect 338038 626634 338094 626668
rect 338128 626634 338184 626668
rect 338218 626634 338349 626668
rect 337387 626615 338349 626634
rect 338675 627558 339637 627577
rect 338675 627524 338786 627558
rect 338820 627524 338876 627558
rect 338910 627524 338966 627558
rect 339000 627524 339056 627558
rect 339090 627524 339146 627558
rect 339180 627524 339236 627558
rect 339270 627524 339326 627558
rect 339360 627524 339416 627558
rect 339450 627524 339506 627558
rect 339540 627524 339637 627558
rect 338675 627505 339637 627524
rect 338675 627464 338747 627505
rect 338675 627430 338694 627464
rect 338728 627430 338747 627464
rect 339565 627445 339637 627505
rect 338675 627374 338747 627430
rect 338675 627340 338694 627374
rect 338728 627340 338747 627374
rect 338675 627284 338747 627340
rect 338675 627250 338694 627284
rect 338728 627250 338747 627284
rect 338675 627194 338747 627250
rect 338675 627160 338694 627194
rect 338728 627160 338747 627194
rect 338675 627104 338747 627160
rect 338675 627070 338694 627104
rect 338728 627070 338747 627104
rect 338675 627014 338747 627070
rect 338675 626980 338694 627014
rect 338728 626980 338747 627014
rect 338675 626924 338747 626980
rect 338675 626890 338694 626924
rect 338728 626890 338747 626924
rect 338675 626834 338747 626890
rect 338675 626800 338694 626834
rect 338728 626800 338747 626834
rect 338675 626744 338747 626800
rect 339565 627411 339584 627445
rect 339618 627411 339637 627445
rect 339565 627355 339637 627411
rect 339565 627321 339584 627355
rect 339618 627321 339637 627355
rect 339565 627265 339637 627321
rect 339565 627231 339584 627265
rect 339618 627231 339637 627265
rect 339565 627175 339637 627231
rect 339565 627141 339584 627175
rect 339618 627141 339637 627175
rect 339565 627085 339637 627141
rect 339565 627051 339584 627085
rect 339618 627051 339637 627085
rect 339565 626995 339637 627051
rect 339565 626961 339584 626995
rect 339618 626961 339637 626995
rect 339565 626905 339637 626961
rect 339565 626871 339584 626905
rect 339618 626871 339637 626905
rect 339565 626815 339637 626871
rect 339565 626781 339584 626815
rect 339618 626781 339637 626815
rect 338675 626710 338694 626744
rect 338728 626710 338747 626744
rect 338675 626687 338747 626710
rect 339565 626725 339637 626781
rect 339565 626691 339584 626725
rect 339618 626691 339637 626725
rect 339565 626687 339637 626691
rect 338675 626668 339637 626687
rect 338675 626634 338752 626668
rect 338786 626634 338842 626668
rect 338876 626634 338932 626668
rect 338966 626634 339022 626668
rect 339056 626634 339112 626668
rect 339146 626634 339202 626668
rect 339236 626634 339292 626668
rect 339326 626634 339382 626668
rect 339416 626634 339472 626668
rect 339506 626634 339637 626668
rect 338675 626615 339637 626634
rect 339963 627558 340925 627577
rect 339963 627524 340074 627558
rect 340108 627524 340164 627558
rect 340198 627524 340254 627558
rect 340288 627524 340344 627558
rect 340378 627524 340434 627558
rect 340468 627524 340524 627558
rect 340558 627524 340614 627558
rect 340648 627524 340704 627558
rect 340738 627524 340794 627558
rect 340828 627524 340925 627558
rect 339963 627505 340925 627524
rect 339963 627464 340035 627505
rect 339963 627430 339982 627464
rect 340016 627430 340035 627464
rect 340853 627445 340925 627505
rect 339963 627374 340035 627430
rect 339963 627340 339982 627374
rect 340016 627340 340035 627374
rect 339963 627284 340035 627340
rect 339963 627250 339982 627284
rect 340016 627250 340035 627284
rect 339963 627194 340035 627250
rect 339963 627160 339982 627194
rect 340016 627160 340035 627194
rect 339963 627104 340035 627160
rect 339963 627070 339982 627104
rect 340016 627070 340035 627104
rect 339963 627014 340035 627070
rect 339963 626980 339982 627014
rect 340016 626980 340035 627014
rect 339963 626924 340035 626980
rect 339963 626890 339982 626924
rect 340016 626890 340035 626924
rect 339963 626834 340035 626890
rect 339963 626800 339982 626834
rect 340016 626800 340035 626834
rect 339963 626744 340035 626800
rect 340853 627411 340872 627445
rect 340906 627411 340925 627445
rect 340853 627355 340925 627411
rect 340853 627321 340872 627355
rect 340906 627321 340925 627355
rect 340853 627265 340925 627321
rect 340853 627231 340872 627265
rect 340906 627231 340925 627265
rect 340853 627175 340925 627231
rect 340853 627141 340872 627175
rect 340906 627141 340925 627175
rect 340853 627085 340925 627141
rect 340853 627051 340872 627085
rect 340906 627051 340925 627085
rect 340853 626995 340925 627051
rect 340853 626961 340872 626995
rect 340906 626961 340925 626995
rect 340853 626905 340925 626961
rect 340853 626871 340872 626905
rect 340906 626871 340925 626905
rect 340853 626815 340925 626871
rect 340853 626781 340872 626815
rect 340906 626781 340925 626815
rect 339963 626710 339982 626744
rect 340016 626710 340035 626744
rect 339963 626687 340035 626710
rect 340853 626725 340925 626781
rect 340853 626691 340872 626725
rect 340906 626691 340925 626725
rect 340853 626687 340925 626691
rect 339963 626668 340925 626687
rect 339963 626634 340040 626668
rect 340074 626634 340130 626668
rect 340164 626634 340220 626668
rect 340254 626634 340310 626668
rect 340344 626634 340400 626668
rect 340434 626634 340490 626668
rect 340524 626634 340580 626668
rect 340614 626634 340670 626668
rect 340704 626634 340760 626668
rect 340794 626634 340925 626668
rect 339963 626615 340925 626634
rect 334811 626270 335773 626289
rect 334811 626236 334922 626270
rect 334956 626236 335012 626270
rect 335046 626236 335102 626270
rect 335136 626236 335192 626270
rect 335226 626236 335282 626270
rect 335316 626236 335372 626270
rect 335406 626236 335462 626270
rect 335496 626236 335552 626270
rect 335586 626236 335642 626270
rect 335676 626236 335773 626270
rect 334811 626217 335773 626236
rect 334811 626176 334883 626217
rect 334811 626142 334830 626176
rect 334864 626142 334883 626176
rect 335701 626157 335773 626217
rect 334811 626086 334883 626142
rect 334811 626052 334830 626086
rect 334864 626052 334883 626086
rect 334811 625996 334883 626052
rect 334811 625962 334830 625996
rect 334864 625962 334883 625996
rect 334811 625906 334883 625962
rect 334811 625872 334830 625906
rect 334864 625872 334883 625906
rect 334811 625816 334883 625872
rect 334811 625782 334830 625816
rect 334864 625782 334883 625816
rect 334811 625726 334883 625782
rect 334811 625692 334830 625726
rect 334864 625692 334883 625726
rect 334811 625636 334883 625692
rect 334811 625602 334830 625636
rect 334864 625602 334883 625636
rect 334811 625546 334883 625602
rect 334811 625512 334830 625546
rect 334864 625512 334883 625546
rect 334811 625456 334883 625512
rect 335701 626123 335720 626157
rect 335754 626123 335773 626157
rect 335701 626067 335773 626123
rect 335701 626033 335720 626067
rect 335754 626033 335773 626067
rect 335701 625977 335773 626033
rect 335701 625943 335720 625977
rect 335754 625943 335773 625977
rect 335701 625887 335773 625943
rect 335701 625853 335720 625887
rect 335754 625853 335773 625887
rect 335701 625797 335773 625853
rect 335701 625763 335720 625797
rect 335754 625763 335773 625797
rect 335701 625707 335773 625763
rect 335701 625673 335720 625707
rect 335754 625673 335773 625707
rect 335701 625617 335773 625673
rect 335701 625583 335720 625617
rect 335754 625583 335773 625617
rect 335701 625527 335773 625583
rect 335701 625493 335720 625527
rect 335754 625493 335773 625527
rect 334811 625422 334830 625456
rect 334864 625422 334883 625456
rect 334811 625399 334883 625422
rect 335701 625437 335773 625493
rect 335701 625403 335720 625437
rect 335754 625403 335773 625437
rect 335701 625399 335773 625403
rect 334811 625380 335773 625399
rect 334811 625346 334888 625380
rect 334922 625346 334978 625380
rect 335012 625346 335068 625380
rect 335102 625346 335158 625380
rect 335192 625346 335248 625380
rect 335282 625346 335338 625380
rect 335372 625346 335428 625380
rect 335462 625346 335518 625380
rect 335552 625346 335608 625380
rect 335642 625346 335773 625380
rect 334811 625327 335773 625346
rect 336099 626270 337061 626289
rect 336099 626236 336210 626270
rect 336244 626236 336300 626270
rect 336334 626236 336390 626270
rect 336424 626236 336480 626270
rect 336514 626236 336570 626270
rect 336604 626236 336660 626270
rect 336694 626236 336750 626270
rect 336784 626236 336840 626270
rect 336874 626236 336930 626270
rect 336964 626236 337061 626270
rect 336099 626217 337061 626236
rect 336099 626176 336171 626217
rect 336099 626142 336118 626176
rect 336152 626142 336171 626176
rect 336989 626157 337061 626217
rect 336099 626086 336171 626142
rect 336099 626052 336118 626086
rect 336152 626052 336171 626086
rect 336099 625996 336171 626052
rect 336099 625962 336118 625996
rect 336152 625962 336171 625996
rect 336099 625906 336171 625962
rect 336099 625872 336118 625906
rect 336152 625872 336171 625906
rect 336099 625816 336171 625872
rect 336099 625782 336118 625816
rect 336152 625782 336171 625816
rect 336099 625726 336171 625782
rect 336099 625692 336118 625726
rect 336152 625692 336171 625726
rect 336099 625636 336171 625692
rect 336099 625602 336118 625636
rect 336152 625602 336171 625636
rect 336099 625546 336171 625602
rect 336099 625512 336118 625546
rect 336152 625512 336171 625546
rect 336099 625456 336171 625512
rect 336989 626123 337008 626157
rect 337042 626123 337061 626157
rect 336989 626067 337061 626123
rect 336989 626033 337008 626067
rect 337042 626033 337061 626067
rect 336989 625977 337061 626033
rect 336989 625943 337008 625977
rect 337042 625943 337061 625977
rect 336989 625887 337061 625943
rect 336989 625853 337008 625887
rect 337042 625853 337061 625887
rect 336989 625797 337061 625853
rect 336989 625763 337008 625797
rect 337042 625763 337061 625797
rect 336989 625707 337061 625763
rect 336989 625673 337008 625707
rect 337042 625673 337061 625707
rect 336989 625617 337061 625673
rect 336989 625583 337008 625617
rect 337042 625583 337061 625617
rect 336989 625527 337061 625583
rect 336989 625493 337008 625527
rect 337042 625493 337061 625527
rect 336099 625422 336118 625456
rect 336152 625422 336171 625456
rect 336099 625399 336171 625422
rect 336989 625437 337061 625493
rect 336989 625403 337008 625437
rect 337042 625403 337061 625437
rect 336989 625399 337061 625403
rect 336099 625380 337061 625399
rect 336099 625346 336176 625380
rect 336210 625346 336266 625380
rect 336300 625346 336356 625380
rect 336390 625346 336446 625380
rect 336480 625346 336536 625380
rect 336570 625346 336626 625380
rect 336660 625346 336716 625380
rect 336750 625346 336806 625380
rect 336840 625346 336896 625380
rect 336930 625346 337061 625380
rect 336099 625327 337061 625346
rect 337387 626270 338349 626289
rect 337387 626236 337498 626270
rect 337532 626236 337588 626270
rect 337622 626236 337678 626270
rect 337712 626236 337768 626270
rect 337802 626236 337858 626270
rect 337892 626236 337948 626270
rect 337982 626236 338038 626270
rect 338072 626236 338128 626270
rect 338162 626236 338218 626270
rect 338252 626236 338349 626270
rect 337387 626217 338349 626236
rect 337387 626176 337459 626217
rect 337387 626142 337406 626176
rect 337440 626142 337459 626176
rect 338277 626157 338349 626217
rect 337387 626086 337459 626142
rect 337387 626052 337406 626086
rect 337440 626052 337459 626086
rect 337387 625996 337459 626052
rect 337387 625962 337406 625996
rect 337440 625962 337459 625996
rect 337387 625906 337459 625962
rect 337387 625872 337406 625906
rect 337440 625872 337459 625906
rect 337387 625816 337459 625872
rect 337387 625782 337406 625816
rect 337440 625782 337459 625816
rect 337387 625726 337459 625782
rect 337387 625692 337406 625726
rect 337440 625692 337459 625726
rect 337387 625636 337459 625692
rect 337387 625602 337406 625636
rect 337440 625602 337459 625636
rect 337387 625546 337459 625602
rect 337387 625512 337406 625546
rect 337440 625512 337459 625546
rect 337387 625456 337459 625512
rect 338277 626123 338296 626157
rect 338330 626123 338349 626157
rect 338277 626067 338349 626123
rect 338277 626033 338296 626067
rect 338330 626033 338349 626067
rect 338277 625977 338349 626033
rect 338277 625943 338296 625977
rect 338330 625943 338349 625977
rect 338277 625887 338349 625943
rect 338277 625853 338296 625887
rect 338330 625853 338349 625887
rect 338277 625797 338349 625853
rect 338277 625763 338296 625797
rect 338330 625763 338349 625797
rect 338277 625707 338349 625763
rect 338277 625673 338296 625707
rect 338330 625673 338349 625707
rect 338277 625617 338349 625673
rect 338277 625583 338296 625617
rect 338330 625583 338349 625617
rect 338277 625527 338349 625583
rect 338277 625493 338296 625527
rect 338330 625493 338349 625527
rect 337387 625422 337406 625456
rect 337440 625422 337459 625456
rect 337387 625399 337459 625422
rect 338277 625437 338349 625493
rect 338277 625403 338296 625437
rect 338330 625403 338349 625437
rect 338277 625399 338349 625403
rect 337387 625380 338349 625399
rect 337387 625346 337464 625380
rect 337498 625346 337554 625380
rect 337588 625346 337644 625380
rect 337678 625346 337734 625380
rect 337768 625346 337824 625380
rect 337858 625346 337914 625380
rect 337948 625346 338004 625380
rect 338038 625346 338094 625380
rect 338128 625346 338184 625380
rect 338218 625346 338349 625380
rect 337387 625327 338349 625346
rect 338675 626270 339637 626289
rect 338675 626236 338786 626270
rect 338820 626236 338876 626270
rect 338910 626236 338966 626270
rect 339000 626236 339056 626270
rect 339090 626236 339146 626270
rect 339180 626236 339236 626270
rect 339270 626236 339326 626270
rect 339360 626236 339416 626270
rect 339450 626236 339506 626270
rect 339540 626236 339637 626270
rect 338675 626217 339637 626236
rect 338675 626176 338747 626217
rect 338675 626142 338694 626176
rect 338728 626142 338747 626176
rect 339565 626157 339637 626217
rect 338675 626086 338747 626142
rect 338675 626052 338694 626086
rect 338728 626052 338747 626086
rect 338675 625996 338747 626052
rect 338675 625962 338694 625996
rect 338728 625962 338747 625996
rect 338675 625906 338747 625962
rect 338675 625872 338694 625906
rect 338728 625872 338747 625906
rect 338675 625816 338747 625872
rect 338675 625782 338694 625816
rect 338728 625782 338747 625816
rect 338675 625726 338747 625782
rect 338675 625692 338694 625726
rect 338728 625692 338747 625726
rect 338675 625636 338747 625692
rect 338675 625602 338694 625636
rect 338728 625602 338747 625636
rect 338675 625546 338747 625602
rect 338675 625512 338694 625546
rect 338728 625512 338747 625546
rect 338675 625456 338747 625512
rect 339565 626123 339584 626157
rect 339618 626123 339637 626157
rect 339565 626067 339637 626123
rect 339565 626033 339584 626067
rect 339618 626033 339637 626067
rect 339565 625977 339637 626033
rect 339565 625943 339584 625977
rect 339618 625943 339637 625977
rect 339565 625887 339637 625943
rect 339565 625853 339584 625887
rect 339618 625853 339637 625887
rect 339565 625797 339637 625853
rect 339565 625763 339584 625797
rect 339618 625763 339637 625797
rect 339565 625707 339637 625763
rect 339565 625673 339584 625707
rect 339618 625673 339637 625707
rect 339565 625617 339637 625673
rect 339565 625583 339584 625617
rect 339618 625583 339637 625617
rect 339565 625527 339637 625583
rect 339565 625493 339584 625527
rect 339618 625493 339637 625527
rect 338675 625422 338694 625456
rect 338728 625422 338747 625456
rect 338675 625399 338747 625422
rect 339565 625437 339637 625493
rect 339565 625403 339584 625437
rect 339618 625403 339637 625437
rect 339565 625399 339637 625403
rect 338675 625380 339637 625399
rect 338675 625346 338752 625380
rect 338786 625346 338842 625380
rect 338876 625346 338932 625380
rect 338966 625346 339022 625380
rect 339056 625346 339112 625380
rect 339146 625346 339202 625380
rect 339236 625346 339292 625380
rect 339326 625346 339382 625380
rect 339416 625346 339472 625380
rect 339506 625346 339637 625380
rect 338675 625327 339637 625346
rect 339963 626270 340925 626289
rect 339963 626236 340074 626270
rect 340108 626236 340164 626270
rect 340198 626236 340254 626270
rect 340288 626236 340344 626270
rect 340378 626236 340434 626270
rect 340468 626236 340524 626270
rect 340558 626236 340614 626270
rect 340648 626236 340704 626270
rect 340738 626236 340794 626270
rect 340828 626236 340925 626270
rect 339963 626217 340925 626236
rect 339963 626176 340035 626217
rect 339963 626142 339982 626176
rect 340016 626142 340035 626176
rect 340853 626157 340925 626217
rect 339963 626086 340035 626142
rect 339963 626052 339982 626086
rect 340016 626052 340035 626086
rect 339963 625996 340035 626052
rect 339963 625962 339982 625996
rect 340016 625962 340035 625996
rect 339963 625906 340035 625962
rect 339963 625872 339982 625906
rect 340016 625872 340035 625906
rect 339963 625816 340035 625872
rect 339963 625782 339982 625816
rect 340016 625782 340035 625816
rect 339963 625726 340035 625782
rect 339963 625692 339982 625726
rect 340016 625692 340035 625726
rect 339963 625636 340035 625692
rect 339963 625602 339982 625636
rect 340016 625602 340035 625636
rect 339963 625546 340035 625602
rect 339963 625512 339982 625546
rect 340016 625512 340035 625546
rect 339963 625456 340035 625512
rect 340853 626123 340872 626157
rect 340906 626123 340925 626157
rect 340853 626067 340925 626123
rect 340853 626033 340872 626067
rect 340906 626033 340925 626067
rect 340853 625977 340925 626033
rect 340853 625943 340872 625977
rect 340906 625943 340925 625977
rect 340853 625887 340925 625943
rect 340853 625853 340872 625887
rect 340906 625853 340925 625887
rect 340853 625797 340925 625853
rect 340853 625763 340872 625797
rect 340906 625763 340925 625797
rect 340853 625707 340925 625763
rect 340853 625673 340872 625707
rect 340906 625673 340925 625707
rect 340853 625617 340925 625673
rect 340853 625583 340872 625617
rect 340906 625583 340925 625617
rect 340853 625527 340925 625583
rect 340853 625493 340872 625527
rect 340906 625493 340925 625527
rect 339963 625422 339982 625456
rect 340016 625422 340035 625456
rect 339963 625399 340035 625422
rect 340853 625437 340925 625493
rect 340853 625403 340872 625437
rect 340906 625403 340925 625437
rect 340853 625399 340925 625403
rect 339963 625380 340925 625399
rect 339963 625346 340040 625380
rect 340074 625346 340130 625380
rect 340164 625346 340220 625380
rect 340254 625346 340310 625380
rect 340344 625346 340400 625380
rect 340434 625346 340490 625380
rect 340524 625346 340580 625380
rect 340614 625346 340670 625380
rect 340704 625346 340760 625380
rect 340794 625346 340925 625380
rect 339963 625327 340925 625346
rect 312704 624608 313304 624808
rect 302904 619648 303104 619748
rect 302904 617306 302954 619648
rect 303054 617306 303104 619648
rect 302904 617206 303104 617306
rect 312032 619648 312232 619748
rect 312032 617306 312082 619648
rect 312182 617306 312232 619648
rect 312704 617608 312904 624608
rect 313104 617608 313304 624608
rect 312704 617408 313304 617608
rect 312032 617206 312232 617306
rect 318614 624608 319214 624808
rect 318614 617608 318814 624608
rect 319014 617608 319214 624608
rect 318614 617408 319214 617608
rect 324114 624608 324714 624808
rect 324114 617608 324314 624608
rect 324514 617608 324714 624608
rect 324114 617408 324714 617608
rect 330070 624606 330670 624806
rect 330070 617606 330270 624606
rect 330470 617606 330670 624606
rect 330070 617406 330670 617606
rect 334811 624982 335773 625001
rect 334811 624948 334922 624982
rect 334956 624948 335012 624982
rect 335046 624948 335102 624982
rect 335136 624948 335192 624982
rect 335226 624948 335282 624982
rect 335316 624948 335372 624982
rect 335406 624948 335462 624982
rect 335496 624948 335552 624982
rect 335586 624948 335642 624982
rect 335676 624948 335773 624982
rect 334811 624929 335773 624948
rect 334811 624888 334883 624929
rect 334811 624854 334830 624888
rect 334864 624854 334883 624888
rect 335701 624869 335773 624929
rect 334811 624798 334883 624854
rect 334811 624764 334830 624798
rect 334864 624764 334883 624798
rect 334811 624708 334883 624764
rect 334811 624674 334830 624708
rect 334864 624674 334883 624708
rect 334811 624618 334883 624674
rect 334811 624584 334830 624618
rect 334864 624584 334883 624618
rect 334811 624528 334883 624584
rect 334811 624494 334830 624528
rect 334864 624494 334883 624528
rect 334811 624438 334883 624494
rect 334811 624404 334830 624438
rect 334864 624404 334883 624438
rect 334811 624348 334883 624404
rect 334811 624314 334830 624348
rect 334864 624314 334883 624348
rect 334811 624258 334883 624314
rect 334811 624224 334830 624258
rect 334864 624224 334883 624258
rect 334811 624168 334883 624224
rect 335701 624835 335720 624869
rect 335754 624835 335773 624869
rect 335701 624779 335773 624835
rect 335701 624745 335720 624779
rect 335754 624745 335773 624779
rect 335701 624689 335773 624745
rect 335701 624655 335720 624689
rect 335754 624655 335773 624689
rect 335701 624599 335773 624655
rect 335701 624565 335720 624599
rect 335754 624565 335773 624599
rect 335701 624509 335773 624565
rect 335701 624475 335720 624509
rect 335754 624475 335773 624509
rect 335701 624419 335773 624475
rect 335701 624385 335720 624419
rect 335754 624385 335773 624419
rect 335701 624329 335773 624385
rect 335701 624295 335720 624329
rect 335754 624295 335773 624329
rect 335701 624239 335773 624295
rect 335701 624205 335720 624239
rect 335754 624205 335773 624239
rect 334811 624134 334830 624168
rect 334864 624134 334883 624168
rect 334811 624111 334883 624134
rect 335701 624149 335773 624205
rect 335701 624115 335720 624149
rect 335754 624115 335773 624149
rect 335701 624111 335773 624115
rect 334811 624092 335773 624111
rect 334811 624058 334888 624092
rect 334922 624058 334978 624092
rect 335012 624058 335068 624092
rect 335102 624058 335158 624092
rect 335192 624058 335248 624092
rect 335282 624058 335338 624092
rect 335372 624058 335428 624092
rect 335462 624058 335518 624092
rect 335552 624058 335608 624092
rect 335642 624058 335773 624092
rect 334811 624039 335773 624058
rect 336099 624982 337061 625001
rect 336099 624948 336210 624982
rect 336244 624948 336300 624982
rect 336334 624948 336390 624982
rect 336424 624948 336480 624982
rect 336514 624948 336570 624982
rect 336604 624948 336660 624982
rect 336694 624948 336750 624982
rect 336784 624948 336840 624982
rect 336874 624948 336930 624982
rect 336964 624948 337061 624982
rect 336099 624929 337061 624948
rect 336099 624888 336171 624929
rect 336099 624854 336118 624888
rect 336152 624854 336171 624888
rect 336989 624869 337061 624929
rect 336099 624798 336171 624854
rect 336099 624764 336118 624798
rect 336152 624764 336171 624798
rect 336099 624708 336171 624764
rect 336099 624674 336118 624708
rect 336152 624674 336171 624708
rect 336099 624618 336171 624674
rect 336099 624584 336118 624618
rect 336152 624584 336171 624618
rect 336099 624528 336171 624584
rect 336099 624494 336118 624528
rect 336152 624494 336171 624528
rect 336099 624438 336171 624494
rect 336099 624404 336118 624438
rect 336152 624404 336171 624438
rect 336099 624348 336171 624404
rect 336099 624314 336118 624348
rect 336152 624314 336171 624348
rect 336099 624258 336171 624314
rect 336099 624224 336118 624258
rect 336152 624224 336171 624258
rect 336099 624168 336171 624224
rect 336989 624835 337008 624869
rect 337042 624835 337061 624869
rect 336989 624779 337061 624835
rect 336989 624745 337008 624779
rect 337042 624745 337061 624779
rect 336989 624689 337061 624745
rect 336989 624655 337008 624689
rect 337042 624655 337061 624689
rect 336989 624599 337061 624655
rect 336989 624565 337008 624599
rect 337042 624565 337061 624599
rect 336989 624509 337061 624565
rect 336989 624475 337008 624509
rect 337042 624475 337061 624509
rect 336989 624419 337061 624475
rect 336989 624385 337008 624419
rect 337042 624385 337061 624419
rect 336989 624329 337061 624385
rect 336989 624295 337008 624329
rect 337042 624295 337061 624329
rect 336989 624239 337061 624295
rect 336989 624205 337008 624239
rect 337042 624205 337061 624239
rect 336099 624134 336118 624168
rect 336152 624134 336171 624168
rect 336099 624111 336171 624134
rect 336989 624149 337061 624205
rect 336989 624115 337008 624149
rect 337042 624115 337061 624149
rect 336989 624111 337061 624115
rect 336099 624092 337061 624111
rect 336099 624058 336176 624092
rect 336210 624058 336266 624092
rect 336300 624058 336356 624092
rect 336390 624058 336446 624092
rect 336480 624058 336536 624092
rect 336570 624058 336626 624092
rect 336660 624058 336716 624092
rect 336750 624058 336806 624092
rect 336840 624058 336896 624092
rect 336930 624058 337061 624092
rect 336099 624039 337061 624058
rect 337387 624982 338349 625001
rect 337387 624948 337498 624982
rect 337532 624948 337588 624982
rect 337622 624948 337678 624982
rect 337712 624948 337768 624982
rect 337802 624948 337858 624982
rect 337892 624948 337948 624982
rect 337982 624948 338038 624982
rect 338072 624948 338128 624982
rect 338162 624948 338218 624982
rect 338252 624948 338349 624982
rect 337387 624929 338349 624948
rect 337387 624888 337459 624929
rect 337387 624854 337406 624888
rect 337440 624854 337459 624888
rect 338277 624869 338349 624929
rect 337387 624798 337459 624854
rect 337387 624764 337406 624798
rect 337440 624764 337459 624798
rect 337387 624708 337459 624764
rect 337387 624674 337406 624708
rect 337440 624674 337459 624708
rect 337387 624618 337459 624674
rect 337387 624584 337406 624618
rect 337440 624584 337459 624618
rect 337387 624528 337459 624584
rect 337387 624494 337406 624528
rect 337440 624494 337459 624528
rect 337387 624438 337459 624494
rect 337387 624404 337406 624438
rect 337440 624404 337459 624438
rect 337387 624348 337459 624404
rect 337387 624314 337406 624348
rect 337440 624314 337459 624348
rect 337387 624258 337459 624314
rect 337387 624224 337406 624258
rect 337440 624224 337459 624258
rect 337387 624168 337459 624224
rect 338277 624835 338296 624869
rect 338330 624835 338349 624869
rect 338277 624779 338349 624835
rect 338277 624745 338296 624779
rect 338330 624745 338349 624779
rect 338277 624689 338349 624745
rect 338277 624655 338296 624689
rect 338330 624655 338349 624689
rect 338277 624599 338349 624655
rect 338277 624565 338296 624599
rect 338330 624565 338349 624599
rect 338277 624509 338349 624565
rect 338277 624475 338296 624509
rect 338330 624475 338349 624509
rect 338277 624419 338349 624475
rect 338277 624385 338296 624419
rect 338330 624385 338349 624419
rect 338277 624329 338349 624385
rect 338277 624295 338296 624329
rect 338330 624295 338349 624329
rect 338277 624239 338349 624295
rect 338277 624205 338296 624239
rect 338330 624205 338349 624239
rect 337387 624134 337406 624168
rect 337440 624134 337459 624168
rect 337387 624111 337459 624134
rect 338277 624149 338349 624205
rect 338277 624115 338296 624149
rect 338330 624115 338349 624149
rect 338277 624111 338349 624115
rect 337387 624092 338349 624111
rect 337387 624058 337464 624092
rect 337498 624058 337554 624092
rect 337588 624058 337644 624092
rect 337678 624058 337734 624092
rect 337768 624058 337824 624092
rect 337858 624058 337914 624092
rect 337948 624058 338004 624092
rect 338038 624058 338094 624092
rect 338128 624058 338184 624092
rect 338218 624058 338349 624092
rect 337387 624039 338349 624058
rect 338675 624982 339637 625001
rect 338675 624948 338786 624982
rect 338820 624948 338876 624982
rect 338910 624948 338966 624982
rect 339000 624948 339056 624982
rect 339090 624948 339146 624982
rect 339180 624948 339236 624982
rect 339270 624948 339326 624982
rect 339360 624948 339416 624982
rect 339450 624948 339506 624982
rect 339540 624948 339637 624982
rect 338675 624929 339637 624948
rect 338675 624888 338747 624929
rect 338675 624854 338694 624888
rect 338728 624854 338747 624888
rect 339565 624869 339637 624929
rect 338675 624798 338747 624854
rect 338675 624764 338694 624798
rect 338728 624764 338747 624798
rect 338675 624708 338747 624764
rect 338675 624674 338694 624708
rect 338728 624674 338747 624708
rect 338675 624618 338747 624674
rect 338675 624584 338694 624618
rect 338728 624584 338747 624618
rect 338675 624528 338747 624584
rect 338675 624494 338694 624528
rect 338728 624494 338747 624528
rect 338675 624438 338747 624494
rect 338675 624404 338694 624438
rect 338728 624404 338747 624438
rect 338675 624348 338747 624404
rect 338675 624314 338694 624348
rect 338728 624314 338747 624348
rect 338675 624258 338747 624314
rect 338675 624224 338694 624258
rect 338728 624224 338747 624258
rect 338675 624168 338747 624224
rect 339565 624835 339584 624869
rect 339618 624835 339637 624869
rect 339565 624779 339637 624835
rect 339565 624745 339584 624779
rect 339618 624745 339637 624779
rect 339565 624689 339637 624745
rect 339565 624655 339584 624689
rect 339618 624655 339637 624689
rect 339565 624599 339637 624655
rect 339565 624565 339584 624599
rect 339618 624565 339637 624599
rect 339565 624509 339637 624565
rect 339565 624475 339584 624509
rect 339618 624475 339637 624509
rect 339565 624419 339637 624475
rect 339565 624385 339584 624419
rect 339618 624385 339637 624419
rect 339565 624329 339637 624385
rect 339565 624295 339584 624329
rect 339618 624295 339637 624329
rect 339565 624239 339637 624295
rect 339565 624205 339584 624239
rect 339618 624205 339637 624239
rect 338675 624134 338694 624168
rect 338728 624134 338747 624168
rect 338675 624111 338747 624134
rect 339565 624149 339637 624205
rect 339565 624115 339584 624149
rect 339618 624115 339637 624149
rect 339565 624111 339637 624115
rect 338675 624092 339637 624111
rect 338675 624058 338752 624092
rect 338786 624058 338842 624092
rect 338876 624058 338932 624092
rect 338966 624058 339022 624092
rect 339056 624058 339112 624092
rect 339146 624058 339202 624092
rect 339236 624058 339292 624092
rect 339326 624058 339382 624092
rect 339416 624058 339472 624092
rect 339506 624058 339637 624092
rect 338675 624039 339637 624058
rect 339963 624982 340925 625001
rect 339963 624948 340074 624982
rect 340108 624948 340164 624982
rect 340198 624948 340254 624982
rect 340288 624948 340344 624982
rect 340378 624948 340434 624982
rect 340468 624948 340524 624982
rect 340558 624948 340614 624982
rect 340648 624948 340704 624982
rect 340738 624948 340794 624982
rect 340828 624948 340925 624982
rect 339963 624929 340925 624948
rect 339963 624888 340035 624929
rect 339963 624854 339982 624888
rect 340016 624854 340035 624888
rect 340853 624869 340925 624929
rect 339963 624798 340035 624854
rect 339963 624764 339982 624798
rect 340016 624764 340035 624798
rect 339963 624708 340035 624764
rect 339963 624674 339982 624708
rect 340016 624674 340035 624708
rect 339963 624618 340035 624674
rect 339963 624584 339982 624618
rect 340016 624584 340035 624618
rect 339963 624528 340035 624584
rect 339963 624494 339982 624528
rect 340016 624494 340035 624528
rect 339963 624438 340035 624494
rect 339963 624404 339982 624438
rect 340016 624404 340035 624438
rect 339963 624348 340035 624404
rect 339963 624314 339982 624348
rect 340016 624314 340035 624348
rect 339963 624258 340035 624314
rect 339963 624224 339982 624258
rect 340016 624224 340035 624258
rect 339963 624168 340035 624224
rect 340853 624835 340872 624869
rect 340906 624835 340925 624869
rect 340853 624779 340925 624835
rect 340853 624745 340872 624779
rect 340906 624745 340925 624779
rect 340853 624689 340925 624745
rect 340853 624655 340872 624689
rect 340906 624655 340925 624689
rect 340853 624599 340925 624655
rect 340853 624565 340872 624599
rect 340906 624565 340925 624599
rect 340853 624509 340925 624565
rect 340853 624475 340872 624509
rect 340906 624475 340925 624509
rect 340853 624419 340925 624475
rect 340853 624385 340872 624419
rect 340906 624385 340925 624419
rect 340853 624329 340925 624385
rect 340853 624295 340872 624329
rect 340906 624295 340925 624329
rect 340853 624239 340925 624295
rect 340853 624205 340872 624239
rect 340906 624205 340925 624239
rect 339963 624134 339982 624168
rect 340016 624134 340035 624168
rect 339963 624111 340035 624134
rect 340853 624149 340925 624205
rect 340853 624115 340872 624149
rect 340906 624115 340925 624149
rect 340853 624111 340925 624115
rect 339963 624092 340925 624111
rect 339963 624058 340040 624092
rect 340074 624058 340130 624092
rect 340164 624058 340220 624092
rect 340254 624058 340310 624092
rect 340344 624058 340400 624092
rect 340434 624058 340490 624092
rect 340524 624058 340580 624092
rect 340614 624058 340670 624092
rect 340704 624058 340760 624092
rect 340794 624058 340925 624092
rect 339963 624039 340925 624058
rect 334811 623694 335773 623713
rect 334811 623660 334922 623694
rect 334956 623660 335012 623694
rect 335046 623660 335102 623694
rect 335136 623660 335192 623694
rect 335226 623660 335282 623694
rect 335316 623660 335372 623694
rect 335406 623660 335462 623694
rect 335496 623660 335552 623694
rect 335586 623660 335642 623694
rect 335676 623660 335773 623694
rect 334811 623641 335773 623660
rect 334811 623600 334883 623641
rect 334811 623566 334830 623600
rect 334864 623566 334883 623600
rect 335701 623581 335773 623641
rect 334811 623510 334883 623566
rect 334811 623476 334830 623510
rect 334864 623476 334883 623510
rect 334811 623420 334883 623476
rect 334811 623386 334830 623420
rect 334864 623386 334883 623420
rect 334811 623330 334883 623386
rect 334811 623296 334830 623330
rect 334864 623296 334883 623330
rect 334811 623240 334883 623296
rect 334811 623206 334830 623240
rect 334864 623206 334883 623240
rect 334811 623150 334883 623206
rect 334811 623116 334830 623150
rect 334864 623116 334883 623150
rect 334811 623060 334883 623116
rect 334811 623026 334830 623060
rect 334864 623026 334883 623060
rect 334811 622970 334883 623026
rect 334811 622936 334830 622970
rect 334864 622936 334883 622970
rect 334811 622880 334883 622936
rect 335701 623547 335720 623581
rect 335754 623547 335773 623581
rect 335701 623491 335773 623547
rect 335701 623457 335720 623491
rect 335754 623457 335773 623491
rect 335701 623401 335773 623457
rect 335701 623367 335720 623401
rect 335754 623367 335773 623401
rect 335701 623311 335773 623367
rect 335701 623277 335720 623311
rect 335754 623277 335773 623311
rect 335701 623221 335773 623277
rect 335701 623187 335720 623221
rect 335754 623187 335773 623221
rect 335701 623131 335773 623187
rect 335701 623097 335720 623131
rect 335754 623097 335773 623131
rect 335701 623041 335773 623097
rect 335701 623007 335720 623041
rect 335754 623007 335773 623041
rect 335701 622951 335773 623007
rect 335701 622917 335720 622951
rect 335754 622917 335773 622951
rect 334811 622846 334830 622880
rect 334864 622846 334883 622880
rect 334811 622823 334883 622846
rect 335701 622861 335773 622917
rect 335701 622827 335720 622861
rect 335754 622827 335773 622861
rect 335701 622823 335773 622827
rect 334811 622804 335773 622823
rect 334811 622770 334888 622804
rect 334922 622770 334978 622804
rect 335012 622770 335068 622804
rect 335102 622770 335158 622804
rect 335192 622770 335248 622804
rect 335282 622770 335338 622804
rect 335372 622770 335428 622804
rect 335462 622770 335518 622804
rect 335552 622770 335608 622804
rect 335642 622770 335773 622804
rect 334811 622751 335773 622770
rect 336099 623694 337061 623713
rect 336099 623660 336210 623694
rect 336244 623660 336300 623694
rect 336334 623660 336390 623694
rect 336424 623660 336480 623694
rect 336514 623660 336570 623694
rect 336604 623660 336660 623694
rect 336694 623660 336750 623694
rect 336784 623660 336840 623694
rect 336874 623660 336930 623694
rect 336964 623660 337061 623694
rect 336099 623641 337061 623660
rect 336099 623600 336171 623641
rect 336099 623566 336118 623600
rect 336152 623566 336171 623600
rect 336989 623581 337061 623641
rect 336099 623510 336171 623566
rect 336099 623476 336118 623510
rect 336152 623476 336171 623510
rect 336099 623420 336171 623476
rect 336099 623386 336118 623420
rect 336152 623386 336171 623420
rect 336099 623330 336171 623386
rect 336099 623296 336118 623330
rect 336152 623296 336171 623330
rect 336099 623240 336171 623296
rect 336099 623206 336118 623240
rect 336152 623206 336171 623240
rect 336099 623150 336171 623206
rect 336099 623116 336118 623150
rect 336152 623116 336171 623150
rect 336099 623060 336171 623116
rect 336099 623026 336118 623060
rect 336152 623026 336171 623060
rect 336099 622970 336171 623026
rect 336099 622936 336118 622970
rect 336152 622936 336171 622970
rect 336099 622880 336171 622936
rect 336989 623547 337008 623581
rect 337042 623547 337061 623581
rect 336989 623491 337061 623547
rect 336989 623457 337008 623491
rect 337042 623457 337061 623491
rect 336989 623401 337061 623457
rect 336989 623367 337008 623401
rect 337042 623367 337061 623401
rect 336989 623311 337061 623367
rect 336989 623277 337008 623311
rect 337042 623277 337061 623311
rect 336989 623221 337061 623277
rect 336989 623187 337008 623221
rect 337042 623187 337061 623221
rect 336989 623131 337061 623187
rect 336989 623097 337008 623131
rect 337042 623097 337061 623131
rect 336989 623041 337061 623097
rect 336989 623007 337008 623041
rect 337042 623007 337061 623041
rect 336989 622951 337061 623007
rect 336989 622917 337008 622951
rect 337042 622917 337061 622951
rect 336099 622846 336118 622880
rect 336152 622846 336171 622880
rect 336099 622823 336171 622846
rect 336989 622861 337061 622917
rect 336989 622827 337008 622861
rect 337042 622827 337061 622861
rect 336989 622823 337061 622827
rect 336099 622804 337061 622823
rect 336099 622770 336176 622804
rect 336210 622770 336266 622804
rect 336300 622770 336356 622804
rect 336390 622770 336446 622804
rect 336480 622770 336536 622804
rect 336570 622770 336626 622804
rect 336660 622770 336716 622804
rect 336750 622770 336806 622804
rect 336840 622770 336896 622804
rect 336930 622770 337061 622804
rect 336099 622751 337061 622770
rect 337387 623694 338349 623713
rect 337387 623660 337498 623694
rect 337532 623660 337588 623694
rect 337622 623660 337678 623694
rect 337712 623660 337768 623694
rect 337802 623660 337858 623694
rect 337892 623660 337948 623694
rect 337982 623660 338038 623694
rect 338072 623660 338128 623694
rect 338162 623660 338218 623694
rect 338252 623660 338349 623694
rect 337387 623641 338349 623660
rect 337387 623600 337459 623641
rect 337387 623566 337406 623600
rect 337440 623566 337459 623600
rect 338277 623581 338349 623641
rect 337387 623510 337459 623566
rect 337387 623476 337406 623510
rect 337440 623476 337459 623510
rect 337387 623420 337459 623476
rect 337387 623386 337406 623420
rect 337440 623386 337459 623420
rect 337387 623330 337459 623386
rect 337387 623296 337406 623330
rect 337440 623296 337459 623330
rect 337387 623240 337459 623296
rect 337387 623206 337406 623240
rect 337440 623206 337459 623240
rect 337387 623150 337459 623206
rect 337387 623116 337406 623150
rect 337440 623116 337459 623150
rect 337387 623060 337459 623116
rect 337387 623026 337406 623060
rect 337440 623026 337459 623060
rect 337387 622970 337459 623026
rect 337387 622936 337406 622970
rect 337440 622936 337459 622970
rect 337387 622880 337459 622936
rect 338277 623547 338296 623581
rect 338330 623547 338349 623581
rect 338277 623491 338349 623547
rect 338277 623457 338296 623491
rect 338330 623457 338349 623491
rect 338277 623401 338349 623457
rect 338277 623367 338296 623401
rect 338330 623367 338349 623401
rect 338277 623311 338349 623367
rect 338277 623277 338296 623311
rect 338330 623277 338349 623311
rect 338277 623221 338349 623277
rect 338277 623187 338296 623221
rect 338330 623187 338349 623221
rect 338277 623131 338349 623187
rect 338277 623097 338296 623131
rect 338330 623097 338349 623131
rect 338277 623041 338349 623097
rect 338277 623007 338296 623041
rect 338330 623007 338349 623041
rect 338277 622951 338349 623007
rect 338277 622917 338296 622951
rect 338330 622917 338349 622951
rect 337387 622846 337406 622880
rect 337440 622846 337459 622880
rect 337387 622823 337459 622846
rect 338277 622861 338349 622917
rect 338277 622827 338296 622861
rect 338330 622827 338349 622861
rect 338277 622823 338349 622827
rect 337387 622804 338349 622823
rect 337387 622770 337464 622804
rect 337498 622770 337554 622804
rect 337588 622770 337644 622804
rect 337678 622770 337734 622804
rect 337768 622770 337824 622804
rect 337858 622770 337914 622804
rect 337948 622770 338004 622804
rect 338038 622770 338094 622804
rect 338128 622770 338184 622804
rect 338218 622770 338349 622804
rect 337387 622751 338349 622770
rect 338675 623694 339637 623713
rect 338675 623660 338786 623694
rect 338820 623660 338876 623694
rect 338910 623660 338966 623694
rect 339000 623660 339056 623694
rect 339090 623660 339146 623694
rect 339180 623660 339236 623694
rect 339270 623660 339326 623694
rect 339360 623660 339416 623694
rect 339450 623660 339506 623694
rect 339540 623660 339637 623694
rect 338675 623641 339637 623660
rect 338675 623600 338747 623641
rect 338675 623566 338694 623600
rect 338728 623566 338747 623600
rect 339565 623581 339637 623641
rect 338675 623510 338747 623566
rect 338675 623476 338694 623510
rect 338728 623476 338747 623510
rect 338675 623420 338747 623476
rect 338675 623386 338694 623420
rect 338728 623386 338747 623420
rect 338675 623330 338747 623386
rect 338675 623296 338694 623330
rect 338728 623296 338747 623330
rect 338675 623240 338747 623296
rect 338675 623206 338694 623240
rect 338728 623206 338747 623240
rect 338675 623150 338747 623206
rect 338675 623116 338694 623150
rect 338728 623116 338747 623150
rect 338675 623060 338747 623116
rect 338675 623026 338694 623060
rect 338728 623026 338747 623060
rect 338675 622970 338747 623026
rect 338675 622936 338694 622970
rect 338728 622936 338747 622970
rect 338675 622880 338747 622936
rect 339565 623547 339584 623581
rect 339618 623547 339637 623581
rect 339565 623491 339637 623547
rect 339565 623457 339584 623491
rect 339618 623457 339637 623491
rect 339565 623401 339637 623457
rect 339565 623367 339584 623401
rect 339618 623367 339637 623401
rect 339565 623311 339637 623367
rect 339565 623277 339584 623311
rect 339618 623277 339637 623311
rect 339565 623221 339637 623277
rect 339565 623187 339584 623221
rect 339618 623187 339637 623221
rect 339565 623131 339637 623187
rect 339565 623097 339584 623131
rect 339618 623097 339637 623131
rect 339565 623041 339637 623097
rect 339565 623007 339584 623041
rect 339618 623007 339637 623041
rect 339565 622951 339637 623007
rect 339565 622917 339584 622951
rect 339618 622917 339637 622951
rect 338675 622846 338694 622880
rect 338728 622846 338747 622880
rect 338675 622823 338747 622846
rect 339565 622861 339637 622917
rect 339565 622827 339584 622861
rect 339618 622827 339637 622861
rect 339565 622823 339637 622827
rect 338675 622804 339637 622823
rect 338675 622770 338752 622804
rect 338786 622770 338842 622804
rect 338876 622770 338932 622804
rect 338966 622770 339022 622804
rect 339056 622770 339112 622804
rect 339146 622770 339202 622804
rect 339236 622770 339292 622804
rect 339326 622770 339382 622804
rect 339416 622770 339472 622804
rect 339506 622770 339637 622804
rect 338675 622751 339637 622770
rect 339963 623694 340925 623713
rect 339963 623660 340074 623694
rect 340108 623660 340164 623694
rect 340198 623660 340254 623694
rect 340288 623660 340344 623694
rect 340378 623660 340434 623694
rect 340468 623660 340524 623694
rect 340558 623660 340614 623694
rect 340648 623660 340704 623694
rect 340738 623660 340794 623694
rect 340828 623660 340925 623694
rect 339963 623641 340925 623660
rect 339963 623600 340035 623641
rect 339963 623566 339982 623600
rect 340016 623566 340035 623600
rect 340853 623581 340925 623641
rect 339963 623510 340035 623566
rect 339963 623476 339982 623510
rect 340016 623476 340035 623510
rect 339963 623420 340035 623476
rect 339963 623386 339982 623420
rect 340016 623386 340035 623420
rect 339963 623330 340035 623386
rect 339963 623296 339982 623330
rect 340016 623296 340035 623330
rect 339963 623240 340035 623296
rect 339963 623206 339982 623240
rect 340016 623206 340035 623240
rect 339963 623150 340035 623206
rect 339963 623116 339982 623150
rect 340016 623116 340035 623150
rect 339963 623060 340035 623116
rect 339963 623026 339982 623060
rect 340016 623026 340035 623060
rect 339963 622970 340035 623026
rect 339963 622936 339982 622970
rect 340016 622936 340035 622970
rect 339963 622880 340035 622936
rect 340853 623547 340872 623581
rect 340906 623547 340925 623581
rect 340853 623491 340925 623547
rect 340853 623457 340872 623491
rect 340906 623457 340925 623491
rect 340853 623401 340925 623457
rect 340853 623367 340872 623401
rect 340906 623367 340925 623401
rect 340853 623311 340925 623367
rect 340853 623277 340872 623311
rect 340906 623277 340925 623311
rect 340853 623221 340925 623277
rect 340853 623187 340872 623221
rect 340906 623187 340925 623221
rect 340853 623131 340925 623187
rect 340853 623097 340872 623131
rect 340906 623097 340925 623131
rect 340853 623041 340925 623097
rect 340853 623007 340872 623041
rect 340906 623007 340925 623041
rect 340853 622951 340925 623007
rect 340853 622917 340872 622951
rect 340906 622917 340925 622951
rect 339963 622846 339982 622880
rect 340016 622846 340035 622880
rect 339963 622823 340035 622846
rect 340853 622861 340925 622917
rect 340853 622827 340872 622861
rect 340906 622827 340925 622861
rect 340853 622823 340925 622827
rect 339963 622804 340925 622823
rect 339963 622770 340040 622804
rect 340074 622770 340130 622804
rect 340164 622770 340220 622804
rect 340254 622770 340310 622804
rect 340344 622770 340400 622804
rect 340434 622770 340490 622804
rect 340524 622770 340580 622804
rect 340614 622770 340670 622804
rect 340704 622770 340760 622804
rect 340794 622770 340925 622804
rect 339963 622751 340925 622770
rect 334811 622406 335773 622425
rect 334811 622372 334922 622406
rect 334956 622372 335012 622406
rect 335046 622372 335102 622406
rect 335136 622372 335192 622406
rect 335226 622372 335282 622406
rect 335316 622372 335372 622406
rect 335406 622372 335462 622406
rect 335496 622372 335552 622406
rect 335586 622372 335642 622406
rect 335676 622372 335773 622406
rect 334811 622353 335773 622372
rect 334811 622312 334883 622353
rect 334811 622278 334830 622312
rect 334864 622278 334883 622312
rect 335701 622293 335773 622353
rect 334811 622222 334883 622278
rect 334811 622188 334830 622222
rect 334864 622188 334883 622222
rect 334811 622132 334883 622188
rect 334811 622098 334830 622132
rect 334864 622098 334883 622132
rect 334811 622042 334883 622098
rect 334811 622008 334830 622042
rect 334864 622008 334883 622042
rect 334811 621952 334883 622008
rect 334811 621918 334830 621952
rect 334864 621918 334883 621952
rect 334811 621862 334883 621918
rect 334811 621828 334830 621862
rect 334864 621828 334883 621862
rect 334811 621772 334883 621828
rect 334811 621738 334830 621772
rect 334864 621738 334883 621772
rect 334811 621682 334883 621738
rect 334811 621648 334830 621682
rect 334864 621648 334883 621682
rect 334811 621592 334883 621648
rect 335701 622259 335720 622293
rect 335754 622259 335773 622293
rect 335701 622203 335773 622259
rect 335701 622169 335720 622203
rect 335754 622169 335773 622203
rect 335701 622113 335773 622169
rect 335701 622079 335720 622113
rect 335754 622079 335773 622113
rect 335701 622023 335773 622079
rect 335701 621989 335720 622023
rect 335754 621989 335773 622023
rect 335701 621933 335773 621989
rect 335701 621899 335720 621933
rect 335754 621899 335773 621933
rect 335701 621843 335773 621899
rect 335701 621809 335720 621843
rect 335754 621809 335773 621843
rect 335701 621753 335773 621809
rect 335701 621719 335720 621753
rect 335754 621719 335773 621753
rect 335701 621663 335773 621719
rect 335701 621629 335720 621663
rect 335754 621629 335773 621663
rect 334811 621558 334830 621592
rect 334864 621558 334883 621592
rect 334811 621535 334883 621558
rect 335701 621573 335773 621629
rect 335701 621539 335720 621573
rect 335754 621539 335773 621573
rect 335701 621535 335773 621539
rect 334811 621516 335773 621535
rect 334811 621482 334888 621516
rect 334922 621482 334978 621516
rect 335012 621482 335068 621516
rect 335102 621482 335158 621516
rect 335192 621482 335248 621516
rect 335282 621482 335338 621516
rect 335372 621482 335428 621516
rect 335462 621482 335518 621516
rect 335552 621482 335608 621516
rect 335642 621482 335773 621516
rect 334811 621463 335773 621482
rect 336099 622406 337061 622425
rect 336099 622372 336210 622406
rect 336244 622372 336300 622406
rect 336334 622372 336390 622406
rect 336424 622372 336480 622406
rect 336514 622372 336570 622406
rect 336604 622372 336660 622406
rect 336694 622372 336750 622406
rect 336784 622372 336840 622406
rect 336874 622372 336930 622406
rect 336964 622372 337061 622406
rect 336099 622353 337061 622372
rect 336099 622312 336171 622353
rect 336099 622278 336118 622312
rect 336152 622278 336171 622312
rect 336989 622293 337061 622353
rect 336099 622222 336171 622278
rect 336099 622188 336118 622222
rect 336152 622188 336171 622222
rect 336099 622132 336171 622188
rect 336099 622098 336118 622132
rect 336152 622098 336171 622132
rect 336099 622042 336171 622098
rect 336099 622008 336118 622042
rect 336152 622008 336171 622042
rect 336099 621952 336171 622008
rect 336099 621918 336118 621952
rect 336152 621918 336171 621952
rect 336099 621862 336171 621918
rect 336099 621828 336118 621862
rect 336152 621828 336171 621862
rect 336099 621772 336171 621828
rect 336099 621738 336118 621772
rect 336152 621738 336171 621772
rect 336099 621682 336171 621738
rect 336099 621648 336118 621682
rect 336152 621648 336171 621682
rect 336099 621592 336171 621648
rect 336989 622259 337008 622293
rect 337042 622259 337061 622293
rect 336989 622203 337061 622259
rect 336989 622169 337008 622203
rect 337042 622169 337061 622203
rect 336989 622113 337061 622169
rect 336989 622079 337008 622113
rect 337042 622079 337061 622113
rect 336989 622023 337061 622079
rect 336989 621989 337008 622023
rect 337042 621989 337061 622023
rect 336989 621933 337061 621989
rect 336989 621899 337008 621933
rect 337042 621899 337061 621933
rect 336989 621843 337061 621899
rect 336989 621809 337008 621843
rect 337042 621809 337061 621843
rect 336989 621753 337061 621809
rect 336989 621719 337008 621753
rect 337042 621719 337061 621753
rect 336989 621663 337061 621719
rect 336989 621629 337008 621663
rect 337042 621629 337061 621663
rect 336099 621558 336118 621592
rect 336152 621558 336171 621592
rect 336099 621535 336171 621558
rect 336989 621573 337061 621629
rect 336989 621539 337008 621573
rect 337042 621539 337061 621573
rect 336989 621535 337061 621539
rect 336099 621516 337061 621535
rect 336099 621482 336176 621516
rect 336210 621482 336266 621516
rect 336300 621482 336356 621516
rect 336390 621482 336446 621516
rect 336480 621482 336536 621516
rect 336570 621482 336626 621516
rect 336660 621482 336716 621516
rect 336750 621482 336806 621516
rect 336840 621482 336896 621516
rect 336930 621482 337061 621516
rect 336099 621463 337061 621482
rect 337387 622406 338349 622425
rect 337387 622372 337498 622406
rect 337532 622372 337588 622406
rect 337622 622372 337678 622406
rect 337712 622372 337768 622406
rect 337802 622372 337858 622406
rect 337892 622372 337948 622406
rect 337982 622372 338038 622406
rect 338072 622372 338128 622406
rect 338162 622372 338218 622406
rect 338252 622372 338349 622406
rect 337387 622353 338349 622372
rect 337387 622312 337459 622353
rect 337387 622278 337406 622312
rect 337440 622278 337459 622312
rect 338277 622293 338349 622353
rect 337387 622222 337459 622278
rect 337387 622188 337406 622222
rect 337440 622188 337459 622222
rect 337387 622132 337459 622188
rect 337387 622098 337406 622132
rect 337440 622098 337459 622132
rect 337387 622042 337459 622098
rect 337387 622008 337406 622042
rect 337440 622008 337459 622042
rect 337387 621952 337459 622008
rect 337387 621918 337406 621952
rect 337440 621918 337459 621952
rect 337387 621862 337459 621918
rect 337387 621828 337406 621862
rect 337440 621828 337459 621862
rect 337387 621772 337459 621828
rect 337387 621738 337406 621772
rect 337440 621738 337459 621772
rect 337387 621682 337459 621738
rect 337387 621648 337406 621682
rect 337440 621648 337459 621682
rect 337387 621592 337459 621648
rect 338277 622259 338296 622293
rect 338330 622259 338349 622293
rect 338277 622203 338349 622259
rect 338277 622169 338296 622203
rect 338330 622169 338349 622203
rect 338277 622113 338349 622169
rect 338277 622079 338296 622113
rect 338330 622079 338349 622113
rect 338277 622023 338349 622079
rect 338277 621989 338296 622023
rect 338330 621989 338349 622023
rect 338277 621933 338349 621989
rect 338277 621899 338296 621933
rect 338330 621899 338349 621933
rect 338277 621843 338349 621899
rect 338277 621809 338296 621843
rect 338330 621809 338349 621843
rect 338277 621753 338349 621809
rect 338277 621719 338296 621753
rect 338330 621719 338349 621753
rect 338277 621663 338349 621719
rect 338277 621629 338296 621663
rect 338330 621629 338349 621663
rect 337387 621558 337406 621592
rect 337440 621558 337459 621592
rect 337387 621535 337459 621558
rect 338277 621573 338349 621629
rect 338277 621539 338296 621573
rect 338330 621539 338349 621573
rect 338277 621535 338349 621539
rect 337387 621516 338349 621535
rect 337387 621482 337464 621516
rect 337498 621482 337554 621516
rect 337588 621482 337644 621516
rect 337678 621482 337734 621516
rect 337768 621482 337824 621516
rect 337858 621482 337914 621516
rect 337948 621482 338004 621516
rect 338038 621482 338094 621516
rect 338128 621482 338184 621516
rect 338218 621482 338349 621516
rect 337387 621463 338349 621482
rect 338675 622406 339637 622425
rect 338675 622372 338786 622406
rect 338820 622372 338876 622406
rect 338910 622372 338966 622406
rect 339000 622372 339056 622406
rect 339090 622372 339146 622406
rect 339180 622372 339236 622406
rect 339270 622372 339326 622406
rect 339360 622372 339416 622406
rect 339450 622372 339506 622406
rect 339540 622372 339637 622406
rect 338675 622353 339637 622372
rect 338675 622312 338747 622353
rect 338675 622278 338694 622312
rect 338728 622278 338747 622312
rect 339565 622293 339637 622353
rect 338675 622222 338747 622278
rect 338675 622188 338694 622222
rect 338728 622188 338747 622222
rect 338675 622132 338747 622188
rect 338675 622098 338694 622132
rect 338728 622098 338747 622132
rect 338675 622042 338747 622098
rect 338675 622008 338694 622042
rect 338728 622008 338747 622042
rect 338675 621952 338747 622008
rect 338675 621918 338694 621952
rect 338728 621918 338747 621952
rect 338675 621862 338747 621918
rect 338675 621828 338694 621862
rect 338728 621828 338747 621862
rect 338675 621772 338747 621828
rect 338675 621738 338694 621772
rect 338728 621738 338747 621772
rect 338675 621682 338747 621738
rect 338675 621648 338694 621682
rect 338728 621648 338747 621682
rect 338675 621592 338747 621648
rect 339565 622259 339584 622293
rect 339618 622259 339637 622293
rect 339565 622203 339637 622259
rect 339565 622169 339584 622203
rect 339618 622169 339637 622203
rect 339565 622113 339637 622169
rect 339565 622079 339584 622113
rect 339618 622079 339637 622113
rect 339565 622023 339637 622079
rect 339565 621989 339584 622023
rect 339618 621989 339637 622023
rect 339565 621933 339637 621989
rect 339565 621899 339584 621933
rect 339618 621899 339637 621933
rect 339565 621843 339637 621899
rect 339565 621809 339584 621843
rect 339618 621809 339637 621843
rect 339565 621753 339637 621809
rect 339565 621719 339584 621753
rect 339618 621719 339637 621753
rect 339565 621663 339637 621719
rect 339565 621629 339584 621663
rect 339618 621629 339637 621663
rect 338675 621558 338694 621592
rect 338728 621558 338747 621592
rect 338675 621535 338747 621558
rect 339565 621573 339637 621629
rect 339565 621539 339584 621573
rect 339618 621539 339637 621573
rect 339565 621535 339637 621539
rect 338675 621516 339637 621535
rect 338675 621482 338752 621516
rect 338786 621482 338842 621516
rect 338876 621482 338932 621516
rect 338966 621482 339022 621516
rect 339056 621482 339112 621516
rect 339146 621482 339202 621516
rect 339236 621482 339292 621516
rect 339326 621482 339382 621516
rect 339416 621482 339472 621516
rect 339506 621482 339637 621516
rect 338675 621463 339637 621482
rect 339963 622406 340925 622425
rect 339963 622372 340074 622406
rect 340108 622372 340164 622406
rect 340198 622372 340254 622406
rect 340288 622372 340344 622406
rect 340378 622372 340434 622406
rect 340468 622372 340524 622406
rect 340558 622372 340614 622406
rect 340648 622372 340704 622406
rect 340738 622372 340794 622406
rect 340828 622372 340925 622406
rect 339963 622353 340925 622372
rect 339963 622312 340035 622353
rect 339963 622278 339982 622312
rect 340016 622278 340035 622312
rect 340853 622293 340925 622353
rect 339963 622222 340035 622278
rect 339963 622188 339982 622222
rect 340016 622188 340035 622222
rect 339963 622132 340035 622188
rect 339963 622098 339982 622132
rect 340016 622098 340035 622132
rect 339963 622042 340035 622098
rect 339963 622008 339982 622042
rect 340016 622008 340035 622042
rect 339963 621952 340035 622008
rect 339963 621918 339982 621952
rect 340016 621918 340035 621952
rect 339963 621862 340035 621918
rect 339963 621828 339982 621862
rect 340016 621828 340035 621862
rect 339963 621772 340035 621828
rect 339963 621738 339982 621772
rect 340016 621738 340035 621772
rect 339963 621682 340035 621738
rect 339963 621648 339982 621682
rect 340016 621648 340035 621682
rect 339963 621592 340035 621648
rect 340853 622259 340872 622293
rect 340906 622259 340925 622293
rect 340853 622203 340925 622259
rect 340853 622169 340872 622203
rect 340906 622169 340925 622203
rect 340853 622113 340925 622169
rect 340853 622079 340872 622113
rect 340906 622079 340925 622113
rect 340853 622023 340925 622079
rect 340853 621989 340872 622023
rect 340906 621989 340925 622023
rect 340853 621933 340925 621989
rect 340853 621899 340872 621933
rect 340906 621899 340925 621933
rect 340853 621843 340925 621899
rect 340853 621809 340872 621843
rect 340906 621809 340925 621843
rect 340853 621753 340925 621809
rect 340853 621719 340872 621753
rect 340906 621719 340925 621753
rect 340853 621663 340925 621719
rect 340853 621629 340872 621663
rect 340906 621629 340925 621663
rect 339963 621558 339982 621592
rect 340016 621558 340035 621592
rect 339963 621535 340035 621558
rect 340853 621573 340925 621629
rect 340853 621539 340872 621573
rect 340906 621539 340925 621573
rect 340853 621535 340925 621539
rect 339963 621516 340925 621535
rect 339963 621482 340040 621516
rect 340074 621482 340130 621516
rect 340164 621482 340220 621516
rect 340254 621482 340310 621516
rect 340344 621482 340400 621516
rect 340434 621482 340490 621516
rect 340524 621482 340580 621516
rect 340614 621482 340670 621516
rect 340704 621482 340760 621516
rect 340794 621482 340925 621516
rect 339963 621463 340925 621482
rect 334811 621118 335773 621137
rect 334811 621084 334922 621118
rect 334956 621084 335012 621118
rect 335046 621084 335102 621118
rect 335136 621084 335192 621118
rect 335226 621084 335282 621118
rect 335316 621084 335372 621118
rect 335406 621084 335462 621118
rect 335496 621084 335552 621118
rect 335586 621084 335642 621118
rect 335676 621084 335773 621118
rect 334811 621065 335773 621084
rect 334811 621024 334883 621065
rect 334811 620990 334830 621024
rect 334864 620990 334883 621024
rect 335701 621005 335773 621065
rect 334811 620934 334883 620990
rect 334811 620900 334830 620934
rect 334864 620900 334883 620934
rect 334811 620844 334883 620900
rect 334811 620810 334830 620844
rect 334864 620810 334883 620844
rect 334811 620754 334883 620810
rect 334811 620720 334830 620754
rect 334864 620720 334883 620754
rect 334811 620664 334883 620720
rect 334811 620630 334830 620664
rect 334864 620630 334883 620664
rect 334811 620574 334883 620630
rect 334811 620540 334830 620574
rect 334864 620540 334883 620574
rect 334811 620484 334883 620540
rect 334811 620450 334830 620484
rect 334864 620450 334883 620484
rect 334811 620394 334883 620450
rect 334811 620360 334830 620394
rect 334864 620360 334883 620394
rect 334811 620304 334883 620360
rect 335701 620971 335720 621005
rect 335754 620971 335773 621005
rect 335701 620915 335773 620971
rect 335701 620881 335720 620915
rect 335754 620881 335773 620915
rect 335701 620825 335773 620881
rect 335701 620791 335720 620825
rect 335754 620791 335773 620825
rect 335701 620735 335773 620791
rect 335701 620701 335720 620735
rect 335754 620701 335773 620735
rect 335701 620645 335773 620701
rect 335701 620611 335720 620645
rect 335754 620611 335773 620645
rect 335701 620555 335773 620611
rect 335701 620521 335720 620555
rect 335754 620521 335773 620555
rect 335701 620465 335773 620521
rect 335701 620431 335720 620465
rect 335754 620431 335773 620465
rect 335701 620375 335773 620431
rect 335701 620341 335720 620375
rect 335754 620341 335773 620375
rect 334811 620270 334830 620304
rect 334864 620270 334883 620304
rect 334811 620247 334883 620270
rect 335701 620285 335773 620341
rect 335701 620251 335720 620285
rect 335754 620251 335773 620285
rect 335701 620247 335773 620251
rect 334811 620228 335773 620247
rect 334811 620194 334888 620228
rect 334922 620194 334978 620228
rect 335012 620194 335068 620228
rect 335102 620194 335158 620228
rect 335192 620194 335248 620228
rect 335282 620194 335338 620228
rect 335372 620194 335428 620228
rect 335462 620194 335518 620228
rect 335552 620194 335608 620228
rect 335642 620194 335773 620228
rect 334811 620175 335773 620194
rect 336099 621118 337061 621137
rect 336099 621084 336210 621118
rect 336244 621084 336300 621118
rect 336334 621084 336390 621118
rect 336424 621084 336480 621118
rect 336514 621084 336570 621118
rect 336604 621084 336660 621118
rect 336694 621084 336750 621118
rect 336784 621084 336840 621118
rect 336874 621084 336930 621118
rect 336964 621084 337061 621118
rect 336099 621065 337061 621084
rect 336099 621024 336171 621065
rect 336099 620990 336118 621024
rect 336152 620990 336171 621024
rect 336989 621005 337061 621065
rect 336099 620934 336171 620990
rect 336099 620900 336118 620934
rect 336152 620900 336171 620934
rect 336099 620844 336171 620900
rect 336099 620810 336118 620844
rect 336152 620810 336171 620844
rect 336099 620754 336171 620810
rect 336099 620720 336118 620754
rect 336152 620720 336171 620754
rect 336099 620664 336171 620720
rect 336099 620630 336118 620664
rect 336152 620630 336171 620664
rect 336099 620574 336171 620630
rect 336099 620540 336118 620574
rect 336152 620540 336171 620574
rect 336099 620484 336171 620540
rect 336099 620450 336118 620484
rect 336152 620450 336171 620484
rect 336099 620394 336171 620450
rect 336099 620360 336118 620394
rect 336152 620360 336171 620394
rect 336099 620304 336171 620360
rect 336989 620971 337008 621005
rect 337042 620971 337061 621005
rect 336989 620915 337061 620971
rect 336989 620881 337008 620915
rect 337042 620881 337061 620915
rect 336989 620825 337061 620881
rect 336989 620791 337008 620825
rect 337042 620791 337061 620825
rect 336989 620735 337061 620791
rect 336989 620701 337008 620735
rect 337042 620701 337061 620735
rect 336989 620645 337061 620701
rect 336989 620611 337008 620645
rect 337042 620611 337061 620645
rect 336989 620555 337061 620611
rect 336989 620521 337008 620555
rect 337042 620521 337061 620555
rect 336989 620465 337061 620521
rect 336989 620431 337008 620465
rect 337042 620431 337061 620465
rect 336989 620375 337061 620431
rect 336989 620341 337008 620375
rect 337042 620341 337061 620375
rect 336099 620270 336118 620304
rect 336152 620270 336171 620304
rect 336099 620247 336171 620270
rect 336989 620285 337061 620341
rect 336989 620251 337008 620285
rect 337042 620251 337061 620285
rect 336989 620247 337061 620251
rect 336099 620228 337061 620247
rect 336099 620194 336176 620228
rect 336210 620194 336266 620228
rect 336300 620194 336356 620228
rect 336390 620194 336446 620228
rect 336480 620194 336536 620228
rect 336570 620194 336626 620228
rect 336660 620194 336716 620228
rect 336750 620194 336806 620228
rect 336840 620194 336896 620228
rect 336930 620194 337061 620228
rect 336099 620175 337061 620194
rect 337387 621118 338349 621137
rect 337387 621084 337498 621118
rect 337532 621084 337588 621118
rect 337622 621084 337678 621118
rect 337712 621084 337768 621118
rect 337802 621084 337858 621118
rect 337892 621084 337948 621118
rect 337982 621084 338038 621118
rect 338072 621084 338128 621118
rect 338162 621084 338218 621118
rect 338252 621084 338349 621118
rect 337387 621065 338349 621084
rect 337387 621024 337459 621065
rect 337387 620990 337406 621024
rect 337440 620990 337459 621024
rect 338277 621005 338349 621065
rect 337387 620934 337459 620990
rect 337387 620900 337406 620934
rect 337440 620900 337459 620934
rect 337387 620844 337459 620900
rect 337387 620810 337406 620844
rect 337440 620810 337459 620844
rect 337387 620754 337459 620810
rect 337387 620720 337406 620754
rect 337440 620720 337459 620754
rect 337387 620664 337459 620720
rect 337387 620630 337406 620664
rect 337440 620630 337459 620664
rect 337387 620574 337459 620630
rect 337387 620540 337406 620574
rect 337440 620540 337459 620574
rect 337387 620484 337459 620540
rect 337387 620450 337406 620484
rect 337440 620450 337459 620484
rect 337387 620394 337459 620450
rect 337387 620360 337406 620394
rect 337440 620360 337459 620394
rect 337387 620304 337459 620360
rect 338277 620971 338296 621005
rect 338330 620971 338349 621005
rect 338277 620915 338349 620971
rect 338277 620881 338296 620915
rect 338330 620881 338349 620915
rect 338277 620825 338349 620881
rect 338277 620791 338296 620825
rect 338330 620791 338349 620825
rect 338277 620735 338349 620791
rect 338277 620701 338296 620735
rect 338330 620701 338349 620735
rect 338277 620645 338349 620701
rect 338277 620611 338296 620645
rect 338330 620611 338349 620645
rect 338277 620555 338349 620611
rect 338277 620521 338296 620555
rect 338330 620521 338349 620555
rect 338277 620465 338349 620521
rect 338277 620431 338296 620465
rect 338330 620431 338349 620465
rect 338277 620375 338349 620431
rect 338277 620341 338296 620375
rect 338330 620341 338349 620375
rect 337387 620270 337406 620304
rect 337440 620270 337459 620304
rect 337387 620247 337459 620270
rect 338277 620285 338349 620341
rect 338277 620251 338296 620285
rect 338330 620251 338349 620285
rect 338277 620247 338349 620251
rect 337387 620228 338349 620247
rect 337387 620194 337464 620228
rect 337498 620194 337554 620228
rect 337588 620194 337644 620228
rect 337678 620194 337734 620228
rect 337768 620194 337824 620228
rect 337858 620194 337914 620228
rect 337948 620194 338004 620228
rect 338038 620194 338094 620228
rect 338128 620194 338184 620228
rect 338218 620194 338349 620228
rect 337387 620175 338349 620194
rect 338675 621118 339637 621137
rect 338675 621084 338786 621118
rect 338820 621084 338876 621118
rect 338910 621084 338966 621118
rect 339000 621084 339056 621118
rect 339090 621084 339146 621118
rect 339180 621084 339236 621118
rect 339270 621084 339326 621118
rect 339360 621084 339416 621118
rect 339450 621084 339506 621118
rect 339540 621084 339637 621118
rect 338675 621065 339637 621084
rect 338675 621024 338747 621065
rect 338675 620990 338694 621024
rect 338728 620990 338747 621024
rect 339565 621005 339637 621065
rect 338675 620934 338747 620990
rect 338675 620900 338694 620934
rect 338728 620900 338747 620934
rect 338675 620844 338747 620900
rect 338675 620810 338694 620844
rect 338728 620810 338747 620844
rect 338675 620754 338747 620810
rect 338675 620720 338694 620754
rect 338728 620720 338747 620754
rect 338675 620664 338747 620720
rect 338675 620630 338694 620664
rect 338728 620630 338747 620664
rect 338675 620574 338747 620630
rect 338675 620540 338694 620574
rect 338728 620540 338747 620574
rect 338675 620484 338747 620540
rect 338675 620450 338694 620484
rect 338728 620450 338747 620484
rect 338675 620394 338747 620450
rect 338675 620360 338694 620394
rect 338728 620360 338747 620394
rect 338675 620304 338747 620360
rect 339565 620971 339584 621005
rect 339618 620971 339637 621005
rect 339565 620915 339637 620971
rect 339565 620881 339584 620915
rect 339618 620881 339637 620915
rect 339565 620825 339637 620881
rect 339565 620791 339584 620825
rect 339618 620791 339637 620825
rect 339565 620735 339637 620791
rect 339565 620701 339584 620735
rect 339618 620701 339637 620735
rect 339565 620645 339637 620701
rect 339565 620611 339584 620645
rect 339618 620611 339637 620645
rect 339565 620555 339637 620611
rect 339565 620521 339584 620555
rect 339618 620521 339637 620555
rect 339565 620465 339637 620521
rect 339565 620431 339584 620465
rect 339618 620431 339637 620465
rect 339565 620375 339637 620431
rect 339565 620341 339584 620375
rect 339618 620341 339637 620375
rect 338675 620270 338694 620304
rect 338728 620270 338747 620304
rect 338675 620247 338747 620270
rect 339565 620285 339637 620341
rect 339565 620251 339584 620285
rect 339618 620251 339637 620285
rect 339565 620247 339637 620251
rect 338675 620228 339637 620247
rect 338675 620194 338752 620228
rect 338786 620194 338842 620228
rect 338876 620194 338932 620228
rect 338966 620194 339022 620228
rect 339056 620194 339112 620228
rect 339146 620194 339202 620228
rect 339236 620194 339292 620228
rect 339326 620194 339382 620228
rect 339416 620194 339472 620228
rect 339506 620194 339637 620228
rect 338675 620175 339637 620194
rect 339963 621118 340925 621137
rect 339963 621084 340074 621118
rect 340108 621084 340164 621118
rect 340198 621084 340254 621118
rect 340288 621084 340344 621118
rect 340378 621084 340434 621118
rect 340468 621084 340524 621118
rect 340558 621084 340614 621118
rect 340648 621084 340704 621118
rect 340738 621084 340794 621118
rect 340828 621084 340925 621118
rect 339963 621065 340925 621084
rect 339963 621024 340035 621065
rect 339963 620990 339982 621024
rect 340016 620990 340035 621024
rect 340853 621005 340925 621065
rect 339963 620934 340035 620990
rect 339963 620900 339982 620934
rect 340016 620900 340035 620934
rect 339963 620844 340035 620900
rect 339963 620810 339982 620844
rect 340016 620810 340035 620844
rect 339963 620754 340035 620810
rect 339963 620720 339982 620754
rect 340016 620720 340035 620754
rect 339963 620664 340035 620720
rect 339963 620630 339982 620664
rect 340016 620630 340035 620664
rect 339963 620574 340035 620630
rect 339963 620540 339982 620574
rect 340016 620540 340035 620574
rect 339963 620484 340035 620540
rect 339963 620450 339982 620484
rect 340016 620450 340035 620484
rect 339963 620394 340035 620450
rect 339963 620360 339982 620394
rect 340016 620360 340035 620394
rect 339963 620304 340035 620360
rect 340853 620971 340872 621005
rect 340906 620971 340925 621005
rect 340853 620915 340925 620971
rect 340853 620881 340872 620915
rect 340906 620881 340925 620915
rect 340853 620825 340925 620881
rect 340853 620791 340872 620825
rect 340906 620791 340925 620825
rect 340853 620735 340925 620791
rect 340853 620701 340872 620735
rect 340906 620701 340925 620735
rect 340853 620645 340925 620701
rect 340853 620611 340872 620645
rect 340906 620611 340925 620645
rect 340853 620555 340925 620611
rect 340853 620521 340872 620555
rect 340906 620521 340925 620555
rect 340853 620465 340925 620521
rect 340853 620431 340872 620465
rect 340906 620431 340925 620465
rect 340853 620375 340925 620431
rect 340853 620341 340872 620375
rect 340906 620341 340925 620375
rect 339963 620270 339982 620304
rect 340016 620270 340035 620304
rect 339963 620247 340035 620270
rect 340853 620285 340925 620341
rect 340853 620251 340872 620285
rect 340906 620251 340925 620285
rect 340853 620247 340925 620251
rect 339963 620228 340925 620247
rect 339963 620194 340040 620228
rect 340074 620194 340130 620228
rect 340164 620194 340220 620228
rect 340254 620194 340310 620228
rect 340344 620194 340400 620228
rect 340434 620194 340490 620228
rect 340524 620194 340580 620228
rect 340614 620194 340670 620228
rect 340704 620194 340760 620228
rect 340794 620194 340925 620228
rect 339963 620175 340925 620194
rect 334811 619830 335773 619849
rect 334811 619796 334922 619830
rect 334956 619796 335012 619830
rect 335046 619796 335102 619830
rect 335136 619796 335192 619830
rect 335226 619796 335282 619830
rect 335316 619796 335372 619830
rect 335406 619796 335462 619830
rect 335496 619796 335552 619830
rect 335586 619796 335642 619830
rect 335676 619796 335773 619830
rect 334811 619777 335773 619796
rect 334811 619736 334883 619777
rect 334811 619702 334830 619736
rect 334864 619702 334883 619736
rect 335701 619717 335773 619777
rect 334811 619646 334883 619702
rect 334811 619612 334830 619646
rect 334864 619612 334883 619646
rect 334811 619556 334883 619612
rect 334811 619522 334830 619556
rect 334864 619522 334883 619556
rect 334811 619466 334883 619522
rect 334811 619432 334830 619466
rect 334864 619432 334883 619466
rect 334811 619376 334883 619432
rect 334811 619342 334830 619376
rect 334864 619342 334883 619376
rect 334811 619286 334883 619342
rect 334811 619252 334830 619286
rect 334864 619252 334883 619286
rect 334811 619196 334883 619252
rect 334811 619162 334830 619196
rect 334864 619162 334883 619196
rect 334811 619106 334883 619162
rect 334811 619072 334830 619106
rect 334864 619072 334883 619106
rect 334811 619016 334883 619072
rect 335701 619683 335720 619717
rect 335754 619683 335773 619717
rect 335701 619627 335773 619683
rect 335701 619593 335720 619627
rect 335754 619593 335773 619627
rect 335701 619537 335773 619593
rect 335701 619503 335720 619537
rect 335754 619503 335773 619537
rect 335701 619447 335773 619503
rect 335701 619413 335720 619447
rect 335754 619413 335773 619447
rect 335701 619357 335773 619413
rect 335701 619323 335720 619357
rect 335754 619323 335773 619357
rect 335701 619267 335773 619323
rect 335701 619233 335720 619267
rect 335754 619233 335773 619267
rect 335701 619177 335773 619233
rect 335701 619143 335720 619177
rect 335754 619143 335773 619177
rect 335701 619087 335773 619143
rect 335701 619053 335720 619087
rect 335754 619053 335773 619087
rect 334811 618982 334830 619016
rect 334864 618982 334883 619016
rect 334811 618959 334883 618982
rect 335701 618997 335773 619053
rect 335701 618963 335720 618997
rect 335754 618963 335773 618997
rect 335701 618959 335773 618963
rect 334811 618940 335773 618959
rect 334811 618906 334888 618940
rect 334922 618906 334978 618940
rect 335012 618906 335068 618940
rect 335102 618906 335158 618940
rect 335192 618906 335248 618940
rect 335282 618906 335338 618940
rect 335372 618906 335428 618940
rect 335462 618906 335518 618940
rect 335552 618906 335608 618940
rect 335642 618906 335773 618940
rect 334811 618887 335773 618906
rect 336099 619830 337061 619849
rect 336099 619796 336210 619830
rect 336244 619796 336300 619830
rect 336334 619796 336390 619830
rect 336424 619796 336480 619830
rect 336514 619796 336570 619830
rect 336604 619796 336660 619830
rect 336694 619796 336750 619830
rect 336784 619796 336840 619830
rect 336874 619796 336930 619830
rect 336964 619796 337061 619830
rect 336099 619777 337061 619796
rect 336099 619736 336171 619777
rect 336099 619702 336118 619736
rect 336152 619702 336171 619736
rect 336989 619717 337061 619777
rect 336099 619646 336171 619702
rect 336099 619612 336118 619646
rect 336152 619612 336171 619646
rect 336099 619556 336171 619612
rect 336099 619522 336118 619556
rect 336152 619522 336171 619556
rect 336099 619466 336171 619522
rect 336099 619432 336118 619466
rect 336152 619432 336171 619466
rect 336099 619376 336171 619432
rect 336099 619342 336118 619376
rect 336152 619342 336171 619376
rect 336099 619286 336171 619342
rect 336099 619252 336118 619286
rect 336152 619252 336171 619286
rect 336099 619196 336171 619252
rect 336099 619162 336118 619196
rect 336152 619162 336171 619196
rect 336099 619106 336171 619162
rect 336099 619072 336118 619106
rect 336152 619072 336171 619106
rect 336099 619016 336171 619072
rect 336989 619683 337008 619717
rect 337042 619683 337061 619717
rect 336989 619627 337061 619683
rect 336989 619593 337008 619627
rect 337042 619593 337061 619627
rect 336989 619537 337061 619593
rect 336989 619503 337008 619537
rect 337042 619503 337061 619537
rect 336989 619447 337061 619503
rect 336989 619413 337008 619447
rect 337042 619413 337061 619447
rect 336989 619357 337061 619413
rect 336989 619323 337008 619357
rect 337042 619323 337061 619357
rect 336989 619267 337061 619323
rect 336989 619233 337008 619267
rect 337042 619233 337061 619267
rect 336989 619177 337061 619233
rect 336989 619143 337008 619177
rect 337042 619143 337061 619177
rect 336989 619087 337061 619143
rect 336989 619053 337008 619087
rect 337042 619053 337061 619087
rect 336099 618982 336118 619016
rect 336152 618982 336171 619016
rect 336099 618959 336171 618982
rect 336989 618997 337061 619053
rect 336989 618963 337008 618997
rect 337042 618963 337061 618997
rect 336989 618959 337061 618963
rect 336099 618940 337061 618959
rect 336099 618906 336176 618940
rect 336210 618906 336266 618940
rect 336300 618906 336356 618940
rect 336390 618906 336446 618940
rect 336480 618906 336536 618940
rect 336570 618906 336626 618940
rect 336660 618906 336716 618940
rect 336750 618906 336806 618940
rect 336840 618906 336896 618940
rect 336930 618906 337061 618940
rect 336099 618887 337061 618906
rect 337387 619830 338349 619849
rect 337387 619796 337498 619830
rect 337532 619796 337588 619830
rect 337622 619796 337678 619830
rect 337712 619796 337768 619830
rect 337802 619796 337858 619830
rect 337892 619796 337948 619830
rect 337982 619796 338038 619830
rect 338072 619796 338128 619830
rect 338162 619796 338218 619830
rect 338252 619796 338349 619830
rect 337387 619777 338349 619796
rect 337387 619736 337459 619777
rect 337387 619702 337406 619736
rect 337440 619702 337459 619736
rect 338277 619717 338349 619777
rect 337387 619646 337459 619702
rect 337387 619612 337406 619646
rect 337440 619612 337459 619646
rect 337387 619556 337459 619612
rect 337387 619522 337406 619556
rect 337440 619522 337459 619556
rect 337387 619466 337459 619522
rect 337387 619432 337406 619466
rect 337440 619432 337459 619466
rect 337387 619376 337459 619432
rect 337387 619342 337406 619376
rect 337440 619342 337459 619376
rect 337387 619286 337459 619342
rect 337387 619252 337406 619286
rect 337440 619252 337459 619286
rect 337387 619196 337459 619252
rect 337387 619162 337406 619196
rect 337440 619162 337459 619196
rect 337387 619106 337459 619162
rect 337387 619072 337406 619106
rect 337440 619072 337459 619106
rect 337387 619016 337459 619072
rect 338277 619683 338296 619717
rect 338330 619683 338349 619717
rect 338277 619627 338349 619683
rect 338277 619593 338296 619627
rect 338330 619593 338349 619627
rect 338277 619537 338349 619593
rect 338277 619503 338296 619537
rect 338330 619503 338349 619537
rect 338277 619447 338349 619503
rect 338277 619413 338296 619447
rect 338330 619413 338349 619447
rect 338277 619357 338349 619413
rect 338277 619323 338296 619357
rect 338330 619323 338349 619357
rect 338277 619267 338349 619323
rect 338277 619233 338296 619267
rect 338330 619233 338349 619267
rect 338277 619177 338349 619233
rect 338277 619143 338296 619177
rect 338330 619143 338349 619177
rect 338277 619087 338349 619143
rect 338277 619053 338296 619087
rect 338330 619053 338349 619087
rect 337387 618982 337406 619016
rect 337440 618982 337459 619016
rect 337387 618959 337459 618982
rect 338277 618997 338349 619053
rect 338277 618963 338296 618997
rect 338330 618963 338349 618997
rect 338277 618959 338349 618963
rect 337387 618940 338349 618959
rect 337387 618906 337464 618940
rect 337498 618906 337554 618940
rect 337588 618906 337644 618940
rect 337678 618906 337734 618940
rect 337768 618906 337824 618940
rect 337858 618906 337914 618940
rect 337948 618906 338004 618940
rect 338038 618906 338094 618940
rect 338128 618906 338184 618940
rect 338218 618906 338349 618940
rect 337387 618887 338349 618906
rect 338675 619830 339637 619849
rect 338675 619796 338786 619830
rect 338820 619796 338876 619830
rect 338910 619796 338966 619830
rect 339000 619796 339056 619830
rect 339090 619796 339146 619830
rect 339180 619796 339236 619830
rect 339270 619796 339326 619830
rect 339360 619796 339416 619830
rect 339450 619796 339506 619830
rect 339540 619796 339637 619830
rect 338675 619777 339637 619796
rect 338675 619736 338747 619777
rect 338675 619702 338694 619736
rect 338728 619702 338747 619736
rect 339565 619717 339637 619777
rect 338675 619646 338747 619702
rect 338675 619612 338694 619646
rect 338728 619612 338747 619646
rect 338675 619556 338747 619612
rect 338675 619522 338694 619556
rect 338728 619522 338747 619556
rect 338675 619466 338747 619522
rect 338675 619432 338694 619466
rect 338728 619432 338747 619466
rect 338675 619376 338747 619432
rect 338675 619342 338694 619376
rect 338728 619342 338747 619376
rect 338675 619286 338747 619342
rect 338675 619252 338694 619286
rect 338728 619252 338747 619286
rect 338675 619196 338747 619252
rect 338675 619162 338694 619196
rect 338728 619162 338747 619196
rect 338675 619106 338747 619162
rect 338675 619072 338694 619106
rect 338728 619072 338747 619106
rect 338675 619016 338747 619072
rect 339565 619683 339584 619717
rect 339618 619683 339637 619717
rect 339565 619627 339637 619683
rect 339565 619593 339584 619627
rect 339618 619593 339637 619627
rect 339565 619537 339637 619593
rect 339565 619503 339584 619537
rect 339618 619503 339637 619537
rect 339565 619447 339637 619503
rect 339565 619413 339584 619447
rect 339618 619413 339637 619447
rect 339565 619357 339637 619413
rect 339565 619323 339584 619357
rect 339618 619323 339637 619357
rect 339565 619267 339637 619323
rect 339565 619233 339584 619267
rect 339618 619233 339637 619267
rect 339565 619177 339637 619233
rect 339565 619143 339584 619177
rect 339618 619143 339637 619177
rect 339565 619087 339637 619143
rect 339565 619053 339584 619087
rect 339618 619053 339637 619087
rect 338675 618982 338694 619016
rect 338728 618982 338747 619016
rect 338675 618959 338747 618982
rect 339565 618997 339637 619053
rect 339565 618963 339584 618997
rect 339618 618963 339637 618997
rect 339565 618959 339637 618963
rect 338675 618940 339637 618959
rect 338675 618906 338752 618940
rect 338786 618906 338842 618940
rect 338876 618906 338932 618940
rect 338966 618906 339022 618940
rect 339056 618906 339112 618940
rect 339146 618906 339202 618940
rect 339236 618906 339292 618940
rect 339326 618906 339382 618940
rect 339416 618906 339472 618940
rect 339506 618906 339637 618940
rect 338675 618887 339637 618906
rect 339963 619830 340925 619849
rect 339963 619796 340074 619830
rect 340108 619796 340164 619830
rect 340198 619796 340254 619830
rect 340288 619796 340344 619830
rect 340378 619796 340434 619830
rect 340468 619796 340524 619830
rect 340558 619796 340614 619830
rect 340648 619796 340704 619830
rect 340738 619796 340794 619830
rect 340828 619796 340925 619830
rect 339963 619777 340925 619796
rect 339963 619736 340035 619777
rect 339963 619702 339982 619736
rect 340016 619702 340035 619736
rect 340853 619717 340925 619777
rect 339963 619646 340035 619702
rect 339963 619612 339982 619646
rect 340016 619612 340035 619646
rect 339963 619556 340035 619612
rect 339963 619522 339982 619556
rect 340016 619522 340035 619556
rect 339963 619466 340035 619522
rect 339963 619432 339982 619466
rect 340016 619432 340035 619466
rect 339963 619376 340035 619432
rect 339963 619342 339982 619376
rect 340016 619342 340035 619376
rect 339963 619286 340035 619342
rect 339963 619252 339982 619286
rect 340016 619252 340035 619286
rect 339963 619196 340035 619252
rect 339963 619162 339982 619196
rect 340016 619162 340035 619196
rect 339963 619106 340035 619162
rect 339963 619072 339982 619106
rect 340016 619072 340035 619106
rect 339963 619016 340035 619072
rect 340853 619683 340872 619717
rect 340906 619683 340925 619717
rect 340853 619627 340925 619683
rect 340853 619593 340872 619627
rect 340906 619593 340925 619627
rect 340853 619537 340925 619593
rect 340853 619503 340872 619537
rect 340906 619503 340925 619537
rect 340853 619447 340925 619503
rect 340853 619413 340872 619447
rect 340906 619413 340925 619447
rect 340853 619357 340925 619413
rect 340853 619323 340872 619357
rect 340906 619323 340925 619357
rect 340853 619267 340925 619323
rect 340853 619233 340872 619267
rect 340906 619233 340925 619267
rect 340853 619177 340925 619233
rect 340853 619143 340872 619177
rect 340906 619143 340925 619177
rect 340853 619087 340925 619143
rect 340853 619053 340872 619087
rect 340906 619053 340925 619087
rect 339963 618982 339982 619016
rect 340016 618982 340035 619016
rect 339963 618959 340035 618982
rect 340853 618997 340925 619053
rect 340853 618963 340872 618997
rect 340906 618963 340925 618997
rect 340853 618959 340925 618963
rect 339963 618940 340925 618959
rect 339963 618906 340040 618940
rect 340074 618906 340130 618940
rect 340164 618906 340220 618940
rect 340254 618906 340310 618940
rect 340344 618906 340400 618940
rect 340434 618906 340490 618940
rect 340524 618906 340580 618940
rect 340614 618906 340670 618940
rect 340704 618906 340760 618940
rect 340794 618906 340925 618940
rect 339963 618887 340925 618906
rect 334811 618542 335773 618561
rect 334811 618508 334922 618542
rect 334956 618508 335012 618542
rect 335046 618508 335102 618542
rect 335136 618508 335192 618542
rect 335226 618508 335282 618542
rect 335316 618508 335372 618542
rect 335406 618508 335462 618542
rect 335496 618508 335552 618542
rect 335586 618508 335642 618542
rect 335676 618508 335773 618542
rect 334811 618489 335773 618508
rect 334811 618448 334883 618489
rect 334811 618414 334830 618448
rect 334864 618414 334883 618448
rect 335701 618429 335773 618489
rect 334811 618358 334883 618414
rect 334811 618324 334830 618358
rect 334864 618324 334883 618358
rect 334811 618268 334883 618324
rect 334811 618234 334830 618268
rect 334864 618234 334883 618268
rect 334811 618178 334883 618234
rect 334811 618144 334830 618178
rect 334864 618144 334883 618178
rect 334811 618088 334883 618144
rect 334811 618054 334830 618088
rect 334864 618054 334883 618088
rect 334811 617998 334883 618054
rect 334811 617964 334830 617998
rect 334864 617964 334883 617998
rect 334811 617908 334883 617964
rect 334811 617874 334830 617908
rect 334864 617874 334883 617908
rect 334811 617818 334883 617874
rect 334811 617784 334830 617818
rect 334864 617784 334883 617818
rect 334811 617728 334883 617784
rect 335701 618395 335720 618429
rect 335754 618395 335773 618429
rect 335701 618339 335773 618395
rect 335701 618305 335720 618339
rect 335754 618305 335773 618339
rect 335701 618249 335773 618305
rect 335701 618215 335720 618249
rect 335754 618215 335773 618249
rect 335701 618159 335773 618215
rect 335701 618125 335720 618159
rect 335754 618125 335773 618159
rect 335701 618069 335773 618125
rect 335701 618035 335720 618069
rect 335754 618035 335773 618069
rect 335701 617979 335773 618035
rect 335701 617945 335720 617979
rect 335754 617945 335773 617979
rect 335701 617889 335773 617945
rect 335701 617855 335720 617889
rect 335754 617855 335773 617889
rect 335701 617799 335773 617855
rect 335701 617765 335720 617799
rect 335754 617765 335773 617799
rect 334811 617694 334830 617728
rect 334864 617694 334883 617728
rect 334811 617671 334883 617694
rect 335701 617709 335773 617765
rect 335701 617675 335720 617709
rect 335754 617675 335773 617709
rect 335701 617671 335773 617675
rect 334811 617652 335773 617671
rect 334811 617618 334888 617652
rect 334922 617618 334978 617652
rect 335012 617618 335068 617652
rect 335102 617618 335158 617652
rect 335192 617618 335248 617652
rect 335282 617618 335338 617652
rect 335372 617618 335428 617652
rect 335462 617618 335518 617652
rect 335552 617618 335608 617652
rect 335642 617618 335773 617652
rect 334811 617599 335773 617618
rect 336099 618542 337061 618561
rect 336099 618508 336210 618542
rect 336244 618508 336300 618542
rect 336334 618508 336390 618542
rect 336424 618508 336480 618542
rect 336514 618508 336570 618542
rect 336604 618508 336660 618542
rect 336694 618508 336750 618542
rect 336784 618508 336840 618542
rect 336874 618508 336930 618542
rect 336964 618508 337061 618542
rect 336099 618489 337061 618508
rect 336099 618448 336171 618489
rect 336099 618414 336118 618448
rect 336152 618414 336171 618448
rect 336989 618429 337061 618489
rect 336099 618358 336171 618414
rect 336099 618324 336118 618358
rect 336152 618324 336171 618358
rect 336099 618268 336171 618324
rect 336099 618234 336118 618268
rect 336152 618234 336171 618268
rect 336099 618178 336171 618234
rect 336099 618144 336118 618178
rect 336152 618144 336171 618178
rect 336099 618088 336171 618144
rect 336099 618054 336118 618088
rect 336152 618054 336171 618088
rect 336099 617998 336171 618054
rect 336099 617964 336118 617998
rect 336152 617964 336171 617998
rect 336099 617908 336171 617964
rect 336099 617874 336118 617908
rect 336152 617874 336171 617908
rect 336099 617818 336171 617874
rect 336099 617784 336118 617818
rect 336152 617784 336171 617818
rect 336099 617728 336171 617784
rect 336989 618395 337008 618429
rect 337042 618395 337061 618429
rect 336989 618339 337061 618395
rect 336989 618305 337008 618339
rect 337042 618305 337061 618339
rect 336989 618249 337061 618305
rect 336989 618215 337008 618249
rect 337042 618215 337061 618249
rect 336989 618159 337061 618215
rect 336989 618125 337008 618159
rect 337042 618125 337061 618159
rect 336989 618069 337061 618125
rect 336989 618035 337008 618069
rect 337042 618035 337061 618069
rect 336989 617979 337061 618035
rect 336989 617945 337008 617979
rect 337042 617945 337061 617979
rect 336989 617889 337061 617945
rect 336989 617855 337008 617889
rect 337042 617855 337061 617889
rect 336989 617799 337061 617855
rect 336989 617765 337008 617799
rect 337042 617765 337061 617799
rect 336099 617694 336118 617728
rect 336152 617694 336171 617728
rect 336099 617671 336171 617694
rect 336989 617709 337061 617765
rect 336989 617675 337008 617709
rect 337042 617675 337061 617709
rect 336989 617671 337061 617675
rect 336099 617652 337061 617671
rect 336099 617618 336176 617652
rect 336210 617618 336266 617652
rect 336300 617618 336356 617652
rect 336390 617618 336446 617652
rect 336480 617618 336536 617652
rect 336570 617618 336626 617652
rect 336660 617618 336716 617652
rect 336750 617618 336806 617652
rect 336840 617618 336896 617652
rect 336930 617618 337061 617652
rect 336099 617599 337061 617618
rect 337387 618542 338349 618561
rect 337387 618508 337498 618542
rect 337532 618508 337588 618542
rect 337622 618508 337678 618542
rect 337712 618508 337768 618542
rect 337802 618508 337858 618542
rect 337892 618508 337948 618542
rect 337982 618508 338038 618542
rect 338072 618508 338128 618542
rect 338162 618508 338218 618542
rect 338252 618508 338349 618542
rect 337387 618489 338349 618508
rect 337387 618448 337459 618489
rect 337387 618414 337406 618448
rect 337440 618414 337459 618448
rect 338277 618429 338349 618489
rect 337387 618358 337459 618414
rect 337387 618324 337406 618358
rect 337440 618324 337459 618358
rect 337387 618268 337459 618324
rect 337387 618234 337406 618268
rect 337440 618234 337459 618268
rect 337387 618178 337459 618234
rect 337387 618144 337406 618178
rect 337440 618144 337459 618178
rect 337387 618088 337459 618144
rect 337387 618054 337406 618088
rect 337440 618054 337459 618088
rect 337387 617998 337459 618054
rect 337387 617964 337406 617998
rect 337440 617964 337459 617998
rect 337387 617908 337459 617964
rect 337387 617874 337406 617908
rect 337440 617874 337459 617908
rect 337387 617818 337459 617874
rect 337387 617784 337406 617818
rect 337440 617784 337459 617818
rect 337387 617728 337459 617784
rect 338277 618395 338296 618429
rect 338330 618395 338349 618429
rect 338277 618339 338349 618395
rect 338277 618305 338296 618339
rect 338330 618305 338349 618339
rect 338277 618249 338349 618305
rect 338277 618215 338296 618249
rect 338330 618215 338349 618249
rect 338277 618159 338349 618215
rect 338277 618125 338296 618159
rect 338330 618125 338349 618159
rect 338277 618069 338349 618125
rect 338277 618035 338296 618069
rect 338330 618035 338349 618069
rect 338277 617979 338349 618035
rect 338277 617945 338296 617979
rect 338330 617945 338349 617979
rect 338277 617889 338349 617945
rect 338277 617855 338296 617889
rect 338330 617855 338349 617889
rect 338277 617799 338349 617855
rect 338277 617765 338296 617799
rect 338330 617765 338349 617799
rect 337387 617694 337406 617728
rect 337440 617694 337459 617728
rect 337387 617671 337459 617694
rect 338277 617709 338349 617765
rect 338277 617675 338296 617709
rect 338330 617675 338349 617709
rect 338277 617671 338349 617675
rect 337387 617652 338349 617671
rect 337387 617618 337464 617652
rect 337498 617618 337554 617652
rect 337588 617618 337644 617652
rect 337678 617618 337734 617652
rect 337768 617618 337824 617652
rect 337858 617618 337914 617652
rect 337948 617618 338004 617652
rect 338038 617618 338094 617652
rect 338128 617618 338184 617652
rect 338218 617618 338349 617652
rect 337387 617599 338349 617618
rect 338675 618542 339637 618561
rect 338675 618508 338786 618542
rect 338820 618508 338876 618542
rect 338910 618508 338966 618542
rect 339000 618508 339056 618542
rect 339090 618508 339146 618542
rect 339180 618508 339236 618542
rect 339270 618508 339326 618542
rect 339360 618508 339416 618542
rect 339450 618508 339506 618542
rect 339540 618508 339637 618542
rect 338675 618489 339637 618508
rect 338675 618448 338747 618489
rect 338675 618414 338694 618448
rect 338728 618414 338747 618448
rect 339565 618429 339637 618489
rect 338675 618358 338747 618414
rect 338675 618324 338694 618358
rect 338728 618324 338747 618358
rect 338675 618268 338747 618324
rect 338675 618234 338694 618268
rect 338728 618234 338747 618268
rect 338675 618178 338747 618234
rect 338675 618144 338694 618178
rect 338728 618144 338747 618178
rect 338675 618088 338747 618144
rect 338675 618054 338694 618088
rect 338728 618054 338747 618088
rect 338675 617998 338747 618054
rect 338675 617964 338694 617998
rect 338728 617964 338747 617998
rect 338675 617908 338747 617964
rect 338675 617874 338694 617908
rect 338728 617874 338747 617908
rect 338675 617818 338747 617874
rect 338675 617784 338694 617818
rect 338728 617784 338747 617818
rect 338675 617728 338747 617784
rect 339565 618395 339584 618429
rect 339618 618395 339637 618429
rect 339565 618339 339637 618395
rect 339565 618305 339584 618339
rect 339618 618305 339637 618339
rect 339565 618249 339637 618305
rect 339565 618215 339584 618249
rect 339618 618215 339637 618249
rect 339565 618159 339637 618215
rect 339565 618125 339584 618159
rect 339618 618125 339637 618159
rect 339565 618069 339637 618125
rect 339565 618035 339584 618069
rect 339618 618035 339637 618069
rect 339565 617979 339637 618035
rect 339565 617945 339584 617979
rect 339618 617945 339637 617979
rect 339565 617889 339637 617945
rect 339565 617855 339584 617889
rect 339618 617855 339637 617889
rect 339565 617799 339637 617855
rect 339565 617765 339584 617799
rect 339618 617765 339637 617799
rect 338675 617694 338694 617728
rect 338728 617694 338747 617728
rect 338675 617671 338747 617694
rect 339565 617709 339637 617765
rect 339565 617675 339584 617709
rect 339618 617675 339637 617709
rect 339565 617671 339637 617675
rect 338675 617652 339637 617671
rect 338675 617618 338752 617652
rect 338786 617618 338842 617652
rect 338876 617618 338932 617652
rect 338966 617618 339022 617652
rect 339056 617618 339112 617652
rect 339146 617618 339202 617652
rect 339236 617618 339292 617652
rect 339326 617618 339382 617652
rect 339416 617618 339472 617652
rect 339506 617618 339637 617652
rect 338675 617599 339637 617618
rect 339963 618542 340925 618561
rect 339963 618508 340074 618542
rect 340108 618508 340164 618542
rect 340198 618508 340254 618542
rect 340288 618508 340344 618542
rect 340378 618508 340434 618542
rect 340468 618508 340524 618542
rect 340558 618508 340614 618542
rect 340648 618508 340704 618542
rect 340738 618508 340794 618542
rect 340828 618508 340925 618542
rect 339963 618489 340925 618508
rect 339963 618448 340035 618489
rect 339963 618414 339982 618448
rect 340016 618414 340035 618448
rect 340853 618429 340925 618489
rect 339963 618358 340035 618414
rect 339963 618324 339982 618358
rect 340016 618324 340035 618358
rect 339963 618268 340035 618324
rect 339963 618234 339982 618268
rect 340016 618234 340035 618268
rect 339963 618178 340035 618234
rect 339963 618144 339982 618178
rect 340016 618144 340035 618178
rect 339963 618088 340035 618144
rect 339963 618054 339982 618088
rect 340016 618054 340035 618088
rect 339963 617998 340035 618054
rect 339963 617964 339982 617998
rect 340016 617964 340035 617998
rect 339963 617908 340035 617964
rect 339963 617874 339982 617908
rect 340016 617874 340035 617908
rect 339963 617818 340035 617874
rect 339963 617784 339982 617818
rect 340016 617784 340035 617818
rect 339963 617728 340035 617784
rect 340853 618395 340872 618429
rect 340906 618395 340925 618429
rect 340853 618339 340925 618395
rect 340853 618305 340872 618339
rect 340906 618305 340925 618339
rect 340853 618249 340925 618305
rect 340853 618215 340872 618249
rect 340906 618215 340925 618249
rect 340853 618159 340925 618215
rect 340853 618125 340872 618159
rect 340906 618125 340925 618159
rect 340853 618069 340925 618125
rect 340853 618035 340872 618069
rect 340906 618035 340925 618069
rect 340853 617979 340925 618035
rect 340853 617945 340872 617979
rect 340906 617945 340925 617979
rect 340853 617889 340925 617945
rect 340853 617855 340872 617889
rect 340906 617855 340925 617889
rect 340853 617799 340925 617855
rect 340853 617765 340872 617799
rect 340906 617765 340925 617799
rect 339963 617694 339982 617728
rect 340016 617694 340035 617728
rect 339963 617671 340035 617694
rect 340853 617709 340925 617765
rect 340853 617675 340872 617709
rect 340906 617675 340925 617709
rect 340853 617671 340925 617675
rect 339963 617652 340925 617671
rect 339963 617618 340040 617652
rect 340074 617618 340130 617652
rect 340164 617618 340220 617652
rect 340254 617618 340310 617652
rect 340344 617618 340400 617652
rect 340434 617618 340490 617652
rect 340524 617618 340580 617652
rect 340614 617618 340670 617652
rect 340704 617618 340760 617652
rect 340794 617618 340925 617652
rect 339963 617599 340925 617618
rect 306436 616802 308978 616852
rect 306436 616702 306536 616802
rect 308878 616702 308978 616802
rect 306436 616652 308978 616702
<< psubdiffcont >>
rect 297824 641672 343136 642672
rect 297872 616472 298872 640624
rect 300688 639776 311872 640542
rect 312448 630702 313018 637006
rect 315692 630702 316262 637006
rect 320652 630702 321222 637006
rect 335340 630702 335910 637006
rect 334782 627674 334816 627708
rect 334872 627674 334906 627708
rect 334962 627674 334996 627708
rect 335052 627674 335086 627708
rect 335142 627674 335176 627708
rect 335232 627674 335266 627708
rect 335322 627674 335356 627708
rect 335412 627674 335446 627708
rect 335502 627674 335536 627708
rect 335592 627674 335626 627708
rect 335682 627674 335716 627708
rect 335772 627674 335806 627708
rect 336070 627674 336104 627708
rect 336160 627674 336194 627708
rect 336250 627674 336284 627708
rect 336340 627674 336374 627708
rect 336430 627674 336464 627708
rect 336520 627674 336554 627708
rect 336610 627674 336644 627708
rect 336700 627674 336734 627708
rect 336790 627674 336824 627708
rect 336880 627674 336914 627708
rect 336970 627674 337004 627708
rect 337060 627674 337094 627708
rect 337358 627674 337392 627708
rect 337448 627674 337482 627708
rect 337538 627674 337572 627708
rect 337628 627674 337662 627708
rect 337718 627674 337752 627708
rect 337808 627674 337842 627708
rect 337898 627674 337932 627708
rect 337988 627674 338022 627708
rect 338078 627674 338112 627708
rect 338168 627674 338202 627708
rect 338258 627674 338292 627708
rect 338348 627674 338382 627708
rect 338646 627674 338680 627708
rect 338736 627674 338770 627708
rect 338826 627674 338860 627708
rect 338916 627674 338950 627708
rect 339006 627674 339040 627708
rect 339096 627674 339130 627708
rect 339186 627674 339220 627708
rect 339276 627674 339310 627708
rect 339366 627674 339400 627708
rect 339456 627674 339490 627708
rect 339546 627674 339580 627708
rect 339636 627674 339670 627708
rect 339934 627674 339968 627708
rect 340024 627674 340058 627708
rect 340114 627674 340148 627708
rect 340204 627674 340238 627708
rect 340294 627674 340328 627708
rect 340384 627674 340418 627708
rect 340474 627674 340508 627708
rect 340564 627674 340598 627708
rect 340654 627674 340688 627708
rect 340744 627674 340778 627708
rect 340834 627674 340868 627708
rect 340924 627674 340958 627708
rect 334681 627590 334715 627624
rect 335868 627590 335902 627624
rect 335969 627590 336003 627624
rect 334681 627500 334715 627534
rect 334681 627410 334715 627444
rect 334681 627320 334715 627354
rect 334681 627230 334715 627264
rect 334681 627140 334715 627174
rect 334681 627050 334715 627084
rect 334681 626960 334715 626994
rect 334681 626870 334715 626904
rect 334681 626780 334715 626814
rect 334681 626690 334715 626724
rect 334681 626600 334715 626634
rect 337156 627590 337190 627624
rect 337257 627590 337291 627624
rect 335868 627500 335902 627534
rect 335969 627500 336003 627534
rect 335868 627410 335902 627444
rect 335969 627410 336003 627444
rect 335868 627320 335902 627354
rect 335969 627320 336003 627354
rect 335868 627230 335902 627264
rect 335969 627230 336003 627264
rect 335868 627140 335902 627174
rect 335969 627140 336003 627174
rect 335868 627050 335902 627084
rect 335969 627050 336003 627084
rect 335868 626960 335902 626994
rect 335969 626960 336003 626994
rect 335868 626870 335902 626904
rect 335969 626870 336003 626904
rect 335868 626780 335902 626814
rect 335969 626780 336003 626814
rect 335868 626690 335902 626724
rect 335969 626690 336003 626724
rect 335868 626600 335902 626634
rect 335969 626600 336003 626634
rect 338444 627590 338478 627624
rect 338545 627590 338579 627624
rect 337156 627500 337190 627534
rect 337257 627500 337291 627534
rect 337156 627410 337190 627444
rect 337257 627410 337291 627444
rect 337156 627320 337190 627354
rect 337257 627320 337291 627354
rect 337156 627230 337190 627264
rect 337257 627230 337291 627264
rect 337156 627140 337190 627174
rect 337257 627140 337291 627174
rect 337156 627050 337190 627084
rect 337257 627050 337291 627084
rect 337156 626960 337190 626994
rect 337257 626960 337291 626994
rect 337156 626870 337190 626904
rect 337257 626870 337291 626904
rect 337156 626780 337190 626814
rect 337257 626780 337291 626814
rect 337156 626690 337190 626724
rect 337257 626690 337291 626724
rect 337156 626600 337190 626634
rect 337257 626600 337291 626634
rect 339732 627590 339766 627624
rect 339833 627590 339867 627624
rect 338444 627500 338478 627534
rect 338545 627500 338579 627534
rect 338444 627410 338478 627444
rect 338545 627410 338579 627444
rect 338444 627320 338478 627354
rect 338545 627320 338579 627354
rect 338444 627230 338478 627264
rect 338545 627230 338579 627264
rect 338444 627140 338478 627174
rect 338545 627140 338579 627174
rect 338444 627050 338478 627084
rect 338545 627050 338579 627084
rect 338444 626960 338478 626994
rect 338545 626960 338579 626994
rect 338444 626870 338478 626904
rect 338545 626870 338579 626904
rect 338444 626780 338478 626814
rect 338545 626780 338579 626814
rect 338444 626690 338478 626724
rect 338545 626690 338579 626724
rect 338444 626600 338478 626634
rect 338545 626600 338579 626634
rect 341020 627590 341054 627624
rect 339732 627500 339766 627534
rect 339833 627500 339867 627534
rect 339732 627410 339766 627444
rect 339833 627410 339867 627444
rect 339732 627320 339766 627354
rect 339833 627320 339867 627354
rect 339732 627230 339766 627264
rect 339833 627230 339867 627264
rect 339732 627140 339766 627174
rect 339833 627140 339867 627174
rect 339732 627050 339766 627084
rect 339833 627050 339867 627084
rect 339732 626960 339766 626994
rect 339833 626960 339867 626994
rect 339732 626870 339766 626904
rect 339833 626870 339867 626904
rect 339732 626780 339766 626814
rect 339833 626780 339867 626814
rect 339732 626690 339766 626724
rect 339833 626690 339867 626724
rect 339732 626600 339766 626634
rect 339833 626600 339867 626634
rect 341020 627500 341054 627534
rect 341020 627410 341054 627444
rect 341020 627320 341054 627354
rect 341020 627230 341054 627264
rect 341020 627140 341054 627174
rect 341020 627050 341054 627084
rect 341020 626960 341054 626994
rect 341020 626870 341054 626904
rect 341020 626780 341054 626814
rect 341020 626690 341054 626724
rect 341020 626600 341054 626634
rect 334681 626510 334715 626544
rect 334782 626487 334816 626521
rect 334872 626487 334906 626521
rect 334962 626487 334996 626521
rect 335052 626487 335086 626521
rect 335142 626487 335176 626521
rect 335232 626487 335266 626521
rect 335322 626487 335356 626521
rect 335412 626487 335446 626521
rect 335502 626487 335536 626521
rect 335592 626487 335626 626521
rect 335682 626487 335716 626521
rect 335772 626487 335806 626521
rect 335868 626510 335902 626544
rect 335969 626510 336003 626544
rect 336070 626487 336104 626521
rect 336160 626487 336194 626521
rect 336250 626487 336284 626521
rect 336340 626487 336374 626521
rect 336430 626487 336464 626521
rect 336520 626487 336554 626521
rect 336610 626487 336644 626521
rect 336700 626487 336734 626521
rect 336790 626487 336824 626521
rect 336880 626487 336914 626521
rect 336970 626487 337004 626521
rect 337060 626487 337094 626521
rect 337156 626510 337190 626544
rect 337257 626510 337291 626544
rect 337358 626487 337392 626521
rect 337448 626487 337482 626521
rect 337538 626487 337572 626521
rect 337628 626487 337662 626521
rect 337718 626487 337752 626521
rect 337808 626487 337842 626521
rect 337898 626487 337932 626521
rect 337988 626487 338022 626521
rect 338078 626487 338112 626521
rect 338168 626487 338202 626521
rect 338258 626487 338292 626521
rect 338348 626487 338382 626521
rect 338444 626510 338478 626544
rect 338545 626510 338579 626544
rect 338646 626487 338680 626521
rect 338736 626487 338770 626521
rect 338826 626487 338860 626521
rect 338916 626487 338950 626521
rect 339006 626487 339040 626521
rect 339096 626487 339130 626521
rect 339186 626487 339220 626521
rect 339276 626487 339310 626521
rect 339366 626487 339400 626521
rect 339456 626487 339490 626521
rect 339546 626487 339580 626521
rect 339636 626487 339670 626521
rect 339732 626510 339766 626544
rect 339833 626510 339867 626544
rect 339934 626487 339968 626521
rect 340024 626487 340058 626521
rect 340114 626487 340148 626521
rect 340204 626487 340238 626521
rect 340294 626487 340328 626521
rect 340384 626487 340418 626521
rect 340474 626487 340508 626521
rect 340564 626487 340598 626521
rect 340654 626487 340688 626521
rect 340744 626487 340778 626521
rect 340834 626487 340868 626521
rect 340924 626487 340958 626521
rect 341020 626510 341054 626544
rect 334782 626386 334816 626420
rect 334872 626386 334906 626420
rect 334962 626386 334996 626420
rect 335052 626386 335086 626420
rect 335142 626386 335176 626420
rect 335232 626386 335266 626420
rect 335322 626386 335356 626420
rect 335412 626386 335446 626420
rect 335502 626386 335536 626420
rect 335592 626386 335626 626420
rect 335682 626386 335716 626420
rect 335772 626386 335806 626420
rect 336070 626386 336104 626420
rect 336160 626386 336194 626420
rect 336250 626386 336284 626420
rect 336340 626386 336374 626420
rect 336430 626386 336464 626420
rect 336520 626386 336554 626420
rect 336610 626386 336644 626420
rect 336700 626386 336734 626420
rect 336790 626386 336824 626420
rect 336880 626386 336914 626420
rect 336970 626386 337004 626420
rect 337060 626386 337094 626420
rect 337358 626386 337392 626420
rect 337448 626386 337482 626420
rect 337538 626386 337572 626420
rect 337628 626386 337662 626420
rect 337718 626386 337752 626420
rect 337808 626386 337842 626420
rect 337898 626386 337932 626420
rect 337988 626386 338022 626420
rect 338078 626386 338112 626420
rect 338168 626386 338202 626420
rect 338258 626386 338292 626420
rect 338348 626386 338382 626420
rect 338646 626386 338680 626420
rect 338736 626386 338770 626420
rect 338826 626386 338860 626420
rect 338916 626386 338950 626420
rect 339006 626386 339040 626420
rect 339096 626386 339130 626420
rect 339186 626386 339220 626420
rect 339276 626386 339310 626420
rect 339366 626386 339400 626420
rect 339456 626386 339490 626420
rect 339546 626386 339580 626420
rect 339636 626386 339670 626420
rect 339934 626386 339968 626420
rect 340024 626386 340058 626420
rect 340114 626386 340148 626420
rect 340204 626386 340238 626420
rect 340294 626386 340328 626420
rect 340384 626386 340418 626420
rect 340474 626386 340508 626420
rect 340564 626386 340598 626420
rect 340654 626386 340688 626420
rect 340744 626386 340778 626420
rect 340834 626386 340868 626420
rect 340924 626386 340958 626420
rect 334681 626302 334715 626336
rect 335868 626302 335902 626336
rect 335969 626302 336003 626336
rect 334681 626212 334715 626246
rect 334681 626122 334715 626156
rect 334681 626032 334715 626066
rect 334681 625942 334715 625976
rect 334681 625852 334715 625886
rect 334681 625762 334715 625796
rect 334681 625672 334715 625706
rect 334681 625582 334715 625616
rect 334681 625492 334715 625526
rect 334681 625402 334715 625436
rect 334681 625312 334715 625346
rect 337156 626302 337190 626336
rect 337257 626302 337291 626336
rect 335868 626212 335902 626246
rect 335969 626212 336003 626246
rect 335868 626122 335902 626156
rect 335969 626122 336003 626156
rect 335868 626032 335902 626066
rect 335969 626032 336003 626066
rect 335868 625942 335902 625976
rect 335969 625942 336003 625976
rect 335868 625852 335902 625886
rect 335969 625852 336003 625886
rect 335868 625762 335902 625796
rect 335969 625762 336003 625796
rect 335868 625672 335902 625706
rect 335969 625672 336003 625706
rect 335868 625582 335902 625616
rect 335969 625582 336003 625616
rect 335868 625492 335902 625526
rect 335969 625492 336003 625526
rect 335868 625402 335902 625436
rect 335969 625402 336003 625436
rect 335868 625312 335902 625346
rect 335969 625312 336003 625346
rect 338444 626302 338478 626336
rect 338545 626302 338579 626336
rect 337156 626212 337190 626246
rect 337257 626212 337291 626246
rect 337156 626122 337190 626156
rect 337257 626122 337291 626156
rect 337156 626032 337190 626066
rect 337257 626032 337291 626066
rect 337156 625942 337190 625976
rect 337257 625942 337291 625976
rect 337156 625852 337190 625886
rect 337257 625852 337291 625886
rect 337156 625762 337190 625796
rect 337257 625762 337291 625796
rect 337156 625672 337190 625706
rect 337257 625672 337291 625706
rect 337156 625582 337190 625616
rect 337257 625582 337291 625616
rect 337156 625492 337190 625526
rect 337257 625492 337291 625526
rect 337156 625402 337190 625436
rect 337257 625402 337291 625436
rect 337156 625312 337190 625346
rect 337257 625312 337291 625346
rect 339732 626302 339766 626336
rect 339833 626302 339867 626336
rect 338444 626212 338478 626246
rect 338545 626212 338579 626246
rect 338444 626122 338478 626156
rect 338545 626122 338579 626156
rect 338444 626032 338478 626066
rect 338545 626032 338579 626066
rect 338444 625942 338478 625976
rect 338545 625942 338579 625976
rect 338444 625852 338478 625886
rect 338545 625852 338579 625886
rect 338444 625762 338478 625796
rect 338545 625762 338579 625796
rect 338444 625672 338478 625706
rect 338545 625672 338579 625706
rect 338444 625582 338478 625616
rect 338545 625582 338579 625616
rect 338444 625492 338478 625526
rect 338545 625492 338579 625526
rect 338444 625402 338478 625436
rect 338545 625402 338579 625436
rect 338444 625312 338478 625346
rect 338545 625312 338579 625346
rect 341020 626302 341054 626336
rect 339732 626212 339766 626246
rect 339833 626212 339867 626246
rect 339732 626122 339766 626156
rect 339833 626122 339867 626156
rect 339732 626032 339766 626066
rect 339833 626032 339867 626066
rect 339732 625942 339766 625976
rect 339833 625942 339867 625976
rect 339732 625852 339766 625886
rect 339833 625852 339867 625886
rect 339732 625762 339766 625796
rect 339833 625762 339867 625796
rect 339732 625672 339766 625706
rect 339833 625672 339867 625706
rect 339732 625582 339766 625616
rect 339833 625582 339867 625616
rect 339732 625492 339766 625526
rect 339833 625492 339867 625526
rect 339732 625402 339766 625436
rect 339833 625402 339867 625436
rect 339732 625312 339766 625346
rect 339833 625312 339867 625346
rect 341020 626212 341054 626246
rect 341020 626122 341054 626156
rect 341020 626032 341054 626066
rect 341020 625942 341054 625976
rect 341020 625852 341054 625886
rect 341020 625762 341054 625796
rect 341020 625672 341054 625706
rect 341020 625582 341054 625616
rect 341020 625492 341054 625526
rect 341020 625402 341054 625436
rect 341020 625312 341054 625346
rect 334681 625222 334715 625256
rect 334782 625199 334816 625233
rect 334872 625199 334906 625233
rect 334962 625199 334996 625233
rect 335052 625199 335086 625233
rect 335142 625199 335176 625233
rect 335232 625199 335266 625233
rect 335322 625199 335356 625233
rect 335412 625199 335446 625233
rect 335502 625199 335536 625233
rect 335592 625199 335626 625233
rect 335682 625199 335716 625233
rect 335772 625199 335806 625233
rect 335868 625222 335902 625256
rect 335969 625222 336003 625256
rect 336070 625199 336104 625233
rect 336160 625199 336194 625233
rect 336250 625199 336284 625233
rect 336340 625199 336374 625233
rect 336430 625199 336464 625233
rect 336520 625199 336554 625233
rect 336610 625199 336644 625233
rect 336700 625199 336734 625233
rect 336790 625199 336824 625233
rect 336880 625199 336914 625233
rect 336970 625199 337004 625233
rect 337060 625199 337094 625233
rect 337156 625222 337190 625256
rect 337257 625222 337291 625256
rect 337358 625199 337392 625233
rect 337448 625199 337482 625233
rect 337538 625199 337572 625233
rect 337628 625199 337662 625233
rect 337718 625199 337752 625233
rect 337808 625199 337842 625233
rect 337898 625199 337932 625233
rect 337988 625199 338022 625233
rect 338078 625199 338112 625233
rect 338168 625199 338202 625233
rect 338258 625199 338292 625233
rect 338348 625199 338382 625233
rect 338444 625222 338478 625256
rect 338545 625222 338579 625256
rect 338646 625199 338680 625233
rect 338736 625199 338770 625233
rect 338826 625199 338860 625233
rect 338916 625199 338950 625233
rect 339006 625199 339040 625233
rect 339096 625199 339130 625233
rect 339186 625199 339220 625233
rect 339276 625199 339310 625233
rect 339366 625199 339400 625233
rect 339456 625199 339490 625233
rect 339546 625199 339580 625233
rect 339636 625199 339670 625233
rect 339732 625222 339766 625256
rect 339833 625222 339867 625256
rect 339934 625199 339968 625233
rect 340024 625199 340058 625233
rect 340114 625199 340148 625233
rect 340204 625199 340238 625233
rect 340294 625199 340328 625233
rect 340384 625199 340418 625233
rect 340474 625199 340508 625233
rect 340564 625199 340598 625233
rect 340654 625199 340688 625233
rect 340744 625199 340778 625233
rect 340834 625199 340868 625233
rect 340924 625199 340958 625233
rect 341020 625222 341054 625256
rect 334782 625098 334816 625132
rect 334872 625098 334906 625132
rect 334962 625098 334996 625132
rect 335052 625098 335086 625132
rect 335142 625098 335176 625132
rect 335232 625098 335266 625132
rect 335322 625098 335356 625132
rect 335412 625098 335446 625132
rect 335502 625098 335536 625132
rect 335592 625098 335626 625132
rect 335682 625098 335716 625132
rect 335772 625098 335806 625132
rect 336070 625098 336104 625132
rect 336160 625098 336194 625132
rect 336250 625098 336284 625132
rect 336340 625098 336374 625132
rect 336430 625098 336464 625132
rect 336520 625098 336554 625132
rect 336610 625098 336644 625132
rect 336700 625098 336734 625132
rect 336790 625098 336824 625132
rect 336880 625098 336914 625132
rect 336970 625098 337004 625132
rect 337060 625098 337094 625132
rect 337358 625098 337392 625132
rect 337448 625098 337482 625132
rect 337538 625098 337572 625132
rect 337628 625098 337662 625132
rect 337718 625098 337752 625132
rect 337808 625098 337842 625132
rect 337898 625098 337932 625132
rect 337988 625098 338022 625132
rect 338078 625098 338112 625132
rect 338168 625098 338202 625132
rect 338258 625098 338292 625132
rect 338348 625098 338382 625132
rect 338646 625098 338680 625132
rect 338736 625098 338770 625132
rect 338826 625098 338860 625132
rect 338916 625098 338950 625132
rect 339006 625098 339040 625132
rect 339096 625098 339130 625132
rect 339186 625098 339220 625132
rect 339276 625098 339310 625132
rect 339366 625098 339400 625132
rect 339456 625098 339490 625132
rect 339546 625098 339580 625132
rect 339636 625098 339670 625132
rect 339934 625098 339968 625132
rect 340024 625098 340058 625132
rect 340114 625098 340148 625132
rect 340204 625098 340238 625132
rect 340294 625098 340328 625132
rect 340384 625098 340418 625132
rect 340474 625098 340508 625132
rect 340564 625098 340598 625132
rect 340654 625098 340688 625132
rect 340744 625098 340778 625132
rect 340834 625098 340868 625132
rect 340924 625098 340958 625132
rect 334681 625014 334715 625048
rect 335868 625014 335902 625048
rect 335969 625014 336003 625048
rect 304322 624556 310774 624888
rect 301286 621266 302278 621342
rect 299900 620612 300300 621188
rect 303266 620612 303666 621188
rect 304770 620548 304870 622148
rect 310270 620548 310370 622148
rect 334681 624924 334715 624958
rect 334681 624834 334715 624868
rect 334681 624744 334715 624778
rect 334681 624654 334715 624688
rect 334681 624564 334715 624598
rect 334681 624474 334715 624508
rect 334681 624384 334715 624418
rect 334681 624294 334715 624328
rect 334681 624204 334715 624238
rect 334681 624114 334715 624148
rect 334681 624024 334715 624058
rect 337156 625014 337190 625048
rect 337257 625014 337291 625048
rect 335868 624924 335902 624958
rect 335969 624924 336003 624958
rect 335868 624834 335902 624868
rect 335969 624834 336003 624868
rect 335868 624744 335902 624778
rect 335969 624744 336003 624778
rect 335868 624654 335902 624688
rect 335969 624654 336003 624688
rect 335868 624564 335902 624598
rect 335969 624564 336003 624598
rect 335868 624474 335902 624508
rect 335969 624474 336003 624508
rect 335868 624384 335902 624418
rect 335969 624384 336003 624418
rect 335868 624294 335902 624328
rect 335969 624294 336003 624328
rect 335868 624204 335902 624238
rect 335969 624204 336003 624238
rect 335868 624114 335902 624148
rect 335969 624114 336003 624148
rect 335868 624024 335902 624058
rect 335969 624024 336003 624058
rect 338444 625014 338478 625048
rect 338545 625014 338579 625048
rect 337156 624924 337190 624958
rect 337257 624924 337291 624958
rect 337156 624834 337190 624868
rect 337257 624834 337291 624868
rect 337156 624744 337190 624778
rect 337257 624744 337291 624778
rect 337156 624654 337190 624688
rect 337257 624654 337291 624688
rect 337156 624564 337190 624598
rect 337257 624564 337291 624598
rect 337156 624474 337190 624508
rect 337257 624474 337291 624508
rect 337156 624384 337190 624418
rect 337257 624384 337291 624418
rect 337156 624294 337190 624328
rect 337257 624294 337291 624328
rect 337156 624204 337190 624238
rect 337257 624204 337291 624238
rect 337156 624114 337190 624148
rect 337257 624114 337291 624148
rect 337156 624024 337190 624058
rect 337257 624024 337291 624058
rect 339732 625014 339766 625048
rect 339833 625014 339867 625048
rect 338444 624924 338478 624958
rect 338545 624924 338579 624958
rect 338444 624834 338478 624868
rect 338545 624834 338579 624868
rect 338444 624744 338478 624778
rect 338545 624744 338579 624778
rect 338444 624654 338478 624688
rect 338545 624654 338579 624688
rect 338444 624564 338478 624598
rect 338545 624564 338579 624598
rect 338444 624474 338478 624508
rect 338545 624474 338579 624508
rect 338444 624384 338478 624418
rect 338545 624384 338579 624418
rect 338444 624294 338478 624328
rect 338545 624294 338579 624328
rect 338444 624204 338478 624238
rect 338545 624204 338579 624238
rect 338444 624114 338478 624148
rect 338545 624114 338579 624148
rect 338444 624024 338478 624058
rect 338545 624024 338579 624058
rect 341020 625014 341054 625048
rect 339732 624924 339766 624958
rect 339833 624924 339867 624958
rect 339732 624834 339766 624868
rect 339833 624834 339867 624868
rect 339732 624744 339766 624778
rect 339833 624744 339867 624778
rect 339732 624654 339766 624688
rect 339833 624654 339867 624688
rect 339732 624564 339766 624598
rect 339833 624564 339867 624598
rect 339732 624474 339766 624508
rect 339833 624474 339867 624508
rect 339732 624384 339766 624418
rect 339833 624384 339867 624418
rect 339732 624294 339766 624328
rect 339833 624294 339867 624328
rect 339732 624204 339766 624238
rect 339833 624204 339867 624238
rect 339732 624114 339766 624148
rect 339833 624114 339867 624148
rect 339732 624024 339766 624058
rect 339833 624024 339867 624058
rect 341020 624924 341054 624958
rect 341020 624834 341054 624868
rect 341020 624744 341054 624778
rect 341020 624654 341054 624688
rect 341020 624564 341054 624598
rect 341020 624474 341054 624508
rect 341020 624384 341054 624418
rect 341020 624294 341054 624328
rect 341020 624204 341054 624238
rect 341020 624114 341054 624148
rect 341020 624024 341054 624058
rect 334681 623934 334715 623968
rect 334782 623911 334816 623945
rect 334872 623911 334906 623945
rect 334962 623911 334996 623945
rect 335052 623911 335086 623945
rect 335142 623911 335176 623945
rect 335232 623911 335266 623945
rect 335322 623911 335356 623945
rect 335412 623911 335446 623945
rect 335502 623911 335536 623945
rect 335592 623911 335626 623945
rect 335682 623911 335716 623945
rect 335772 623911 335806 623945
rect 335868 623934 335902 623968
rect 335969 623934 336003 623968
rect 336070 623911 336104 623945
rect 336160 623911 336194 623945
rect 336250 623911 336284 623945
rect 336340 623911 336374 623945
rect 336430 623911 336464 623945
rect 336520 623911 336554 623945
rect 336610 623911 336644 623945
rect 336700 623911 336734 623945
rect 336790 623911 336824 623945
rect 336880 623911 336914 623945
rect 336970 623911 337004 623945
rect 337060 623911 337094 623945
rect 337156 623934 337190 623968
rect 337257 623934 337291 623968
rect 337358 623911 337392 623945
rect 337448 623911 337482 623945
rect 337538 623911 337572 623945
rect 337628 623911 337662 623945
rect 337718 623911 337752 623945
rect 337808 623911 337842 623945
rect 337898 623911 337932 623945
rect 337988 623911 338022 623945
rect 338078 623911 338112 623945
rect 338168 623911 338202 623945
rect 338258 623911 338292 623945
rect 338348 623911 338382 623945
rect 338444 623934 338478 623968
rect 338545 623934 338579 623968
rect 338646 623911 338680 623945
rect 338736 623911 338770 623945
rect 338826 623911 338860 623945
rect 338916 623911 338950 623945
rect 339006 623911 339040 623945
rect 339096 623911 339130 623945
rect 339186 623911 339220 623945
rect 339276 623911 339310 623945
rect 339366 623911 339400 623945
rect 339456 623911 339490 623945
rect 339546 623911 339580 623945
rect 339636 623911 339670 623945
rect 339732 623934 339766 623968
rect 339833 623934 339867 623968
rect 339934 623911 339968 623945
rect 340024 623911 340058 623945
rect 340114 623911 340148 623945
rect 340204 623911 340238 623945
rect 340294 623911 340328 623945
rect 340384 623911 340418 623945
rect 340474 623911 340508 623945
rect 340564 623911 340598 623945
rect 340654 623911 340688 623945
rect 340744 623911 340778 623945
rect 340834 623911 340868 623945
rect 340924 623911 340958 623945
rect 341020 623934 341054 623968
rect 334782 623810 334816 623844
rect 334872 623810 334906 623844
rect 334962 623810 334996 623844
rect 335052 623810 335086 623844
rect 335142 623810 335176 623844
rect 335232 623810 335266 623844
rect 335322 623810 335356 623844
rect 335412 623810 335446 623844
rect 335502 623810 335536 623844
rect 335592 623810 335626 623844
rect 335682 623810 335716 623844
rect 335772 623810 335806 623844
rect 336070 623810 336104 623844
rect 336160 623810 336194 623844
rect 336250 623810 336284 623844
rect 336340 623810 336374 623844
rect 336430 623810 336464 623844
rect 336520 623810 336554 623844
rect 336610 623810 336644 623844
rect 336700 623810 336734 623844
rect 336790 623810 336824 623844
rect 336880 623810 336914 623844
rect 336970 623810 337004 623844
rect 337060 623810 337094 623844
rect 337358 623810 337392 623844
rect 337448 623810 337482 623844
rect 337538 623810 337572 623844
rect 337628 623810 337662 623844
rect 337718 623810 337752 623844
rect 337808 623810 337842 623844
rect 337898 623810 337932 623844
rect 337988 623810 338022 623844
rect 338078 623810 338112 623844
rect 338168 623810 338202 623844
rect 338258 623810 338292 623844
rect 338348 623810 338382 623844
rect 338646 623810 338680 623844
rect 338736 623810 338770 623844
rect 338826 623810 338860 623844
rect 338916 623810 338950 623844
rect 339006 623810 339040 623844
rect 339096 623810 339130 623844
rect 339186 623810 339220 623844
rect 339276 623810 339310 623844
rect 339366 623810 339400 623844
rect 339456 623810 339490 623844
rect 339546 623810 339580 623844
rect 339636 623810 339670 623844
rect 339934 623810 339968 623844
rect 340024 623810 340058 623844
rect 340114 623810 340148 623844
rect 340204 623810 340238 623844
rect 340294 623810 340328 623844
rect 340384 623810 340418 623844
rect 340474 623810 340508 623844
rect 340564 623810 340598 623844
rect 340654 623810 340688 623844
rect 340744 623810 340778 623844
rect 340834 623810 340868 623844
rect 340924 623810 340958 623844
rect 334681 623726 334715 623760
rect 335868 623726 335902 623760
rect 335969 623726 336003 623760
rect 334681 623636 334715 623670
rect 334681 623546 334715 623580
rect 334681 623456 334715 623490
rect 334681 623366 334715 623400
rect 334681 623276 334715 623310
rect 334681 623186 334715 623220
rect 334681 623096 334715 623130
rect 334681 623006 334715 623040
rect 334681 622916 334715 622950
rect 334681 622826 334715 622860
rect 334681 622736 334715 622770
rect 337156 623726 337190 623760
rect 337257 623726 337291 623760
rect 335868 623636 335902 623670
rect 335969 623636 336003 623670
rect 335868 623546 335902 623580
rect 335969 623546 336003 623580
rect 335868 623456 335902 623490
rect 335969 623456 336003 623490
rect 335868 623366 335902 623400
rect 335969 623366 336003 623400
rect 335868 623276 335902 623310
rect 335969 623276 336003 623310
rect 335868 623186 335902 623220
rect 335969 623186 336003 623220
rect 335868 623096 335902 623130
rect 335969 623096 336003 623130
rect 335868 623006 335902 623040
rect 335969 623006 336003 623040
rect 335868 622916 335902 622950
rect 335969 622916 336003 622950
rect 335868 622826 335902 622860
rect 335969 622826 336003 622860
rect 335868 622736 335902 622770
rect 335969 622736 336003 622770
rect 338444 623726 338478 623760
rect 338545 623726 338579 623760
rect 337156 623636 337190 623670
rect 337257 623636 337291 623670
rect 337156 623546 337190 623580
rect 337257 623546 337291 623580
rect 337156 623456 337190 623490
rect 337257 623456 337291 623490
rect 337156 623366 337190 623400
rect 337257 623366 337291 623400
rect 337156 623276 337190 623310
rect 337257 623276 337291 623310
rect 337156 623186 337190 623220
rect 337257 623186 337291 623220
rect 337156 623096 337190 623130
rect 337257 623096 337291 623130
rect 337156 623006 337190 623040
rect 337257 623006 337291 623040
rect 337156 622916 337190 622950
rect 337257 622916 337291 622950
rect 337156 622826 337190 622860
rect 337257 622826 337291 622860
rect 337156 622736 337190 622770
rect 337257 622736 337291 622770
rect 339732 623726 339766 623760
rect 339833 623726 339867 623760
rect 338444 623636 338478 623670
rect 338545 623636 338579 623670
rect 338444 623546 338478 623580
rect 338545 623546 338579 623580
rect 338444 623456 338478 623490
rect 338545 623456 338579 623490
rect 338444 623366 338478 623400
rect 338545 623366 338579 623400
rect 338444 623276 338478 623310
rect 338545 623276 338579 623310
rect 338444 623186 338478 623220
rect 338545 623186 338579 623220
rect 338444 623096 338478 623130
rect 338545 623096 338579 623130
rect 338444 623006 338478 623040
rect 338545 623006 338579 623040
rect 338444 622916 338478 622950
rect 338545 622916 338579 622950
rect 338444 622826 338478 622860
rect 338545 622826 338579 622860
rect 338444 622736 338478 622770
rect 338545 622736 338579 622770
rect 341020 623726 341054 623760
rect 339732 623636 339766 623670
rect 339833 623636 339867 623670
rect 339732 623546 339766 623580
rect 339833 623546 339867 623580
rect 339732 623456 339766 623490
rect 339833 623456 339867 623490
rect 339732 623366 339766 623400
rect 339833 623366 339867 623400
rect 339732 623276 339766 623310
rect 339833 623276 339867 623310
rect 339732 623186 339766 623220
rect 339833 623186 339867 623220
rect 339732 623096 339766 623130
rect 339833 623096 339867 623130
rect 339732 623006 339766 623040
rect 339833 623006 339867 623040
rect 339732 622916 339766 622950
rect 339833 622916 339867 622950
rect 339732 622826 339766 622860
rect 339833 622826 339867 622860
rect 339732 622736 339766 622770
rect 339833 622736 339867 622770
rect 341020 623636 341054 623670
rect 341020 623546 341054 623580
rect 341020 623456 341054 623490
rect 341020 623366 341054 623400
rect 341020 623276 341054 623310
rect 341020 623186 341054 623220
rect 341020 623096 341054 623130
rect 341020 623006 341054 623040
rect 341020 622916 341054 622950
rect 341020 622826 341054 622860
rect 341020 622736 341054 622770
rect 334681 622646 334715 622680
rect 334782 622623 334816 622657
rect 334872 622623 334906 622657
rect 334962 622623 334996 622657
rect 335052 622623 335086 622657
rect 335142 622623 335176 622657
rect 335232 622623 335266 622657
rect 335322 622623 335356 622657
rect 335412 622623 335446 622657
rect 335502 622623 335536 622657
rect 335592 622623 335626 622657
rect 335682 622623 335716 622657
rect 335772 622623 335806 622657
rect 335868 622646 335902 622680
rect 335969 622646 336003 622680
rect 336070 622623 336104 622657
rect 336160 622623 336194 622657
rect 336250 622623 336284 622657
rect 336340 622623 336374 622657
rect 336430 622623 336464 622657
rect 336520 622623 336554 622657
rect 336610 622623 336644 622657
rect 336700 622623 336734 622657
rect 336790 622623 336824 622657
rect 336880 622623 336914 622657
rect 336970 622623 337004 622657
rect 337060 622623 337094 622657
rect 337156 622646 337190 622680
rect 337257 622646 337291 622680
rect 337358 622623 337392 622657
rect 337448 622623 337482 622657
rect 337538 622623 337572 622657
rect 337628 622623 337662 622657
rect 337718 622623 337752 622657
rect 337808 622623 337842 622657
rect 337898 622623 337932 622657
rect 337988 622623 338022 622657
rect 338078 622623 338112 622657
rect 338168 622623 338202 622657
rect 338258 622623 338292 622657
rect 338348 622623 338382 622657
rect 338444 622646 338478 622680
rect 338545 622646 338579 622680
rect 338646 622623 338680 622657
rect 338736 622623 338770 622657
rect 338826 622623 338860 622657
rect 338916 622623 338950 622657
rect 339006 622623 339040 622657
rect 339096 622623 339130 622657
rect 339186 622623 339220 622657
rect 339276 622623 339310 622657
rect 339366 622623 339400 622657
rect 339456 622623 339490 622657
rect 339546 622623 339580 622657
rect 339636 622623 339670 622657
rect 339732 622646 339766 622680
rect 339833 622646 339867 622680
rect 339934 622623 339968 622657
rect 340024 622623 340058 622657
rect 340114 622623 340148 622657
rect 340204 622623 340238 622657
rect 340294 622623 340328 622657
rect 340384 622623 340418 622657
rect 340474 622623 340508 622657
rect 340564 622623 340598 622657
rect 340654 622623 340688 622657
rect 340744 622623 340778 622657
rect 340834 622623 340868 622657
rect 340924 622623 340958 622657
rect 341020 622646 341054 622680
rect 334782 622522 334816 622556
rect 334872 622522 334906 622556
rect 334962 622522 334996 622556
rect 335052 622522 335086 622556
rect 335142 622522 335176 622556
rect 335232 622522 335266 622556
rect 335322 622522 335356 622556
rect 335412 622522 335446 622556
rect 335502 622522 335536 622556
rect 335592 622522 335626 622556
rect 335682 622522 335716 622556
rect 335772 622522 335806 622556
rect 336070 622522 336104 622556
rect 336160 622522 336194 622556
rect 336250 622522 336284 622556
rect 336340 622522 336374 622556
rect 336430 622522 336464 622556
rect 336520 622522 336554 622556
rect 336610 622522 336644 622556
rect 336700 622522 336734 622556
rect 336790 622522 336824 622556
rect 336880 622522 336914 622556
rect 336970 622522 337004 622556
rect 337060 622522 337094 622556
rect 337358 622522 337392 622556
rect 337448 622522 337482 622556
rect 337538 622522 337572 622556
rect 337628 622522 337662 622556
rect 337718 622522 337752 622556
rect 337808 622522 337842 622556
rect 337898 622522 337932 622556
rect 337988 622522 338022 622556
rect 338078 622522 338112 622556
rect 338168 622522 338202 622556
rect 338258 622522 338292 622556
rect 338348 622522 338382 622556
rect 338646 622522 338680 622556
rect 338736 622522 338770 622556
rect 338826 622522 338860 622556
rect 338916 622522 338950 622556
rect 339006 622522 339040 622556
rect 339096 622522 339130 622556
rect 339186 622522 339220 622556
rect 339276 622522 339310 622556
rect 339366 622522 339400 622556
rect 339456 622522 339490 622556
rect 339546 622522 339580 622556
rect 339636 622522 339670 622556
rect 339934 622522 339968 622556
rect 340024 622522 340058 622556
rect 340114 622522 340148 622556
rect 340204 622522 340238 622556
rect 340294 622522 340328 622556
rect 340384 622522 340418 622556
rect 340474 622522 340508 622556
rect 340564 622522 340598 622556
rect 340654 622522 340688 622556
rect 340744 622522 340778 622556
rect 340834 622522 340868 622556
rect 340924 622522 340958 622556
rect 334681 622438 334715 622472
rect 335868 622438 335902 622472
rect 335969 622438 336003 622472
rect 334681 622348 334715 622382
rect 334681 622258 334715 622292
rect 334681 622168 334715 622202
rect 334681 622078 334715 622112
rect 334681 621988 334715 622022
rect 334681 621898 334715 621932
rect 334681 621808 334715 621842
rect 334681 621718 334715 621752
rect 334681 621628 334715 621662
rect 334681 621538 334715 621572
rect 334681 621448 334715 621482
rect 337156 622438 337190 622472
rect 337257 622438 337291 622472
rect 335868 622348 335902 622382
rect 335969 622348 336003 622382
rect 335868 622258 335902 622292
rect 335969 622258 336003 622292
rect 335868 622168 335902 622202
rect 335969 622168 336003 622202
rect 335868 622078 335902 622112
rect 335969 622078 336003 622112
rect 335868 621988 335902 622022
rect 335969 621988 336003 622022
rect 335868 621898 335902 621932
rect 335969 621898 336003 621932
rect 335868 621808 335902 621842
rect 335969 621808 336003 621842
rect 335868 621718 335902 621752
rect 335969 621718 336003 621752
rect 335868 621628 335902 621662
rect 335969 621628 336003 621662
rect 335868 621538 335902 621572
rect 335969 621538 336003 621572
rect 335868 621448 335902 621482
rect 335969 621448 336003 621482
rect 338444 622438 338478 622472
rect 338545 622438 338579 622472
rect 337156 622348 337190 622382
rect 337257 622348 337291 622382
rect 337156 622258 337190 622292
rect 337257 622258 337291 622292
rect 337156 622168 337190 622202
rect 337257 622168 337291 622202
rect 337156 622078 337190 622112
rect 337257 622078 337291 622112
rect 337156 621988 337190 622022
rect 337257 621988 337291 622022
rect 337156 621898 337190 621932
rect 337257 621898 337291 621932
rect 337156 621808 337190 621842
rect 337257 621808 337291 621842
rect 337156 621718 337190 621752
rect 337257 621718 337291 621752
rect 337156 621628 337190 621662
rect 337257 621628 337291 621662
rect 337156 621538 337190 621572
rect 337257 621538 337291 621572
rect 337156 621448 337190 621482
rect 337257 621448 337291 621482
rect 339732 622438 339766 622472
rect 339833 622438 339867 622472
rect 338444 622348 338478 622382
rect 338545 622348 338579 622382
rect 338444 622258 338478 622292
rect 338545 622258 338579 622292
rect 338444 622168 338478 622202
rect 338545 622168 338579 622202
rect 338444 622078 338478 622112
rect 338545 622078 338579 622112
rect 338444 621988 338478 622022
rect 338545 621988 338579 622022
rect 338444 621898 338478 621932
rect 338545 621898 338579 621932
rect 338444 621808 338478 621842
rect 338545 621808 338579 621842
rect 338444 621718 338478 621752
rect 338545 621718 338579 621752
rect 338444 621628 338478 621662
rect 338545 621628 338579 621662
rect 338444 621538 338478 621572
rect 338545 621538 338579 621572
rect 338444 621448 338478 621482
rect 338545 621448 338579 621482
rect 341020 622438 341054 622472
rect 339732 622348 339766 622382
rect 339833 622348 339867 622382
rect 339732 622258 339766 622292
rect 339833 622258 339867 622292
rect 339732 622168 339766 622202
rect 339833 622168 339867 622202
rect 339732 622078 339766 622112
rect 339833 622078 339867 622112
rect 339732 621988 339766 622022
rect 339833 621988 339867 622022
rect 339732 621898 339766 621932
rect 339833 621898 339867 621932
rect 339732 621808 339766 621842
rect 339833 621808 339867 621842
rect 339732 621718 339766 621752
rect 339833 621718 339867 621752
rect 339732 621628 339766 621662
rect 339833 621628 339867 621662
rect 339732 621538 339766 621572
rect 339833 621538 339867 621572
rect 339732 621448 339766 621482
rect 339833 621448 339867 621482
rect 341020 622348 341054 622382
rect 341020 622258 341054 622292
rect 341020 622168 341054 622202
rect 341020 622078 341054 622112
rect 341020 621988 341054 622022
rect 341020 621898 341054 621932
rect 341020 621808 341054 621842
rect 341020 621718 341054 621752
rect 341020 621628 341054 621662
rect 341020 621538 341054 621572
rect 341020 621448 341054 621482
rect 334681 621358 334715 621392
rect 334782 621335 334816 621369
rect 334872 621335 334906 621369
rect 334962 621335 334996 621369
rect 335052 621335 335086 621369
rect 335142 621335 335176 621369
rect 335232 621335 335266 621369
rect 335322 621335 335356 621369
rect 335412 621335 335446 621369
rect 335502 621335 335536 621369
rect 335592 621335 335626 621369
rect 335682 621335 335716 621369
rect 335772 621335 335806 621369
rect 335868 621358 335902 621392
rect 335969 621358 336003 621392
rect 336070 621335 336104 621369
rect 336160 621335 336194 621369
rect 336250 621335 336284 621369
rect 336340 621335 336374 621369
rect 336430 621335 336464 621369
rect 336520 621335 336554 621369
rect 336610 621335 336644 621369
rect 336700 621335 336734 621369
rect 336790 621335 336824 621369
rect 336880 621335 336914 621369
rect 336970 621335 337004 621369
rect 337060 621335 337094 621369
rect 337156 621358 337190 621392
rect 337257 621358 337291 621392
rect 337358 621335 337392 621369
rect 337448 621335 337482 621369
rect 337538 621335 337572 621369
rect 337628 621335 337662 621369
rect 337718 621335 337752 621369
rect 337808 621335 337842 621369
rect 337898 621335 337932 621369
rect 337988 621335 338022 621369
rect 338078 621335 338112 621369
rect 338168 621335 338202 621369
rect 338258 621335 338292 621369
rect 338348 621335 338382 621369
rect 338444 621358 338478 621392
rect 338545 621358 338579 621392
rect 338646 621335 338680 621369
rect 338736 621335 338770 621369
rect 338826 621335 338860 621369
rect 338916 621335 338950 621369
rect 339006 621335 339040 621369
rect 339096 621335 339130 621369
rect 339186 621335 339220 621369
rect 339276 621335 339310 621369
rect 339366 621335 339400 621369
rect 339456 621335 339490 621369
rect 339546 621335 339580 621369
rect 339636 621335 339670 621369
rect 339732 621358 339766 621392
rect 339833 621358 339867 621392
rect 339934 621335 339968 621369
rect 340024 621335 340058 621369
rect 340114 621335 340148 621369
rect 340204 621335 340238 621369
rect 340294 621335 340328 621369
rect 340384 621335 340418 621369
rect 340474 621335 340508 621369
rect 340564 621335 340598 621369
rect 340654 621335 340688 621369
rect 340744 621335 340778 621369
rect 340834 621335 340868 621369
rect 340924 621335 340958 621369
rect 341020 621358 341054 621392
rect 334782 621234 334816 621268
rect 334872 621234 334906 621268
rect 334962 621234 334996 621268
rect 335052 621234 335086 621268
rect 335142 621234 335176 621268
rect 335232 621234 335266 621268
rect 335322 621234 335356 621268
rect 335412 621234 335446 621268
rect 335502 621234 335536 621268
rect 335592 621234 335626 621268
rect 335682 621234 335716 621268
rect 335772 621234 335806 621268
rect 336070 621234 336104 621268
rect 336160 621234 336194 621268
rect 336250 621234 336284 621268
rect 336340 621234 336374 621268
rect 336430 621234 336464 621268
rect 336520 621234 336554 621268
rect 336610 621234 336644 621268
rect 336700 621234 336734 621268
rect 336790 621234 336824 621268
rect 336880 621234 336914 621268
rect 336970 621234 337004 621268
rect 337060 621234 337094 621268
rect 337358 621234 337392 621268
rect 337448 621234 337482 621268
rect 337538 621234 337572 621268
rect 337628 621234 337662 621268
rect 337718 621234 337752 621268
rect 337808 621234 337842 621268
rect 337898 621234 337932 621268
rect 337988 621234 338022 621268
rect 338078 621234 338112 621268
rect 338168 621234 338202 621268
rect 338258 621234 338292 621268
rect 338348 621234 338382 621268
rect 338646 621234 338680 621268
rect 338736 621234 338770 621268
rect 338826 621234 338860 621268
rect 338916 621234 338950 621268
rect 339006 621234 339040 621268
rect 339096 621234 339130 621268
rect 339186 621234 339220 621268
rect 339276 621234 339310 621268
rect 339366 621234 339400 621268
rect 339456 621234 339490 621268
rect 339546 621234 339580 621268
rect 339636 621234 339670 621268
rect 339934 621234 339968 621268
rect 340024 621234 340058 621268
rect 340114 621234 340148 621268
rect 340204 621234 340238 621268
rect 340294 621234 340328 621268
rect 340384 621234 340418 621268
rect 340474 621234 340508 621268
rect 340564 621234 340598 621268
rect 340654 621234 340688 621268
rect 340744 621234 340778 621268
rect 340834 621234 340868 621268
rect 340924 621234 340958 621268
rect 334681 621150 334715 621184
rect 335868 621150 335902 621184
rect 335969 621150 336003 621184
rect 334681 621060 334715 621094
rect 334681 620970 334715 621004
rect 334681 620880 334715 620914
rect 334681 620790 334715 620824
rect 334681 620700 334715 620734
rect 334681 620610 334715 620644
rect 334681 620520 334715 620554
rect 334681 620430 334715 620464
rect 334681 620340 334715 620374
rect 334681 620250 334715 620284
rect 334681 620160 334715 620194
rect 337156 621150 337190 621184
rect 337257 621150 337291 621184
rect 335868 621060 335902 621094
rect 335969 621060 336003 621094
rect 335868 620970 335902 621004
rect 335969 620970 336003 621004
rect 335868 620880 335902 620914
rect 335969 620880 336003 620914
rect 335868 620790 335902 620824
rect 335969 620790 336003 620824
rect 335868 620700 335902 620734
rect 335969 620700 336003 620734
rect 335868 620610 335902 620644
rect 335969 620610 336003 620644
rect 335868 620520 335902 620554
rect 335969 620520 336003 620554
rect 335868 620430 335902 620464
rect 335969 620430 336003 620464
rect 335868 620340 335902 620374
rect 335969 620340 336003 620374
rect 335868 620250 335902 620284
rect 335969 620250 336003 620284
rect 335868 620160 335902 620194
rect 335969 620160 336003 620194
rect 338444 621150 338478 621184
rect 338545 621150 338579 621184
rect 337156 621060 337190 621094
rect 337257 621060 337291 621094
rect 337156 620970 337190 621004
rect 337257 620970 337291 621004
rect 337156 620880 337190 620914
rect 337257 620880 337291 620914
rect 337156 620790 337190 620824
rect 337257 620790 337291 620824
rect 337156 620700 337190 620734
rect 337257 620700 337291 620734
rect 337156 620610 337190 620644
rect 337257 620610 337291 620644
rect 337156 620520 337190 620554
rect 337257 620520 337291 620554
rect 337156 620430 337190 620464
rect 337257 620430 337291 620464
rect 337156 620340 337190 620374
rect 337257 620340 337291 620374
rect 337156 620250 337190 620284
rect 337257 620250 337291 620284
rect 337156 620160 337190 620194
rect 337257 620160 337291 620194
rect 339732 621150 339766 621184
rect 339833 621150 339867 621184
rect 338444 621060 338478 621094
rect 338545 621060 338579 621094
rect 338444 620970 338478 621004
rect 338545 620970 338579 621004
rect 338444 620880 338478 620914
rect 338545 620880 338579 620914
rect 338444 620790 338478 620824
rect 338545 620790 338579 620824
rect 338444 620700 338478 620734
rect 338545 620700 338579 620734
rect 338444 620610 338478 620644
rect 338545 620610 338579 620644
rect 338444 620520 338478 620554
rect 338545 620520 338579 620554
rect 338444 620430 338478 620464
rect 338545 620430 338579 620464
rect 338444 620340 338478 620374
rect 338545 620340 338579 620374
rect 338444 620250 338478 620284
rect 338545 620250 338579 620284
rect 338444 620160 338478 620194
rect 338545 620160 338579 620194
rect 341020 621150 341054 621184
rect 339732 621060 339766 621094
rect 339833 621060 339867 621094
rect 339732 620970 339766 621004
rect 339833 620970 339867 621004
rect 339732 620880 339766 620914
rect 339833 620880 339867 620914
rect 339732 620790 339766 620824
rect 339833 620790 339867 620824
rect 339732 620700 339766 620734
rect 339833 620700 339867 620734
rect 339732 620610 339766 620644
rect 339833 620610 339867 620644
rect 339732 620520 339766 620554
rect 339833 620520 339867 620554
rect 339732 620430 339766 620464
rect 339833 620430 339867 620464
rect 339732 620340 339766 620374
rect 339833 620340 339867 620374
rect 339732 620250 339766 620284
rect 339833 620250 339867 620284
rect 339732 620160 339766 620194
rect 339833 620160 339867 620194
rect 341020 621060 341054 621094
rect 341020 620970 341054 621004
rect 341020 620880 341054 620914
rect 341020 620790 341054 620824
rect 341020 620700 341054 620734
rect 341020 620610 341054 620644
rect 341020 620520 341054 620554
rect 341020 620430 341054 620464
rect 341020 620340 341054 620374
rect 341020 620250 341054 620284
rect 341020 620160 341054 620194
rect 334681 620070 334715 620104
rect 334782 620047 334816 620081
rect 334872 620047 334906 620081
rect 334962 620047 334996 620081
rect 335052 620047 335086 620081
rect 335142 620047 335176 620081
rect 335232 620047 335266 620081
rect 335322 620047 335356 620081
rect 335412 620047 335446 620081
rect 335502 620047 335536 620081
rect 335592 620047 335626 620081
rect 335682 620047 335716 620081
rect 335772 620047 335806 620081
rect 335868 620070 335902 620104
rect 335969 620070 336003 620104
rect 336070 620047 336104 620081
rect 336160 620047 336194 620081
rect 336250 620047 336284 620081
rect 336340 620047 336374 620081
rect 336430 620047 336464 620081
rect 336520 620047 336554 620081
rect 336610 620047 336644 620081
rect 336700 620047 336734 620081
rect 336790 620047 336824 620081
rect 336880 620047 336914 620081
rect 336970 620047 337004 620081
rect 337060 620047 337094 620081
rect 337156 620070 337190 620104
rect 337257 620070 337291 620104
rect 337358 620047 337392 620081
rect 337448 620047 337482 620081
rect 337538 620047 337572 620081
rect 337628 620047 337662 620081
rect 337718 620047 337752 620081
rect 337808 620047 337842 620081
rect 337898 620047 337932 620081
rect 337988 620047 338022 620081
rect 338078 620047 338112 620081
rect 338168 620047 338202 620081
rect 338258 620047 338292 620081
rect 338348 620047 338382 620081
rect 338444 620070 338478 620104
rect 338545 620070 338579 620104
rect 338646 620047 338680 620081
rect 338736 620047 338770 620081
rect 338826 620047 338860 620081
rect 338916 620047 338950 620081
rect 339006 620047 339040 620081
rect 339096 620047 339130 620081
rect 339186 620047 339220 620081
rect 339276 620047 339310 620081
rect 339366 620047 339400 620081
rect 339456 620047 339490 620081
rect 339546 620047 339580 620081
rect 339636 620047 339670 620081
rect 339732 620070 339766 620104
rect 339833 620070 339867 620104
rect 339934 620047 339968 620081
rect 340024 620047 340058 620081
rect 340114 620047 340148 620081
rect 340204 620047 340238 620081
rect 340294 620047 340328 620081
rect 340384 620047 340418 620081
rect 340474 620047 340508 620081
rect 340564 620047 340598 620081
rect 340654 620047 340688 620081
rect 340744 620047 340778 620081
rect 340834 620047 340868 620081
rect 340924 620047 340958 620081
rect 341020 620070 341054 620104
rect 334782 619946 334816 619980
rect 334872 619946 334906 619980
rect 334962 619946 334996 619980
rect 335052 619946 335086 619980
rect 335142 619946 335176 619980
rect 335232 619946 335266 619980
rect 335322 619946 335356 619980
rect 335412 619946 335446 619980
rect 335502 619946 335536 619980
rect 335592 619946 335626 619980
rect 335682 619946 335716 619980
rect 335772 619946 335806 619980
rect 336070 619946 336104 619980
rect 336160 619946 336194 619980
rect 336250 619946 336284 619980
rect 336340 619946 336374 619980
rect 336430 619946 336464 619980
rect 336520 619946 336554 619980
rect 336610 619946 336644 619980
rect 336700 619946 336734 619980
rect 336790 619946 336824 619980
rect 336880 619946 336914 619980
rect 336970 619946 337004 619980
rect 337060 619946 337094 619980
rect 337358 619946 337392 619980
rect 337448 619946 337482 619980
rect 337538 619946 337572 619980
rect 337628 619946 337662 619980
rect 337718 619946 337752 619980
rect 337808 619946 337842 619980
rect 337898 619946 337932 619980
rect 337988 619946 338022 619980
rect 338078 619946 338112 619980
rect 338168 619946 338202 619980
rect 338258 619946 338292 619980
rect 338348 619946 338382 619980
rect 338646 619946 338680 619980
rect 338736 619946 338770 619980
rect 338826 619946 338860 619980
rect 338916 619946 338950 619980
rect 339006 619946 339040 619980
rect 339096 619946 339130 619980
rect 339186 619946 339220 619980
rect 339276 619946 339310 619980
rect 339366 619946 339400 619980
rect 339456 619946 339490 619980
rect 339546 619946 339580 619980
rect 339636 619946 339670 619980
rect 339934 619946 339968 619980
rect 340024 619946 340058 619980
rect 340114 619946 340148 619980
rect 340204 619946 340238 619980
rect 340294 619946 340328 619980
rect 340384 619946 340418 619980
rect 340474 619946 340508 619980
rect 340564 619946 340598 619980
rect 340654 619946 340688 619980
rect 340744 619946 340778 619980
rect 340834 619946 340868 619980
rect 340924 619946 340958 619980
rect 334681 619862 334715 619896
rect 335868 619862 335902 619896
rect 335969 619862 336003 619896
rect 334681 619772 334715 619806
rect 334681 619682 334715 619716
rect 334681 619592 334715 619626
rect 334681 619502 334715 619536
rect 334681 619412 334715 619446
rect 334681 619322 334715 619356
rect 334681 619232 334715 619266
rect 334681 619142 334715 619176
rect 334681 619052 334715 619086
rect 334681 618962 334715 618996
rect 334681 618872 334715 618906
rect 337156 619862 337190 619896
rect 337257 619862 337291 619896
rect 335868 619772 335902 619806
rect 335969 619772 336003 619806
rect 335868 619682 335902 619716
rect 335969 619682 336003 619716
rect 335868 619592 335902 619626
rect 335969 619592 336003 619626
rect 335868 619502 335902 619536
rect 335969 619502 336003 619536
rect 335868 619412 335902 619446
rect 335969 619412 336003 619446
rect 335868 619322 335902 619356
rect 335969 619322 336003 619356
rect 335868 619232 335902 619266
rect 335969 619232 336003 619266
rect 335868 619142 335902 619176
rect 335969 619142 336003 619176
rect 335868 619052 335902 619086
rect 335969 619052 336003 619086
rect 335868 618962 335902 618996
rect 335969 618962 336003 618996
rect 335868 618872 335902 618906
rect 335969 618872 336003 618906
rect 338444 619862 338478 619896
rect 338545 619862 338579 619896
rect 337156 619772 337190 619806
rect 337257 619772 337291 619806
rect 337156 619682 337190 619716
rect 337257 619682 337291 619716
rect 337156 619592 337190 619626
rect 337257 619592 337291 619626
rect 337156 619502 337190 619536
rect 337257 619502 337291 619536
rect 337156 619412 337190 619446
rect 337257 619412 337291 619446
rect 337156 619322 337190 619356
rect 337257 619322 337291 619356
rect 337156 619232 337190 619266
rect 337257 619232 337291 619266
rect 337156 619142 337190 619176
rect 337257 619142 337291 619176
rect 337156 619052 337190 619086
rect 337257 619052 337291 619086
rect 337156 618962 337190 618996
rect 337257 618962 337291 618996
rect 337156 618872 337190 618906
rect 337257 618872 337291 618906
rect 339732 619862 339766 619896
rect 339833 619862 339867 619896
rect 338444 619772 338478 619806
rect 338545 619772 338579 619806
rect 338444 619682 338478 619716
rect 338545 619682 338579 619716
rect 338444 619592 338478 619626
rect 338545 619592 338579 619626
rect 338444 619502 338478 619536
rect 338545 619502 338579 619536
rect 338444 619412 338478 619446
rect 338545 619412 338579 619446
rect 338444 619322 338478 619356
rect 338545 619322 338579 619356
rect 338444 619232 338478 619266
rect 338545 619232 338579 619266
rect 338444 619142 338478 619176
rect 338545 619142 338579 619176
rect 338444 619052 338478 619086
rect 338545 619052 338579 619086
rect 338444 618962 338478 618996
rect 338545 618962 338579 618996
rect 338444 618872 338478 618906
rect 338545 618872 338579 618906
rect 341020 619862 341054 619896
rect 339732 619772 339766 619806
rect 339833 619772 339867 619806
rect 339732 619682 339766 619716
rect 339833 619682 339867 619716
rect 339732 619592 339766 619626
rect 339833 619592 339867 619626
rect 339732 619502 339766 619536
rect 339833 619502 339867 619536
rect 339732 619412 339766 619446
rect 339833 619412 339867 619446
rect 339732 619322 339766 619356
rect 339833 619322 339867 619356
rect 339732 619232 339766 619266
rect 339833 619232 339867 619266
rect 339732 619142 339766 619176
rect 339833 619142 339867 619176
rect 339732 619052 339766 619086
rect 339833 619052 339867 619086
rect 339732 618962 339766 618996
rect 339833 618962 339867 618996
rect 339732 618872 339766 618906
rect 339833 618872 339867 618906
rect 341020 619772 341054 619806
rect 341020 619682 341054 619716
rect 341020 619592 341054 619626
rect 341020 619502 341054 619536
rect 341020 619412 341054 619446
rect 341020 619322 341054 619356
rect 341020 619232 341054 619266
rect 341020 619142 341054 619176
rect 341020 619052 341054 619086
rect 341020 618962 341054 618996
rect 341020 618872 341054 618906
rect 334681 618782 334715 618816
rect 334782 618759 334816 618793
rect 334872 618759 334906 618793
rect 334962 618759 334996 618793
rect 335052 618759 335086 618793
rect 335142 618759 335176 618793
rect 335232 618759 335266 618793
rect 335322 618759 335356 618793
rect 335412 618759 335446 618793
rect 335502 618759 335536 618793
rect 335592 618759 335626 618793
rect 335682 618759 335716 618793
rect 335772 618759 335806 618793
rect 335868 618782 335902 618816
rect 335969 618782 336003 618816
rect 336070 618759 336104 618793
rect 336160 618759 336194 618793
rect 336250 618759 336284 618793
rect 336340 618759 336374 618793
rect 336430 618759 336464 618793
rect 336520 618759 336554 618793
rect 336610 618759 336644 618793
rect 336700 618759 336734 618793
rect 336790 618759 336824 618793
rect 336880 618759 336914 618793
rect 336970 618759 337004 618793
rect 337060 618759 337094 618793
rect 337156 618782 337190 618816
rect 337257 618782 337291 618816
rect 337358 618759 337392 618793
rect 337448 618759 337482 618793
rect 337538 618759 337572 618793
rect 337628 618759 337662 618793
rect 337718 618759 337752 618793
rect 337808 618759 337842 618793
rect 337898 618759 337932 618793
rect 337988 618759 338022 618793
rect 338078 618759 338112 618793
rect 338168 618759 338202 618793
rect 338258 618759 338292 618793
rect 338348 618759 338382 618793
rect 338444 618782 338478 618816
rect 338545 618782 338579 618816
rect 338646 618759 338680 618793
rect 338736 618759 338770 618793
rect 338826 618759 338860 618793
rect 338916 618759 338950 618793
rect 339006 618759 339040 618793
rect 339096 618759 339130 618793
rect 339186 618759 339220 618793
rect 339276 618759 339310 618793
rect 339366 618759 339400 618793
rect 339456 618759 339490 618793
rect 339546 618759 339580 618793
rect 339636 618759 339670 618793
rect 339732 618782 339766 618816
rect 339833 618782 339867 618816
rect 339934 618759 339968 618793
rect 340024 618759 340058 618793
rect 340114 618759 340148 618793
rect 340204 618759 340238 618793
rect 340294 618759 340328 618793
rect 340384 618759 340418 618793
rect 340474 618759 340508 618793
rect 340564 618759 340598 618793
rect 340654 618759 340688 618793
rect 340744 618759 340778 618793
rect 340834 618759 340868 618793
rect 340924 618759 340958 618793
rect 341020 618782 341054 618816
rect 334782 618658 334816 618692
rect 334872 618658 334906 618692
rect 334962 618658 334996 618692
rect 335052 618658 335086 618692
rect 335142 618658 335176 618692
rect 335232 618658 335266 618692
rect 335322 618658 335356 618692
rect 335412 618658 335446 618692
rect 335502 618658 335536 618692
rect 335592 618658 335626 618692
rect 335682 618658 335716 618692
rect 335772 618658 335806 618692
rect 336070 618658 336104 618692
rect 336160 618658 336194 618692
rect 336250 618658 336284 618692
rect 336340 618658 336374 618692
rect 336430 618658 336464 618692
rect 336520 618658 336554 618692
rect 336610 618658 336644 618692
rect 336700 618658 336734 618692
rect 336790 618658 336824 618692
rect 336880 618658 336914 618692
rect 336970 618658 337004 618692
rect 337060 618658 337094 618692
rect 337358 618658 337392 618692
rect 337448 618658 337482 618692
rect 337538 618658 337572 618692
rect 337628 618658 337662 618692
rect 337718 618658 337752 618692
rect 337808 618658 337842 618692
rect 337898 618658 337932 618692
rect 337988 618658 338022 618692
rect 338078 618658 338112 618692
rect 338168 618658 338202 618692
rect 338258 618658 338292 618692
rect 338348 618658 338382 618692
rect 338646 618658 338680 618692
rect 338736 618658 338770 618692
rect 338826 618658 338860 618692
rect 338916 618658 338950 618692
rect 339006 618658 339040 618692
rect 339096 618658 339130 618692
rect 339186 618658 339220 618692
rect 339276 618658 339310 618692
rect 339366 618658 339400 618692
rect 339456 618658 339490 618692
rect 339546 618658 339580 618692
rect 339636 618658 339670 618692
rect 339934 618658 339968 618692
rect 340024 618658 340058 618692
rect 340114 618658 340148 618692
rect 340204 618658 340238 618692
rect 340294 618658 340328 618692
rect 340384 618658 340418 618692
rect 340474 618658 340508 618692
rect 340564 618658 340598 618692
rect 340654 618658 340688 618692
rect 340744 618658 340778 618692
rect 340834 618658 340868 618692
rect 340924 618658 340958 618692
rect 334681 618574 334715 618608
rect 335868 618574 335902 618608
rect 335969 618574 336003 618608
rect 334681 618484 334715 618518
rect 334681 618394 334715 618428
rect 334681 618304 334715 618338
rect 334681 618214 334715 618248
rect 334681 618124 334715 618158
rect 334681 618034 334715 618068
rect 334681 617944 334715 617978
rect 334681 617854 334715 617888
rect 334681 617764 334715 617798
rect 334681 617674 334715 617708
rect 334681 617584 334715 617618
rect 337156 618574 337190 618608
rect 337257 618574 337291 618608
rect 335868 618484 335902 618518
rect 335969 618484 336003 618518
rect 335868 618394 335902 618428
rect 335969 618394 336003 618428
rect 335868 618304 335902 618338
rect 335969 618304 336003 618338
rect 335868 618214 335902 618248
rect 335969 618214 336003 618248
rect 335868 618124 335902 618158
rect 335969 618124 336003 618158
rect 335868 618034 335902 618068
rect 335969 618034 336003 618068
rect 335868 617944 335902 617978
rect 335969 617944 336003 617978
rect 335868 617854 335902 617888
rect 335969 617854 336003 617888
rect 335868 617764 335902 617798
rect 335969 617764 336003 617798
rect 335868 617674 335902 617708
rect 335969 617674 336003 617708
rect 335868 617584 335902 617618
rect 335969 617584 336003 617618
rect 338444 618574 338478 618608
rect 338545 618574 338579 618608
rect 337156 618484 337190 618518
rect 337257 618484 337291 618518
rect 337156 618394 337190 618428
rect 337257 618394 337291 618428
rect 337156 618304 337190 618338
rect 337257 618304 337291 618338
rect 337156 618214 337190 618248
rect 337257 618214 337291 618248
rect 337156 618124 337190 618158
rect 337257 618124 337291 618158
rect 337156 618034 337190 618068
rect 337257 618034 337291 618068
rect 337156 617944 337190 617978
rect 337257 617944 337291 617978
rect 337156 617854 337190 617888
rect 337257 617854 337291 617888
rect 337156 617764 337190 617798
rect 337257 617764 337291 617798
rect 337156 617674 337190 617708
rect 337257 617674 337291 617708
rect 337156 617584 337190 617618
rect 337257 617584 337291 617618
rect 339732 618574 339766 618608
rect 339833 618574 339867 618608
rect 338444 618484 338478 618518
rect 338545 618484 338579 618518
rect 338444 618394 338478 618428
rect 338545 618394 338579 618428
rect 338444 618304 338478 618338
rect 338545 618304 338579 618338
rect 338444 618214 338478 618248
rect 338545 618214 338579 618248
rect 338444 618124 338478 618158
rect 338545 618124 338579 618158
rect 338444 618034 338478 618068
rect 338545 618034 338579 618068
rect 338444 617944 338478 617978
rect 338545 617944 338579 617978
rect 338444 617854 338478 617888
rect 338545 617854 338579 617888
rect 338444 617764 338478 617798
rect 338545 617764 338579 617798
rect 338444 617674 338478 617708
rect 338545 617674 338579 617708
rect 338444 617584 338478 617618
rect 338545 617584 338579 617618
rect 341020 618574 341054 618608
rect 339732 618484 339766 618518
rect 339833 618484 339867 618518
rect 339732 618394 339766 618428
rect 339833 618394 339867 618428
rect 339732 618304 339766 618338
rect 339833 618304 339867 618338
rect 339732 618214 339766 618248
rect 339833 618214 339867 618248
rect 339732 618124 339766 618158
rect 339833 618124 339867 618158
rect 339732 618034 339766 618068
rect 339833 618034 339867 618068
rect 339732 617944 339766 617978
rect 339833 617944 339867 617978
rect 339732 617854 339766 617888
rect 339833 617854 339867 617888
rect 339732 617764 339766 617798
rect 339833 617764 339867 617798
rect 339732 617674 339766 617708
rect 339833 617674 339867 617708
rect 339732 617584 339766 617618
rect 339833 617584 339867 617618
rect 341020 618484 341054 618518
rect 341020 618394 341054 618428
rect 341020 618304 341054 618338
rect 341020 618214 341054 618248
rect 341020 618124 341054 618158
rect 341020 618034 341054 618068
rect 341020 617944 341054 617978
rect 341020 617854 341054 617888
rect 341020 617764 341054 617798
rect 341020 617674 341054 617708
rect 341020 617584 341054 617618
rect 334681 617494 334715 617528
rect 334782 617471 334816 617505
rect 334872 617471 334906 617505
rect 334962 617471 334996 617505
rect 335052 617471 335086 617505
rect 335142 617471 335176 617505
rect 335232 617471 335266 617505
rect 335322 617471 335356 617505
rect 335412 617471 335446 617505
rect 335502 617471 335536 617505
rect 335592 617471 335626 617505
rect 335682 617471 335716 617505
rect 335772 617471 335806 617505
rect 335868 617494 335902 617528
rect 335969 617494 336003 617528
rect 336070 617471 336104 617505
rect 336160 617471 336194 617505
rect 336250 617471 336284 617505
rect 336340 617471 336374 617505
rect 336430 617471 336464 617505
rect 336520 617471 336554 617505
rect 336610 617471 336644 617505
rect 336700 617471 336734 617505
rect 336790 617471 336824 617505
rect 336880 617471 336914 617505
rect 336970 617471 337004 617505
rect 337060 617471 337094 617505
rect 337156 617494 337190 617528
rect 337257 617494 337291 617528
rect 337358 617471 337392 617505
rect 337448 617471 337482 617505
rect 337538 617471 337572 617505
rect 337628 617471 337662 617505
rect 337718 617471 337752 617505
rect 337808 617471 337842 617505
rect 337898 617471 337932 617505
rect 337988 617471 338022 617505
rect 338078 617471 338112 617505
rect 338168 617471 338202 617505
rect 338258 617471 338292 617505
rect 338348 617471 338382 617505
rect 338444 617494 338478 617528
rect 338545 617494 338579 617528
rect 338646 617471 338680 617505
rect 338736 617471 338770 617505
rect 338826 617471 338860 617505
rect 338916 617471 338950 617505
rect 339006 617471 339040 617505
rect 339096 617471 339130 617505
rect 339186 617471 339220 617505
rect 339276 617471 339310 617505
rect 339366 617471 339400 617505
rect 339456 617471 339490 617505
rect 339546 617471 339580 617505
rect 339636 617471 339670 617505
rect 339732 617494 339766 617528
rect 339833 617494 339867 617528
rect 339934 617471 339968 617505
rect 340024 617471 340058 617505
rect 340114 617471 340148 617505
rect 340204 617471 340238 617505
rect 340294 617471 340328 617505
rect 340384 617471 340418 617505
rect 340474 617471 340508 617505
rect 340564 617471 340598 617505
rect 340654 617471 340688 617505
rect 340744 617471 340778 617505
rect 340834 617471 340868 617505
rect 340924 617471 340958 617505
rect 341020 617494 341054 617528
rect 297848 614448 341088 615448
rect 342112 614424 343112 640648
<< nsubdiffcont >>
rect 334922 627524 334956 627558
rect 335012 627524 335046 627558
rect 335102 627524 335136 627558
rect 335192 627524 335226 627558
rect 335282 627524 335316 627558
rect 335372 627524 335406 627558
rect 335462 627524 335496 627558
rect 335552 627524 335586 627558
rect 335642 627524 335676 627558
rect 334830 627430 334864 627464
rect 334830 627340 334864 627374
rect 334830 627250 334864 627284
rect 334830 627160 334864 627194
rect 334830 627070 334864 627104
rect 334830 626980 334864 627014
rect 334830 626890 334864 626924
rect 334830 626800 334864 626834
rect 335720 627411 335754 627445
rect 335720 627321 335754 627355
rect 335720 627231 335754 627265
rect 335720 627141 335754 627175
rect 335720 627051 335754 627085
rect 335720 626961 335754 626995
rect 335720 626871 335754 626905
rect 335720 626781 335754 626815
rect 334830 626710 334864 626744
rect 335720 626691 335754 626725
rect 334888 626634 334922 626668
rect 334978 626634 335012 626668
rect 335068 626634 335102 626668
rect 335158 626634 335192 626668
rect 335248 626634 335282 626668
rect 335338 626634 335372 626668
rect 335428 626634 335462 626668
rect 335518 626634 335552 626668
rect 335608 626634 335642 626668
rect 336210 627524 336244 627558
rect 336300 627524 336334 627558
rect 336390 627524 336424 627558
rect 336480 627524 336514 627558
rect 336570 627524 336604 627558
rect 336660 627524 336694 627558
rect 336750 627524 336784 627558
rect 336840 627524 336874 627558
rect 336930 627524 336964 627558
rect 336118 627430 336152 627464
rect 336118 627340 336152 627374
rect 336118 627250 336152 627284
rect 336118 627160 336152 627194
rect 336118 627070 336152 627104
rect 336118 626980 336152 627014
rect 336118 626890 336152 626924
rect 336118 626800 336152 626834
rect 337008 627411 337042 627445
rect 337008 627321 337042 627355
rect 337008 627231 337042 627265
rect 337008 627141 337042 627175
rect 337008 627051 337042 627085
rect 337008 626961 337042 626995
rect 337008 626871 337042 626905
rect 337008 626781 337042 626815
rect 336118 626710 336152 626744
rect 337008 626691 337042 626725
rect 336176 626634 336210 626668
rect 336266 626634 336300 626668
rect 336356 626634 336390 626668
rect 336446 626634 336480 626668
rect 336536 626634 336570 626668
rect 336626 626634 336660 626668
rect 336716 626634 336750 626668
rect 336806 626634 336840 626668
rect 336896 626634 336930 626668
rect 337498 627524 337532 627558
rect 337588 627524 337622 627558
rect 337678 627524 337712 627558
rect 337768 627524 337802 627558
rect 337858 627524 337892 627558
rect 337948 627524 337982 627558
rect 338038 627524 338072 627558
rect 338128 627524 338162 627558
rect 338218 627524 338252 627558
rect 337406 627430 337440 627464
rect 337406 627340 337440 627374
rect 337406 627250 337440 627284
rect 337406 627160 337440 627194
rect 337406 627070 337440 627104
rect 337406 626980 337440 627014
rect 337406 626890 337440 626924
rect 337406 626800 337440 626834
rect 338296 627411 338330 627445
rect 338296 627321 338330 627355
rect 338296 627231 338330 627265
rect 338296 627141 338330 627175
rect 338296 627051 338330 627085
rect 338296 626961 338330 626995
rect 338296 626871 338330 626905
rect 338296 626781 338330 626815
rect 337406 626710 337440 626744
rect 338296 626691 338330 626725
rect 337464 626634 337498 626668
rect 337554 626634 337588 626668
rect 337644 626634 337678 626668
rect 337734 626634 337768 626668
rect 337824 626634 337858 626668
rect 337914 626634 337948 626668
rect 338004 626634 338038 626668
rect 338094 626634 338128 626668
rect 338184 626634 338218 626668
rect 338786 627524 338820 627558
rect 338876 627524 338910 627558
rect 338966 627524 339000 627558
rect 339056 627524 339090 627558
rect 339146 627524 339180 627558
rect 339236 627524 339270 627558
rect 339326 627524 339360 627558
rect 339416 627524 339450 627558
rect 339506 627524 339540 627558
rect 338694 627430 338728 627464
rect 338694 627340 338728 627374
rect 338694 627250 338728 627284
rect 338694 627160 338728 627194
rect 338694 627070 338728 627104
rect 338694 626980 338728 627014
rect 338694 626890 338728 626924
rect 338694 626800 338728 626834
rect 339584 627411 339618 627445
rect 339584 627321 339618 627355
rect 339584 627231 339618 627265
rect 339584 627141 339618 627175
rect 339584 627051 339618 627085
rect 339584 626961 339618 626995
rect 339584 626871 339618 626905
rect 339584 626781 339618 626815
rect 338694 626710 338728 626744
rect 339584 626691 339618 626725
rect 338752 626634 338786 626668
rect 338842 626634 338876 626668
rect 338932 626634 338966 626668
rect 339022 626634 339056 626668
rect 339112 626634 339146 626668
rect 339202 626634 339236 626668
rect 339292 626634 339326 626668
rect 339382 626634 339416 626668
rect 339472 626634 339506 626668
rect 340074 627524 340108 627558
rect 340164 627524 340198 627558
rect 340254 627524 340288 627558
rect 340344 627524 340378 627558
rect 340434 627524 340468 627558
rect 340524 627524 340558 627558
rect 340614 627524 340648 627558
rect 340704 627524 340738 627558
rect 340794 627524 340828 627558
rect 339982 627430 340016 627464
rect 339982 627340 340016 627374
rect 339982 627250 340016 627284
rect 339982 627160 340016 627194
rect 339982 627070 340016 627104
rect 339982 626980 340016 627014
rect 339982 626890 340016 626924
rect 339982 626800 340016 626834
rect 340872 627411 340906 627445
rect 340872 627321 340906 627355
rect 340872 627231 340906 627265
rect 340872 627141 340906 627175
rect 340872 627051 340906 627085
rect 340872 626961 340906 626995
rect 340872 626871 340906 626905
rect 340872 626781 340906 626815
rect 339982 626710 340016 626744
rect 340872 626691 340906 626725
rect 340040 626634 340074 626668
rect 340130 626634 340164 626668
rect 340220 626634 340254 626668
rect 340310 626634 340344 626668
rect 340400 626634 340434 626668
rect 340490 626634 340524 626668
rect 340580 626634 340614 626668
rect 340670 626634 340704 626668
rect 340760 626634 340794 626668
rect 334922 626236 334956 626270
rect 335012 626236 335046 626270
rect 335102 626236 335136 626270
rect 335192 626236 335226 626270
rect 335282 626236 335316 626270
rect 335372 626236 335406 626270
rect 335462 626236 335496 626270
rect 335552 626236 335586 626270
rect 335642 626236 335676 626270
rect 334830 626142 334864 626176
rect 334830 626052 334864 626086
rect 334830 625962 334864 625996
rect 334830 625872 334864 625906
rect 334830 625782 334864 625816
rect 334830 625692 334864 625726
rect 334830 625602 334864 625636
rect 334830 625512 334864 625546
rect 335720 626123 335754 626157
rect 335720 626033 335754 626067
rect 335720 625943 335754 625977
rect 335720 625853 335754 625887
rect 335720 625763 335754 625797
rect 335720 625673 335754 625707
rect 335720 625583 335754 625617
rect 335720 625493 335754 625527
rect 334830 625422 334864 625456
rect 335720 625403 335754 625437
rect 334888 625346 334922 625380
rect 334978 625346 335012 625380
rect 335068 625346 335102 625380
rect 335158 625346 335192 625380
rect 335248 625346 335282 625380
rect 335338 625346 335372 625380
rect 335428 625346 335462 625380
rect 335518 625346 335552 625380
rect 335608 625346 335642 625380
rect 336210 626236 336244 626270
rect 336300 626236 336334 626270
rect 336390 626236 336424 626270
rect 336480 626236 336514 626270
rect 336570 626236 336604 626270
rect 336660 626236 336694 626270
rect 336750 626236 336784 626270
rect 336840 626236 336874 626270
rect 336930 626236 336964 626270
rect 336118 626142 336152 626176
rect 336118 626052 336152 626086
rect 336118 625962 336152 625996
rect 336118 625872 336152 625906
rect 336118 625782 336152 625816
rect 336118 625692 336152 625726
rect 336118 625602 336152 625636
rect 336118 625512 336152 625546
rect 337008 626123 337042 626157
rect 337008 626033 337042 626067
rect 337008 625943 337042 625977
rect 337008 625853 337042 625887
rect 337008 625763 337042 625797
rect 337008 625673 337042 625707
rect 337008 625583 337042 625617
rect 337008 625493 337042 625527
rect 336118 625422 336152 625456
rect 337008 625403 337042 625437
rect 336176 625346 336210 625380
rect 336266 625346 336300 625380
rect 336356 625346 336390 625380
rect 336446 625346 336480 625380
rect 336536 625346 336570 625380
rect 336626 625346 336660 625380
rect 336716 625346 336750 625380
rect 336806 625346 336840 625380
rect 336896 625346 336930 625380
rect 337498 626236 337532 626270
rect 337588 626236 337622 626270
rect 337678 626236 337712 626270
rect 337768 626236 337802 626270
rect 337858 626236 337892 626270
rect 337948 626236 337982 626270
rect 338038 626236 338072 626270
rect 338128 626236 338162 626270
rect 338218 626236 338252 626270
rect 337406 626142 337440 626176
rect 337406 626052 337440 626086
rect 337406 625962 337440 625996
rect 337406 625872 337440 625906
rect 337406 625782 337440 625816
rect 337406 625692 337440 625726
rect 337406 625602 337440 625636
rect 337406 625512 337440 625546
rect 338296 626123 338330 626157
rect 338296 626033 338330 626067
rect 338296 625943 338330 625977
rect 338296 625853 338330 625887
rect 338296 625763 338330 625797
rect 338296 625673 338330 625707
rect 338296 625583 338330 625617
rect 338296 625493 338330 625527
rect 337406 625422 337440 625456
rect 338296 625403 338330 625437
rect 337464 625346 337498 625380
rect 337554 625346 337588 625380
rect 337644 625346 337678 625380
rect 337734 625346 337768 625380
rect 337824 625346 337858 625380
rect 337914 625346 337948 625380
rect 338004 625346 338038 625380
rect 338094 625346 338128 625380
rect 338184 625346 338218 625380
rect 338786 626236 338820 626270
rect 338876 626236 338910 626270
rect 338966 626236 339000 626270
rect 339056 626236 339090 626270
rect 339146 626236 339180 626270
rect 339236 626236 339270 626270
rect 339326 626236 339360 626270
rect 339416 626236 339450 626270
rect 339506 626236 339540 626270
rect 338694 626142 338728 626176
rect 338694 626052 338728 626086
rect 338694 625962 338728 625996
rect 338694 625872 338728 625906
rect 338694 625782 338728 625816
rect 338694 625692 338728 625726
rect 338694 625602 338728 625636
rect 338694 625512 338728 625546
rect 339584 626123 339618 626157
rect 339584 626033 339618 626067
rect 339584 625943 339618 625977
rect 339584 625853 339618 625887
rect 339584 625763 339618 625797
rect 339584 625673 339618 625707
rect 339584 625583 339618 625617
rect 339584 625493 339618 625527
rect 338694 625422 338728 625456
rect 339584 625403 339618 625437
rect 338752 625346 338786 625380
rect 338842 625346 338876 625380
rect 338932 625346 338966 625380
rect 339022 625346 339056 625380
rect 339112 625346 339146 625380
rect 339202 625346 339236 625380
rect 339292 625346 339326 625380
rect 339382 625346 339416 625380
rect 339472 625346 339506 625380
rect 340074 626236 340108 626270
rect 340164 626236 340198 626270
rect 340254 626236 340288 626270
rect 340344 626236 340378 626270
rect 340434 626236 340468 626270
rect 340524 626236 340558 626270
rect 340614 626236 340648 626270
rect 340704 626236 340738 626270
rect 340794 626236 340828 626270
rect 339982 626142 340016 626176
rect 339982 626052 340016 626086
rect 339982 625962 340016 625996
rect 339982 625872 340016 625906
rect 339982 625782 340016 625816
rect 339982 625692 340016 625726
rect 339982 625602 340016 625636
rect 339982 625512 340016 625546
rect 340872 626123 340906 626157
rect 340872 626033 340906 626067
rect 340872 625943 340906 625977
rect 340872 625853 340906 625887
rect 340872 625763 340906 625797
rect 340872 625673 340906 625707
rect 340872 625583 340906 625617
rect 340872 625493 340906 625527
rect 339982 625422 340016 625456
rect 340872 625403 340906 625437
rect 340040 625346 340074 625380
rect 340130 625346 340164 625380
rect 340220 625346 340254 625380
rect 340310 625346 340344 625380
rect 340400 625346 340434 625380
rect 340490 625346 340524 625380
rect 340580 625346 340614 625380
rect 340670 625346 340704 625380
rect 340760 625346 340794 625380
rect 302954 617306 303054 619648
rect 312082 617306 312182 619648
rect 312904 617608 313104 624608
rect 318814 617608 319014 624608
rect 324314 617608 324514 624608
rect 330270 617606 330470 624606
rect 334922 624948 334956 624982
rect 335012 624948 335046 624982
rect 335102 624948 335136 624982
rect 335192 624948 335226 624982
rect 335282 624948 335316 624982
rect 335372 624948 335406 624982
rect 335462 624948 335496 624982
rect 335552 624948 335586 624982
rect 335642 624948 335676 624982
rect 334830 624854 334864 624888
rect 334830 624764 334864 624798
rect 334830 624674 334864 624708
rect 334830 624584 334864 624618
rect 334830 624494 334864 624528
rect 334830 624404 334864 624438
rect 334830 624314 334864 624348
rect 334830 624224 334864 624258
rect 335720 624835 335754 624869
rect 335720 624745 335754 624779
rect 335720 624655 335754 624689
rect 335720 624565 335754 624599
rect 335720 624475 335754 624509
rect 335720 624385 335754 624419
rect 335720 624295 335754 624329
rect 335720 624205 335754 624239
rect 334830 624134 334864 624168
rect 335720 624115 335754 624149
rect 334888 624058 334922 624092
rect 334978 624058 335012 624092
rect 335068 624058 335102 624092
rect 335158 624058 335192 624092
rect 335248 624058 335282 624092
rect 335338 624058 335372 624092
rect 335428 624058 335462 624092
rect 335518 624058 335552 624092
rect 335608 624058 335642 624092
rect 336210 624948 336244 624982
rect 336300 624948 336334 624982
rect 336390 624948 336424 624982
rect 336480 624948 336514 624982
rect 336570 624948 336604 624982
rect 336660 624948 336694 624982
rect 336750 624948 336784 624982
rect 336840 624948 336874 624982
rect 336930 624948 336964 624982
rect 336118 624854 336152 624888
rect 336118 624764 336152 624798
rect 336118 624674 336152 624708
rect 336118 624584 336152 624618
rect 336118 624494 336152 624528
rect 336118 624404 336152 624438
rect 336118 624314 336152 624348
rect 336118 624224 336152 624258
rect 337008 624835 337042 624869
rect 337008 624745 337042 624779
rect 337008 624655 337042 624689
rect 337008 624565 337042 624599
rect 337008 624475 337042 624509
rect 337008 624385 337042 624419
rect 337008 624295 337042 624329
rect 337008 624205 337042 624239
rect 336118 624134 336152 624168
rect 337008 624115 337042 624149
rect 336176 624058 336210 624092
rect 336266 624058 336300 624092
rect 336356 624058 336390 624092
rect 336446 624058 336480 624092
rect 336536 624058 336570 624092
rect 336626 624058 336660 624092
rect 336716 624058 336750 624092
rect 336806 624058 336840 624092
rect 336896 624058 336930 624092
rect 337498 624948 337532 624982
rect 337588 624948 337622 624982
rect 337678 624948 337712 624982
rect 337768 624948 337802 624982
rect 337858 624948 337892 624982
rect 337948 624948 337982 624982
rect 338038 624948 338072 624982
rect 338128 624948 338162 624982
rect 338218 624948 338252 624982
rect 337406 624854 337440 624888
rect 337406 624764 337440 624798
rect 337406 624674 337440 624708
rect 337406 624584 337440 624618
rect 337406 624494 337440 624528
rect 337406 624404 337440 624438
rect 337406 624314 337440 624348
rect 337406 624224 337440 624258
rect 338296 624835 338330 624869
rect 338296 624745 338330 624779
rect 338296 624655 338330 624689
rect 338296 624565 338330 624599
rect 338296 624475 338330 624509
rect 338296 624385 338330 624419
rect 338296 624295 338330 624329
rect 338296 624205 338330 624239
rect 337406 624134 337440 624168
rect 338296 624115 338330 624149
rect 337464 624058 337498 624092
rect 337554 624058 337588 624092
rect 337644 624058 337678 624092
rect 337734 624058 337768 624092
rect 337824 624058 337858 624092
rect 337914 624058 337948 624092
rect 338004 624058 338038 624092
rect 338094 624058 338128 624092
rect 338184 624058 338218 624092
rect 338786 624948 338820 624982
rect 338876 624948 338910 624982
rect 338966 624948 339000 624982
rect 339056 624948 339090 624982
rect 339146 624948 339180 624982
rect 339236 624948 339270 624982
rect 339326 624948 339360 624982
rect 339416 624948 339450 624982
rect 339506 624948 339540 624982
rect 338694 624854 338728 624888
rect 338694 624764 338728 624798
rect 338694 624674 338728 624708
rect 338694 624584 338728 624618
rect 338694 624494 338728 624528
rect 338694 624404 338728 624438
rect 338694 624314 338728 624348
rect 338694 624224 338728 624258
rect 339584 624835 339618 624869
rect 339584 624745 339618 624779
rect 339584 624655 339618 624689
rect 339584 624565 339618 624599
rect 339584 624475 339618 624509
rect 339584 624385 339618 624419
rect 339584 624295 339618 624329
rect 339584 624205 339618 624239
rect 338694 624134 338728 624168
rect 339584 624115 339618 624149
rect 338752 624058 338786 624092
rect 338842 624058 338876 624092
rect 338932 624058 338966 624092
rect 339022 624058 339056 624092
rect 339112 624058 339146 624092
rect 339202 624058 339236 624092
rect 339292 624058 339326 624092
rect 339382 624058 339416 624092
rect 339472 624058 339506 624092
rect 340074 624948 340108 624982
rect 340164 624948 340198 624982
rect 340254 624948 340288 624982
rect 340344 624948 340378 624982
rect 340434 624948 340468 624982
rect 340524 624948 340558 624982
rect 340614 624948 340648 624982
rect 340704 624948 340738 624982
rect 340794 624948 340828 624982
rect 339982 624854 340016 624888
rect 339982 624764 340016 624798
rect 339982 624674 340016 624708
rect 339982 624584 340016 624618
rect 339982 624494 340016 624528
rect 339982 624404 340016 624438
rect 339982 624314 340016 624348
rect 339982 624224 340016 624258
rect 340872 624835 340906 624869
rect 340872 624745 340906 624779
rect 340872 624655 340906 624689
rect 340872 624565 340906 624599
rect 340872 624475 340906 624509
rect 340872 624385 340906 624419
rect 340872 624295 340906 624329
rect 340872 624205 340906 624239
rect 339982 624134 340016 624168
rect 340872 624115 340906 624149
rect 340040 624058 340074 624092
rect 340130 624058 340164 624092
rect 340220 624058 340254 624092
rect 340310 624058 340344 624092
rect 340400 624058 340434 624092
rect 340490 624058 340524 624092
rect 340580 624058 340614 624092
rect 340670 624058 340704 624092
rect 340760 624058 340794 624092
rect 334922 623660 334956 623694
rect 335012 623660 335046 623694
rect 335102 623660 335136 623694
rect 335192 623660 335226 623694
rect 335282 623660 335316 623694
rect 335372 623660 335406 623694
rect 335462 623660 335496 623694
rect 335552 623660 335586 623694
rect 335642 623660 335676 623694
rect 334830 623566 334864 623600
rect 334830 623476 334864 623510
rect 334830 623386 334864 623420
rect 334830 623296 334864 623330
rect 334830 623206 334864 623240
rect 334830 623116 334864 623150
rect 334830 623026 334864 623060
rect 334830 622936 334864 622970
rect 335720 623547 335754 623581
rect 335720 623457 335754 623491
rect 335720 623367 335754 623401
rect 335720 623277 335754 623311
rect 335720 623187 335754 623221
rect 335720 623097 335754 623131
rect 335720 623007 335754 623041
rect 335720 622917 335754 622951
rect 334830 622846 334864 622880
rect 335720 622827 335754 622861
rect 334888 622770 334922 622804
rect 334978 622770 335012 622804
rect 335068 622770 335102 622804
rect 335158 622770 335192 622804
rect 335248 622770 335282 622804
rect 335338 622770 335372 622804
rect 335428 622770 335462 622804
rect 335518 622770 335552 622804
rect 335608 622770 335642 622804
rect 336210 623660 336244 623694
rect 336300 623660 336334 623694
rect 336390 623660 336424 623694
rect 336480 623660 336514 623694
rect 336570 623660 336604 623694
rect 336660 623660 336694 623694
rect 336750 623660 336784 623694
rect 336840 623660 336874 623694
rect 336930 623660 336964 623694
rect 336118 623566 336152 623600
rect 336118 623476 336152 623510
rect 336118 623386 336152 623420
rect 336118 623296 336152 623330
rect 336118 623206 336152 623240
rect 336118 623116 336152 623150
rect 336118 623026 336152 623060
rect 336118 622936 336152 622970
rect 337008 623547 337042 623581
rect 337008 623457 337042 623491
rect 337008 623367 337042 623401
rect 337008 623277 337042 623311
rect 337008 623187 337042 623221
rect 337008 623097 337042 623131
rect 337008 623007 337042 623041
rect 337008 622917 337042 622951
rect 336118 622846 336152 622880
rect 337008 622827 337042 622861
rect 336176 622770 336210 622804
rect 336266 622770 336300 622804
rect 336356 622770 336390 622804
rect 336446 622770 336480 622804
rect 336536 622770 336570 622804
rect 336626 622770 336660 622804
rect 336716 622770 336750 622804
rect 336806 622770 336840 622804
rect 336896 622770 336930 622804
rect 337498 623660 337532 623694
rect 337588 623660 337622 623694
rect 337678 623660 337712 623694
rect 337768 623660 337802 623694
rect 337858 623660 337892 623694
rect 337948 623660 337982 623694
rect 338038 623660 338072 623694
rect 338128 623660 338162 623694
rect 338218 623660 338252 623694
rect 337406 623566 337440 623600
rect 337406 623476 337440 623510
rect 337406 623386 337440 623420
rect 337406 623296 337440 623330
rect 337406 623206 337440 623240
rect 337406 623116 337440 623150
rect 337406 623026 337440 623060
rect 337406 622936 337440 622970
rect 338296 623547 338330 623581
rect 338296 623457 338330 623491
rect 338296 623367 338330 623401
rect 338296 623277 338330 623311
rect 338296 623187 338330 623221
rect 338296 623097 338330 623131
rect 338296 623007 338330 623041
rect 338296 622917 338330 622951
rect 337406 622846 337440 622880
rect 338296 622827 338330 622861
rect 337464 622770 337498 622804
rect 337554 622770 337588 622804
rect 337644 622770 337678 622804
rect 337734 622770 337768 622804
rect 337824 622770 337858 622804
rect 337914 622770 337948 622804
rect 338004 622770 338038 622804
rect 338094 622770 338128 622804
rect 338184 622770 338218 622804
rect 338786 623660 338820 623694
rect 338876 623660 338910 623694
rect 338966 623660 339000 623694
rect 339056 623660 339090 623694
rect 339146 623660 339180 623694
rect 339236 623660 339270 623694
rect 339326 623660 339360 623694
rect 339416 623660 339450 623694
rect 339506 623660 339540 623694
rect 338694 623566 338728 623600
rect 338694 623476 338728 623510
rect 338694 623386 338728 623420
rect 338694 623296 338728 623330
rect 338694 623206 338728 623240
rect 338694 623116 338728 623150
rect 338694 623026 338728 623060
rect 338694 622936 338728 622970
rect 339584 623547 339618 623581
rect 339584 623457 339618 623491
rect 339584 623367 339618 623401
rect 339584 623277 339618 623311
rect 339584 623187 339618 623221
rect 339584 623097 339618 623131
rect 339584 623007 339618 623041
rect 339584 622917 339618 622951
rect 338694 622846 338728 622880
rect 339584 622827 339618 622861
rect 338752 622770 338786 622804
rect 338842 622770 338876 622804
rect 338932 622770 338966 622804
rect 339022 622770 339056 622804
rect 339112 622770 339146 622804
rect 339202 622770 339236 622804
rect 339292 622770 339326 622804
rect 339382 622770 339416 622804
rect 339472 622770 339506 622804
rect 340074 623660 340108 623694
rect 340164 623660 340198 623694
rect 340254 623660 340288 623694
rect 340344 623660 340378 623694
rect 340434 623660 340468 623694
rect 340524 623660 340558 623694
rect 340614 623660 340648 623694
rect 340704 623660 340738 623694
rect 340794 623660 340828 623694
rect 339982 623566 340016 623600
rect 339982 623476 340016 623510
rect 339982 623386 340016 623420
rect 339982 623296 340016 623330
rect 339982 623206 340016 623240
rect 339982 623116 340016 623150
rect 339982 623026 340016 623060
rect 339982 622936 340016 622970
rect 340872 623547 340906 623581
rect 340872 623457 340906 623491
rect 340872 623367 340906 623401
rect 340872 623277 340906 623311
rect 340872 623187 340906 623221
rect 340872 623097 340906 623131
rect 340872 623007 340906 623041
rect 340872 622917 340906 622951
rect 339982 622846 340016 622880
rect 340872 622827 340906 622861
rect 340040 622770 340074 622804
rect 340130 622770 340164 622804
rect 340220 622770 340254 622804
rect 340310 622770 340344 622804
rect 340400 622770 340434 622804
rect 340490 622770 340524 622804
rect 340580 622770 340614 622804
rect 340670 622770 340704 622804
rect 340760 622770 340794 622804
rect 334922 622372 334956 622406
rect 335012 622372 335046 622406
rect 335102 622372 335136 622406
rect 335192 622372 335226 622406
rect 335282 622372 335316 622406
rect 335372 622372 335406 622406
rect 335462 622372 335496 622406
rect 335552 622372 335586 622406
rect 335642 622372 335676 622406
rect 334830 622278 334864 622312
rect 334830 622188 334864 622222
rect 334830 622098 334864 622132
rect 334830 622008 334864 622042
rect 334830 621918 334864 621952
rect 334830 621828 334864 621862
rect 334830 621738 334864 621772
rect 334830 621648 334864 621682
rect 335720 622259 335754 622293
rect 335720 622169 335754 622203
rect 335720 622079 335754 622113
rect 335720 621989 335754 622023
rect 335720 621899 335754 621933
rect 335720 621809 335754 621843
rect 335720 621719 335754 621753
rect 335720 621629 335754 621663
rect 334830 621558 334864 621592
rect 335720 621539 335754 621573
rect 334888 621482 334922 621516
rect 334978 621482 335012 621516
rect 335068 621482 335102 621516
rect 335158 621482 335192 621516
rect 335248 621482 335282 621516
rect 335338 621482 335372 621516
rect 335428 621482 335462 621516
rect 335518 621482 335552 621516
rect 335608 621482 335642 621516
rect 336210 622372 336244 622406
rect 336300 622372 336334 622406
rect 336390 622372 336424 622406
rect 336480 622372 336514 622406
rect 336570 622372 336604 622406
rect 336660 622372 336694 622406
rect 336750 622372 336784 622406
rect 336840 622372 336874 622406
rect 336930 622372 336964 622406
rect 336118 622278 336152 622312
rect 336118 622188 336152 622222
rect 336118 622098 336152 622132
rect 336118 622008 336152 622042
rect 336118 621918 336152 621952
rect 336118 621828 336152 621862
rect 336118 621738 336152 621772
rect 336118 621648 336152 621682
rect 337008 622259 337042 622293
rect 337008 622169 337042 622203
rect 337008 622079 337042 622113
rect 337008 621989 337042 622023
rect 337008 621899 337042 621933
rect 337008 621809 337042 621843
rect 337008 621719 337042 621753
rect 337008 621629 337042 621663
rect 336118 621558 336152 621592
rect 337008 621539 337042 621573
rect 336176 621482 336210 621516
rect 336266 621482 336300 621516
rect 336356 621482 336390 621516
rect 336446 621482 336480 621516
rect 336536 621482 336570 621516
rect 336626 621482 336660 621516
rect 336716 621482 336750 621516
rect 336806 621482 336840 621516
rect 336896 621482 336930 621516
rect 337498 622372 337532 622406
rect 337588 622372 337622 622406
rect 337678 622372 337712 622406
rect 337768 622372 337802 622406
rect 337858 622372 337892 622406
rect 337948 622372 337982 622406
rect 338038 622372 338072 622406
rect 338128 622372 338162 622406
rect 338218 622372 338252 622406
rect 337406 622278 337440 622312
rect 337406 622188 337440 622222
rect 337406 622098 337440 622132
rect 337406 622008 337440 622042
rect 337406 621918 337440 621952
rect 337406 621828 337440 621862
rect 337406 621738 337440 621772
rect 337406 621648 337440 621682
rect 338296 622259 338330 622293
rect 338296 622169 338330 622203
rect 338296 622079 338330 622113
rect 338296 621989 338330 622023
rect 338296 621899 338330 621933
rect 338296 621809 338330 621843
rect 338296 621719 338330 621753
rect 338296 621629 338330 621663
rect 337406 621558 337440 621592
rect 338296 621539 338330 621573
rect 337464 621482 337498 621516
rect 337554 621482 337588 621516
rect 337644 621482 337678 621516
rect 337734 621482 337768 621516
rect 337824 621482 337858 621516
rect 337914 621482 337948 621516
rect 338004 621482 338038 621516
rect 338094 621482 338128 621516
rect 338184 621482 338218 621516
rect 338786 622372 338820 622406
rect 338876 622372 338910 622406
rect 338966 622372 339000 622406
rect 339056 622372 339090 622406
rect 339146 622372 339180 622406
rect 339236 622372 339270 622406
rect 339326 622372 339360 622406
rect 339416 622372 339450 622406
rect 339506 622372 339540 622406
rect 338694 622278 338728 622312
rect 338694 622188 338728 622222
rect 338694 622098 338728 622132
rect 338694 622008 338728 622042
rect 338694 621918 338728 621952
rect 338694 621828 338728 621862
rect 338694 621738 338728 621772
rect 338694 621648 338728 621682
rect 339584 622259 339618 622293
rect 339584 622169 339618 622203
rect 339584 622079 339618 622113
rect 339584 621989 339618 622023
rect 339584 621899 339618 621933
rect 339584 621809 339618 621843
rect 339584 621719 339618 621753
rect 339584 621629 339618 621663
rect 338694 621558 338728 621592
rect 339584 621539 339618 621573
rect 338752 621482 338786 621516
rect 338842 621482 338876 621516
rect 338932 621482 338966 621516
rect 339022 621482 339056 621516
rect 339112 621482 339146 621516
rect 339202 621482 339236 621516
rect 339292 621482 339326 621516
rect 339382 621482 339416 621516
rect 339472 621482 339506 621516
rect 340074 622372 340108 622406
rect 340164 622372 340198 622406
rect 340254 622372 340288 622406
rect 340344 622372 340378 622406
rect 340434 622372 340468 622406
rect 340524 622372 340558 622406
rect 340614 622372 340648 622406
rect 340704 622372 340738 622406
rect 340794 622372 340828 622406
rect 339982 622278 340016 622312
rect 339982 622188 340016 622222
rect 339982 622098 340016 622132
rect 339982 622008 340016 622042
rect 339982 621918 340016 621952
rect 339982 621828 340016 621862
rect 339982 621738 340016 621772
rect 339982 621648 340016 621682
rect 340872 622259 340906 622293
rect 340872 622169 340906 622203
rect 340872 622079 340906 622113
rect 340872 621989 340906 622023
rect 340872 621899 340906 621933
rect 340872 621809 340906 621843
rect 340872 621719 340906 621753
rect 340872 621629 340906 621663
rect 339982 621558 340016 621592
rect 340872 621539 340906 621573
rect 340040 621482 340074 621516
rect 340130 621482 340164 621516
rect 340220 621482 340254 621516
rect 340310 621482 340344 621516
rect 340400 621482 340434 621516
rect 340490 621482 340524 621516
rect 340580 621482 340614 621516
rect 340670 621482 340704 621516
rect 340760 621482 340794 621516
rect 334922 621084 334956 621118
rect 335012 621084 335046 621118
rect 335102 621084 335136 621118
rect 335192 621084 335226 621118
rect 335282 621084 335316 621118
rect 335372 621084 335406 621118
rect 335462 621084 335496 621118
rect 335552 621084 335586 621118
rect 335642 621084 335676 621118
rect 334830 620990 334864 621024
rect 334830 620900 334864 620934
rect 334830 620810 334864 620844
rect 334830 620720 334864 620754
rect 334830 620630 334864 620664
rect 334830 620540 334864 620574
rect 334830 620450 334864 620484
rect 334830 620360 334864 620394
rect 335720 620971 335754 621005
rect 335720 620881 335754 620915
rect 335720 620791 335754 620825
rect 335720 620701 335754 620735
rect 335720 620611 335754 620645
rect 335720 620521 335754 620555
rect 335720 620431 335754 620465
rect 335720 620341 335754 620375
rect 334830 620270 334864 620304
rect 335720 620251 335754 620285
rect 334888 620194 334922 620228
rect 334978 620194 335012 620228
rect 335068 620194 335102 620228
rect 335158 620194 335192 620228
rect 335248 620194 335282 620228
rect 335338 620194 335372 620228
rect 335428 620194 335462 620228
rect 335518 620194 335552 620228
rect 335608 620194 335642 620228
rect 336210 621084 336244 621118
rect 336300 621084 336334 621118
rect 336390 621084 336424 621118
rect 336480 621084 336514 621118
rect 336570 621084 336604 621118
rect 336660 621084 336694 621118
rect 336750 621084 336784 621118
rect 336840 621084 336874 621118
rect 336930 621084 336964 621118
rect 336118 620990 336152 621024
rect 336118 620900 336152 620934
rect 336118 620810 336152 620844
rect 336118 620720 336152 620754
rect 336118 620630 336152 620664
rect 336118 620540 336152 620574
rect 336118 620450 336152 620484
rect 336118 620360 336152 620394
rect 337008 620971 337042 621005
rect 337008 620881 337042 620915
rect 337008 620791 337042 620825
rect 337008 620701 337042 620735
rect 337008 620611 337042 620645
rect 337008 620521 337042 620555
rect 337008 620431 337042 620465
rect 337008 620341 337042 620375
rect 336118 620270 336152 620304
rect 337008 620251 337042 620285
rect 336176 620194 336210 620228
rect 336266 620194 336300 620228
rect 336356 620194 336390 620228
rect 336446 620194 336480 620228
rect 336536 620194 336570 620228
rect 336626 620194 336660 620228
rect 336716 620194 336750 620228
rect 336806 620194 336840 620228
rect 336896 620194 336930 620228
rect 337498 621084 337532 621118
rect 337588 621084 337622 621118
rect 337678 621084 337712 621118
rect 337768 621084 337802 621118
rect 337858 621084 337892 621118
rect 337948 621084 337982 621118
rect 338038 621084 338072 621118
rect 338128 621084 338162 621118
rect 338218 621084 338252 621118
rect 337406 620990 337440 621024
rect 337406 620900 337440 620934
rect 337406 620810 337440 620844
rect 337406 620720 337440 620754
rect 337406 620630 337440 620664
rect 337406 620540 337440 620574
rect 337406 620450 337440 620484
rect 337406 620360 337440 620394
rect 338296 620971 338330 621005
rect 338296 620881 338330 620915
rect 338296 620791 338330 620825
rect 338296 620701 338330 620735
rect 338296 620611 338330 620645
rect 338296 620521 338330 620555
rect 338296 620431 338330 620465
rect 338296 620341 338330 620375
rect 337406 620270 337440 620304
rect 338296 620251 338330 620285
rect 337464 620194 337498 620228
rect 337554 620194 337588 620228
rect 337644 620194 337678 620228
rect 337734 620194 337768 620228
rect 337824 620194 337858 620228
rect 337914 620194 337948 620228
rect 338004 620194 338038 620228
rect 338094 620194 338128 620228
rect 338184 620194 338218 620228
rect 338786 621084 338820 621118
rect 338876 621084 338910 621118
rect 338966 621084 339000 621118
rect 339056 621084 339090 621118
rect 339146 621084 339180 621118
rect 339236 621084 339270 621118
rect 339326 621084 339360 621118
rect 339416 621084 339450 621118
rect 339506 621084 339540 621118
rect 338694 620990 338728 621024
rect 338694 620900 338728 620934
rect 338694 620810 338728 620844
rect 338694 620720 338728 620754
rect 338694 620630 338728 620664
rect 338694 620540 338728 620574
rect 338694 620450 338728 620484
rect 338694 620360 338728 620394
rect 339584 620971 339618 621005
rect 339584 620881 339618 620915
rect 339584 620791 339618 620825
rect 339584 620701 339618 620735
rect 339584 620611 339618 620645
rect 339584 620521 339618 620555
rect 339584 620431 339618 620465
rect 339584 620341 339618 620375
rect 338694 620270 338728 620304
rect 339584 620251 339618 620285
rect 338752 620194 338786 620228
rect 338842 620194 338876 620228
rect 338932 620194 338966 620228
rect 339022 620194 339056 620228
rect 339112 620194 339146 620228
rect 339202 620194 339236 620228
rect 339292 620194 339326 620228
rect 339382 620194 339416 620228
rect 339472 620194 339506 620228
rect 340074 621084 340108 621118
rect 340164 621084 340198 621118
rect 340254 621084 340288 621118
rect 340344 621084 340378 621118
rect 340434 621084 340468 621118
rect 340524 621084 340558 621118
rect 340614 621084 340648 621118
rect 340704 621084 340738 621118
rect 340794 621084 340828 621118
rect 339982 620990 340016 621024
rect 339982 620900 340016 620934
rect 339982 620810 340016 620844
rect 339982 620720 340016 620754
rect 339982 620630 340016 620664
rect 339982 620540 340016 620574
rect 339982 620450 340016 620484
rect 339982 620360 340016 620394
rect 340872 620971 340906 621005
rect 340872 620881 340906 620915
rect 340872 620791 340906 620825
rect 340872 620701 340906 620735
rect 340872 620611 340906 620645
rect 340872 620521 340906 620555
rect 340872 620431 340906 620465
rect 340872 620341 340906 620375
rect 339982 620270 340016 620304
rect 340872 620251 340906 620285
rect 340040 620194 340074 620228
rect 340130 620194 340164 620228
rect 340220 620194 340254 620228
rect 340310 620194 340344 620228
rect 340400 620194 340434 620228
rect 340490 620194 340524 620228
rect 340580 620194 340614 620228
rect 340670 620194 340704 620228
rect 340760 620194 340794 620228
rect 334922 619796 334956 619830
rect 335012 619796 335046 619830
rect 335102 619796 335136 619830
rect 335192 619796 335226 619830
rect 335282 619796 335316 619830
rect 335372 619796 335406 619830
rect 335462 619796 335496 619830
rect 335552 619796 335586 619830
rect 335642 619796 335676 619830
rect 334830 619702 334864 619736
rect 334830 619612 334864 619646
rect 334830 619522 334864 619556
rect 334830 619432 334864 619466
rect 334830 619342 334864 619376
rect 334830 619252 334864 619286
rect 334830 619162 334864 619196
rect 334830 619072 334864 619106
rect 335720 619683 335754 619717
rect 335720 619593 335754 619627
rect 335720 619503 335754 619537
rect 335720 619413 335754 619447
rect 335720 619323 335754 619357
rect 335720 619233 335754 619267
rect 335720 619143 335754 619177
rect 335720 619053 335754 619087
rect 334830 618982 334864 619016
rect 335720 618963 335754 618997
rect 334888 618906 334922 618940
rect 334978 618906 335012 618940
rect 335068 618906 335102 618940
rect 335158 618906 335192 618940
rect 335248 618906 335282 618940
rect 335338 618906 335372 618940
rect 335428 618906 335462 618940
rect 335518 618906 335552 618940
rect 335608 618906 335642 618940
rect 336210 619796 336244 619830
rect 336300 619796 336334 619830
rect 336390 619796 336424 619830
rect 336480 619796 336514 619830
rect 336570 619796 336604 619830
rect 336660 619796 336694 619830
rect 336750 619796 336784 619830
rect 336840 619796 336874 619830
rect 336930 619796 336964 619830
rect 336118 619702 336152 619736
rect 336118 619612 336152 619646
rect 336118 619522 336152 619556
rect 336118 619432 336152 619466
rect 336118 619342 336152 619376
rect 336118 619252 336152 619286
rect 336118 619162 336152 619196
rect 336118 619072 336152 619106
rect 337008 619683 337042 619717
rect 337008 619593 337042 619627
rect 337008 619503 337042 619537
rect 337008 619413 337042 619447
rect 337008 619323 337042 619357
rect 337008 619233 337042 619267
rect 337008 619143 337042 619177
rect 337008 619053 337042 619087
rect 336118 618982 336152 619016
rect 337008 618963 337042 618997
rect 336176 618906 336210 618940
rect 336266 618906 336300 618940
rect 336356 618906 336390 618940
rect 336446 618906 336480 618940
rect 336536 618906 336570 618940
rect 336626 618906 336660 618940
rect 336716 618906 336750 618940
rect 336806 618906 336840 618940
rect 336896 618906 336930 618940
rect 337498 619796 337532 619830
rect 337588 619796 337622 619830
rect 337678 619796 337712 619830
rect 337768 619796 337802 619830
rect 337858 619796 337892 619830
rect 337948 619796 337982 619830
rect 338038 619796 338072 619830
rect 338128 619796 338162 619830
rect 338218 619796 338252 619830
rect 337406 619702 337440 619736
rect 337406 619612 337440 619646
rect 337406 619522 337440 619556
rect 337406 619432 337440 619466
rect 337406 619342 337440 619376
rect 337406 619252 337440 619286
rect 337406 619162 337440 619196
rect 337406 619072 337440 619106
rect 338296 619683 338330 619717
rect 338296 619593 338330 619627
rect 338296 619503 338330 619537
rect 338296 619413 338330 619447
rect 338296 619323 338330 619357
rect 338296 619233 338330 619267
rect 338296 619143 338330 619177
rect 338296 619053 338330 619087
rect 337406 618982 337440 619016
rect 338296 618963 338330 618997
rect 337464 618906 337498 618940
rect 337554 618906 337588 618940
rect 337644 618906 337678 618940
rect 337734 618906 337768 618940
rect 337824 618906 337858 618940
rect 337914 618906 337948 618940
rect 338004 618906 338038 618940
rect 338094 618906 338128 618940
rect 338184 618906 338218 618940
rect 338786 619796 338820 619830
rect 338876 619796 338910 619830
rect 338966 619796 339000 619830
rect 339056 619796 339090 619830
rect 339146 619796 339180 619830
rect 339236 619796 339270 619830
rect 339326 619796 339360 619830
rect 339416 619796 339450 619830
rect 339506 619796 339540 619830
rect 338694 619702 338728 619736
rect 338694 619612 338728 619646
rect 338694 619522 338728 619556
rect 338694 619432 338728 619466
rect 338694 619342 338728 619376
rect 338694 619252 338728 619286
rect 338694 619162 338728 619196
rect 338694 619072 338728 619106
rect 339584 619683 339618 619717
rect 339584 619593 339618 619627
rect 339584 619503 339618 619537
rect 339584 619413 339618 619447
rect 339584 619323 339618 619357
rect 339584 619233 339618 619267
rect 339584 619143 339618 619177
rect 339584 619053 339618 619087
rect 338694 618982 338728 619016
rect 339584 618963 339618 618997
rect 338752 618906 338786 618940
rect 338842 618906 338876 618940
rect 338932 618906 338966 618940
rect 339022 618906 339056 618940
rect 339112 618906 339146 618940
rect 339202 618906 339236 618940
rect 339292 618906 339326 618940
rect 339382 618906 339416 618940
rect 339472 618906 339506 618940
rect 340074 619796 340108 619830
rect 340164 619796 340198 619830
rect 340254 619796 340288 619830
rect 340344 619796 340378 619830
rect 340434 619796 340468 619830
rect 340524 619796 340558 619830
rect 340614 619796 340648 619830
rect 340704 619796 340738 619830
rect 340794 619796 340828 619830
rect 339982 619702 340016 619736
rect 339982 619612 340016 619646
rect 339982 619522 340016 619556
rect 339982 619432 340016 619466
rect 339982 619342 340016 619376
rect 339982 619252 340016 619286
rect 339982 619162 340016 619196
rect 339982 619072 340016 619106
rect 340872 619683 340906 619717
rect 340872 619593 340906 619627
rect 340872 619503 340906 619537
rect 340872 619413 340906 619447
rect 340872 619323 340906 619357
rect 340872 619233 340906 619267
rect 340872 619143 340906 619177
rect 340872 619053 340906 619087
rect 339982 618982 340016 619016
rect 340872 618963 340906 618997
rect 340040 618906 340074 618940
rect 340130 618906 340164 618940
rect 340220 618906 340254 618940
rect 340310 618906 340344 618940
rect 340400 618906 340434 618940
rect 340490 618906 340524 618940
rect 340580 618906 340614 618940
rect 340670 618906 340704 618940
rect 340760 618906 340794 618940
rect 334922 618508 334956 618542
rect 335012 618508 335046 618542
rect 335102 618508 335136 618542
rect 335192 618508 335226 618542
rect 335282 618508 335316 618542
rect 335372 618508 335406 618542
rect 335462 618508 335496 618542
rect 335552 618508 335586 618542
rect 335642 618508 335676 618542
rect 334830 618414 334864 618448
rect 334830 618324 334864 618358
rect 334830 618234 334864 618268
rect 334830 618144 334864 618178
rect 334830 618054 334864 618088
rect 334830 617964 334864 617998
rect 334830 617874 334864 617908
rect 334830 617784 334864 617818
rect 335720 618395 335754 618429
rect 335720 618305 335754 618339
rect 335720 618215 335754 618249
rect 335720 618125 335754 618159
rect 335720 618035 335754 618069
rect 335720 617945 335754 617979
rect 335720 617855 335754 617889
rect 335720 617765 335754 617799
rect 334830 617694 334864 617728
rect 335720 617675 335754 617709
rect 334888 617618 334922 617652
rect 334978 617618 335012 617652
rect 335068 617618 335102 617652
rect 335158 617618 335192 617652
rect 335248 617618 335282 617652
rect 335338 617618 335372 617652
rect 335428 617618 335462 617652
rect 335518 617618 335552 617652
rect 335608 617618 335642 617652
rect 336210 618508 336244 618542
rect 336300 618508 336334 618542
rect 336390 618508 336424 618542
rect 336480 618508 336514 618542
rect 336570 618508 336604 618542
rect 336660 618508 336694 618542
rect 336750 618508 336784 618542
rect 336840 618508 336874 618542
rect 336930 618508 336964 618542
rect 336118 618414 336152 618448
rect 336118 618324 336152 618358
rect 336118 618234 336152 618268
rect 336118 618144 336152 618178
rect 336118 618054 336152 618088
rect 336118 617964 336152 617998
rect 336118 617874 336152 617908
rect 336118 617784 336152 617818
rect 337008 618395 337042 618429
rect 337008 618305 337042 618339
rect 337008 618215 337042 618249
rect 337008 618125 337042 618159
rect 337008 618035 337042 618069
rect 337008 617945 337042 617979
rect 337008 617855 337042 617889
rect 337008 617765 337042 617799
rect 336118 617694 336152 617728
rect 337008 617675 337042 617709
rect 336176 617618 336210 617652
rect 336266 617618 336300 617652
rect 336356 617618 336390 617652
rect 336446 617618 336480 617652
rect 336536 617618 336570 617652
rect 336626 617618 336660 617652
rect 336716 617618 336750 617652
rect 336806 617618 336840 617652
rect 336896 617618 336930 617652
rect 337498 618508 337532 618542
rect 337588 618508 337622 618542
rect 337678 618508 337712 618542
rect 337768 618508 337802 618542
rect 337858 618508 337892 618542
rect 337948 618508 337982 618542
rect 338038 618508 338072 618542
rect 338128 618508 338162 618542
rect 338218 618508 338252 618542
rect 337406 618414 337440 618448
rect 337406 618324 337440 618358
rect 337406 618234 337440 618268
rect 337406 618144 337440 618178
rect 337406 618054 337440 618088
rect 337406 617964 337440 617998
rect 337406 617874 337440 617908
rect 337406 617784 337440 617818
rect 338296 618395 338330 618429
rect 338296 618305 338330 618339
rect 338296 618215 338330 618249
rect 338296 618125 338330 618159
rect 338296 618035 338330 618069
rect 338296 617945 338330 617979
rect 338296 617855 338330 617889
rect 338296 617765 338330 617799
rect 337406 617694 337440 617728
rect 338296 617675 338330 617709
rect 337464 617618 337498 617652
rect 337554 617618 337588 617652
rect 337644 617618 337678 617652
rect 337734 617618 337768 617652
rect 337824 617618 337858 617652
rect 337914 617618 337948 617652
rect 338004 617618 338038 617652
rect 338094 617618 338128 617652
rect 338184 617618 338218 617652
rect 338786 618508 338820 618542
rect 338876 618508 338910 618542
rect 338966 618508 339000 618542
rect 339056 618508 339090 618542
rect 339146 618508 339180 618542
rect 339236 618508 339270 618542
rect 339326 618508 339360 618542
rect 339416 618508 339450 618542
rect 339506 618508 339540 618542
rect 338694 618414 338728 618448
rect 338694 618324 338728 618358
rect 338694 618234 338728 618268
rect 338694 618144 338728 618178
rect 338694 618054 338728 618088
rect 338694 617964 338728 617998
rect 338694 617874 338728 617908
rect 338694 617784 338728 617818
rect 339584 618395 339618 618429
rect 339584 618305 339618 618339
rect 339584 618215 339618 618249
rect 339584 618125 339618 618159
rect 339584 618035 339618 618069
rect 339584 617945 339618 617979
rect 339584 617855 339618 617889
rect 339584 617765 339618 617799
rect 338694 617694 338728 617728
rect 339584 617675 339618 617709
rect 338752 617618 338786 617652
rect 338842 617618 338876 617652
rect 338932 617618 338966 617652
rect 339022 617618 339056 617652
rect 339112 617618 339146 617652
rect 339202 617618 339236 617652
rect 339292 617618 339326 617652
rect 339382 617618 339416 617652
rect 339472 617618 339506 617652
rect 340074 618508 340108 618542
rect 340164 618508 340198 618542
rect 340254 618508 340288 618542
rect 340344 618508 340378 618542
rect 340434 618508 340468 618542
rect 340524 618508 340558 618542
rect 340614 618508 340648 618542
rect 340704 618508 340738 618542
rect 340794 618508 340828 618542
rect 339982 618414 340016 618448
rect 339982 618324 340016 618358
rect 339982 618234 340016 618268
rect 339982 618144 340016 618178
rect 339982 618054 340016 618088
rect 339982 617964 340016 617998
rect 339982 617874 340016 617908
rect 339982 617784 340016 617818
rect 340872 618395 340906 618429
rect 340872 618305 340906 618339
rect 340872 618215 340906 618249
rect 340872 618125 340906 618159
rect 340872 618035 340906 618069
rect 340872 617945 340906 617979
rect 340872 617855 340906 617889
rect 340872 617765 340906 617799
rect 339982 617694 340016 617728
rect 340872 617675 340906 617709
rect 340040 617618 340074 617652
rect 340130 617618 340164 617652
rect 340220 617618 340254 617652
rect 340310 617618 340344 617652
rect 340400 617618 340434 617652
rect 340490 617618 340524 617652
rect 340580 617618 340614 617652
rect 340670 617618 340704 617652
rect 340760 617618 340794 617652
rect 306536 616702 308878 616802
<< poly >>
rect 313450 624946 313850 624972
rect 313908 624946 314308 624972
rect 314366 624946 314766 624972
rect 314824 624946 315224 624972
rect 315282 624946 315682 624972
rect 315740 624946 316140 624972
rect 316198 624946 316598 624972
rect 316656 624946 317056 624972
rect 317114 624946 317514 624972
rect 317572 624946 317972 624972
rect 318030 624946 318430 624972
rect 319408 624946 319808 624972
rect 319866 624946 320266 624972
rect 320324 624946 320724 624972
rect 320782 624946 321182 624972
rect 321240 624946 321640 624972
rect 321698 624946 322098 624972
rect 322156 624946 322556 624972
rect 322614 624946 323014 624972
rect 323072 624946 323472 624972
rect 323530 624946 323930 624972
rect 324908 624946 325308 624972
rect 325366 624946 325766 624972
rect 325824 624946 326224 624972
rect 326282 624946 326682 624972
rect 326740 624946 327140 624972
rect 327198 624946 327598 624972
rect 327656 624946 328056 624972
rect 328114 624946 328514 624972
rect 328572 624946 328972 624972
rect 329030 624946 329430 624972
rect 329488 624946 329888 624972
rect 304940 624296 305028 624312
rect 304940 623928 304956 624296
rect 304990 623928 305028 624296
rect 304940 623912 305028 623928
rect 310428 623912 310454 624312
rect 305368 622232 305768 622248
rect 305368 622198 305384 622232
rect 305752 622198 305768 622232
rect 305368 622160 305768 622198
rect 305940 622232 306340 622248
rect 305940 622198 305956 622232
rect 306324 622198 306340 622232
rect 305940 622160 306340 622198
rect 306512 622232 306912 622248
rect 306512 622198 306528 622232
rect 306896 622198 306912 622232
rect 306512 622160 306912 622198
rect 307084 622232 307484 622248
rect 307084 622198 307100 622232
rect 307468 622198 307484 622232
rect 307084 622160 307484 622198
rect 307656 622232 308056 622248
rect 307656 622198 307672 622232
rect 308040 622198 308056 622232
rect 307656 622160 308056 622198
rect 308228 622232 308628 622248
rect 308228 622198 308244 622232
rect 308612 622198 308628 622232
rect 308228 622160 308628 622198
rect 308800 622232 309200 622248
rect 308800 622198 308816 622232
rect 309184 622198 309200 622232
rect 308800 622160 309200 622198
rect 309372 622232 309772 622248
rect 309372 622198 309388 622232
rect 309756 622198 309772 622232
rect 309372 622160 309772 622198
rect 300438 621110 300838 621126
rect 300438 621076 300454 621110
rect 300822 621076 300838 621110
rect 300438 621038 300838 621076
rect 300896 621110 301296 621126
rect 300896 621076 300912 621110
rect 301280 621076 301296 621110
rect 300896 621038 301296 621076
rect 301354 621110 301754 621126
rect 301354 621076 301370 621110
rect 301738 621076 301754 621110
rect 301354 621038 301754 621076
rect 301812 621110 302212 621126
rect 301812 621076 301828 621110
rect 302196 621076 302212 621110
rect 301812 621038 302212 621076
rect 302270 621110 302670 621126
rect 302270 621076 302286 621110
rect 302654 621076 302670 621110
rect 302270 621038 302670 621076
rect 302728 621110 303128 621126
rect 302728 621076 302744 621110
rect 303112 621076 303128 621110
rect 302728 621038 303128 621076
rect 300438 620612 300838 620638
rect 300896 620612 301296 620638
rect 301354 620612 301754 620638
rect 301812 620612 302212 620638
rect 302270 620612 302670 620638
rect 302728 620612 303128 620638
rect 305368 620334 305768 620360
rect 305940 620334 306340 620360
rect 306512 620334 306912 620360
rect 307084 620334 307484 620360
rect 307656 620334 308056 620360
rect 308228 620334 308628 620360
rect 308800 620334 309200 620360
rect 309372 620334 309772 620360
rect 303642 619829 304042 619845
rect 303642 619795 303658 619829
rect 304026 619795 304042 619829
rect 303642 619748 304042 619795
rect 304214 619829 304614 619845
rect 304214 619795 304230 619829
rect 304598 619795 304614 619829
rect 304214 619748 304614 619795
rect 304786 619829 305186 619845
rect 304786 619795 304802 619829
rect 305170 619795 305186 619829
rect 304786 619748 305186 619795
rect 305358 619829 305758 619845
rect 305358 619795 305374 619829
rect 305742 619795 305758 619829
rect 305358 619748 305758 619795
rect 305930 619829 306330 619845
rect 305930 619795 305946 619829
rect 306314 619795 306330 619829
rect 305930 619748 306330 619795
rect 306502 619829 306902 619845
rect 306502 619795 306518 619829
rect 306886 619795 306902 619829
rect 306502 619748 306902 619795
rect 307074 619829 307474 619845
rect 307074 619795 307090 619829
rect 307458 619795 307474 619829
rect 307074 619748 307474 619795
rect 307646 619829 308046 619845
rect 307646 619795 307662 619829
rect 308030 619795 308046 619829
rect 307646 619748 308046 619795
rect 308218 619829 308618 619845
rect 308218 619795 308234 619829
rect 308602 619795 308618 619829
rect 308218 619748 308618 619795
rect 308790 619829 309190 619845
rect 308790 619795 308806 619829
rect 309174 619795 309190 619829
rect 308790 619748 309190 619795
rect 309362 619829 309762 619845
rect 309362 619795 309378 619829
rect 309746 619795 309762 619829
rect 309362 619748 309762 619795
rect 309934 619829 310334 619845
rect 309934 619795 309950 619829
rect 310318 619795 310334 619829
rect 309934 619748 310334 619795
rect 310506 619829 310906 619845
rect 310506 619795 310522 619829
rect 310890 619795 310906 619829
rect 310506 619748 310906 619795
rect 311078 619829 311478 619845
rect 311078 619795 311094 619829
rect 311462 619795 311478 619829
rect 311078 619748 311478 619795
rect 303642 617142 304042 617168
rect 304214 617142 304614 617168
rect 304786 617142 305186 617168
rect 305358 617142 305758 617168
rect 305930 617142 306330 617168
rect 306502 617142 306902 617168
rect 307074 617142 307474 617168
rect 307646 617142 308046 617168
rect 308218 617142 308618 617168
rect 308790 617142 309190 617168
rect 309362 617142 309762 617168
rect 309934 617142 310334 617168
rect 310506 617142 310906 617168
rect 311078 617142 311478 617168
rect 313450 617159 313850 617206
rect 313450 617125 313466 617159
rect 313834 617125 313850 617159
rect 313450 617109 313850 617125
rect 313908 617159 314308 617206
rect 313908 617125 313924 617159
rect 314292 617125 314308 617159
rect 313908 617109 314308 617125
rect 314366 617159 314766 617206
rect 314366 617125 314382 617159
rect 314750 617125 314766 617159
rect 314366 617109 314766 617125
rect 314824 617159 315224 617206
rect 314824 617125 314840 617159
rect 315208 617125 315224 617159
rect 314824 617109 315224 617125
rect 315282 617159 315682 617206
rect 315282 617125 315298 617159
rect 315666 617125 315682 617159
rect 315282 617109 315682 617125
rect 315740 617159 316140 617206
rect 315740 617125 315756 617159
rect 316124 617125 316140 617159
rect 315740 617109 316140 617125
rect 316198 617159 316598 617206
rect 316198 617125 316214 617159
rect 316582 617125 316598 617159
rect 316198 617109 316598 617125
rect 316656 617159 317056 617206
rect 316656 617125 316672 617159
rect 317040 617125 317056 617159
rect 316656 617109 317056 617125
rect 317114 617159 317514 617206
rect 317114 617125 317130 617159
rect 317498 617125 317514 617159
rect 317114 617109 317514 617125
rect 317572 617159 317972 617206
rect 317572 617125 317588 617159
rect 317956 617125 317972 617159
rect 317572 617109 317972 617125
rect 318030 617159 318430 617206
rect 318030 617125 318046 617159
rect 318414 617125 318430 617159
rect 318030 617109 318430 617125
rect 319408 617159 319808 617206
rect 319408 617125 319424 617159
rect 319792 617125 319808 617159
rect 319408 617109 319808 617125
rect 319866 617159 320266 617206
rect 319866 617125 319882 617159
rect 320250 617125 320266 617159
rect 319866 617109 320266 617125
rect 320324 617159 320724 617206
rect 320324 617125 320340 617159
rect 320708 617125 320724 617159
rect 320324 617109 320724 617125
rect 320782 617159 321182 617206
rect 320782 617125 320798 617159
rect 321166 617125 321182 617159
rect 320782 617109 321182 617125
rect 321240 617159 321640 617206
rect 321240 617125 321256 617159
rect 321624 617125 321640 617159
rect 321240 617109 321640 617125
rect 321698 617159 322098 617206
rect 321698 617125 321714 617159
rect 322082 617125 322098 617159
rect 321698 617109 322098 617125
rect 322156 617159 322556 617206
rect 322156 617125 322172 617159
rect 322540 617125 322556 617159
rect 322156 617109 322556 617125
rect 322614 617159 323014 617206
rect 322614 617125 322630 617159
rect 322998 617125 323014 617159
rect 322614 617109 323014 617125
rect 323072 617159 323472 617206
rect 323072 617125 323088 617159
rect 323456 617125 323472 617159
rect 323072 617109 323472 617125
rect 323530 617159 323930 617206
rect 323530 617125 323546 617159
rect 323914 617125 323930 617159
rect 323530 617109 323930 617125
rect 324908 617159 325308 617206
rect 324908 617125 324924 617159
rect 325292 617125 325308 617159
rect 324908 617109 325308 617125
rect 325366 617159 325766 617206
rect 325366 617125 325382 617159
rect 325750 617125 325766 617159
rect 325366 617109 325766 617125
rect 325824 617159 326224 617206
rect 325824 617125 325840 617159
rect 326208 617125 326224 617159
rect 325824 617109 326224 617125
rect 326282 617159 326682 617206
rect 326282 617125 326298 617159
rect 326666 617125 326682 617159
rect 326282 617109 326682 617125
rect 326740 617159 327140 617206
rect 326740 617125 326756 617159
rect 327124 617125 327140 617159
rect 326740 617109 327140 617125
rect 327198 617159 327598 617206
rect 327198 617125 327214 617159
rect 327582 617125 327598 617159
rect 327198 617109 327598 617125
rect 327656 617159 328056 617206
rect 327656 617125 327672 617159
rect 328040 617125 328056 617159
rect 327656 617109 328056 617125
rect 328114 617159 328514 617206
rect 328114 617125 328130 617159
rect 328498 617125 328514 617159
rect 328114 617109 328514 617125
rect 328572 617159 328972 617206
rect 328572 617125 328588 617159
rect 328956 617125 328972 617159
rect 328572 617109 328972 617125
rect 329030 617159 329430 617206
rect 329030 617125 329046 617159
rect 329414 617125 329430 617159
rect 329030 617109 329430 617125
rect 329488 617159 329888 617206
rect 329488 617125 329504 617159
rect 329872 617125 329888 617159
rect 329488 617109 329888 617125
<< polycont >>
rect 304956 623928 304990 624296
rect 305384 622198 305752 622232
rect 305956 622198 306324 622232
rect 306528 622198 306896 622232
rect 307100 622198 307468 622232
rect 307672 622198 308040 622232
rect 308244 622198 308612 622232
rect 308816 622198 309184 622232
rect 309388 622198 309756 622232
rect 300454 621076 300822 621110
rect 300912 621076 301280 621110
rect 301370 621076 301738 621110
rect 301828 621076 302196 621110
rect 302286 621076 302654 621110
rect 302744 621076 303112 621110
rect 303658 619795 304026 619829
rect 304230 619795 304598 619829
rect 304802 619795 305170 619829
rect 305374 619795 305742 619829
rect 305946 619795 306314 619829
rect 306518 619795 306886 619829
rect 307090 619795 307458 619829
rect 307662 619795 308030 619829
rect 308234 619795 308602 619829
rect 308806 619795 309174 619829
rect 309378 619795 309746 619829
rect 309950 619795 310318 619829
rect 310522 619795 310890 619829
rect 311094 619795 311462 619829
rect 313466 617125 313834 617159
rect 313924 617125 314292 617159
rect 314382 617125 314750 617159
rect 314840 617125 315208 617159
rect 315298 617125 315666 617159
rect 315756 617125 316124 617159
rect 316214 617125 316582 617159
rect 316672 617125 317040 617159
rect 317130 617125 317498 617159
rect 317588 617125 317956 617159
rect 318046 617125 318414 617159
rect 319424 617125 319792 617159
rect 319882 617125 320250 617159
rect 320340 617125 320708 617159
rect 320798 617125 321166 617159
rect 321256 617125 321624 617159
rect 321714 617125 322082 617159
rect 322172 617125 322540 617159
rect 322630 617125 322998 617159
rect 323088 617125 323456 617159
rect 323546 617125 323914 617159
rect 324924 617125 325292 617159
rect 325382 617125 325750 617159
rect 325840 617125 326208 617159
rect 326298 617125 326666 617159
rect 326756 617125 327124 617159
rect 327214 617125 327582 617159
rect 327672 617125 328040 617159
rect 328130 617125 328498 617159
rect 328588 617125 328956 617159
rect 329046 617125 329414 617159
rect 329504 617125 329872 617159
<< xpolycontact >>
rect 316544 637068 317114 637500
rect 313272 635682 313842 636114
rect 313272 631926 313842 632358
rect 314090 635682 314660 636114
rect 314090 631926 314660 632358
rect 314908 635682 315478 636114
rect 314908 631926 315478 632358
rect 316544 632336 317114 632768
rect 317362 637068 317932 637500
rect 317362 632336 317932 632768
rect 318180 637068 318750 637500
rect 318180 632336 318750 632768
rect 318998 637068 319568 637500
rect 318998 632336 319568 632768
rect 321452 637006 322022 637438
rect 321452 630270 322022 630702
rect 322270 637006 322840 637438
rect 322270 630270 322840 630702
rect 323088 637006 323658 637438
rect 323088 630270 323658 630702
rect 323906 637006 324476 637438
rect 323906 630270 324476 630702
rect 324724 637006 325294 637438
rect 324724 630270 325294 630702
rect 325542 637006 326112 637438
rect 325542 630270 326112 630702
rect 326360 637006 326930 637438
rect 326360 630270 326930 630702
rect 327178 637006 327748 637438
rect 327178 630270 327748 630702
rect 327996 637006 328566 637438
rect 327996 630270 328566 630702
rect 328814 637006 329384 637438
rect 328814 630270 329384 630702
rect 329632 637006 330202 637438
rect 329632 630270 330202 630702
rect 330450 637006 331020 637438
rect 330450 630270 331020 630702
rect 331268 637006 331838 637438
rect 331268 630270 331838 630702
rect 332086 637006 332656 637438
rect 332086 630270 332656 630702
rect 332904 637006 333474 637438
rect 332904 630270 333474 630702
rect 333722 637006 334292 637438
rect 333722 630270 334292 630702
rect 334540 637006 335110 637438
rect 334540 630270 335110 630702
<< xpolyres >>
rect 313272 632358 313842 635682
rect 314090 632358 314660 635682
rect 314908 632358 315478 635682
rect 316544 632768 317114 637068
rect 317362 632768 317932 637068
rect 318180 632768 318750 637068
rect 318998 632768 319568 637068
rect 321452 630702 322022 637006
rect 322270 630702 322840 637006
rect 323088 630702 323658 637006
rect 323906 630702 324476 637006
rect 324724 630702 325294 637006
rect 325542 630702 326112 637006
rect 326360 630702 326930 637006
rect 327178 630702 327748 637006
rect 327996 630702 328566 637006
rect 328814 630702 329384 637006
rect 329632 630702 330202 637006
rect 330450 630702 331020 637006
rect 331268 630702 331838 637006
rect 332086 630702 332656 637006
rect 332904 630702 333474 637006
rect 333722 630702 334292 637006
rect 334540 630702 335110 637006
<< locali >>
rect 297800 642688 298824 642696
rect 297800 642672 298876 642688
rect 298976 642672 299100 642688
rect 299200 642672 299324 642688
rect 299424 642672 299548 642688
rect 299648 642672 299772 642688
rect 299872 642672 299996 642688
rect 300096 642672 300220 642688
rect 300320 642672 300444 642688
rect 300544 642672 300668 642688
rect 300768 642672 300892 642688
rect 300992 642672 301116 642688
rect 301216 642672 301340 642688
rect 301440 642672 301564 642688
rect 301664 642672 301788 642688
rect 301888 642672 302012 642688
rect 302112 642672 302236 642688
rect 302336 642672 302460 642688
rect 302560 642672 302684 642688
rect 302784 642672 302908 642688
rect 303008 642672 303132 642688
rect 303232 642672 303356 642688
rect 303456 642672 303580 642688
rect 303680 642672 303804 642688
rect 303904 642672 304028 642688
rect 304128 642672 304252 642688
rect 304352 642672 304476 642688
rect 304576 642672 304700 642688
rect 304800 642672 304924 642688
rect 305024 642672 305148 642688
rect 305248 642672 305372 642688
rect 305472 642672 309346 642688
rect 309446 642672 309570 642688
rect 309670 642672 309794 642688
rect 309894 642672 310018 642688
rect 310118 642672 310242 642688
rect 310342 642672 310466 642688
rect 310566 642672 310690 642688
rect 310790 642672 310914 642688
rect 311014 642672 311138 642688
rect 311238 642672 311362 642688
rect 311462 642672 311586 642688
rect 311686 642672 311810 642688
rect 311910 642672 312034 642688
rect 312134 642672 312258 642688
rect 312358 642672 312482 642688
rect 312582 642672 312706 642688
rect 312806 642672 312930 642688
rect 313030 642672 313154 642688
rect 313254 642672 313378 642688
rect 313478 642672 313602 642688
rect 313702 642672 313826 642688
rect 313926 642672 314050 642688
rect 314150 642672 314274 642688
rect 314374 642672 314498 642688
rect 314598 642672 314722 642688
rect 314822 642672 314946 642688
rect 315046 642672 315170 642688
rect 315270 642672 315394 642688
rect 315494 642672 315618 642688
rect 315718 642672 315842 642688
rect 315942 642672 335616 642688
rect 335716 642672 335840 642688
rect 335940 642672 336064 642688
rect 336164 642672 336288 642688
rect 336388 642672 336512 642688
rect 336612 642672 336736 642688
rect 336836 642672 336960 642688
rect 337060 642672 337184 642688
rect 337284 642672 337408 642688
rect 337508 642672 337632 642688
rect 337732 642672 337856 642688
rect 337956 642672 338080 642688
rect 338180 642672 338304 642688
rect 338404 642672 338528 642688
rect 338628 642672 338752 642688
rect 338852 642672 338976 642688
rect 339076 642672 339200 642688
rect 339300 642672 339424 642688
rect 339524 642672 339648 642688
rect 339748 642672 339872 642688
rect 339972 642672 340096 642688
rect 340196 642672 340320 642688
rect 340420 642672 340544 642688
rect 340644 642672 340768 642688
rect 340868 642672 340992 642688
rect 341092 642672 341216 642688
rect 341316 642672 341440 642688
rect 341540 642672 341664 642688
rect 341764 642672 341888 642688
rect 341988 642672 342112 642688
rect 342212 642672 343160 642696
rect 297800 641672 297824 642672
rect 343136 641672 343160 642672
rect 297800 641656 343160 641672
rect 297800 640640 298824 641656
rect 342160 640664 343160 641656
rect 342096 640648 343160 640664
rect 297800 640624 298888 640640
rect 297800 637996 297872 640624
rect 297800 637896 297850 637996
rect 297800 637772 297872 637896
rect 297800 637672 297850 637772
rect 297800 637548 297872 637672
rect 297800 637448 297850 637548
rect 297800 637324 297872 637448
rect 297800 637224 297850 637324
rect 297800 637100 297872 637224
rect 297800 637000 297850 637100
rect 297800 636876 297872 637000
rect 297800 636776 297850 636876
rect 297800 636652 297872 636776
rect 297800 636552 297850 636652
rect 297800 636428 297872 636552
rect 297800 636328 297850 636428
rect 297800 636204 297872 636328
rect 297800 636104 297850 636204
rect 297800 635980 297872 636104
rect 297800 635880 297850 635980
rect 297800 635756 297872 635880
rect 297800 635656 297850 635756
rect 297800 635532 297872 635656
rect 297800 635432 297850 635532
rect 297800 635308 297872 635432
rect 297800 635208 297850 635308
rect 297800 635084 297872 635208
rect 297800 634984 297850 635084
rect 297800 634860 297872 634984
rect 297800 634760 297850 634860
rect 297800 634636 297872 634760
rect 297800 634536 297850 634636
rect 297800 634412 297872 634536
rect 297800 634312 297850 634412
rect 297800 634188 297872 634312
rect 297800 634088 297850 634188
rect 297800 633964 297872 634088
rect 297800 633864 297850 633964
rect 297800 633740 297872 633864
rect 297800 633640 297850 633740
rect 297800 633516 297872 633640
rect 297800 633416 297850 633516
rect 297800 633292 297872 633416
rect 297800 633192 297850 633292
rect 297800 633068 297872 633192
rect 297800 632968 297850 633068
rect 297800 632844 297872 632968
rect 297800 632744 297850 632844
rect 297800 632620 297872 632744
rect 297800 632520 297850 632620
rect 297800 632396 297872 632520
rect 297800 632296 297850 632396
rect 297800 632172 297872 632296
rect 297800 632072 297850 632172
rect 297800 631948 297872 632072
rect 297800 631848 297850 631948
rect 297800 631724 297872 631848
rect 297800 631624 297850 631724
rect 297800 631500 297872 631624
rect 297800 631400 297850 631500
rect 297800 624596 297872 631400
rect 297800 624496 297850 624596
rect 297800 624372 297872 624496
rect 297800 624272 297850 624372
rect 297800 624148 297872 624272
rect 297800 624048 297850 624148
rect 297800 623924 297872 624048
rect 297800 623824 297850 623924
rect 297800 623700 297872 623824
rect 297800 623600 297850 623700
rect 297800 623476 297872 623600
rect 297800 623376 297850 623476
rect 297800 623252 297872 623376
rect 297800 623152 297850 623252
rect 297800 623028 297872 623152
rect 297800 622928 297850 623028
rect 297800 622804 297872 622928
rect 297800 622704 297850 622804
rect 297800 622580 297872 622704
rect 297800 622480 297850 622580
rect 297800 622356 297872 622480
rect 297800 622256 297850 622356
rect 297800 622132 297872 622256
rect 297800 622032 297850 622132
rect 297800 621908 297872 622032
rect 297800 621808 297850 621908
rect 297800 621684 297872 621808
rect 297800 621584 297850 621684
rect 297800 621460 297872 621584
rect 297800 621360 297850 621460
rect 297800 621236 297872 621360
rect 297800 621136 297850 621236
rect 297800 621012 297872 621136
rect 297800 620912 297850 621012
rect 297800 620788 297872 620912
rect 297800 620688 297850 620788
rect 297800 620564 297872 620688
rect 297800 620464 297850 620564
rect 297800 620340 297872 620464
rect 297800 620240 297850 620340
rect 297800 620116 297872 620240
rect 297800 620016 297850 620116
rect 297800 619892 297872 620016
rect 297800 619792 297850 619892
rect 297800 619668 297872 619792
rect 297800 619568 297850 619668
rect 297800 619444 297872 619568
rect 297800 619344 297850 619444
rect 297800 619220 297872 619344
rect 297800 619120 297850 619220
rect 297800 618996 297872 619120
rect 297800 618896 297850 618996
rect 297800 618772 297872 618896
rect 297800 618672 297850 618772
rect 297800 618548 297872 618672
rect 297800 618448 297850 618548
rect 297800 618324 297872 618448
rect 297800 618224 297850 618324
rect 297800 618100 297872 618224
rect 297800 618000 297850 618100
rect 297800 616472 297872 618000
rect 298872 616472 298888 640624
rect 315670 637068 316544 637500
rect 319568 637438 322022 637500
rect 319568 637068 321452 637438
rect 315670 637022 316274 637068
rect 312432 637006 313034 637022
rect 312432 636114 312448 637006
rect 312422 635672 312448 636114
rect 312432 631612 312448 635672
rect 312428 631108 312448 631612
rect 312432 630702 312448 631108
rect 313018 636114 313034 637006
rect 315670 637006 316278 637022
rect 318998 637006 321452 637068
rect 335110 637006 335934 637438
rect 315670 636510 315692 637006
rect 315676 636114 315692 636510
rect 313018 635682 313272 636114
rect 313842 635682 314090 636114
rect 314660 635682 314908 636114
rect 315478 635682 315692 636114
rect 313018 635672 315692 635682
rect 313018 631612 313034 635672
rect 315676 632358 315692 635672
rect 316262 632764 316278 637006
rect 320636 632768 320652 637006
rect 315478 631926 315692 632358
rect 313272 631616 313842 631926
rect 315676 631616 315692 631926
rect 316262 632336 316544 632764
rect 317114 632336 317220 632768
rect 318882 632336 318998 632768
rect 319568 632336 320652 632768
rect 316262 632238 317220 632336
rect 318882 632238 320652 632336
rect 313272 631612 315692 631616
rect 313018 631108 315692 631612
rect 313018 630702 313034 631108
rect 312432 630686 313034 630702
rect 315676 630702 315692 631108
rect 316262 631616 316278 632238
rect 316262 631108 316288 631616
rect 316262 630702 316278 631108
rect 320636 630702 320652 632238
rect 321222 630702 321238 637006
rect 335324 630702 335340 637006
rect 335910 630702 335926 637006
rect 315676 630686 316278 630702
rect 320628 630270 321452 630702
rect 335110 630270 335934 630702
rect 334648 627708 341088 627740
rect 334648 627674 334782 627708
rect 334816 627674 334872 627708
rect 334906 627674 334962 627708
rect 334996 627674 335052 627708
rect 335086 627674 335142 627708
rect 335176 627674 335232 627708
rect 335266 627674 335322 627708
rect 335356 627674 335412 627708
rect 335446 627674 335502 627708
rect 335536 627674 335592 627708
rect 335626 627674 335682 627708
rect 335716 627674 335772 627708
rect 335806 627674 336070 627708
rect 336104 627674 336160 627708
rect 336194 627674 336250 627708
rect 336284 627674 336340 627708
rect 336374 627674 336430 627708
rect 336464 627674 336520 627708
rect 336554 627674 336610 627708
rect 336644 627674 336700 627708
rect 336734 627674 336790 627708
rect 336824 627674 336880 627708
rect 336914 627674 336970 627708
rect 337004 627674 337060 627708
rect 337094 627674 337358 627708
rect 337392 627674 337448 627708
rect 337482 627674 337538 627708
rect 337572 627674 337628 627708
rect 337662 627674 337718 627708
rect 337752 627674 337808 627708
rect 337842 627674 337898 627708
rect 337932 627674 337988 627708
rect 338022 627674 338078 627708
rect 338112 627674 338168 627708
rect 338202 627674 338258 627708
rect 338292 627674 338348 627708
rect 338382 627674 338646 627708
rect 338680 627674 338736 627708
rect 338770 627674 338826 627708
rect 338860 627674 338916 627708
rect 338950 627674 339006 627708
rect 339040 627674 339096 627708
rect 339130 627674 339186 627708
rect 339220 627674 339276 627708
rect 339310 627674 339366 627708
rect 339400 627674 339456 627708
rect 339490 627674 339546 627708
rect 339580 627674 339636 627708
rect 339670 627674 339934 627708
rect 339968 627674 340024 627708
rect 340058 627674 340114 627708
rect 340148 627674 340204 627708
rect 340238 627674 340294 627708
rect 340328 627674 340384 627708
rect 340418 627674 340474 627708
rect 340508 627674 340564 627708
rect 340598 627674 340654 627708
rect 340688 627674 340744 627708
rect 340778 627674 340834 627708
rect 340868 627674 340924 627708
rect 340958 627674 341088 627708
rect 334648 627641 341088 627674
rect 334648 627624 334888 627641
rect 334648 627590 334681 627624
rect 334715 627590 334888 627624
rect 334648 627577 334888 627590
rect 335688 627624 336188 627641
rect 335688 627590 335868 627624
rect 335902 627590 335969 627624
rect 336003 627590 336188 627624
rect 335688 627577 336188 627590
rect 336988 627624 337388 627641
rect 336988 627590 337156 627624
rect 337190 627590 337257 627624
rect 337291 627590 337388 627624
rect 336988 627577 337388 627590
rect 338288 627624 338688 627641
rect 338288 627590 338444 627624
rect 338478 627590 338545 627624
rect 338579 627590 338688 627624
rect 338288 627577 338688 627590
rect 339588 627624 339988 627641
rect 339588 627590 339732 627624
rect 339766 627590 339833 627624
rect 339867 627590 339988 627624
rect 339588 627577 339988 627590
rect 340888 627624 341088 627641
rect 340888 627590 341020 627624
rect 341054 627590 341088 627624
rect 340888 627577 341088 627590
rect 334648 627558 341088 627577
rect 334648 627534 334922 627558
rect 334648 627500 334681 627534
rect 334715 627524 334922 627534
rect 334956 627524 335012 627558
rect 335046 627524 335102 627558
rect 335136 627524 335192 627558
rect 335226 627524 335282 627558
rect 335316 627524 335372 627558
rect 335406 627524 335462 627558
rect 335496 627524 335552 627558
rect 335586 627524 335642 627558
rect 335676 627534 336210 627558
rect 335676 627524 335868 627534
rect 334715 627505 335868 627524
rect 334715 627500 334888 627505
rect 334648 627464 334888 627500
rect 334648 627444 334830 627464
rect 334648 627410 334681 627444
rect 334715 627430 334830 627444
rect 334864 627430 334888 627464
rect 335688 627500 335868 627505
rect 335902 627500 335969 627534
rect 336003 627524 336210 627534
rect 336244 627524 336300 627558
rect 336334 627524 336390 627558
rect 336424 627524 336480 627558
rect 336514 627524 336570 627558
rect 336604 627524 336660 627558
rect 336694 627524 336750 627558
rect 336784 627524 336840 627558
rect 336874 627524 336930 627558
rect 336964 627534 337498 627558
rect 336964 627524 337156 627534
rect 336003 627505 337156 627524
rect 336003 627500 336188 627505
rect 335688 627464 336188 627500
rect 335688 627445 336118 627464
rect 334715 627410 334888 627430
rect 334648 627374 334888 627410
rect 334648 627354 334830 627374
rect 334648 627320 334681 627354
rect 334715 627340 334830 627354
rect 334864 627340 334888 627374
rect 334715 627320 334888 627340
rect 334648 627284 334888 627320
rect 334648 627264 334830 627284
rect 334648 627230 334681 627264
rect 334715 627250 334830 627264
rect 334864 627250 334888 627284
rect 334715 627230 334888 627250
rect 334648 627194 334888 627230
rect 334648 627174 334830 627194
rect 334648 627140 334681 627174
rect 334715 627160 334830 627174
rect 334864 627160 334888 627194
rect 334715 627140 334888 627160
rect 334648 627104 334888 627140
rect 334648 627084 334830 627104
rect 334648 627050 334681 627084
rect 334715 627070 334830 627084
rect 334864 627070 334888 627104
rect 334715 627050 334888 627070
rect 334648 627014 334888 627050
rect 334648 626994 334830 627014
rect 334648 626960 334681 626994
rect 334715 626980 334830 626994
rect 334864 626980 334888 627014
rect 334715 626960 334888 626980
rect 334648 626924 334888 626960
rect 334648 626904 334830 626924
rect 334648 626870 334681 626904
rect 334715 626890 334830 626904
rect 334864 626890 334888 626924
rect 334715 626870 334888 626890
rect 334648 626834 334888 626870
rect 334648 626814 334830 626834
rect 334648 626780 334681 626814
rect 334715 626800 334830 626814
rect 334864 626800 334888 626834
rect 334715 626780 334888 626800
rect 334648 626744 334888 626780
rect 334945 627382 335639 627443
rect 334945 627348 335004 627382
rect 335038 627370 335094 627382
rect 335066 627348 335094 627370
rect 335128 627370 335184 627382
rect 335128 627348 335132 627370
rect 334945 627336 335032 627348
rect 335066 627336 335132 627348
rect 335166 627348 335184 627370
rect 335218 627370 335274 627382
rect 335218 627348 335232 627370
rect 335166 627336 335232 627348
rect 335266 627348 335274 627370
rect 335308 627370 335364 627382
rect 335398 627370 335454 627382
rect 335488 627370 335544 627382
rect 335308 627348 335332 627370
rect 335398 627348 335432 627370
rect 335488 627348 335532 627370
rect 335578 627348 335639 627382
rect 335266 627336 335332 627348
rect 335366 627336 335432 627348
rect 335466 627336 335532 627348
rect 335566 627336 335639 627348
rect 334945 627292 335639 627336
rect 334945 627258 335004 627292
rect 335038 627270 335094 627292
rect 335066 627258 335094 627270
rect 335128 627270 335184 627292
rect 335128 627258 335132 627270
rect 334945 627236 335032 627258
rect 335066 627236 335132 627258
rect 335166 627258 335184 627270
rect 335218 627270 335274 627292
rect 335218 627258 335232 627270
rect 335166 627236 335232 627258
rect 335266 627258 335274 627270
rect 335308 627270 335364 627292
rect 335398 627270 335454 627292
rect 335488 627270 335544 627292
rect 335308 627258 335332 627270
rect 335398 627258 335432 627270
rect 335488 627258 335532 627270
rect 335578 627258 335639 627292
rect 335266 627236 335332 627258
rect 335366 627236 335432 627258
rect 335466 627236 335532 627258
rect 335566 627236 335639 627258
rect 334945 627202 335639 627236
rect 334945 627168 335004 627202
rect 335038 627170 335094 627202
rect 335066 627168 335094 627170
rect 335128 627170 335184 627202
rect 335128 627168 335132 627170
rect 334945 627136 335032 627168
rect 335066 627136 335132 627168
rect 335166 627168 335184 627170
rect 335218 627170 335274 627202
rect 335218 627168 335232 627170
rect 335166 627136 335232 627168
rect 335266 627168 335274 627170
rect 335308 627170 335364 627202
rect 335398 627170 335454 627202
rect 335488 627170 335544 627202
rect 335308 627168 335332 627170
rect 335398 627168 335432 627170
rect 335488 627168 335532 627170
rect 335578 627168 335639 627202
rect 335266 627136 335332 627168
rect 335366 627136 335432 627168
rect 335466 627136 335532 627168
rect 335566 627136 335639 627168
rect 334945 627112 335639 627136
rect 334945 627078 335004 627112
rect 335038 627078 335094 627112
rect 335128 627078 335184 627112
rect 335218 627078 335274 627112
rect 335308 627078 335364 627112
rect 335398 627078 335454 627112
rect 335488 627078 335544 627112
rect 335578 627078 335639 627112
rect 334945 627070 335639 627078
rect 334945 627036 335032 627070
rect 335066 627036 335132 627070
rect 335166 627036 335232 627070
rect 335266 627036 335332 627070
rect 335366 627036 335432 627070
rect 335466 627036 335532 627070
rect 335566 627036 335639 627070
rect 334945 627022 335639 627036
rect 334945 626988 335004 627022
rect 335038 626988 335094 627022
rect 335128 626988 335184 627022
rect 335218 626988 335274 627022
rect 335308 626988 335364 627022
rect 335398 626988 335454 627022
rect 335488 626988 335544 627022
rect 335578 626988 335639 627022
rect 334945 626970 335639 626988
rect 334945 626936 335032 626970
rect 335066 626936 335132 626970
rect 335166 626936 335232 626970
rect 335266 626936 335332 626970
rect 335366 626936 335432 626970
rect 335466 626936 335532 626970
rect 335566 626936 335639 626970
rect 334945 626932 335639 626936
rect 334945 626898 335004 626932
rect 335038 626898 335094 626932
rect 335128 626898 335184 626932
rect 335218 626898 335274 626932
rect 335308 626898 335364 626932
rect 335398 626898 335454 626932
rect 335488 626898 335544 626932
rect 335578 626898 335639 626932
rect 334945 626870 335639 626898
rect 334945 626842 335032 626870
rect 335066 626842 335132 626870
rect 334945 626808 335004 626842
rect 335066 626836 335094 626842
rect 335038 626808 335094 626836
rect 335128 626836 335132 626842
rect 335166 626842 335232 626870
rect 335166 626836 335184 626842
rect 335128 626808 335184 626836
rect 335218 626836 335232 626842
rect 335266 626842 335332 626870
rect 335366 626842 335432 626870
rect 335466 626842 335532 626870
rect 335566 626842 335639 626870
rect 335266 626836 335274 626842
rect 335218 626808 335274 626836
rect 335308 626836 335332 626842
rect 335398 626836 335432 626842
rect 335488 626836 335532 626842
rect 335308 626808 335364 626836
rect 335398 626808 335454 626836
rect 335488 626808 335544 626836
rect 335578 626808 335639 626842
rect 334945 626749 335639 626808
rect 335688 627411 335720 627445
rect 335754 627444 336118 627445
rect 335754 627411 335868 627444
rect 335688 627410 335868 627411
rect 335902 627410 335969 627444
rect 336003 627430 336118 627444
rect 336152 627430 336188 627464
rect 336988 627500 337156 627505
rect 337190 627500 337257 627534
rect 337291 627524 337498 627534
rect 337532 627524 337588 627558
rect 337622 627524 337678 627558
rect 337712 627524 337768 627558
rect 337802 627524 337858 627558
rect 337892 627524 337948 627558
rect 337982 627524 338038 627558
rect 338072 627524 338128 627558
rect 338162 627524 338218 627558
rect 338252 627534 338786 627558
rect 338252 627524 338444 627534
rect 337291 627505 338444 627524
rect 337291 627500 337459 627505
rect 336988 627464 337459 627500
rect 336988 627445 337406 627464
rect 336003 627410 336188 627430
rect 335688 627374 336188 627410
rect 335688 627355 336118 627374
rect 335688 627321 335720 627355
rect 335754 627354 336118 627355
rect 335754 627321 335868 627354
rect 335688 627320 335868 627321
rect 335902 627320 335969 627354
rect 336003 627340 336118 627354
rect 336152 627340 336188 627374
rect 336003 627320 336188 627340
rect 335688 627284 336188 627320
rect 335688 627265 336118 627284
rect 335688 627231 335720 627265
rect 335754 627264 336118 627265
rect 335754 627231 335868 627264
rect 335688 627230 335868 627231
rect 335902 627230 335969 627264
rect 336003 627250 336118 627264
rect 336152 627250 336188 627284
rect 336003 627230 336188 627250
rect 335688 627194 336188 627230
rect 335688 627175 336118 627194
rect 335688 627141 335720 627175
rect 335754 627174 336118 627175
rect 335754 627141 335868 627174
rect 335688 627140 335868 627141
rect 335902 627140 335969 627174
rect 336003 627160 336118 627174
rect 336152 627160 336188 627194
rect 336003 627140 336188 627160
rect 335688 627104 336188 627140
rect 335688 627085 336118 627104
rect 335688 627051 335720 627085
rect 335754 627084 336118 627085
rect 335754 627051 335868 627084
rect 335688 627050 335868 627051
rect 335902 627050 335969 627084
rect 336003 627070 336118 627084
rect 336152 627070 336188 627104
rect 336003 627050 336188 627070
rect 335688 627014 336188 627050
rect 335688 626995 336118 627014
rect 335688 626961 335720 626995
rect 335754 626994 336118 626995
rect 335754 626961 335868 626994
rect 335688 626960 335868 626961
rect 335902 626960 335969 626994
rect 336003 626980 336118 626994
rect 336152 626980 336188 627014
rect 336003 626960 336188 626980
rect 335688 626924 336188 626960
rect 335688 626905 336118 626924
rect 335688 626871 335720 626905
rect 335754 626904 336118 626905
rect 335754 626871 335868 626904
rect 335688 626870 335868 626871
rect 335902 626870 335969 626904
rect 336003 626890 336118 626904
rect 336152 626890 336188 626924
rect 336003 626870 336188 626890
rect 335688 626834 336188 626870
rect 335688 626815 336118 626834
rect 335688 626781 335720 626815
rect 335754 626814 336118 626815
rect 335754 626781 335868 626814
rect 335688 626780 335868 626781
rect 335902 626780 335969 626814
rect 336003 626800 336118 626814
rect 336152 626800 336188 626834
rect 336003 626780 336188 626800
rect 334648 626724 334830 626744
rect 334648 626690 334681 626724
rect 334715 626710 334830 626724
rect 334864 626710 334888 626744
rect 334715 626690 334888 626710
rect 334648 626687 334888 626690
rect 335688 626744 336188 626780
rect 336233 627382 336927 627443
rect 336233 627348 336292 627382
rect 336326 627370 336382 627382
rect 336354 627348 336382 627370
rect 336416 627370 336472 627382
rect 336416 627348 336420 627370
rect 336233 627336 336320 627348
rect 336354 627336 336420 627348
rect 336454 627348 336472 627370
rect 336506 627370 336562 627382
rect 336506 627348 336520 627370
rect 336454 627336 336520 627348
rect 336554 627348 336562 627370
rect 336596 627370 336652 627382
rect 336686 627370 336742 627382
rect 336776 627370 336832 627382
rect 336596 627348 336620 627370
rect 336686 627348 336720 627370
rect 336776 627348 336820 627370
rect 336866 627348 336927 627382
rect 336554 627336 336620 627348
rect 336654 627336 336720 627348
rect 336754 627336 336820 627348
rect 336854 627336 336927 627348
rect 336233 627292 336927 627336
rect 336233 627258 336292 627292
rect 336326 627270 336382 627292
rect 336354 627258 336382 627270
rect 336416 627270 336472 627292
rect 336416 627258 336420 627270
rect 336233 627236 336320 627258
rect 336354 627236 336420 627258
rect 336454 627258 336472 627270
rect 336506 627270 336562 627292
rect 336506 627258 336520 627270
rect 336454 627236 336520 627258
rect 336554 627258 336562 627270
rect 336596 627270 336652 627292
rect 336686 627270 336742 627292
rect 336776 627270 336832 627292
rect 336596 627258 336620 627270
rect 336686 627258 336720 627270
rect 336776 627258 336820 627270
rect 336866 627258 336927 627292
rect 336554 627236 336620 627258
rect 336654 627236 336720 627258
rect 336754 627236 336820 627258
rect 336854 627236 336927 627258
rect 336233 627202 336927 627236
rect 336233 627168 336292 627202
rect 336326 627170 336382 627202
rect 336354 627168 336382 627170
rect 336416 627170 336472 627202
rect 336416 627168 336420 627170
rect 336233 627136 336320 627168
rect 336354 627136 336420 627168
rect 336454 627168 336472 627170
rect 336506 627170 336562 627202
rect 336506 627168 336520 627170
rect 336454 627136 336520 627168
rect 336554 627168 336562 627170
rect 336596 627170 336652 627202
rect 336686 627170 336742 627202
rect 336776 627170 336832 627202
rect 336596 627168 336620 627170
rect 336686 627168 336720 627170
rect 336776 627168 336820 627170
rect 336866 627168 336927 627202
rect 336554 627136 336620 627168
rect 336654 627136 336720 627168
rect 336754 627136 336820 627168
rect 336854 627136 336927 627168
rect 336233 627112 336927 627136
rect 336233 627078 336292 627112
rect 336326 627078 336382 627112
rect 336416 627078 336472 627112
rect 336506 627078 336562 627112
rect 336596 627078 336652 627112
rect 336686 627078 336742 627112
rect 336776 627078 336832 627112
rect 336866 627078 336927 627112
rect 336233 627070 336927 627078
rect 336233 627036 336320 627070
rect 336354 627036 336420 627070
rect 336454 627036 336520 627070
rect 336554 627036 336620 627070
rect 336654 627036 336720 627070
rect 336754 627036 336820 627070
rect 336854 627036 336927 627070
rect 336233 627022 336927 627036
rect 336233 626988 336292 627022
rect 336326 626988 336382 627022
rect 336416 626988 336472 627022
rect 336506 626988 336562 627022
rect 336596 626988 336652 627022
rect 336686 626988 336742 627022
rect 336776 626988 336832 627022
rect 336866 626988 336927 627022
rect 336233 626970 336927 626988
rect 336233 626936 336320 626970
rect 336354 626936 336420 626970
rect 336454 626936 336520 626970
rect 336554 626936 336620 626970
rect 336654 626936 336720 626970
rect 336754 626936 336820 626970
rect 336854 626936 336927 626970
rect 336233 626932 336927 626936
rect 336233 626898 336292 626932
rect 336326 626898 336382 626932
rect 336416 626898 336472 626932
rect 336506 626898 336562 626932
rect 336596 626898 336652 626932
rect 336686 626898 336742 626932
rect 336776 626898 336832 626932
rect 336866 626898 336927 626932
rect 336233 626870 336927 626898
rect 336233 626842 336320 626870
rect 336354 626842 336420 626870
rect 336233 626808 336292 626842
rect 336354 626836 336382 626842
rect 336326 626808 336382 626836
rect 336416 626836 336420 626842
rect 336454 626842 336520 626870
rect 336454 626836 336472 626842
rect 336416 626808 336472 626836
rect 336506 626836 336520 626842
rect 336554 626842 336620 626870
rect 336654 626842 336720 626870
rect 336754 626842 336820 626870
rect 336854 626842 336927 626870
rect 336554 626836 336562 626842
rect 336506 626808 336562 626836
rect 336596 626836 336620 626842
rect 336686 626836 336720 626842
rect 336776 626836 336820 626842
rect 336596 626808 336652 626836
rect 336686 626808 336742 626836
rect 336776 626808 336832 626836
rect 336866 626808 336927 626842
rect 336233 626749 336927 626808
rect 336988 627411 337008 627445
rect 337042 627444 337406 627445
rect 337042 627411 337156 627444
rect 336988 627410 337156 627411
rect 337190 627410 337257 627444
rect 337291 627430 337406 627444
rect 337440 627430 337459 627464
rect 338277 627500 338444 627505
rect 338478 627500 338545 627534
rect 338579 627524 338786 627534
rect 338820 627524 338876 627558
rect 338910 627524 338966 627558
rect 339000 627524 339056 627558
rect 339090 627524 339146 627558
rect 339180 627524 339236 627558
rect 339270 627524 339326 627558
rect 339360 627524 339416 627558
rect 339450 627524 339506 627558
rect 339540 627534 340074 627558
rect 339540 627524 339732 627534
rect 338579 627505 339732 627524
rect 338579 627500 338747 627505
rect 338277 627464 338747 627500
rect 338277 627445 338694 627464
rect 337291 627410 337459 627430
rect 336988 627374 337459 627410
rect 336988 627355 337406 627374
rect 336988 627321 337008 627355
rect 337042 627354 337406 627355
rect 337042 627321 337156 627354
rect 336988 627320 337156 627321
rect 337190 627320 337257 627354
rect 337291 627340 337406 627354
rect 337440 627340 337459 627374
rect 337291 627320 337459 627340
rect 336988 627284 337459 627320
rect 336988 627265 337406 627284
rect 336988 627231 337008 627265
rect 337042 627264 337406 627265
rect 337042 627231 337156 627264
rect 336988 627230 337156 627231
rect 337190 627230 337257 627264
rect 337291 627250 337406 627264
rect 337440 627250 337459 627284
rect 337291 627230 337459 627250
rect 336988 627194 337459 627230
rect 336988 627175 337406 627194
rect 336988 627141 337008 627175
rect 337042 627174 337406 627175
rect 337042 627141 337156 627174
rect 336988 627140 337156 627141
rect 337190 627140 337257 627174
rect 337291 627160 337406 627174
rect 337440 627160 337459 627194
rect 337291 627140 337459 627160
rect 336988 627104 337459 627140
rect 336988 627085 337406 627104
rect 336988 627051 337008 627085
rect 337042 627084 337406 627085
rect 337042 627051 337156 627084
rect 336988 627050 337156 627051
rect 337190 627050 337257 627084
rect 337291 627070 337406 627084
rect 337440 627070 337459 627104
rect 337291 627050 337459 627070
rect 336988 627014 337459 627050
rect 336988 626995 337406 627014
rect 336988 626961 337008 626995
rect 337042 626994 337406 626995
rect 337042 626961 337156 626994
rect 336988 626960 337156 626961
rect 337190 626960 337257 626994
rect 337291 626980 337406 626994
rect 337440 626980 337459 627014
rect 337291 626960 337459 626980
rect 336988 626924 337459 626960
rect 336988 626905 337406 626924
rect 336988 626871 337008 626905
rect 337042 626904 337406 626905
rect 337042 626871 337156 626904
rect 336988 626870 337156 626871
rect 337190 626870 337257 626904
rect 337291 626890 337406 626904
rect 337440 626890 337459 626924
rect 337291 626870 337459 626890
rect 336988 626834 337459 626870
rect 336988 626815 337406 626834
rect 336988 626781 337008 626815
rect 337042 626814 337406 626815
rect 337042 626781 337156 626814
rect 336988 626780 337156 626781
rect 337190 626780 337257 626814
rect 337291 626800 337406 626814
rect 337440 626800 337459 626834
rect 337291 626780 337459 626800
rect 335688 626725 336118 626744
rect 335688 626691 335720 626725
rect 335754 626724 336118 626725
rect 335754 626691 335868 626724
rect 335688 626690 335868 626691
rect 335902 626690 335969 626724
rect 336003 626710 336118 626724
rect 336152 626710 336188 626744
rect 336003 626690 336188 626710
rect 335688 626687 336188 626690
rect 336988 626744 337459 626780
rect 337521 627382 338215 627443
rect 337521 627348 337580 627382
rect 337614 627370 337670 627382
rect 337642 627348 337670 627370
rect 337704 627370 337760 627382
rect 337704 627348 337708 627370
rect 337521 627336 337608 627348
rect 337642 627336 337708 627348
rect 337742 627348 337760 627370
rect 337794 627370 337850 627382
rect 337794 627348 337808 627370
rect 337742 627336 337808 627348
rect 337842 627348 337850 627370
rect 337884 627370 337940 627382
rect 337974 627370 338030 627382
rect 338064 627370 338120 627382
rect 337884 627348 337908 627370
rect 337974 627348 338008 627370
rect 338064 627348 338108 627370
rect 338154 627348 338215 627382
rect 337842 627336 337908 627348
rect 337942 627336 338008 627348
rect 338042 627336 338108 627348
rect 338142 627336 338215 627348
rect 337521 627292 338215 627336
rect 337521 627258 337580 627292
rect 337614 627270 337670 627292
rect 337642 627258 337670 627270
rect 337704 627270 337760 627292
rect 337704 627258 337708 627270
rect 337521 627236 337608 627258
rect 337642 627236 337708 627258
rect 337742 627258 337760 627270
rect 337794 627270 337850 627292
rect 337794 627258 337808 627270
rect 337742 627236 337808 627258
rect 337842 627258 337850 627270
rect 337884 627270 337940 627292
rect 337974 627270 338030 627292
rect 338064 627270 338120 627292
rect 337884 627258 337908 627270
rect 337974 627258 338008 627270
rect 338064 627258 338108 627270
rect 338154 627258 338215 627292
rect 337842 627236 337908 627258
rect 337942 627236 338008 627258
rect 338042 627236 338108 627258
rect 338142 627236 338215 627258
rect 337521 627202 338215 627236
rect 337521 627168 337580 627202
rect 337614 627170 337670 627202
rect 337642 627168 337670 627170
rect 337704 627170 337760 627202
rect 337704 627168 337708 627170
rect 337521 627136 337608 627168
rect 337642 627136 337708 627168
rect 337742 627168 337760 627170
rect 337794 627170 337850 627202
rect 337794 627168 337808 627170
rect 337742 627136 337808 627168
rect 337842 627168 337850 627170
rect 337884 627170 337940 627202
rect 337974 627170 338030 627202
rect 338064 627170 338120 627202
rect 337884 627168 337908 627170
rect 337974 627168 338008 627170
rect 338064 627168 338108 627170
rect 338154 627168 338215 627202
rect 337842 627136 337908 627168
rect 337942 627136 338008 627168
rect 338042 627136 338108 627168
rect 338142 627136 338215 627168
rect 337521 627112 338215 627136
rect 337521 627078 337580 627112
rect 337614 627078 337670 627112
rect 337704 627078 337760 627112
rect 337794 627078 337850 627112
rect 337884 627078 337940 627112
rect 337974 627078 338030 627112
rect 338064 627078 338120 627112
rect 338154 627078 338215 627112
rect 337521 627070 338215 627078
rect 337521 627036 337608 627070
rect 337642 627036 337708 627070
rect 337742 627036 337808 627070
rect 337842 627036 337908 627070
rect 337942 627036 338008 627070
rect 338042 627036 338108 627070
rect 338142 627036 338215 627070
rect 337521 627022 338215 627036
rect 337521 626988 337580 627022
rect 337614 626988 337670 627022
rect 337704 626988 337760 627022
rect 337794 626988 337850 627022
rect 337884 626988 337940 627022
rect 337974 626988 338030 627022
rect 338064 626988 338120 627022
rect 338154 626988 338215 627022
rect 337521 626970 338215 626988
rect 337521 626936 337608 626970
rect 337642 626936 337708 626970
rect 337742 626936 337808 626970
rect 337842 626936 337908 626970
rect 337942 626936 338008 626970
rect 338042 626936 338108 626970
rect 338142 626936 338215 626970
rect 337521 626932 338215 626936
rect 337521 626898 337580 626932
rect 337614 626898 337670 626932
rect 337704 626898 337760 626932
rect 337794 626898 337850 626932
rect 337884 626898 337940 626932
rect 337974 626898 338030 626932
rect 338064 626898 338120 626932
rect 338154 626898 338215 626932
rect 337521 626870 338215 626898
rect 337521 626842 337608 626870
rect 337642 626842 337708 626870
rect 337521 626808 337580 626842
rect 337642 626836 337670 626842
rect 337614 626808 337670 626836
rect 337704 626836 337708 626842
rect 337742 626842 337808 626870
rect 337742 626836 337760 626842
rect 337704 626808 337760 626836
rect 337794 626836 337808 626842
rect 337842 626842 337908 626870
rect 337942 626842 338008 626870
rect 338042 626842 338108 626870
rect 338142 626842 338215 626870
rect 337842 626836 337850 626842
rect 337794 626808 337850 626836
rect 337884 626836 337908 626842
rect 337974 626836 338008 626842
rect 338064 626836 338108 626842
rect 337884 626808 337940 626836
rect 337974 626808 338030 626836
rect 338064 626808 338120 626836
rect 338154 626808 338215 626842
rect 337521 626749 338215 626808
rect 338277 627411 338296 627445
rect 338330 627444 338694 627445
rect 338330 627411 338444 627444
rect 338277 627410 338444 627411
rect 338478 627410 338545 627444
rect 338579 627430 338694 627444
rect 338728 627430 338747 627464
rect 339565 627500 339732 627505
rect 339766 627500 339833 627534
rect 339867 627524 340074 627534
rect 340108 627524 340164 627558
rect 340198 627524 340254 627558
rect 340288 627524 340344 627558
rect 340378 627524 340434 627558
rect 340468 627524 340524 627558
rect 340558 627524 340614 627558
rect 340648 627524 340704 627558
rect 340738 627524 340794 627558
rect 340828 627534 341088 627558
rect 340828 627524 341020 627534
rect 339867 627505 341020 627524
rect 339867 627500 340035 627505
rect 339565 627464 340035 627500
rect 339565 627445 339982 627464
rect 338579 627410 338747 627430
rect 338277 627374 338747 627410
rect 338277 627355 338694 627374
rect 338277 627321 338296 627355
rect 338330 627354 338694 627355
rect 338330 627321 338444 627354
rect 338277 627320 338444 627321
rect 338478 627320 338545 627354
rect 338579 627340 338694 627354
rect 338728 627340 338747 627374
rect 338579 627320 338747 627340
rect 338277 627284 338747 627320
rect 338277 627265 338694 627284
rect 338277 627231 338296 627265
rect 338330 627264 338694 627265
rect 338330 627231 338444 627264
rect 338277 627230 338444 627231
rect 338478 627230 338545 627264
rect 338579 627250 338694 627264
rect 338728 627250 338747 627284
rect 338579 627230 338747 627250
rect 338277 627194 338747 627230
rect 338277 627175 338694 627194
rect 338277 627141 338296 627175
rect 338330 627174 338694 627175
rect 338330 627141 338444 627174
rect 338277 627140 338444 627141
rect 338478 627140 338545 627174
rect 338579 627160 338694 627174
rect 338728 627160 338747 627194
rect 338579 627140 338747 627160
rect 338277 627104 338747 627140
rect 338277 627085 338694 627104
rect 338277 627051 338296 627085
rect 338330 627084 338694 627085
rect 338330 627051 338444 627084
rect 338277 627050 338444 627051
rect 338478 627050 338545 627084
rect 338579 627070 338694 627084
rect 338728 627070 338747 627104
rect 338579 627050 338747 627070
rect 338277 627014 338747 627050
rect 338277 626995 338694 627014
rect 338277 626961 338296 626995
rect 338330 626994 338694 626995
rect 338330 626961 338444 626994
rect 338277 626960 338444 626961
rect 338478 626960 338545 626994
rect 338579 626980 338694 626994
rect 338728 626980 338747 627014
rect 338579 626960 338747 626980
rect 338277 626924 338747 626960
rect 338277 626905 338694 626924
rect 338277 626871 338296 626905
rect 338330 626904 338694 626905
rect 338330 626871 338444 626904
rect 338277 626870 338444 626871
rect 338478 626870 338545 626904
rect 338579 626890 338694 626904
rect 338728 626890 338747 626924
rect 338579 626870 338747 626890
rect 338277 626834 338747 626870
rect 338277 626815 338694 626834
rect 338277 626781 338296 626815
rect 338330 626814 338694 626815
rect 338330 626781 338444 626814
rect 338277 626780 338444 626781
rect 338478 626780 338545 626814
rect 338579 626800 338694 626814
rect 338728 626800 338747 626834
rect 338579 626780 338747 626800
rect 336988 626725 337406 626744
rect 336988 626691 337008 626725
rect 337042 626724 337406 626725
rect 337042 626691 337156 626724
rect 336988 626690 337156 626691
rect 337190 626690 337257 626724
rect 337291 626710 337406 626724
rect 337440 626710 337459 626744
rect 337291 626690 337459 626710
rect 336988 626687 337459 626690
rect 338277 626744 338747 626780
rect 338809 627382 339503 627443
rect 338809 627348 338868 627382
rect 338902 627370 338958 627382
rect 338930 627348 338958 627370
rect 338992 627370 339048 627382
rect 338992 627348 338996 627370
rect 338809 627336 338896 627348
rect 338930 627336 338996 627348
rect 339030 627348 339048 627370
rect 339082 627370 339138 627382
rect 339082 627348 339096 627370
rect 339030 627336 339096 627348
rect 339130 627348 339138 627370
rect 339172 627370 339228 627382
rect 339262 627370 339318 627382
rect 339352 627370 339408 627382
rect 339172 627348 339196 627370
rect 339262 627348 339296 627370
rect 339352 627348 339396 627370
rect 339442 627348 339503 627382
rect 339130 627336 339196 627348
rect 339230 627336 339296 627348
rect 339330 627336 339396 627348
rect 339430 627336 339503 627348
rect 338809 627292 339503 627336
rect 338809 627258 338868 627292
rect 338902 627270 338958 627292
rect 338930 627258 338958 627270
rect 338992 627270 339048 627292
rect 338992 627258 338996 627270
rect 338809 627236 338896 627258
rect 338930 627236 338996 627258
rect 339030 627258 339048 627270
rect 339082 627270 339138 627292
rect 339082 627258 339096 627270
rect 339030 627236 339096 627258
rect 339130 627258 339138 627270
rect 339172 627270 339228 627292
rect 339262 627270 339318 627292
rect 339352 627270 339408 627292
rect 339172 627258 339196 627270
rect 339262 627258 339296 627270
rect 339352 627258 339396 627270
rect 339442 627258 339503 627292
rect 339130 627236 339196 627258
rect 339230 627236 339296 627258
rect 339330 627236 339396 627258
rect 339430 627236 339503 627258
rect 338809 627202 339503 627236
rect 338809 627168 338868 627202
rect 338902 627170 338958 627202
rect 338930 627168 338958 627170
rect 338992 627170 339048 627202
rect 338992 627168 338996 627170
rect 338809 627136 338896 627168
rect 338930 627136 338996 627168
rect 339030 627168 339048 627170
rect 339082 627170 339138 627202
rect 339082 627168 339096 627170
rect 339030 627136 339096 627168
rect 339130 627168 339138 627170
rect 339172 627170 339228 627202
rect 339262 627170 339318 627202
rect 339352 627170 339408 627202
rect 339172 627168 339196 627170
rect 339262 627168 339296 627170
rect 339352 627168 339396 627170
rect 339442 627168 339503 627202
rect 339130 627136 339196 627168
rect 339230 627136 339296 627168
rect 339330 627136 339396 627168
rect 339430 627136 339503 627168
rect 338809 627112 339503 627136
rect 338809 627078 338868 627112
rect 338902 627078 338958 627112
rect 338992 627078 339048 627112
rect 339082 627078 339138 627112
rect 339172 627078 339228 627112
rect 339262 627078 339318 627112
rect 339352 627078 339408 627112
rect 339442 627078 339503 627112
rect 338809 627070 339503 627078
rect 338809 627036 338896 627070
rect 338930 627036 338996 627070
rect 339030 627036 339096 627070
rect 339130 627036 339196 627070
rect 339230 627036 339296 627070
rect 339330 627036 339396 627070
rect 339430 627036 339503 627070
rect 338809 627022 339503 627036
rect 338809 626988 338868 627022
rect 338902 626988 338958 627022
rect 338992 626988 339048 627022
rect 339082 626988 339138 627022
rect 339172 626988 339228 627022
rect 339262 626988 339318 627022
rect 339352 626988 339408 627022
rect 339442 626988 339503 627022
rect 338809 626970 339503 626988
rect 338809 626936 338896 626970
rect 338930 626936 338996 626970
rect 339030 626936 339096 626970
rect 339130 626936 339196 626970
rect 339230 626936 339296 626970
rect 339330 626936 339396 626970
rect 339430 626936 339503 626970
rect 338809 626932 339503 626936
rect 338809 626898 338868 626932
rect 338902 626898 338958 626932
rect 338992 626898 339048 626932
rect 339082 626898 339138 626932
rect 339172 626898 339228 626932
rect 339262 626898 339318 626932
rect 339352 626898 339408 626932
rect 339442 626898 339503 626932
rect 338809 626870 339503 626898
rect 338809 626842 338896 626870
rect 338930 626842 338996 626870
rect 338809 626808 338868 626842
rect 338930 626836 338958 626842
rect 338902 626808 338958 626836
rect 338992 626836 338996 626842
rect 339030 626842 339096 626870
rect 339030 626836 339048 626842
rect 338992 626808 339048 626836
rect 339082 626836 339096 626842
rect 339130 626842 339196 626870
rect 339230 626842 339296 626870
rect 339330 626842 339396 626870
rect 339430 626842 339503 626870
rect 339130 626836 339138 626842
rect 339082 626808 339138 626836
rect 339172 626836 339196 626842
rect 339262 626836 339296 626842
rect 339352 626836 339396 626842
rect 339172 626808 339228 626836
rect 339262 626808 339318 626836
rect 339352 626808 339408 626836
rect 339442 626808 339503 626842
rect 338809 626749 339503 626808
rect 339565 627411 339584 627445
rect 339618 627444 339982 627445
rect 339618 627411 339732 627444
rect 339565 627410 339732 627411
rect 339766 627410 339833 627444
rect 339867 627430 339982 627444
rect 340016 627430 340035 627464
rect 340853 627500 341020 627505
rect 341054 627500 341088 627534
rect 340853 627445 341088 627500
rect 339867 627410 340035 627430
rect 339565 627374 340035 627410
rect 339565 627355 339982 627374
rect 339565 627321 339584 627355
rect 339618 627354 339982 627355
rect 339618 627321 339732 627354
rect 339565 627320 339732 627321
rect 339766 627320 339833 627354
rect 339867 627340 339982 627354
rect 340016 627340 340035 627374
rect 339867 627320 340035 627340
rect 339565 627284 340035 627320
rect 339565 627265 339982 627284
rect 339565 627231 339584 627265
rect 339618 627264 339982 627265
rect 339618 627231 339732 627264
rect 339565 627230 339732 627231
rect 339766 627230 339833 627264
rect 339867 627250 339982 627264
rect 340016 627250 340035 627284
rect 339867 627230 340035 627250
rect 339565 627194 340035 627230
rect 339565 627175 339982 627194
rect 339565 627141 339584 627175
rect 339618 627174 339982 627175
rect 339618 627141 339732 627174
rect 339565 627140 339732 627141
rect 339766 627140 339833 627174
rect 339867 627160 339982 627174
rect 340016 627160 340035 627194
rect 339867 627140 340035 627160
rect 339565 627104 340035 627140
rect 339565 627085 339982 627104
rect 339565 627051 339584 627085
rect 339618 627084 339982 627085
rect 339618 627051 339732 627084
rect 339565 627050 339732 627051
rect 339766 627050 339833 627084
rect 339867 627070 339982 627084
rect 340016 627070 340035 627104
rect 339867 627050 340035 627070
rect 339565 627014 340035 627050
rect 339565 626995 339982 627014
rect 339565 626961 339584 626995
rect 339618 626994 339982 626995
rect 339618 626961 339732 626994
rect 339565 626960 339732 626961
rect 339766 626960 339833 626994
rect 339867 626980 339982 626994
rect 340016 626980 340035 627014
rect 339867 626960 340035 626980
rect 339565 626924 340035 626960
rect 339565 626905 339982 626924
rect 339565 626871 339584 626905
rect 339618 626904 339982 626905
rect 339618 626871 339732 626904
rect 339565 626870 339732 626871
rect 339766 626870 339833 626904
rect 339867 626890 339982 626904
rect 340016 626890 340035 626924
rect 339867 626870 340035 626890
rect 339565 626834 340035 626870
rect 339565 626815 339982 626834
rect 339565 626781 339584 626815
rect 339618 626814 339982 626815
rect 339618 626781 339732 626814
rect 339565 626780 339732 626781
rect 339766 626780 339833 626814
rect 339867 626800 339982 626814
rect 340016 626800 340035 626834
rect 339867 626780 340035 626800
rect 338277 626725 338694 626744
rect 338277 626691 338296 626725
rect 338330 626724 338694 626725
rect 338330 626691 338444 626724
rect 338277 626690 338444 626691
rect 338478 626690 338545 626724
rect 338579 626710 338694 626724
rect 338728 626710 338747 626744
rect 338579 626690 338747 626710
rect 338277 626687 338747 626690
rect 339565 626744 340035 626780
rect 340097 627382 340791 627443
rect 340097 627348 340156 627382
rect 340190 627370 340246 627382
rect 340218 627348 340246 627370
rect 340280 627370 340336 627382
rect 340280 627348 340284 627370
rect 340097 627336 340184 627348
rect 340218 627336 340284 627348
rect 340318 627348 340336 627370
rect 340370 627370 340426 627382
rect 340370 627348 340384 627370
rect 340318 627336 340384 627348
rect 340418 627348 340426 627370
rect 340460 627370 340516 627382
rect 340550 627370 340606 627382
rect 340640 627370 340696 627382
rect 340460 627348 340484 627370
rect 340550 627348 340584 627370
rect 340640 627348 340684 627370
rect 340730 627348 340791 627382
rect 340418 627336 340484 627348
rect 340518 627336 340584 627348
rect 340618 627336 340684 627348
rect 340718 627336 340791 627348
rect 340097 627292 340791 627336
rect 340097 627258 340156 627292
rect 340190 627270 340246 627292
rect 340218 627258 340246 627270
rect 340280 627270 340336 627292
rect 340280 627258 340284 627270
rect 340097 627236 340184 627258
rect 340218 627236 340284 627258
rect 340318 627258 340336 627270
rect 340370 627270 340426 627292
rect 340370 627258 340384 627270
rect 340318 627236 340384 627258
rect 340418 627258 340426 627270
rect 340460 627270 340516 627292
rect 340550 627270 340606 627292
rect 340640 627270 340696 627292
rect 340460 627258 340484 627270
rect 340550 627258 340584 627270
rect 340640 627258 340684 627270
rect 340730 627258 340791 627292
rect 340418 627236 340484 627258
rect 340518 627236 340584 627258
rect 340618 627236 340684 627258
rect 340718 627236 340791 627258
rect 340097 627202 340791 627236
rect 340097 627168 340156 627202
rect 340190 627170 340246 627202
rect 340218 627168 340246 627170
rect 340280 627170 340336 627202
rect 340280 627168 340284 627170
rect 340097 627136 340184 627168
rect 340218 627136 340284 627168
rect 340318 627168 340336 627170
rect 340370 627170 340426 627202
rect 340370 627168 340384 627170
rect 340318 627136 340384 627168
rect 340418 627168 340426 627170
rect 340460 627170 340516 627202
rect 340550 627170 340606 627202
rect 340640 627170 340696 627202
rect 340460 627168 340484 627170
rect 340550 627168 340584 627170
rect 340640 627168 340684 627170
rect 340730 627168 340791 627202
rect 340418 627136 340484 627168
rect 340518 627136 340584 627168
rect 340618 627136 340684 627168
rect 340718 627136 340791 627168
rect 340097 627112 340791 627136
rect 340097 627078 340156 627112
rect 340190 627078 340246 627112
rect 340280 627078 340336 627112
rect 340370 627078 340426 627112
rect 340460 627078 340516 627112
rect 340550 627078 340606 627112
rect 340640 627078 340696 627112
rect 340730 627078 340791 627112
rect 340097 627070 340791 627078
rect 340097 627036 340184 627070
rect 340218 627036 340284 627070
rect 340318 627036 340384 627070
rect 340418 627036 340484 627070
rect 340518 627036 340584 627070
rect 340618 627036 340684 627070
rect 340718 627036 340791 627070
rect 340097 627022 340791 627036
rect 340097 626988 340156 627022
rect 340190 626988 340246 627022
rect 340280 626988 340336 627022
rect 340370 626988 340426 627022
rect 340460 626988 340516 627022
rect 340550 626988 340606 627022
rect 340640 626988 340696 627022
rect 340730 626988 340791 627022
rect 340097 626970 340791 626988
rect 340097 626936 340184 626970
rect 340218 626936 340284 626970
rect 340318 626936 340384 626970
rect 340418 626936 340484 626970
rect 340518 626936 340584 626970
rect 340618 626936 340684 626970
rect 340718 626936 340791 626970
rect 340097 626932 340791 626936
rect 340097 626898 340156 626932
rect 340190 626898 340246 626932
rect 340280 626898 340336 626932
rect 340370 626898 340426 626932
rect 340460 626898 340516 626932
rect 340550 626898 340606 626932
rect 340640 626898 340696 626932
rect 340730 626898 340791 626932
rect 340097 626870 340791 626898
rect 340097 626842 340184 626870
rect 340218 626842 340284 626870
rect 340097 626808 340156 626842
rect 340218 626836 340246 626842
rect 340190 626808 340246 626836
rect 340280 626836 340284 626842
rect 340318 626842 340384 626870
rect 340318 626836 340336 626842
rect 340280 626808 340336 626836
rect 340370 626836 340384 626842
rect 340418 626842 340484 626870
rect 340518 626842 340584 626870
rect 340618 626842 340684 626870
rect 340718 626842 340791 626870
rect 340418 626836 340426 626842
rect 340370 626808 340426 626836
rect 340460 626836 340484 626842
rect 340550 626836 340584 626842
rect 340640 626836 340684 626842
rect 340460 626808 340516 626836
rect 340550 626808 340606 626836
rect 340640 626808 340696 626836
rect 340730 626808 340791 626842
rect 340097 626749 340791 626808
rect 340853 627411 340872 627445
rect 340906 627444 341088 627445
rect 340906 627411 341020 627444
rect 340853 627410 341020 627411
rect 341054 627410 341088 627444
rect 340853 627355 341088 627410
rect 340853 627321 340872 627355
rect 340906 627354 341088 627355
rect 340906 627321 341020 627354
rect 340853 627320 341020 627321
rect 341054 627320 341088 627354
rect 340853 627265 341088 627320
rect 340853 627231 340872 627265
rect 340906 627264 341088 627265
rect 340906 627231 341020 627264
rect 340853 627230 341020 627231
rect 341054 627230 341088 627264
rect 340853 627175 341088 627230
rect 340853 627141 340872 627175
rect 340906 627174 341088 627175
rect 340906 627141 341020 627174
rect 340853 627140 341020 627141
rect 341054 627140 341088 627174
rect 340853 627085 341088 627140
rect 340853 627051 340872 627085
rect 340906 627084 341088 627085
rect 340906 627051 341020 627084
rect 340853 627050 341020 627051
rect 341054 627050 341088 627084
rect 340853 626995 341088 627050
rect 340853 626961 340872 626995
rect 340906 626994 341088 626995
rect 340906 626961 341020 626994
rect 340853 626960 341020 626961
rect 341054 626960 341088 626994
rect 340853 626905 341088 626960
rect 340853 626871 340872 626905
rect 340906 626904 341088 626905
rect 340906 626871 341020 626904
rect 340853 626870 341020 626871
rect 341054 626870 341088 626904
rect 340853 626815 341088 626870
rect 340853 626781 340872 626815
rect 340906 626814 341088 626815
rect 340906 626781 341020 626814
rect 340853 626780 341020 626781
rect 341054 626780 341088 626814
rect 339565 626725 339982 626744
rect 339565 626691 339584 626725
rect 339618 626724 339982 626725
rect 339618 626691 339732 626724
rect 339565 626690 339732 626691
rect 339766 626690 339833 626724
rect 339867 626710 339982 626724
rect 340016 626710 340035 626744
rect 339867 626690 340035 626710
rect 339565 626687 340035 626690
rect 340853 626725 341088 626780
rect 340853 626691 340872 626725
rect 340906 626724 341088 626725
rect 340906 626691 341020 626724
rect 340853 626690 341020 626691
rect 341054 626690 341088 626724
rect 340853 626687 341088 626690
rect 334648 626668 341088 626687
rect 334648 626634 334888 626668
rect 334922 626634 334978 626668
rect 335012 626634 335068 626668
rect 335102 626634 335158 626668
rect 335192 626634 335248 626668
rect 335282 626634 335338 626668
rect 335372 626634 335428 626668
rect 335462 626634 335518 626668
rect 335552 626634 335608 626668
rect 335642 626634 336176 626668
rect 336210 626634 336266 626668
rect 336300 626634 336356 626668
rect 336390 626634 336446 626668
rect 336480 626634 336536 626668
rect 336570 626634 336626 626668
rect 336660 626634 336716 626668
rect 336750 626634 336806 626668
rect 336840 626634 336896 626668
rect 336930 626634 337464 626668
rect 337498 626634 337554 626668
rect 337588 626634 337644 626668
rect 337678 626634 337734 626668
rect 337768 626634 337824 626668
rect 337858 626634 337914 626668
rect 337948 626634 338004 626668
rect 338038 626634 338094 626668
rect 338128 626634 338184 626668
rect 338218 626634 338752 626668
rect 338786 626634 338842 626668
rect 338876 626634 338932 626668
rect 338966 626634 339022 626668
rect 339056 626634 339112 626668
rect 339146 626634 339202 626668
rect 339236 626634 339292 626668
rect 339326 626634 339382 626668
rect 339416 626634 339472 626668
rect 339506 626634 340040 626668
rect 340074 626634 340130 626668
rect 340164 626634 340220 626668
rect 340254 626634 340310 626668
rect 340344 626634 340400 626668
rect 340434 626634 340490 626668
rect 340524 626634 340580 626668
rect 340614 626634 340670 626668
rect 340704 626634 340760 626668
rect 340794 626634 341088 626668
rect 334648 626600 334681 626634
rect 334715 626615 335868 626634
rect 334715 626600 334888 626615
rect 334648 626551 334888 626600
rect 335688 626600 335868 626615
rect 335902 626600 335969 626634
rect 336003 626615 337156 626634
rect 336003 626600 336188 626615
rect 335688 626551 336188 626600
rect 336988 626600 337156 626615
rect 337190 626600 337257 626634
rect 337291 626615 338444 626634
rect 337291 626600 337388 626615
rect 336988 626551 337388 626600
rect 338288 626600 338444 626615
rect 338478 626600 338545 626634
rect 338579 626615 339732 626634
rect 338579 626600 338688 626615
rect 338288 626551 338688 626600
rect 339588 626600 339732 626615
rect 339766 626600 339833 626634
rect 339867 626615 341020 626634
rect 339867 626600 339988 626615
rect 339588 626551 339988 626600
rect 340888 626600 341020 626615
rect 341054 626600 341088 626634
rect 340888 626551 341088 626600
rect 334648 626544 341088 626551
rect 334648 626510 334681 626544
rect 334715 626521 335868 626544
rect 334715 626510 334782 626521
rect 334648 626487 334782 626510
rect 334816 626487 334872 626521
rect 334906 626487 334962 626521
rect 334996 626487 335052 626521
rect 335086 626487 335142 626521
rect 335176 626487 335232 626521
rect 335266 626487 335322 626521
rect 335356 626487 335412 626521
rect 335446 626487 335502 626521
rect 335536 626487 335592 626521
rect 335626 626487 335682 626521
rect 335716 626487 335772 626521
rect 335806 626510 335868 626521
rect 335902 626510 335969 626544
rect 336003 626521 337156 626544
rect 336003 626510 336070 626521
rect 335806 626487 336070 626510
rect 336104 626487 336160 626521
rect 336194 626487 336250 626521
rect 336284 626487 336340 626521
rect 336374 626487 336430 626521
rect 336464 626487 336520 626521
rect 336554 626487 336610 626521
rect 336644 626487 336700 626521
rect 336734 626487 336790 626521
rect 336824 626487 336880 626521
rect 336914 626487 336970 626521
rect 337004 626487 337060 626521
rect 337094 626510 337156 626521
rect 337190 626510 337257 626544
rect 337291 626521 338444 626544
rect 337291 626510 337358 626521
rect 337094 626487 337358 626510
rect 337392 626487 337448 626521
rect 337482 626487 337538 626521
rect 337572 626487 337628 626521
rect 337662 626487 337718 626521
rect 337752 626487 337808 626521
rect 337842 626487 337898 626521
rect 337932 626487 337988 626521
rect 338022 626487 338078 626521
rect 338112 626487 338168 626521
rect 338202 626487 338258 626521
rect 338292 626487 338348 626521
rect 338382 626510 338444 626521
rect 338478 626510 338545 626544
rect 338579 626521 339732 626544
rect 338579 626510 338646 626521
rect 338382 626487 338646 626510
rect 338680 626487 338736 626521
rect 338770 626487 338826 626521
rect 338860 626487 338916 626521
rect 338950 626487 339006 626521
rect 339040 626487 339096 626521
rect 339130 626487 339186 626521
rect 339220 626487 339276 626521
rect 339310 626487 339366 626521
rect 339400 626487 339456 626521
rect 339490 626487 339546 626521
rect 339580 626487 339636 626521
rect 339670 626510 339732 626521
rect 339766 626510 339833 626544
rect 339867 626521 341020 626544
rect 339867 626510 339934 626521
rect 339670 626487 339934 626510
rect 339968 626487 340024 626521
rect 340058 626487 340114 626521
rect 340148 626487 340204 626521
rect 340238 626487 340294 626521
rect 340328 626487 340384 626521
rect 340418 626487 340474 626521
rect 340508 626487 340564 626521
rect 340598 626487 340654 626521
rect 340688 626487 340744 626521
rect 340778 626487 340834 626521
rect 340868 626487 340924 626521
rect 340958 626510 341020 626521
rect 341054 626510 341088 626544
rect 340958 626487 341088 626510
rect 334648 626420 341088 626487
rect 334648 626386 334782 626420
rect 334816 626386 334872 626420
rect 334906 626386 334962 626420
rect 334996 626386 335052 626420
rect 335086 626386 335142 626420
rect 335176 626386 335232 626420
rect 335266 626386 335322 626420
rect 335356 626386 335412 626420
rect 335446 626386 335502 626420
rect 335536 626386 335592 626420
rect 335626 626386 335682 626420
rect 335716 626386 335772 626420
rect 335806 626386 336070 626420
rect 336104 626386 336160 626420
rect 336194 626386 336250 626420
rect 336284 626386 336340 626420
rect 336374 626386 336430 626420
rect 336464 626386 336520 626420
rect 336554 626386 336610 626420
rect 336644 626386 336700 626420
rect 336734 626386 336790 626420
rect 336824 626386 336880 626420
rect 336914 626386 336970 626420
rect 337004 626386 337060 626420
rect 337094 626386 337358 626420
rect 337392 626386 337448 626420
rect 337482 626386 337538 626420
rect 337572 626386 337628 626420
rect 337662 626386 337718 626420
rect 337752 626386 337808 626420
rect 337842 626386 337898 626420
rect 337932 626386 337988 626420
rect 338022 626386 338078 626420
rect 338112 626386 338168 626420
rect 338202 626386 338258 626420
rect 338292 626386 338348 626420
rect 338382 626386 338646 626420
rect 338680 626386 338736 626420
rect 338770 626386 338826 626420
rect 338860 626386 338916 626420
rect 338950 626386 339006 626420
rect 339040 626386 339096 626420
rect 339130 626386 339186 626420
rect 339220 626386 339276 626420
rect 339310 626386 339366 626420
rect 339400 626386 339456 626420
rect 339490 626386 339546 626420
rect 339580 626386 339636 626420
rect 339670 626386 339934 626420
rect 339968 626386 340024 626420
rect 340058 626386 340114 626420
rect 340148 626386 340204 626420
rect 340238 626386 340294 626420
rect 340328 626386 340384 626420
rect 340418 626386 340474 626420
rect 340508 626386 340564 626420
rect 340598 626386 340654 626420
rect 340688 626386 340744 626420
rect 340778 626386 340834 626420
rect 340868 626386 340924 626420
rect 340958 626386 341088 626420
rect 334648 626353 341088 626386
rect 334648 626336 334888 626353
rect 334648 626302 334681 626336
rect 334715 626302 334888 626336
rect 334648 626289 334888 626302
rect 335688 626336 336188 626353
rect 335688 626302 335868 626336
rect 335902 626302 335969 626336
rect 336003 626302 336188 626336
rect 335688 626289 336188 626302
rect 336988 626336 337388 626353
rect 336988 626302 337156 626336
rect 337190 626302 337257 626336
rect 337291 626302 337388 626336
rect 336988 626289 337388 626302
rect 338288 626336 338688 626353
rect 338288 626302 338444 626336
rect 338478 626302 338545 626336
rect 338579 626302 338688 626336
rect 338288 626289 338688 626302
rect 339588 626336 339988 626353
rect 339588 626302 339732 626336
rect 339766 626302 339833 626336
rect 339867 626302 339988 626336
rect 339588 626289 339988 626302
rect 340888 626336 341088 626353
rect 340888 626302 341020 626336
rect 341054 626302 341088 626336
rect 340888 626289 341088 626302
rect 334648 626270 341088 626289
rect 334648 626246 334922 626270
rect 334648 626212 334681 626246
rect 334715 626236 334922 626246
rect 334956 626236 335012 626270
rect 335046 626236 335102 626270
rect 335136 626236 335192 626270
rect 335226 626236 335282 626270
rect 335316 626236 335372 626270
rect 335406 626236 335462 626270
rect 335496 626236 335552 626270
rect 335586 626236 335642 626270
rect 335676 626246 336210 626270
rect 335676 626236 335868 626246
rect 334715 626217 335868 626236
rect 334715 626212 334888 626217
rect 334648 626176 334888 626212
rect 334648 626156 334830 626176
rect 334648 626122 334681 626156
rect 334715 626142 334830 626156
rect 334864 626142 334888 626176
rect 335688 626212 335868 626217
rect 335902 626212 335969 626246
rect 336003 626236 336210 626246
rect 336244 626236 336300 626270
rect 336334 626236 336390 626270
rect 336424 626236 336480 626270
rect 336514 626236 336570 626270
rect 336604 626236 336660 626270
rect 336694 626236 336750 626270
rect 336784 626236 336840 626270
rect 336874 626236 336930 626270
rect 336964 626246 337498 626270
rect 336964 626236 337156 626246
rect 336003 626217 337156 626236
rect 336003 626212 336188 626217
rect 335688 626176 336188 626212
rect 335688 626157 336118 626176
rect 334715 626122 334888 626142
rect 334648 626086 334888 626122
rect 334648 626066 334830 626086
rect 334648 626032 334681 626066
rect 334715 626052 334830 626066
rect 334864 626052 334888 626086
rect 334715 626032 334888 626052
rect 334648 625996 334888 626032
rect 334648 625976 334830 625996
rect 334648 625942 334681 625976
rect 334715 625962 334830 625976
rect 334864 625962 334888 625996
rect 334715 625942 334888 625962
rect 334648 625906 334888 625942
rect 334648 625886 334830 625906
rect 334648 625852 334681 625886
rect 334715 625872 334830 625886
rect 334864 625872 334888 625906
rect 334715 625852 334888 625872
rect 334648 625816 334888 625852
rect 334648 625796 334830 625816
rect 334648 625762 334681 625796
rect 334715 625782 334830 625796
rect 334864 625782 334888 625816
rect 334715 625762 334888 625782
rect 334648 625726 334888 625762
rect 334648 625706 334830 625726
rect 334648 625672 334681 625706
rect 334715 625692 334830 625706
rect 334864 625692 334888 625726
rect 334715 625672 334888 625692
rect 334648 625636 334888 625672
rect 334648 625616 334830 625636
rect 334648 625582 334681 625616
rect 334715 625602 334830 625616
rect 334864 625602 334888 625636
rect 334715 625582 334888 625602
rect 334648 625546 334888 625582
rect 334648 625526 334830 625546
rect 334648 625492 334681 625526
rect 334715 625512 334830 625526
rect 334864 625512 334888 625546
rect 334715 625492 334888 625512
rect 334648 625456 334888 625492
rect 334945 626094 335639 626155
rect 334945 626060 335004 626094
rect 335038 626082 335094 626094
rect 335066 626060 335094 626082
rect 335128 626082 335184 626094
rect 335128 626060 335132 626082
rect 334945 626048 335032 626060
rect 335066 626048 335132 626060
rect 335166 626060 335184 626082
rect 335218 626082 335274 626094
rect 335218 626060 335232 626082
rect 335166 626048 335232 626060
rect 335266 626060 335274 626082
rect 335308 626082 335364 626094
rect 335398 626082 335454 626094
rect 335488 626082 335544 626094
rect 335308 626060 335332 626082
rect 335398 626060 335432 626082
rect 335488 626060 335532 626082
rect 335578 626060 335639 626094
rect 335266 626048 335332 626060
rect 335366 626048 335432 626060
rect 335466 626048 335532 626060
rect 335566 626048 335639 626060
rect 334945 626004 335639 626048
rect 334945 625970 335004 626004
rect 335038 625982 335094 626004
rect 335066 625970 335094 625982
rect 335128 625982 335184 626004
rect 335128 625970 335132 625982
rect 334945 625948 335032 625970
rect 335066 625948 335132 625970
rect 335166 625970 335184 625982
rect 335218 625982 335274 626004
rect 335218 625970 335232 625982
rect 335166 625948 335232 625970
rect 335266 625970 335274 625982
rect 335308 625982 335364 626004
rect 335398 625982 335454 626004
rect 335488 625982 335544 626004
rect 335308 625970 335332 625982
rect 335398 625970 335432 625982
rect 335488 625970 335532 625982
rect 335578 625970 335639 626004
rect 335266 625948 335332 625970
rect 335366 625948 335432 625970
rect 335466 625948 335532 625970
rect 335566 625948 335639 625970
rect 334945 625914 335639 625948
rect 334945 625880 335004 625914
rect 335038 625882 335094 625914
rect 335066 625880 335094 625882
rect 335128 625882 335184 625914
rect 335128 625880 335132 625882
rect 334945 625848 335032 625880
rect 335066 625848 335132 625880
rect 335166 625880 335184 625882
rect 335218 625882 335274 625914
rect 335218 625880 335232 625882
rect 335166 625848 335232 625880
rect 335266 625880 335274 625882
rect 335308 625882 335364 625914
rect 335398 625882 335454 625914
rect 335488 625882 335544 625914
rect 335308 625880 335332 625882
rect 335398 625880 335432 625882
rect 335488 625880 335532 625882
rect 335578 625880 335639 625914
rect 335266 625848 335332 625880
rect 335366 625848 335432 625880
rect 335466 625848 335532 625880
rect 335566 625848 335639 625880
rect 334945 625824 335639 625848
rect 334945 625790 335004 625824
rect 335038 625790 335094 625824
rect 335128 625790 335184 625824
rect 335218 625790 335274 625824
rect 335308 625790 335364 625824
rect 335398 625790 335454 625824
rect 335488 625790 335544 625824
rect 335578 625790 335639 625824
rect 334945 625782 335639 625790
rect 334945 625748 335032 625782
rect 335066 625748 335132 625782
rect 335166 625748 335232 625782
rect 335266 625748 335332 625782
rect 335366 625748 335432 625782
rect 335466 625748 335532 625782
rect 335566 625748 335639 625782
rect 334945 625734 335639 625748
rect 334945 625700 335004 625734
rect 335038 625700 335094 625734
rect 335128 625700 335184 625734
rect 335218 625700 335274 625734
rect 335308 625700 335364 625734
rect 335398 625700 335454 625734
rect 335488 625700 335544 625734
rect 335578 625700 335639 625734
rect 334945 625682 335639 625700
rect 334945 625648 335032 625682
rect 335066 625648 335132 625682
rect 335166 625648 335232 625682
rect 335266 625648 335332 625682
rect 335366 625648 335432 625682
rect 335466 625648 335532 625682
rect 335566 625648 335639 625682
rect 334945 625644 335639 625648
rect 334945 625610 335004 625644
rect 335038 625610 335094 625644
rect 335128 625610 335184 625644
rect 335218 625610 335274 625644
rect 335308 625610 335364 625644
rect 335398 625610 335454 625644
rect 335488 625610 335544 625644
rect 335578 625610 335639 625644
rect 334945 625582 335639 625610
rect 334945 625554 335032 625582
rect 335066 625554 335132 625582
rect 334945 625520 335004 625554
rect 335066 625548 335094 625554
rect 335038 625520 335094 625548
rect 335128 625548 335132 625554
rect 335166 625554 335232 625582
rect 335166 625548 335184 625554
rect 335128 625520 335184 625548
rect 335218 625548 335232 625554
rect 335266 625554 335332 625582
rect 335366 625554 335432 625582
rect 335466 625554 335532 625582
rect 335566 625554 335639 625582
rect 335266 625548 335274 625554
rect 335218 625520 335274 625548
rect 335308 625548 335332 625554
rect 335398 625548 335432 625554
rect 335488 625548 335532 625554
rect 335308 625520 335364 625548
rect 335398 625520 335454 625548
rect 335488 625520 335544 625548
rect 335578 625520 335639 625554
rect 334945 625461 335639 625520
rect 335688 626123 335720 626157
rect 335754 626156 336118 626157
rect 335754 626123 335868 626156
rect 335688 626122 335868 626123
rect 335902 626122 335969 626156
rect 336003 626142 336118 626156
rect 336152 626142 336188 626176
rect 336988 626212 337156 626217
rect 337190 626212 337257 626246
rect 337291 626236 337498 626246
rect 337532 626236 337588 626270
rect 337622 626236 337678 626270
rect 337712 626236 337768 626270
rect 337802 626236 337858 626270
rect 337892 626236 337948 626270
rect 337982 626236 338038 626270
rect 338072 626236 338128 626270
rect 338162 626236 338218 626270
rect 338252 626246 338786 626270
rect 338252 626236 338444 626246
rect 337291 626217 338444 626236
rect 337291 626212 337459 626217
rect 336988 626176 337459 626212
rect 336988 626157 337406 626176
rect 336003 626122 336188 626142
rect 335688 626086 336188 626122
rect 335688 626067 336118 626086
rect 335688 626033 335720 626067
rect 335754 626066 336118 626067
rect 335754 626033 335868 626066
rect 335688 626032 335868 626033
rect 335902 626032 335969 626066
rect 336003 626052 336118 626066
rect 336152 626052 336188 626086
rect 336003 626032 336188 626052
rect 335688 625996 336188 626032
rect 335688 625977 336118 625996
rect 335688 625943 335720 625977
rect 335754 625976 336118 625977
rect 335754 625943 335868 625976
rect 335688 625942 335868 625943
rect 335902 625942 335969 625976
rect 336003 625962 336118 625976
rect 336152 625962 336188 625996
rect 336003 625942 336188 625962
rect 335688 625906 336188 625942
rect 335688 625887 336118 625906
rect 335688 625853 335720 625887
rect 335754 625886 336118 625887
rect 335754 625853 335868 625886
rect 335688 625852 335868 625853
rect 335902 625852 335969 625886
rect 336003 625872 336118 625886
rect 336152 625872 336188 625906
rect 336003 625852 336188 625872
rect 335688 625816 336188 625852
rect 335688 625797 336118 625816
rect 335688 625763 335720 625797
rect 335754 625796 336118 625797
rect 335754 625763 335868 625796
rect 335688 625762 335868 625763
rect 335902 625762 335969 625796
rect 336003 625782 336118 625796
rect 336152 625782 336188 625816
rect 336003 625762 336188 625782
rect 335688 625726 336188 625762
rect 335688 625707 336118 625726
rect 335688 625673 335720 625707
rect 335754 625706 336118 625707
rect 335754 625673 335868 625706
rect 335688 625672 335868 625673
rect 335902 625672 335969 625706
rect 336003 625692 336118 625706
rect 336152 625692 336188 625726
rect 336003 625672 336188 625692
rect 335688 625636 336188 625672
rect 335688 625617 336118 625636
rect 335688 625583 335720 625617
rect 335754 625616 336118 625617
rect 335754 625583 335868 625616
rect 335688 625582 335868 625583
rect 335902 625582 335969 625616
rect 336003 625602 336118 625616
rect 336152 625602 336188 625636
rect 336003 625582 336188 625602
rect 335688 625546 336188 625582
rect 335688 625527 336118 625546
rect 335688 625493 335720 625527
rect 335754 625526 336118 625527
rect 335754 625493 335868 625526
rect 335688 625492 335868 625493
rect 335902 625492 335969 625526
rect 336003 625512 336118 625526
rect 336152 625512 336188 625546
rect 336003 625492 336188 625512
rect 334648 625436 334830 625456
rect 334648 625402 334681 625436
rect 334715 625422 334830 625436
rect 334864 625422 334888 625456
rect 334715 625402 334888 625422
rect 334648 625399 334888 625402
rect 335688 625456 336188 625492
rect 336233 626094 336927 626155
rect 336233 626060 336292 626094
rect 336326 626082 336382 626094
rect 336354 626060 336382 626082
rect 336416 626082 336472 626094
rect 336416 626060 336420 626082
rect 336233 626048 336320 626060
rect 336354 626048 336420 626060
rect 336454 626060 336472 626082
rect 336506 626082 336562 626094
rect 336506 626060 336520 626082
rect 336454 626048 336520 626060
rect 336554 626060 336562 626082
rect 336596 626082 336652 626094
rect 336686 626082 336742 626094
rect 336776 626082 336832 626094
rect 336596 626060 336620 626082
rect 336686 626060 336720 626082
rect 336776 626060 336820 626082
rect 336866 626060 336927 626094
rect 336554 626048 336620 626060
rect 336654 626048 336720 626060
rect 336754 626048 336820 626060
rect 336854 626048 336927 626060
rect 336233 626004 336927 626048
rect 336233 625970 336292 626004
rect 336326 625982 336382 626004
rect 336354 625970 336382 625982
rect 336416 625982 336472 626004
rect 336416 625970 336420 625982
rect 336233 625948 336320 625970
rect 336354 625948 336420 625970
rect 336454 625970 336472 625982
rect 336506 625982 336562 626004
rect 336506 625970 336520 625982
rect 336454 625948 336520 625970
rect 336554 625970 336562 625982
rect 336596 625982 336652 626004
rect 336686 625982 336742 626004
rect 336776 625982 336832 626004
rect 336596 625970 336620 625982
rect 336686 625970 336720 625982
rect 336776 625970 336820 625982
rect 336866 625970 336927 626004
rect 336554 625948 336620 625970
rect 336654 625948 336720 625970
rect 336754 625948 336820 625970
rect 336854 625948 336927 625970
rect 336233 625914 336927 625948
rect 336233 625880 336292 625914
rect 336326 625882 336382 625914
rect 336354 625880 336382 625882
rect 336416 625882 336472 625914
rect 336416 625880 336420 625882
rect 336233 625848 336320 625880
rect 336354 625848 336420 625880
rect 336454 625880 336472 625882
rect 336506 625882 336562 625914
rect 336506 625880 336520 625882
rect 336454 625848 336520 625880
rect 336554 625880 336562 625882
rect 336596 625882 336652 625914
rect 336686 625882 336742 625914
rect 336776 625882 336832 625914
rect 336596 625880 336620 625882
rect 336686 625880 336720 625882
rect 336776 625880 336820 625882
rect 336866 625880 336927 625914
rect 336554 625848 336620 625880
rect 336654 625848 336720 625880
rect 336754 625848 336820 625880
rect 336854 625848 336927 625880
rect 336233 625824 336927 625848
rect 336233 625790 336292 625824
rect 336326 625790 336382 625824
rect 336416 625790 336472 625824
rect 336506 625790 336562 625824
rect 336596 625790 336652 625824
rect 336686 625790 336742 625824
rect 336776 625790 336832 625824
rect 336866 625790 336927 625824
rect 336233 625782 336927 625790
rect 336233 625748 336320 625782
rect 336354 625748 336420 625782
rect 336454 625748 336520 625782
rect 336554 625748 336620 625782
rect 336654 625748 336720 625782
rect 336754 625748 336820 625782
rect 336854 625748 336927 625782
rect 336233 625734 336927 625748
rect 336233 625700 336292 625734
rect 336326 625700 336382 625734
rect 336416 625700 336472 625734
rect 336506 625700 336562 625734
rect 336596 625700 336652 625734
rect 336686 625700 336742 625734
rect 336776 625700 336832 625734
rect 336866 625700 336927 625734
rect 336233 625682 336927 625700
rect 336233 625648 336320 625682
rect 336354 625648 336420 625682
rect 336454 625648 336520 625682
rect 336554 625648 336620 625682
rect 336654 625648 336720 625682
rect 336754 625648 336820 625682
rect 336854 625648 336927 625682
rect 336233 625644 336927 625648
rect 336233 625610 336292 625644
rect 336326 625610 336382 625644
rect 336416 625610 336472 625644
rect 336506 625610 336562 625644
rect 336596 625610 336652 625644
rect 336686 625610 336742 625644
rect 336776 625610 336832 625644
rect 336866 625610 336927 625644
rect 336233 625582 336927 625610
rect 336233 625554 336320 625582
rect 336354 625554 336420 625582
rect 336233 625520 336292 625554
rect 336354 625548 336382 625554
rect 336326 625520 336382 625548
rect 336416 625548 336420 625554
rect 336454 625554 336520 625582
rect 336454 625548 336472 625554
rect 336416 625520 336472 625548
rect 336506 625548 336520 625554
rect 336554 625554 336620 625582
rect 336654 625554 336720 625582
rect 336754 625554 336820 625582
rect 336854 625554 336927 625582
rect 336554 625548 336562 625554
rect 336506 625520 336562 625548
rect 336596 625548 336620 625554
rect 336686 625548 336720 625554
rect 336776 625548 336820 625554
rect 336596 625520 336652 625548
rect 336686 625520 336742 625548
rect 336776 625520 336832 625548
rect 336866 625520 336927 625554
rect 336233 625461 336927 625520
rect 336988 626123 337008 626157
rect 337042 626156 337406 626157
rect 337042 626123 337156 626156
rect 336988 626122 337156 626123
rect 337190 626122 337257 626156
rect 337291 626142 337406 626156
rect 337440 626142 337459 626176
rect 338277 626212 338444 626217
rect 338478 626212 338545 626246
rect 338579 626236 338786 626246
rect 338820 626236 338876 626270
rect 338910 626236 338966 626270
rect 339000 626236 339056 626270
rect 339090 626236 339146 626270
rect 339180 626236 339236 626270
rect 339270 626236 339326 626270
rect 339360 626236 339416 626270
rect 339450 626236 339506 626270
rect 339540 626246 340074 626270
rect 339540 626236 339732 626246
rect 338579 626217 339732 626236
rect 338579 626212 338747 626217
rect 338277 626176 338747 626212
rect 338277 626157 338694 626176
rect 337291 626122 337459 626142
rect 336988 626086 337459 626122
rect 336988 626067 337406 626086
rect 336988 626033 337008 626067
rect 337042 626066 337406 626067
rect 337042 626033 337156 626066
rect 336988 626032 337156 626033
rect 337190 626032 337257 626066
rect 337291 626052 337406 626066
rect 337440 626052 337459 626086
rect 337291 626032 337459 626052
rect 336988 625996 337459 626032
rect 336988 625977 337406 625996
rect 336988 625943 337008 625977
rect 337042 625976 337406 625977
rect 337042 625943 337156 625976
rect 336988 625942 337156 625943
rect 337190 625942 337257 625976
rect 337291 625962 337406 625976
rect 337440 625962 337459 625996
rect 337291 625942 337459 625962
rect 336988 625906 337459 625942
rect 336988 625887 337406 625906
rect 336988 625853 337008 625887
rect 337042 625886 337406 625887
rect 337042 625853 337156 625886
rect 336988 625852 337156 625853
rect 337190 625852 337257 625886
rect 337291 625872 337406 625886
rect 337440 625872 337459 625906
rect 337291 625852 337459 625872
rect 336988 625816 337459 625852
rect 336988 625797 337406 625816
rect 336988 625763 337008 625797
rect 337042 625796 337406 625797
rect 337042 625763 337156 625796
rect 336988 625762 337156 625763
rect 337190 625762 337257 625796
rect 337291 625782 337406 625796
rect 337440 625782 337459 625816
rect 337291 625762 337459 625782
rect 336988 625726 337459 625762
rect 336988 625707 337406 625726
rect 336988 625673 337008 625707
rect 337042 625706 337406 625707
rect 337042 625673 337156 625706
rect 336988 625672 337156 625673
rect 337190 625672 337257 625706
rect 337291 625692 337406 625706
rect 337440 625692 337459 625726
rect 337291 625672 337459 625692
rect 336988 625636 337459 625672
rect 336988 625617 337406 625636
rect 336988 625583 337008 625617
rect 337042 625616 337406 625617
rect 337042 625583 337156 625616
rect 336988 625582 337156 625583
rect 337190 625582 337257 625616
rect 337291 625602 337406 625616
rect 337440 625602 337459 625636
rect 337291 625582 337459 625602
rect 336988 625546 337459 625582
rect 336988 625527 337406 625546
rect 336988 625493 337008 625527
rect 337042 625526 337406 625527
rect 337042 625493 337156 625526
rect 336988 625492 337156 625493
rect 337190 625492 337257 625526
rect 337291 625512 337406 625526
rect 337440 625512 337459 625546
rect 337291 625492 337459 625512
rect 335688 625437 336118 625456
rect 335688 625403 335720 625437
rect 335754 625436 336118 625437
rect 335754 625403 335868 625436
rect 335688 625402 335868 625403
rect 335902 625402 335969 625436
rect 336003 625422 336118 625436
rect 336152 625422 336188 625456
rect 336003 625402 336188 625422
rect 335688 625399 336188 625402
rect 336988 625456 337459 625492
rect 337521 626094 338215 626155
rect 337521 626060 337580 626094
rect 337614 626082 337670 626094
rect 337642 626060 337670 626082
rect 337704 626082 337760 626094
rect 337704 626060 337708 626082
rect 337521 626048 337608 626060
rect 337642 626048 337708 626060
rect 337742 626060 337760 626082
rect 337794 626082 337850 626094
rect 337794 626060 337808 626082
rect 337742 626048 337808 626060
rect 337842 626060 337850 626082
rect 337884 626082 337940 626094
rect 337974 626082 338030 626094
rect 338064 626082 338120 626094
rect 337884 626060 337908 626082
rect 337974 626060 338008 626082
rect 338064 626060 338108 626082
rect 338154 626060 338215 626094
rect 337842 626048 337908 626060
rect 337942 626048 338008 626060
rect 338042 626048 338108 626060
rect 338142 626048 338215 626060
rect 337521 626004 338215 626048
rect 337521 625970 337580 626004
rect 337614 625982 337670 626004
rect 337642 625970 337670 625982
rect 337704 625982 337760 626004
rect 337704 625970 337708 625982
rect 337521 625948 337608 625970
rect 337642 625948 337708 625970
rect 337742 625970 337760 625982
rect 337794 625982 337850 626004
rect 337794 625970 337808 625982
rect 337742 625948 337808 625970
rect 337842 625970 337850 625982
rect 337884 625982 337940 626004
rect 337974 625982 338030 626004
rect 338064 625982 338120 626004
rect 337884 625970 337908 625982
rect 337974 625970 338008 625982
rect 338064 625970 338108 625982
rect 338154 625970 338215 626004
rect 337842 625948 337908 625970
rect 337942 625948 338008 625970
rect 338042 625948 338108 625970
rect 338142 625948 338215 625970
rect 337521 625914 338215 625948
rect 337521 625880 337580 625914
rect 337614 625882 337670 625914
rect 337642 625880 337670 625882
rect 337704 625882 337760 625914
rect 337704 625880 337708 625882
rect 337521 625848 337608 625880
rect 337642 625848 337708 625880
rect 337742 625880 337760 625882
rect 337794 625882 337850 625914
rect 337794 625880 337808 625882
rect 337742 625848 337808 625880
rect 337842 625880 337850 625882
rect 337884 625882 337940 625914
rect 337974 625882 338030 625914
rect 338064 625882 338120 625914
rect 337884 625880 337908 625882
rect 337974 625880 338008 625882
rect 338064 625880 338108 625882
rect 338154 625880 338215 625914
rect 337842 625848 337908 625880
rect 337942 625848 338008 625880
rect 338042 625848 338108 625880
rect 338142 625848 338215 625880
rect 337521 625824 338215 625848
rect 337521 625790 337580 625824
rect 337614 625790 337670 625824
rect 337704 625790 337760 625824
rect 337794 625790 337850 625824
rect 337884 625790 337940 625824
rect 337974 625790 338030 625824
rect 338064 625790 338120 625824
rect 338154 625790 338215 625824
rect 337521 625782 338215 625790
rect 337521 625748 337608 625782
rect 337642 625748 337708 625782
rect 337742 625748 337808 625782
rect 337842 625748 337908 625782
rect 337942 625748 338008 625782
rect 338042 625748 338108 625782
rect 338142 625748 338215 625782
rect 337521 625734 338215 625748
rect 337521 625700 337580 625734
rect 337614 625700 337670 625734
rect 337704 625700 337760 625734
rect 337794 625700 337850 625734
rect 337884 625700 337940 625734
rect 337974 625700 338030 625734
rect 338064 625700 338120 625734
rect 338154 625700 338215 625734
rect 337521 625682 338215 625700
rect 337521 625648 337608 625682
rect 337642 625648 337708 625682
rect 337742 625648 337808 625682
rect 337842 625648 337908 625682
rect 337942 625648 338008 625682
rect 338042 625648 338108 625682
rect 338142 625648 338215 625682
rect 337521 625644 338215 625648
rect 337521 625610 337580 625644
rect 337614 625610 337670 625644
rect 337704 625610 337760 625644
rect 337794 625610 337850 625644
rect 337884 625610 337940 625644
rect 337974 625610 338030 625644
rect 338064 625610 338120 625644
rect 338154 625610 338215 625644
rect 337521 625582 338215 625610
rect 337521 625554 337608 625582
rect 337642 625554 337708 625582
rect 337521 625520 337580 625554
rect 337642 625548 337670 625554
rect 337614 625520 337670 625548
rect 337704 625548 337708 625554
rect 337742 625554 337808 625582
rect 337742 625548 337760 625554
rect 337704 625520 337760 625548
rect 337794 625548 337808 625554
rect 337842 625554 337908 625582
rect 337942 625554 338008 625582
rect 338042 625554 338108 625582
rect 338142 625554 338215 625582
rect 337842 625548 337850 625554
rect 337794 625520 337850 625548
rect 337884 625548 337908 625554
rect 337974 625548 338008 625554
rect 338064 625548 338108 625554
rect 337884 625520 337940 625548
rect 337974 625520 338030 625548
rect 338064 625520 338120 625548
rect 338154 625520 338215 625554
rect 337521 625461 338215 625520
rect 338277 626123 338296 626157
rect 338330 626156 338694 626157
rect 338330 626123 338444 626156
rect 338277 626122 338444 626123
rect 338478 626122 338545 626156
rect 338579 626142 338694 626156
rect 338728 626142 338747 626176
rect 339565 626212 339732 626217
rect 339766 626212 339833 626246
rect 339867 626236 340074 626246
rect 340108 626236 340164 626270
rect 340198 626236 340254 626270
rect 340288 626236 340344 626270
rect 340378 626236 340434 626270
rect 340468 626236 340524 626270
rect 340558 626236 340614 626270
rect 340648 626236 340704 626270
rect 340738 626236 340794 626270
rect 340828 626246 341088 626270
rect 340828 626236 341020 626246
rect 339867 626217 341020 626236
rect 339867 626212 340035 626217
rect 339565 626176 340035 626212
rect 339565 626157 339982 626176
rect 338579 626122 338747 626142
rect 338277 626086 338747 626122
rect 338277 626067 338694 626086
rect 338277 626033 338296 626067
rect 338330 626066 338694 626067
rect 338330 626033 338444 626066
rect 338277 626032 338444 626033
rect 338478 626032 338545 626066
rect 338579 626052 338694 626066
rect 338728 626052 338747 626086
rect 338579 626032 338747 626052
rect 338277 625996 338747 626032
rect 338277 625977 338694 625996
rect 338277 625943 338296 625977
rect 338330 625976 338694 625977
rect 338330 625943 338444 625976
rect 338277 625942 338444 625943
rect 338478 625942 338545 625976
rect 338579 625962 338694 625976
rect 338728 625962 338747 625996
rect 338579 625942 338747 625962
rect 338277 625906 338747 625942
rect 338277 625887 338694 625906
rect 338277 625853 338296 625887
rect 338330 625886 338694 625887
rect 338330 625853 338444 625886
rect 338277 625852 338444 625853
rect 338478 625852 338545 625886
rect 338579 625872 338694 625886
rect 338728 625872 338747 625906
rect 338579 625852 338747 625872
rect 338277 625816 338747 625852
rect 338277 625797 338694 625816
rect 338277 625763 338296 625797
rect 338330 625796 338694 625797
rect 338330 625763 338444 625796
rect 338277 625762 338444 625763
rect 338478 625762 338545 625796
rect 338579 625782 338694 625796
rect 338728 625782 338747 625816
rect 338579 625762 338747 625782
rect 338277 625726 338747 625762
rect 338277 625707 338694 625726
rect 338277 625673 338296 625707
rect 338330 625706 338694 625707
rect 338330 625673 338444 625706
rect 338277 625672 338444 625673
rect 338478 625672 338545 625706
rect 338579 625692 338694 625706
rect 338728 625692 338747 625726
rect 338579 625672 338747 625692
rect 338277 625636 338747 625672
rect 338277 625617 338694 625636
rect 338277 625583 338296 625617
rect 338330 625616 338694 625617
rect 338330 625583 338444 625616
rect 338277 625582 338444 625583
rect 338478 625582 338545 625616
rect 338579 625602 338694 625616
rect 338728 625602 338747 625636
rect 338579 625582 338747 625602
rect 338277 625546 338747 625582
rect 338277 625527 338694 625546
rect 338277 625493 338296 625527
rect 338330 625526 338694 625527
rect 338330 625493 338444 625526
rect 338277 625492 338444 625493
rect 338478 625492 338545 625526
rect 338579 625512 338694 625526
rect 338728 625512 338747 625546
rect 338579 625492 338747 625512
rect 336988 625437 337406 625456
rect 336988 625403 337008 625437
rect 337042 625436 337406 625437
rect 337042 625403 337156 625436
rect 336988 625402 337156 625403
rect 337190 625402 337257 625436
rect 337291 625422 337406 625436
rect 337440 625422 337459 625456
rect 337291 625402 337459 625422
rect 336988 625399 337459 625402
rect 338277 625456 338747 625492
rect 338809 626094 339503 626155
rect 338809 626060 338868 626094
rect 338902 626082 338958 626094
rect 338930 626060 338958 626082
rect 338992 626082 339048 626094
rect 338992 626060 338996 626082
rect 338809 626048 338896 626060
rect 338930 626048 338996 626060
rect 339030 626060 339048 626082
rect 339082 626082 339138 626094
rect 339082 626060 339096 626082
rect 339030 626048 339096 626060
rect 339130 626060 339138 626082
rect 339172 626082 339228 626094
rect 339262 626082 339318 626094
rect 339352 626082 339408 626094
rect 339172 626060 339196 626082
rect 339262 626060 339296 626082
rect 339352 626060 339396 626082
rect 339442 626060 339503 626094
rect 339130 626048 339196 626060
rect 339230 626048 339296 626060
rect 339330 626048 339396 626060
rect 339430 626048 339503 626060
rect 338809 626004 339503 626048
rect 338809 625970 338868 626004
rect 338902 625982 338958 626004
rect 338930 625970 338958 625982
rect 338992 625982 339048 626004
rect 338992 625970 338996 625982
rect 338809 625948 338896 625970
rect 338930 625948 338996 625970
rect 339030 625970 339048 625982
rect 339082 625982 339138 626004
rect 339082 625970 339096 625982
rect 339030 625948 339096 625970
rect 339130 625970 339138 625982
rect 339172 625982 339228 626004
rect 339262 625982 339318 626004
rect 339352 625982 339408 626004
rect 339172 625970 339196 625982
rect 339262 625970 339296 625982
rect 339352 625970 339396 625982
rect 339442 625970 339503 626004
rect 339130 625948 339196 625970
rect 339230 625948 339296 625970
rect 339330 625948 339396 625970
rect 339430 625948 339503 625970
rect 338809 625914 339503 625948
rect 338809 625880 338868 625914
rect 338902 625882 338958 625914
rect 338930 625880 338958 625882
rect 338992 625882 339048 625914
rect 338992 625880 338996 625882
rect 338809 625848 338896 625880
rect 338930 625848 338996 625880
rect 339030 625880 339048 625882
rect 339082 625882 339138 625914
rect 339082 625880 339096 625882
rect 339030 625848 339096 625880
rect 339130 625880 339138 625882
rect 339172 625882 339228 625914
rect 339262 625882 339318 625914
rect 339352 625882 339408 625914
rect 339172 625880 339196 625882
rect 339262 625880 339296 625882
rect 339352 625880 339396 625882
rect 339442 625880 339503 625914
rect 339130 625848 339196 625880
rect 339230 625848 339296 625880
rect 339330 625848 339396 625880
rect 339430 625848 339503 625880
rect 338809 625824 339503 625848
rect 338809 625790 338868 625824
rect 338902 625790 338958 625824
rect 338992 625790 339048 625824
rect 339082 625790 339138 625824
rect 339172 625790 339228 625824
rect 339262 625790 339318 625824
rect 339352 625790 339408 625824
rect 339442 625790 339503 625824
rect 338809 625782 339503 625790
rect 338809 625748 338896 625782
rect 338930 625748 338996 625782
rect 339030 625748 339096 625782
rect 339130 625748 339196 625782
rect 339230 625748 339296 625782
rect 339330 625748 339396 625782
rect 339430 625748 339503 625782
rect 338809 625734 339503 625748
rect 338809 625700 338868 625734
rect 338902 625700 338958 625734
rect 338992 625700 339048 625734
rect 339082 625700 339138 625734
rect 339172 625700 339228 625734
rect 339262 625700 339318 625734
rect 339352 625700 339408 625734
rect 339442 625700 339503 625734
rect 338809 625682 339503 625700
rect 338809 625648 338896 625682
rect 338930 625648 338996 625682
rect 339030 625648 339096 625682
rect 339130 625648 339196 625682
rect 339230 625648 339296 625682
rect 339330 625648 339396 625682
rect 339430 625648 339503 625682
rect 338809 625644 339503 625648
rect 338809 625610 338868 625644
rect 338902 625610 338958 625644
rect 338992 625610 339048 625644
rect 339082 625610 339138 625644
rect 339172 625610 339228 625644
rect 339262 625610 339318 625644
rect 339352 625610 339408 625644
rect 339442 625610 339503 625644
rect 338809 625582 339503 625610
rect 338809 625554 338896 625582
rect 338930 625554 338996 625582
rect 338809 625520 338868 625554
rect 338930 625548 338958 625554
rect 338902 625520 338958 625548
rect 338992 625548 338996 625554
rect 339030 625554 339096 625582
rect 339030 625548 339048 625554
rect 338992 625520 339048 625548
rect 339082 625548 339096 625554
rect 339130 625554 339196 625582
rect 339230 625554 339296 625582
rect 339330 625554 339396 625582
rect 339430 625554 339503 625582
rect 339130 625548 339138 625554
rect 339082 625520 339138 625548
rect 339172 625548 339196 625554
rect 339262 625548 339296 625554
rect 339352 625548 339396 625554
rect 339172 625520 339228 625548
rect 339262 625520 339318 625548
rect 339352 625520 339408 625548
rect 339442 625520 339503 625554
rect 338809 625461 339503 625520
rect 339565 626123 339584 626157
rect 339618 626156 339982 626157
rect 339618 626123 339732 626156
rect 339565 626122 339732 626123
rect 339766 626122 339833 626156
rect 339867 626142 339982 626156
rect 340016 626142 340035 626176
rect 340853 626212 341020 626217
rect 341054 626212 341088 626246
rect 340853 626157 341088 626212
rect 339867 626122 340035 626142
rect 339565 626086 340035 626122
rect 339565 626067 339982 626086
rect 339565 626033 339584 626067
rect 339618 626066 339982 626067
rect 339618 626033 339732 626066
rect 339565 626032 339732 626033
rect 339766 626032 339833 626066
rect 339867 626052 339982 626066
rect 340016 626052 340035 626086
rect 339867 626032 340035 626052
rect 339565 625996 340035 626032
rect 339565 625977 339982 625996
rect 339565 625943 339584 625977
rect 339618 625976 339982 625977
rect 339618 625943 339732 625976
rect 339565 625942 339732 625943
rect 339766 625942 339833 625976
rect 339867 625962 339982 625976
rect 340016 625962 340035 625996
rect 339867 625942 340035 625962
rect 339565 625906 340035 625942
rect 339565 625887 339982 625906
rect 339565 625853 339584 625887
rect 339618 625886 339982 625887
rect 339618 625853 339732 625886
rect 339565 625852 339732 625853
rect 339766 625852 339833 625886
rect 339867 625872 339982 625886
rect 340016 625872 340035 625906
rect 339867 625852 340035 625872
rect 339565 625816 340035 625852
rect 339565 625797 339982 625816
rect 339565 625763 339584 625797
rect 339618 625796 339982 625797
rect 339618 625763 339732 625796
rect 339565 625762 339732 625763
rect 339766 625762 339833 625796
rect 339867 625782 339982 625796
rect 340016 625782 340035 625816
rect 339867 625762 340035 625782
rect 339565 625726 340035 625762
rect 339565 625707 339982 625726
rect 339565 625673 339584 625707
rect 339618 625706 339982 625707
rect 339618 625673 339732 625706
rect 339565 625672 339732 625673
rect 339766 625672 339833 625706
rect 339867 625692 339982 625706
rect 340016 625692 340035 625726
rect 339867 625672 340035 625692
rect 339565 625636 340035 625672
rect 339565 625617 339982 625636
rect 339565 625583 339584 625617
rect 339618 625616 339982 625617
rect 339618 625583 339732 625616
rect 339565 625582 339732 625583
rect 339766 625582 339833 625616
rect 339867 625602 339982 625616
rect 340016 625602 340035 625636
rect 339867 625582 340035 625602
rect 339565 625546 340035 625582
rect 339565 625527 339982 625546
rect 339565 625493 339584 625527
rect 339618 625526 339982 625527
rect 339618 625493 339732 625526
rect 339565 625492 339732 625493
rect 339766 625492 339833 625526
rect 339867 625512 339982 625526
rect 340016 625512 340035 625546
rect 339867 625492 340035 625512
rect 338277 625437 338694 625456
rect 338277 625403 338296 625437
rect 338330 625436 338694 625437
rect 338330 625403 338444 625436
rect 338277 625402 338444 625403
rect 338478 625402 338545 625436
rect 338579 625422 338694 625436
rect 338728 625422 338747 625456
rect 338579 625402 338747 625422
rect 338277 625399 338747 625402
rect 339565 625456 340035 625492
rect 340097 626094 340791 626155
rect 340097 626060 340156 626094
rect 340190 626082 340246 626094
rect 340218 626060 340246 626082
rect 340280 626082 340336 626094
rect 340280 626060 340284 626082
rect 340097 626048 340184 626060
rect 340218 626048 340284 626060
rect 340318 626060 340336 626082
rect 340370 626082 340426 626094
rect 340370 626060 340384 626082
rect 340318 626048 340384 626060
rect 340418 626060 340426 626082
rect 340460 626082 340516 626094
rect 340550 626082 340606 626094
rect 340640 626082 340696 626094
rect 340460 626060 340484 626082
rect 340550 626060 340584 626082
rect 340640 626060 340684 626082
rect 340730 626060 340791 626094
rect 340418 626048 340484 626060
rect 340518 626048 340584 626060
rect 340618 626048 340684 626060
rect 340718 626048 340791 626060
rect 340097 626004 340791 626048
rect 340097 625970 340156 626004
rect 340190 625982 340246 626004
rect 340218 625970 340246 625982
rect 340280 625982 340336 626004
rect 340280 625970 340284 625982
rect 340097 625948 340184 625970
rect 340218 625948 340284 625970
rect 340318 625970 340336 625982
rect 340370 625982 340426 626004
rect 340370 625970 340384 625982
rect 340318 625948 340384 625970
rect 340418 625970 340426 625982
rect 340460 625982 340516 626004
rect 340550 625982 340606 626004
rect 340640 625982 340696 626004
rect 340460 625970 340484 625982
rect 340550 625970 340584 625982
rect 340640 625970 340684 625982
rect 340730 625970 340791 626004
rect 340418 625948 340484 625970
rect 340518 625948 340584 625970
rect 340618 625948 340684 625970
rect 340718 625948 340791 625970
rect 340097 625914 340791 625948
rect 340097 625880 340156 625914
rect 340190 625882 340246 625914
rect 340218 625880 340246 625882
rect 340280 625882 340336 625914
rect 340280 625880 340284 625882
rect 340097 625848 340184 625880
rect 340218 625848 340284 625880
rect 340318 625880 340336 625882
rect 340370 625882 340426 625914
rect 340370 625880 340384 625882
rect 340318 625848 340384 625880
rect 340418 625880 340426 625882
rect 340460 625882 340516 625914
rect 340550 625882 340606 625914
rect 340640 625882 340696 625914
rect 340460 625880 340484 625882
rect 340550 625880 340584 625882
rect 340640 625880 340684 625882
rect 340730 625880 340791 625914
rect 340418 625848 340484 625880
rect 340518 625848 340584 625880
rect 340618 625848 340684 625880
rect 340718 625848 340791 625880
rect 340097 625824 340791 625848
rect 340097 625790 340156 625824
rect 340190 625790 340246 625824
rect 340280 625790 340336 625824
rect 340370 625790 340426 625824
rect 340460 625790 340516 625824
rect 340550 625790 340606 625824
rect 340640 625790 340696 625824
rect 340730 625790 340791 625824
rect 340097 625782 340791 625790
rect 340097 625748 340184 625782
rect 340218 625748 340284 625782
rect 340318 625748 340384 625782
rect 340418 625748 340484 625782
rect 340518 625748 340584 625782
rect 340618 625748 340684 625782
rect 340718 625748 340791 625782
rect 340097 625734 340791 625748
rect 340097 625700 340156 625734
rect 340190 625700 340246 625734
rect 340280 625700 340336 625734
rect 340370 625700 340426 625734
rect 340460 625700 340516 625734
rect 340550 625700 340606 625734
rect 340640 625700 340696 625734
rect 340730 625700 340791 625734
rect 340097 625682 340791 625700
rect 340097 625648 340184 625682
rect 340218 625648 340284 625682
rect 340318 625648 340384 625682
rect 340418 625648 340484 625682
rect 340518 625648 340584 625682
rect 340618 625648 340684 625682
rect 340718 625648 340791 625682
rect 340097 625644 340791 625648
rect 340097 625610 340156 625644
rect 340190 625610 340246 625644
rect 340280 625610 340336 625644
rect 340370 625610 340426 625644
rect 340460 625610 340516 625644
rect 340550 625610 340606 625644
rect 340640 625610 340696 625644
rect 340730 625610 340791 625644
rect 340097 625582 340791 625610
rect 340097 625554 340184 625582
rect 340218 625554 340284 625582
rect 340097 625520 340156 625554
rect 340218 625548 340246 625554
rect 340190 625520 340246 625548
rect 340280 625548 340284 625554
rect 340318 625554 340384 625582
rect 340318 625548 340336 625554
rect 340280 625520 340336 625548
rect 340370 625548 340384 625554
rect 340418 625554 340484 625582
rect 340518 625554 340584 625582
rect 340618 625554 340684 625582
rect 340718 625554 340791 625582
rect 340418 625548 340426 625554
rect 340370 625520 340426 625548
rect 340460 625548 340484 625554
rect 340550 625548 340584 625554
rect 340640 625548 340684 625554
rect 340460 625520 340516 625548
rect 340550 625520 340606 625548
rect 340640 625520 340696 625548
rect 340730 625520 340791 625554
rect 340097 625461 340791 625520
rect 340853 626123 340872 626157
rect 340906 626156 341088 626157
rect 340906 626123 341020 626156
rect 340853 626122 341020 626123
rect 341054 626122 341088 626156
rect 340853 626067 341088 626122
rect 340853 626033 340872 626067
rect 340906 626066 341088 626067
rect 340906 626033 341020 626066
rect 340853 626032 341020 626033
rect 341054 626032 341088 626066
rect 340853 625977 341088 626032
rect 340853 625943 340872 625977
rect 340906 625976 341088 625977
rect 340906 625943 341020 625976
rect 340853 625942 341020 625943
rect 341054 625942 341088 625976
rect 340853 625887 341088 625942
rect 340853 625853 340872 625887
rect 340906 625886 341088 625887
rect 340906 625853 341020 625886
rect 340853 625852 341020 625853
rect 341054 625852 341088 625886
rect 340853 625797 341088 625852
rect 340853 625763 340872 625797
rect 340906 625796 341088 625797
rect 340906 625763 341020 625796
rect 340853 625762 341020 625763
rect 341054 625762 341088 625796
rect 340853 625707 341088 625762
rect 340853 625673 340872 625707
rect 340906 625706 341088 625707
rect 340906 625673 341020 625706
rect 340853 625672 341020 625673
rect 341054 625672 341088 625706
rect 340853 625617 341088 625672
rect 340853 625583 340872 625617
rect 340906 625616 341088 625617
rect 340906 625583 341020 625616
rect 340853 625582 341020 625583
rect 341054 625582 341088 625616
rect 340853 625527 341088 625582
rect 340853 625493 340872 625527
rect 340906 625526 341088 625527
rect 340906 625493 341020 625526
rect 340853 625492 341020 625493
rect 341054 625492 341088 625526
rect 339565 625437 339982 625456
rect 339565 625403 339584 625437
rect 339618 625436 339982 625437
rect 339618 625403 339732 625436
rect 339565 625402 339732 625403
rect 339766 625402 339833 625436
rect 339867 625422 339982 625436
rect 340016 625422 340035 625456
rect 339867 625402 340035 625422
rect 339565 625399 340035 625402
rect 340853 625437 341088 625492
rect 340853 625403 340872 625437
rect 340906 625436 341088 625437
rect 340906 625403 341020 625436
rect 340853 625402 341020 625403
rect 341054 625402 341088 625436
rect 340853 625399 341088 625402
rect 334648 625380 341088 625399
rect 334648 625346 334888 625380
rect 334922 625346 334978 625380
rect 335012 625346 335068 625380
rect 335102 625346 335158 625380
rect 335192 625346 335248 625380
rect 335282 625346 335338 625380
rect 335372 625346 335428 625380
rect 335462 625346 335518 625380
rect 335552 625346 335608 625380
rect 335642 625346 336176 625380
rect 336210 625346 336266 625380
rect 336300 625346 336356 625380
rect 336390 625346 336446 625380
rect 336480 625346 336536 625380
rect 336570 625346 336626 625380
rect 336660 625346 336716 625380
rect 336750 625346 336806 625380
rect 336840 625346 336896 625380
rect 336930 625346 337464 625380
rect 337498 625346 337554 625380
rect 337588 625346 337644 625380
rect 337678 625346 337734 625380
rect 337768 625346 337824 625380
rect 337858 625346 337914 625380
rect 337948 625346 338004 625380
rect 338038 625346 338094 625380
rect 338128 625346 338184 625380
rect 338218 625346 338752 625380
rect 338786 625346 338842 625380
rect 338876 625346 338932 625380
rect 338966 625346 339022 625380
rect 339056 625346 339112 625380
rect 339146 625346 339202 625380
rect 339236 625346 339292 625380
rect 339326 625346 339382 625380
rect 339416 625346 339472 625380
rect 339506 625346 340040 625380
rect 340074 625346 340130 625380
rect 340164 625346 340220 625380
rect 340254 625346 340310 625380
rect 340344 625346 340400 625380
rect 340434 625346 340490 625380
rect 340524 625346 340580 625380
rect 340614 625346 340670 625380
rect 340704 625346 340760 625380
rect 340794 625346 341088 625380
rect 334648 625312 334681 625346
rect 334715 625327 335868 625346
rect 334715 625312 334888 625327
rect 334648 625263 334888 625312
rect 335688 625312 335868 625327
rect 335902 625312 335969 625346
rect 336003 625327 337156 625346
rect 336003 625312 336188 625327
rect 335688 625263 336188 625312
rect 336988 625312 337156 625327
rect 337190 625312 337257 625346
rect 337291 625327 338444 625346
rect 337291 625312 337388 625327
rect 336988 625263 337388 625312
rect 338288 625312 338444 625327
rect 338478 625312 338545 625346
rect 338579 625327 339732 625346
rect 338579 625312 338688 625327
rect 338288 625263 338688 625312
rect 339588 625312 339732 625327
rect 339766 625312 339833 625346
rect 339867 625327 341020 625346
rect 339867 625312 339988 625327
rect 339588 625263 339988 625312
rect 340888 625312 341020 625327
rect 341054 625312 341088 625346
rect 340888 625263 341088 625312
rect 334648 625256 341088 625263
rect 334648 625222 334681 625256
rect 334715 625233 335868 625256
rect 334715 625222 334782 625233
rect 334648 625199 334782 625222
rect 334816 625199 334872 625233
rect 334906 625199 334962 625233
rect 334996 625199 335052 625233
rect 335086 625199 335142 625233
rect 335176 625199 335232 625233
rect 335266 625199 335322 625233
rect 335356 625199 335412 625233
rect 335446 625199 335502 625233
rect 335536 625199 335592 625233
rect 335626 625199 335682 625233
rect 335716 625199 335772 625233
rect 335806 625222 335868 625233
rect 335902 625222 335969 625256
rect 336003 625233 337156 625256
rect 336003 625222 336070 625233
rect 335806 625199 336070 625222
rect 336104 625199 336160 625233
rect 336194 625199 336250 625233
rect 336284 625199 336340 625233
rect 336374 625199 336430 625233
rect 336464 625199 336520 625233
rect 336554 625199 336610 625233
rect 336644 625199 336700 625233
rect 336734 625199 336790 625233
rect 336824 625199 336880 625233
rect 336914 625199 336970 625233
rect 337004 625199 337060 625233
rect 337094 625222 337156 625233
rect 337190 625222 337257 625256
rect 337291 625233 338444 625256
rect 337291 625222 337358 625233
rect 337094 625199 337358 625222
rect 337392 625199 337448 625233
rect 337482 625199 337538 625233
rect 337572 625199 337628 625233
rect 337662 625199 337718 625233
rect 337752 625199 337808 625233
rect 337842 625199 337898 625233
rect 337932 625199 337988 625233
rect 338022 625199 338078 625233
rect 338112 625199 338168 625233
rect 338202 625199 338258 625233
rect 338292 625199 338348 625233
rect 338382 625222 338444 625233
rect 338478 625222 338545 625256
rect 338579 625233 339732 625256
rect 338579 625222 338646 625233
rect 338382 625199 338646 625222
rect 338680 625199 338736 625233
rect 338770 625199 338826 625233
rect 338860 625199 338916 625233
rect 338950 625199 339006 625233
rect 339040 625199 339096 625233
rect 339130 625199 339186 625233
rect 339220 625199 339276 625233
rect 339310 625199 339366 625233
rect 339400 625199 339456 625233
rect 339490 625199 339546 625233
rect 339580 625199 339636 625233
rect 339670 625222 339732 625233
rect 339766 625222 339833 625256
rect 339867 625233 341020 625256
rect 339867 625222 339934 625233
rect 339670 625199 339934 625222
rect 339968 625199 340024 625233
rect 340058 625199 340114 625233
rect 340148 625199 340204 625233
rect 340238 625199 340294 625233
rect 340328 625199 340384 625233
rect 340418 625199 340474 625233
rect 340508 625199 340564 625233
rect 340598 625199 340654 625233
rect 340688 625199 340744 625233
rect 340778 625199 340834 625233
rect 340868 625199 340924 625233
rect 340958 625222 341020 625233
rect 341054 625222 341088 625256
rect 340958 625199 341088 625222
rect 334648 625132 341088 625199
rect 334648 625098 334782 625132
rect 334816 625098 334872 625132
rect 334906 625098 334962 625132
rect 334996 625098 335052 625132
rect 335086 625098 335142 625132
rect 335176 625098 335232 625132
rect 335266 625098 335322 625132
rect 335356 625098 335412 625132
rect 335446 625098 335502 625132
rect 335536 625098 335592 625132
rect 335626 625098 335682 625132
rect 335716 625098 335772 625132
rect 335806 625098 336070 625132
rect 336104 625098 336160 625132
rect 336194 625098 336250 625132
rect 336284 625098 336340 625132
rect 336374 625098 336430 625132
rect 336464 625098 336520 625132
rect 336554 625098 336610 625132
rect 336644 625098 336700 625132
rect 336734 625098 336790 625132
rect 336824 625098 336880 625132
rect 336914 625098 336970 625132
rect 337004 625098 337060 625132
rect 337094 625098 337358 625132
rect 337392 625098 337448 625132
rect 337482 625098 337538 625132
rect 337572 625098 337628 625132
rect 337662 625098 337718 625132
rect 337752 625098 337808 625132
rect 337842 625098 337898 625132
rect 337932 625098 337988 625132
rect 338022 625098 338078 625132
rect 338112 625098 338168 625132
rect 338202 625098 338258 625132
rect 338292 625098 338348 625132
rect 338382 625098 338646 625132
rect 338680 625098 338736 625132
rect 338770 625098 338826 625132
rect 338860 625098 338916 625132
rect 338950 625098 339006 625132
rect 339040 625098 339096 625132
rect 339130 625098 339186 625132
rect 339220 625098 339276 625132
rect 339310 625098 339366 625132
rect 339400 625098 339456 625132
rect 339490 625098 339546 625132
rect 339580 625098 339636 625132
rect 339670 625098 339934 625132
rect 339968 625098 340024 625132
rect 340058 625098 340114 625132
rect 340148 625098 340204 625132
rect 340238 625098 340294 625132
rect 340328 625098 340384 625132
rect 340418 625098 340474 625132
rect 340508 625098 340564 625132
rect 340598 625098 340654 625132
rect 340688 625098 340744 625132
rect 340778 625098 340834 625132
rect 340868 625098 340924 625132
rect 340958 625098 341088 625132
rect 334648 625065 341088 625098
rect 334648 625048 334888 625065
rect 334648 625014 334681 625048
rect 334715 625014 334888 625048
rect 334648 625001 334888 625014
rect 335688 625048 336188 625065
rect 335688 625014 335868 625048
rect 335902 625014 335969 625048
rect 336003 625014 336188 625048
rect 335688 625001 336188 625014
rect 336988 625048 337388 625065
rect 336988 625014 337156 625048
rect 337190 625014 337257 625048
rect 337291 625014 337388 625048
rect 336988 625001 337388 625014
rect 338288 625048 338688 625065
rect 338288 625014 338444 625048
rect 338478 625014 338545 625048
rect 338579 625014 338688 625048
rect 338288 625001 338688 625014
rect 339588 625048 339988 625065
rect 339588 625014 339732 625048
rect 339766 625014 339833 625048
rect 339867 625014 339988 625048
rect 339588 625001 339988 625014
rect 340888 625048 341088 625065
rect 340888 625014 341020 625048
rect 341054 625014 341088 625048
rect 340888 625001 341088 625014
rect 334648 624982 341088 625001
rect 334648 624958 334922 624982
rect 313404 624934 313438 624950
rect 304306 624894 310790 624904
rect 304306 624550 304316 624894
rect 310780 624550 310790 624894
rect 304306 624540 310790 624550
rect 312704 624608 313304 624808
rect 305024 624324 305040 624358
rect 310416 624324 310432 624358
rect 304956 624296 304990 624312
rect 304956 623912 304990 623928
rect 305024 623866 305040 623900
rect 310416 623866 310432 623900
rect 305368 622198 305384 622232
rect 305752 622198 305768 622232
rect 305940 622198 305956 622232
rect 306324 622198 306340 622232
rect 306512 622198 306528 622232
rect 306896 622198 306912 622232
rect 307084 622198 307100 622232
rect 307468 622198 307484 622232
rect 307656 622198 307672 622232
rect 308040 622198 308056 622232
rect 308228 622198 308244 622232
rect 308612 622198 308628 622232
rect 308800 622198 308816 622232
rect 309184 622198 309200 622232
rect 309372 622198 309388 622232
rect 309756 622198 309772 622232
rect 304754 622148 304886 622164
rect 301270 621342 302294 621358
rect 301270 621266 301286 621342
rect 302278 621266 302294 621342
rect 301270 621226 302294 621266
rect 299884 621188 300316 621204
rect 299884 620612 299900 621188
rect 300300 621110 300316 621188
rect 301270 621174 301298 621226
rect 301350 621174 302214 621226
rect 302266 621174 302294 621226
rect 301270 621162 302294 621174
rect 303250 621188 303682 621204
rect 303250 621110 303266 621188
rect 300300 621076 300454 621110
rect 300822 621076 300838 621110
rect 300896 621076 300912 621110
rect 301280 621076 301370 621110
rect 301738 621076 301828 621110
rect 302196 621076 302286 621110
rect 302654 621076 302670 621110
rect 302728 621076 302744 621110
rect 303112 621076 303266 621110
rect 300300 621026 300426 621076
rect 300300 620650 300392 621026
rect 300300 620634 300426 620650
rect 300850 621026 300884 621042
rect 300850 620634 300884 620650
rect 301308 621026 301342 621042
rect 301308 620634 301342 620650
rect 301766 621026 301800 621042
rect 301766 620634 301800 620650
rect 302224 621026 302258 621042
rect 302224 620634 302258 620650
rect 302682 621026 302716 621042
rect 302682 620634 302716 620650
rect 303140 621026 303266 621076
rect 303174 620650 303266 621026
rect 303140 620634 303266 620650
rect 300300 620612 300316 620634
rect 299884 620596 300316 620612
rect 303250 620612 303266 620634
rect 303666 620612 303682 621188
rect 303250 620596 303682 620612
rect 304754 620548 304770 622148
rect 304870 620548 304886 622148
rect 304754 620532 304886 620548
rect 305322 622148 305356 622164
rect 305322 620356 305356 620372
rect 305780 622148 305814 622164
rect 305780 620356 305814 620372
rect 305894 622148 305928 622164
rect 305894 620356 305928 620372
rect 306352 622148 306386 622164
rect 306352 620356 306386 620372
rect 306466 622148 306500 622164
rect 306466 620356 306500 620372
rect 306924 622148 306958 622164
rect 306924 620356 306958 620372
rect 307038 622148 307072 622164
rect 307038 620356 307072 620372
rect 307496 622148 307530 622164
rect 307496 620356 307530 620372
rect 307610 622148 307644 622164
rect 307610 620356 307644 620372
rect 308068 622148 308102 622164
rect 308068 620356 308102 620372
rect 308182 622148 308216 622164
rect 308182 620356 308216 620372
rect 308640 622148 308674 622164
rect 308640 620356 308674 620372
rect 308754 622148 308788 622164
rect 308754 620356 308788 620372
rect 309212 622148 309246 622164
rect 309212 620356 309246 620372
rect 309326 622148 309360 622164
rect 309326 620356 309360 620372
rect 309784 622148 309818 622164
rect 310254 622148 310386 622164
rect 310254 620548 310270 622148
rect 310370 620548 310386 622148
rect 310254 620532 310386 620548
rect 309784 620356 309818 620372
rect 303642 619795 303658 619829
rect 304026 619795 304042 619829
rect 304214 619795 304230 619829
rect 304598 619795 304614 619829
rect 304786 619795 304802 619829
rect 305170 619795 305186 619829
rect 305358 619795 305374 619829
rect 305742 619795 305758 619829
rect 305930 619795 305946 619829
rect 306314 619795 306330 619829
rect 306502 619795 306518 619829
rect 306886 619795 306902 619829
rect 307074 619795 307090 619829
rect 307458 619795 307474 619829
rect 307646 619795 307662 619829
rect 308030 619795 308046 619829
rect 308218 619795 308234 619829
rect 308602 619795 308618 619829
rect 308790 619795 308806 619829
rect 309174 619795 309190 619829
rect 309362 619795 309378 619829
rect 309746 619795 309762 619829
rect 309934 619795 309950 619829
rect 310318 619795 310334 619829
rect 310506 619795 310522 619829
rect 310890 619795 310906 619829
rect 311078 619795 311094 619829
rect 311462 619795 311478 619829
rect 303596 619736 303630 619752
rect 302938 619648 303070 619660
rect 302938 617306 302954 619648
rect 303054 617306 303070 619648
rect 302938 617290 303070 617306
rect 303596 617164 303630 617180
rect 304054 619736 304088 619752
rect 304054 617164 304088 617180
rect 304168 619736 304202 619752
rect 304168 617164 304202 617180
rect 304626 619736 304660 619752
rect 304626 617164 304660 617180
rect 304740 619736 304774 619752
rect 304740 617164 304774 617180
rect 305198 619736 305232 619752
rect 305198 617164 305232 617180
rect 305312 619736 305346 619752
rect 305312 617164 305346 617180
rect 305770 619736 305804 619752
rect 305770 617164 305804 617180
rect 305884 619736 305918 619752
rect 305884 617164 305918 617180
rect 306342 619736 306376 619752
rect 306342 617164 306376 617180
rect 306456 619736 306490 619752
rect 306456 617164 306490 617180
rect 306914 619736 306948 619752
rect 306914 617164 306948 617180
rect 307028 619736 307062 619752
rect 307028 617164 307062 617180
rect 307486 619736 307520 619752
rect 307486 617164 307520 617180
rect 307600 619736 307634 619752
rect 307600 617164 307634 617180
rect 308058 619736 308092 619752
rect 308058 617164 308092 617180
rect 308172 619736 308206 619752
rect 308172 617164 308206 617180
rect 308630 619736 308664 619752
rect 308630 617164 308664 617180
rect 308744 619736 308778 619752
rect 308744 617164 308778 617180
rect 309202 619736 309236 619752
rect 309202 617164 309236 617180
rect 309316 619736 309350 619752
rect 309316 617164 309350 617180
rect 309774 619736 309808 619752
rect 309774 617164 309808 617180
rect 309888 619736 309922 619752
rect 309888 617164 309922 617180
rect 310346 619736 310380 619752
rect 310346 617164 310380 617180
rect 310460 619736 310494 619752
rect 310460 617164 310494 617180
rect 310918 619736 310952 619752
rect 310918 617164 310952 617180
rect 311032 619736 311066 619752
rect 311032 617164 311066 617180
rect 311490 619736 311524 619752
rect 312066 619648 312198 619660
rect 312066 617306 312082 619648
rect 312182 617306 312198 619648
rect 312066 617290 312198 617306
rect 312704 617608 312904 624608
rect 313104 617608 313304 624608
rect 311490 617164 311524 617180
rect 306524 616802 308894 616818
rect 306524 616702 306536 616802
rect 308878 616702 308894 616802
rect 306524 616686 308894 616702
rect 312704 616708 313304 617608
rect 313404 617202 313438 617218
rect 313862 624934 313896 624950
rect 313862 617202 313896 617218
rect 314320 624934 314354 624950
rect 314320 617202 314354 617218
rect 314778 624934 314812 624950
rect 314778 617202 314812 617218
rect 315236 624934 315270 624950
rect 315236 617202 315270 617218
rect 315694 624934 315728 624950
rect 315694 617202 315728 617218
rect 316152 624934 316186 624950
rect 316152 617202 316186 617218
rect 316610 624934 316644 624950
rect 316610 617202 316644 617218
rect 317068 624934 317102 624950
rect 317068 617202 317102 617218
rect 317526 624934 317560 624950
rect 317526 617202 317560 617218
rect 317984 624934 318018 624950
rect 317984 617202 318018 617218
rect 318442 624934 318476 624950
rect 319362 624934 319396 624950
rect 318442 617202 318476 617218
rect 318614 624608 319214 624808
rect 318614 617608 318814 624608
rect 319014 617608 319214 624608
rect 313450 617125 313466 617159
rect 313834 617125 313850 617159
rect 313908 617125 313924 617159
rect 314292 617125 314308 617159
rect 314366 617125 314382 617159
rect 314750 617125 314766 617159
rect 314824 617125 314840 617159
rect 315208 617125 315224 617159
rect 315282 617125 315298 617159
rect 315666 617125 315682 617159
rect 315740 617125 315756 617159
rect 316124 617125 316140 617159
rect 316198 617125 316214 617159
rect 316582 617125 316598 617159
rect 316656 617125 316672 617159
rect 317040 617125 317056 617159
rect 317114 617125 317130 617159
rect 317498 617125 317514 617159
rect 317572 617125 317588 617159
rect 317956 617125 317972 617159
rect 318030 617125 318046 617159
rect 318414 617125 318430 617159
rect 312704 616608 312804 616708
rect 313204 616608 313304 616708
rect 312704 616508 313304 616608
rect 318614 616708 319214 617608
rect 319362 617202 319396 617218
rect 319820 624934 319854 624950
rect 319820 617202 319854 617218
rect 320278 624934 320312 624950
rect 320278 617202 320312 617218
rect 320736 624934 320770 624950
rect 320736 617202 320770 617218
rect 321194 624934 321228 624950
rect 321194 617202 321228 617218
rect 321652 624934 321686 624950
rect 321652 617202 321686 617218
rect 322110 624934 322144 624950
rect 322110 617202 322144 617218
rect 322568 624934 322602 624950
rect 322568 617202 322602 617218
rect 323026 624934 323060 624950
rect 323026 617202 323060 617218
rect 323484 624934 323518 624950
rect 323484 617202 323518 617218
rect 323942 624934 323976 624950
rect 324862 624934 324896 624950
rect 323942 617202 323976 617218
rect 324114 624608 324714 624808
rect 324114 617608 324314 624608
rect 324514 617608 324714 624608
rect 319408 617125 319424 617159
rect 319792 617125 319808 617159
rect 319866 617125 319882 617159
rect 320250 617125 320266 617159
rect 320324 617125 320340 617159
rect 320708 617125 320724 617159
rect 320782 617125 320798 617159
rect 321166 617125 321182 617159
rect 321240 617125 321256 617159
rect 321624 617125 321640 617159
rect 321698 617125 321714 617159
rect 322082 617125 322098 617159
rect 322156 617125 322172 617159
rect 322540 617125 322556 617159
rect 322614 617125 322630 617159
rect 322998 617125 323014 617159
rect 323072 617125 323088 617159
rect 323456 617125 323472 617159
rect 323530 617125 323546 617159
rect 323914 617125 323930 617159
rect 318614 616608 318714 616708
rect 319114 616608 319214 616708
rect 318614 616508 319214 616608
rect 324114 616708 324714 617608
rect 324862 617202 324896 617218
rect 325320 624934 325354 624950
rect 325320 617202 325354 617218
rect 325778 624934 325812 624950
rect 325778 617202 325812 617218
rect 326236 624934 326270 624950
rect 326236 617202 326270 617218
rect 326694 624934 326728 624950
rect 326694 617202 326728 617218
rect 327152 624934 327186 624950
rect 327152 617202 327186 617218
rect 327610 624934 327644 624950
rect 327610 617202 327644 617218
rect 328068 624934 328102 624950
rect 328068 617202 328102 617218
rect 328526 624934 328560 624950
rect 328526 617202 328560 617218
rect 328984 624934 329018 624950
rect 328984 617202 329018 617218
rect 329442 624934 329476 624950
rect 329442 617202 329476 617218
rect 329900 624934 329934 624950
rect 334648 624924 334681 624958
rect 334715 624948 334922 624958
rect 334956 624948 335012 624982
rect 335046 624948 335102 624982
rect 335136 624948 335192 624982
rect 335226 624948 335282 624982
rect 335316 624948 335372 624982
rect 335406 624948 335462 624982
rect 335496 624948 335552 624982
rect 335586 624948 335642 624982
rect 335676 624958 336210 624982
rect 335676 624948 335868 624958
rect 334715 624929 335868 624948
rect 334715 624924 334888 624929
rect 334648 624888 334888 624924
rect 334648 624868 334830 624888
rect 334648 624834 334681 624868
rect 334715 624854 334830 624868
rect 334864 624854 334888 624888
rect 335688 624924 335868 624929
rect 335902 624924 335969 624958
rect 336003 624948 336210 624958
rect 336244 624948 336300 624982
rect 336334 624948 336390 624982
rect 336424 624948 336480 624982
rect 336514 624948 336570 624982
rect 336604 624948 336660 624982
rect 336694 624948 336750 624982
rect 336784 624948 336840 624982
rect 336874 624948 336930 624982
rect 336964 624958 337498 624982
rect 336964 624948 337156 624958
rect 336003 624929 337156 624948
rect 336003 624924 336188 624929
rect 335688 624888 336188 624924
rect 335688 624869 336118 624888
rect 334715 624834 334888 624854
rect 329900 617202 329934 617218
rect 330070 624606 330670 624806
rect 330070 617606 330270 624606
rect 330470 617606 330670 624606
rect 324908 617125 324924 617159
rect 325292 617125 325308 617159
rect 325366 617125 325382 617159
rect 325750 617125 325766 617159
rect 325824 617125 325840 617159
rect 326208 617125 326224 617159
rect 326282 617125 326298 617159
rect 326666 617125 326682 617159
rect 326740 617125 326756 617159
rect 327124 617125 327140 617159
rect 327198 617125 327214 617159
rect 327582 617125 327598 617159
rect 327656 617125 327672 617159
rect 328040 617125 328056 617159
rect 328114 617125 328130 617159
rect 328498 617125 328514 617159
rect 328572 617125 328588 617159
rect 328956 617125 328972 617159
rect 329030 617125 329046 617159
rect 329414 617125 329430 617159
rect 329488 617125 329504 617159
rect 329872 617125 329888 617159
rect 324114 616608 324214 616708
rect 324614 616608 324714 616708
rect 324114 616508 324714 616608
rect 330070 616706 330670 617606
rect 334648 624798 334888 624834
rect 334648 624778 334830 624798
rect 334648 624744 334681 624778
rect 334715 624764 334830 624778
rect 334864 624764 334888 624798
rect 334715 624744 334888 624764
rect 334648 624708 334888 624744
rect 334648 624688 334830 624708
rect 334648 624654 334681 624688
rect 334715 624674 334830 624688
rect 334864 624674 334888 624708
rect 334715 624654 334888 624674
rect 334648 624618 334888 624654
rect 334648 624598 334830 624618
rect 334648 624564 334681 624598
rect 334715 624584 334830 624598
rect 334864 624584 334888 624618
rect 334715 624564 334888 624584
rect 334648 624528 334888 624564
rect 334648 624508 334830 624528
rect 334648 624474 334681 624508
rect 334715 624494 334830 624508
rect 334864 624494 334888 624528
rect 334715 624474 334888 624494
rect 334648 624438 334888 624474
rect 334648 624418 334830 624438
rect 334648 624384 334681 624418
rect 334715 624404 334830 624418
rect 334864 624404 334888 624438
rect 334715 624384 334888 624404
rect 334648 624348 334888 624384
rect 334648 624328 334830 624348
rect 334648 624294 334681 624328
rect 334715 624314 334830 624328
rect 334864 624314 334888 624348
rect 334715 624294 334888 624314
rect 334648 624258 334888 624294
rect 334648 624238 334830 624258
rect 334648 624204 334681 624238
rect 334715 624224 334830 624238
rect 334864 624224 334888 624258
rect 334715 624204 334888 624224
rect 334648 624168 334888 624204
rect 334945 624806 335639 624867
rect 334945 624772 335004 624806
rect 335038 624794 335094 624806
rect 335066 624772 335094 624794
rect 335128 624794 335184 624806
rect 335128 624772 335132 624794
rect 334945 624760 335032 624772
rect 335066 624760 335132 624772
rect 335166 624772 335184 624794
rect 335218 624794 335274 624806
rect 335218 624772 335232 624794
rect 335166 624760 335232 624772
rect 335266 624772 335274 624794
rect 335308 624794 335364 624806
rect 335398 624794 335454 624806
rect 335488 624794 335544 624806
rect 335308 624772 335332 624794
rect 335398 624772 335432 624794
rect 335488 624772 335532 624794
rect 335578 624772 335639 624806
rect 335266 624760 335332 624772
rect 335366 624760 335432 624772
rect 335466 624760 335532 624772
rect 335566 624760 335639 624772
rect 334945 624716 335639 624760
rect 334945 624682 335004 624716
rect 335038 624694 335094 624716
rect 335066 624682 335094 624694
rect 335128 624694 335184 624716
rect 335128 624682 335132 624694
rect 334945 624660 335032 624682
rect 335066 624660 335132 624682
rect 335166 624682 335184 624694
rect 335218 624694 335274 624716
rect 335218 624682 335232 624694
rect 335166 624660 335232 624682
rect 335266 624682 335274 624694
rect 335308 624694 335364 624716
rect 335398 624694 335454 624716
rect 335488 624694 335544 624716
rect 335308 624682 335332 624694
rect 335398 624682 335432 624694
rect 335488 624682 335532 624694
rect 335578 624682 335639 624716
rect 335266 624660 335332 624682
rect 335366 624660 335432 624682
rect 335466 624660 335532 624682
rect 335566 624660 335639 624682
rect 334945 624626 335639 624660
rect 334945 624592 335004 624626
rect 335038 624594 335094 624626
rect 335066 624592 335094 624594
rect 335128 624594 335184 624626
rect 335128 624592 335132 624594
rect 334945 624560 335032 624592
rect 335066 624560 335132 624592
rect 335166 624592 335184 624594
rect 335218 624594 335274 624626
rect 335218 624592 335232 624594
rect 335166 624560 335232 624592
rect 335266 624592 335274 624594
rect 335308 624594 335364 624626
rect 335398 624594 335454 624626
rect 335488 624594 335544 624626
rect 335308 624592 335332 624594
rect 335398 624592 335432 624594
rect 335488 624592 335532 624594
rect 335578 624592 335639 624626
rect 335266 624560 335332 624592
rect 335366 624560 335432 624592
rect 335466 624560 335532 624592
rect 335566 624560 335639 624592
rect 334945 624536 335639 624560
rect 334945 624502 335004 624536
rect 335038 624502 335094 624536
rect 335128 624502 335184 624536
rect 335218 624502 335274 624536
rect 335308 624502 335364 624536
rect 335398 624502 335454 624536
rect 335488 624502 335544 624536
rect 335578 624502 335639 624536
rect 334945 624494 335639 624502
rect 334945 624460 335032 624494
rect 335066 624460 335132 624494
rect 335166 624460 335232 624494
rect 335266 624460 335332 624494
rect 335366 624460 335432 624494
rect 335466 624460 335532 624494
rect 335566 624460 335639 624494
rect 334945 624446 335639 624460
rect 334945 624412 335004 624446
rect 335038 624412 335094 624446
rect 335128 624412 335184 624446
rect 335218 624412 335274 624446
rect 335308 624412 335364 624446
rect 335398 624412 335454 624446
rect 335488 624412 335544 624446
rect 335578 624412 335639 624446
rect 334945 624394 335639 624412
rect 334945 624360 335032 624394
rect 335066 624360 335132 624394
rect 335166 624360 335232 624394
rect 335266 624360 335332 624394
rect 335366 624360 335432 624394
rect 335466 624360 335532 624394
rect 335566 624360 335639 624394
rect 334945 624356 335639 624360
rect 334945 624322 335004 624356
rect 335038 624322 335094 624356
rect 335128 624322 335184 624356
rect 335218 624322 335274 624356
rect 335308 624322 335364 624356
rect 335398 624322 335454 624356
rect 335488 624322 335544 624356
rect 335578 624322 335639 624356
rect 334945 624294 335639 624322
rect 334945 624266 335032 624294
rect 335066 624266 335132 624294
rect 334945 624232 335004 624266
rect 335066 624260 335094 624266
rect 335038 624232 335094 624260
rect 335128 624260 335132 624266
rect 335166 624266 335232 624294
rect 335166 624260 335184 624266
rect 335128 624232 335184 624260
rect 335218 624260 335232 624266
rect 335266 624266 335332 624294
rect 335366 624266 335432 624294
rect 335466 624266 335532 624294
rect 335566 624266 335639 624294
rect 335266 624260 335274 624266
rect 335218 624232 335274 624260
rect 335308 624260 335332 624266
rect 335398 624260 335432 624266
rect 335488 624260 335532 624266
rect 335308 624232 335364 624260
rect 335398 624232 335454 624260
rect 335488 624232 335544 624260
rect 335578 624232 335639 624266
rect 334945 624173 335639 624232
rect 335688 624835 335720 624869
rect 335754 624868 336118 624869
rect 335754 624835 335868 624868
rect 335688 624834 335868 624835
rect 335902 624834 335969 624868
rect 336003 624854 336118 624868
rect 336152 624854 336188 624888
rect 336988 624924 337156 624929
rect 337190 624924 337257 624958
rect 337291 624948 337498 624958
rect 337532 624948 337588 624982
rect 337622 624948 337678 624982
rect 337712 624948 337768 624982
rect 337802 624948 337858 624982
rect 337892 624948 337948 624982
rect 337982 624948 338038 624982
rect 338072 624948 338128 624982
rect 338162 624948 338218 624982
rect 338252 624958 338786 624982
rect 338252 624948 338444 624958
rect 337291 624929 338444 624948
rect 337291 624924 337459 624929
rect 336988 624888 337459 624924
rect 336988 624869 337406 624888
rect 336003 624834 336188 624854
rect 335688 624798 336188 624834
rect 335688 624779 336118 624798
rect 335688 624745 335720 624779
rect 335754 624778 336118 624779
rect 335754 624745 335868 624778
rect 335688 624744 335868 624745
rect 335902 624744 335969 624778
rect 336003 624764 336118 624778
rect 336152 624764 336188 624798
rect 336003 624744 336188 624764
rect 335688 624708 336188 624744
rect 335688 624689 336118 624708
rect 335688 624655 335720 624689
rect 335754 624688 336118 624689
rect 335754 624655 335868 624688
rect 335688 624654 335868 624655
rect 335902 624654 335969 624688
rect 336003 624674 336118 624688
rect 336152 624674 336188 624708
rect 336003 624654 336188 624674
rect 335688 624618 336188 624654
rect 335688 624599 336118 624618
rect 335688 624565 335720 624599
rect 335754 624598 336118 624599
rect 335754 624565 335868 624598
rect 335688 624564 335868 624565
rect 335902 624564 335969 624598
rect 336003 624584 336118 624598
rect 336152 624584 336188 624618
rect 336003 624564 336188 624584
rect 335688 624528 336188 624564
rect 335688 624509 336118 624528
rect 335688 624475 335720 624509
rect 335754 624508 336118 624509
rect 335754 624475 335868 624508
rect 335688 624474 335868 624475
rect 335902 624474 335969 624508
rect 336003 624494 336118 624508
rect 336152 624494 336188 624528
rect 336003 624474 336188 624494
rect 335688 624438 336188 624474
rect 335688 624419 336118 624438
rect 335688 624385 335720 624419
rect 335754 624418 336118 624419
rect 335754 624385 335868 624418
rect 335688 624384 335868 624385
rect 335902 624384 335969 624418
rect 336003 624404 336118 624418
rect 336152 624404 336188 624438
rect 336003 624384 336188 624404
rect 335688 624348 336188 624384
rect 335688 624329 336118 624348
rect 335688 624295 335720 624329
rect 335754 624328 336118 624329
rect 335754 624295 335868 624328
rect 335688 624294 335868 624295
rect 335902 624294 335969 624328
rect 336003 624314 336118 624328
rect 336152 624314 336188 624348
rect 336003 624294 336188 624314
rect 335688 624258 336188 624294
rect 335688 624239 336118 624258
rect 335688 624205 335720 624239
rect 335754 624238 336118 624239
rect 335754 624205 335868 624238
rect 335688 624204 335868 624205
rect 335902 624204 335969 624238
rect 336003 624224 336118 624238
rect 336152 624224 336188 624258
rect 336003 624204 336188 624224
rect 334648 624148 334830 624168
rect 334648 624114 334681 624148
rect 334715 624134 334830 624148
rect 334864 624134 334888 624168
rect 334715 624114 334888 624134
rect 334648 624111 334888 624114
rect 335688 624168 336188 624204
rect 336233 624806 336927 624867
rect 336233 624772 336292 624806
rect 336326 624794 336382 624806
rect 336354 624772 336382 624794
rect 336416 624794 336472 624806
rect 336416 624772 336420 624794
rect 336233 624760 336320 624772
rect 336354 624760 336420 624772
rect 336454 624772 336472 624794
rect 336506 624794 336562 624806
rect 336506 624772 336520 624794
rect 336454 624760 336520 624772
rect 336554 624772 336562 624794
rect 336596 624794 336652 624806
rect 336686 624794 336742 624806
rect 336776 624794 336832 624806
rect 336596 624772 336620 624794
rect 336686 624772 336720 624794
rect 336776 624772 336820 624794
rect 336866 624772 336927 624806
rect 336554 624760 336620 624772
rect 336654 624760 336720 624772
rect 336754 624760 336820 624772
rect 336854 624760 336927 624772
rect 336233 624716 336927 624760
rect 336233 624682 336292 624716
rect 336326 624694 336382 624716
rect 336354 624682 336382 624694
rect 336416 624694 336472 624716
rect 336416 624682 336420 624694
rect 336233 624660 336320 624682
rect 336354 624660 336420 624682
rect 336454 624682 336472 624694
rect 336506 624694 336562 624716
rect 336506 624682 336520 624694
rect 336454 624660 336520 624682
rect 336554 624682 336562 624694
rect 336596 624694 336652 624716
rect 336686 624694 336742 624716
rect 336776 624694 336832 624716
rect 336596 624682 336620 624694
rect 336686 624682 336720 624694
rect 336776 624682 336820 624694
rect 336866 624682 336927 624716
rect 336554 624660 336620 624682
rect 336654 624660 336720 624682
rect 336754 624660 336820 624682
rect 336854 624660 336927 624682
rect 336233 624626 336927 624660
rect 336233 624592 336292 624626
rect 336326 624594 336382 624626
rect 336354 624592 336382 624594
rect 336416 624594 336472 624626
rect 336416 624592 336420 624594
rect 336233 624560 336320 624592
rect 336354 624560 336420 624592
rect 336454 624592 336472 624594
rect 336506 624594 336562 624626
rect 336506 624592 336520 624594
rect 336454 624560 336520 624592
rect 336554 624592 336562 624594
rect 336596 624594 336652 624626
rect 336686 624594 336742 624626
rect 336776 624594 336832 624626
rect 336596 624592 336620 624594
rect 336686 624592 336720 624594
rect 336776 624592 336820 624594
rect 336866 624592 336927 624626
rect 336554 624560 336620 624592
rect 336654 624560 336720 624592
rect 336754 624560 336820 624592
rect 336854 624560 336927 624592
rect 336233 624536 336927 624560
rect 336233 624502 336292 624536
rect 336326 624502 336382 624536
rect 336416 624502 336472 624536
rect 336506 624502 336562 624536
rect 336596 624502 336652 624536
rect 336686 624502 336742 624536
rect 336776 624502 336832 624536
rect 336866 624502 336927 624536
rect 336233 624494 336927 624502
rect 336233 624460 336320 624494
rect 336354 624460 336420 624494
rect 336454 624460 336520 624494
rect 336554 624460 336620 624494
rect 336654 624460 336720 624494
rect 336754 624460 336820 624494
rect 336854 624460 336927 624494
rect 336233 624446 336927 624460
rect 336233 624412 336292 624446
rect 336326 624412 336382 624446
rect 336416 624412 336472 624446
rect 336506 624412 336562 624446
rect 336596 624412 336652 624446
rect 336686 624412 336742 624446
rect 336776 624412 336832 624446
rect 336866 624412 336927 624446
rect 336233 624394 336927 624412
rect 336233 624360 336320 624394
rect 336354 624360 336420 624394
rect 336454 624360 336520 624394
rect 336554 624360 336620 624394
rect 336654 624360 336720 624394
rect 336754 624360 336820 624394
rect 336854 624360 336927 624394
rect 336233 624356 336927 624360
rect 336233 624322 336292 624356
rect 336326 624322 336382 624356
rect 336416 624322 336472 624356
rect 336506 624322 336562 624356
rect 336596 624322 336652 624356
rect 336686 624322 336742 624356
rect 336776 624322 336832 624356
rect 336866 624322 336927 624356
rect 336233 624294 336927 624322
rect 336233 624266 336320 624294
rect 336354 624266 336420 624294
rect 336233 624232 336292 624266
rect 336354 624260 336382 624266
rect 336326 624232 336382 624260
rect 336416 624260 336420 624266
rect 336454 624266 336520 624294
rect 336454 624260 336472 624266
rect 336416 624232 336472 624260
rect 336506 624260 336520 624266
rect 336554 624266 336620 624294
rect 336654 624266 336720 624294
rect 336754 624266 336820 624294
rect 336854 624266 336927 624294
rect 336554 624260 336562 624266
rect 336506 624232 336562 624260
rect 336596 624260 336620 624266
rect 336686 624260 336720 624266
rect 336776 624260 336820 624266
rect 336596 624232 336652 624260
rect 336686 624232 336742 624260
rect 336776 624232 336832 624260
rect 336866 624232 336927 624266
rect 336233 624173 336927 624232
rect 336988 624835 337008 624869
rect 337042 624868 337406 624869
rect 337042 624835 337156 624868
rect 336988 624834 337156 624835
rect 337190 624834 337257 624868
rect 337291 624854 337406 624868
rect 337440 624854 337459 624888
rect 338277 624924 338444 624929
rect 338478 624924 338545 624958
rect 338579 624948 338786 624958
rect 338820 624948 338876 624982
rect 338910 624948 338966 624982
rect 339000 624948 339056 624982
rect 339090 624948 339146 624982
rect 339180 624948 339236 624982
rect 339270 624948 339326 624982
rect 339360 624948 339416 624982
rect 339450 624948 339506 624982
rect 339540 624958 340074 624982
rect 339540 624948 339732 624958
rect 338579 624929 339732 624948
rect 338579 624924 338747 624929
rect 338277 624888 338747 624924
rect 338277 624869 338694 624888
rect 337291 624834 337459 624854
rect 336988 624798 337459 624834
rect 336988 624779 337406 624798
rect 336988 624745 337008 624779
rect 337042 624778 337406 624779
rect 337042 624745 337156 624778
rect 336988 624744 337156 624745
rect 337190 624744 337257 624778
rect 337291 624764 337406 624778
rect 337440 624764 337459 624798
rect 337291 624744 337459 624764
rect 336988 624708 337459 624744
rect 336988 624689 337406 624708
rect 336988 624655 337008 624689
rect 337042 624688 337406 624689
rect 337042 624655 337156 624688
rect 336988 624654 337156 624655
rect 337190 624654 337257 624688
rect 337291 624674 337406 624688
rect 337440 624674 337459 624708
rect 337291 624654 337459 624674
rect 336988 624618 337459 624654
rect 336988 624599 337406 624618
rect 336988 624565 337008 624599
rect 337042 624598 337406 624599
rect 337042 624565 337156 624598
rect 336988 624564 337156 624565
rect 337190 624564 337257 624598
rect 337291 624584 337406 624598
rect 337440 624584 337459 624618
rect 337291 624564 337459 624584
rect 336988 624528 337459 624564
rect 336988 624509 337406 624528
rect 336988 624475 337008 624509
rect 337042 624508 337406 624509
rect 337042 624475 337156 624508
rect 336988 624474 337156 624475
rect 337190 624474 337257 624508
rect 337291 624494 337406 624508
rect 337440 624494 337459 624528
rect 337291 624474 337459 624494
rect 336988 624438 337459 624474
rect 336988 624419 337406 624438
rect 336988 624385 337008 624419
rect 337042 624418 337406 624419
rect 337042 624385 337156 624418
rect 336988 624384 337156 624385
rect 337190 624384 337257 624418
rect 337291 624404 337406 624418
rect 337440 624404 337459 624438
rect 337291 624384 337459 624404
rect 336988 624348 337459 624384
rect 336988 624329 337406 624348
rect 336988 624295 337008 624329
rect 337042 624328 337406 624329
rect 337042 624295 337156 624328
rect 336988 624294 337156 624295
rect 337190 624294 337257 624328
rect 337291 624314 337406 624328
rect 337440 624314 337459 624348
rect 337291 624294 337459 624314
rect 336988 624258 337459 624294
rect 336988 624239 337406 624258
rect 336988 624205 337008 624239
rect 337042 624238 337406 624239
rect 337042 624205 337156 624238
rect 336988 624204 337156 624205
rect 337190 624204 337257 624238
rect 337291 624224 337406 624238
rect 337440 624224 337459 624258
rect 337291 624204 337459 624224
rect 335688 624149 336118 624168
rect 335688 624115 335720 624149
rect 335754 624148 336118 624149
rect 335754 624115 335868 624148
rect 335688 624114 335868 624115
rect 335902 624114 335969 624148
rect 336003 624134 336118 624148
rect 336152 624134 336188 624168
rect 336003 624114 336188 624134
rect 335688 624111 336188 624114
rect 336988 624168 337459 624204
rect 337521 624806 338215 624867
rect 337521 624772 337580 624806
rect 337614 624794 337670 624806
rect 337642 624772 337670 624794
rect 337704 624794 337760 624806
rect 337704 624772 337708 624794
rect 337521 624760 337608 624772
rect 337642 624760 337708 624772
rect 337742 624772 337760 624794
rect 337794 624794 337850 624806
rect 337794 624772 337808 624794
rect 337742 624760 337808 624772
rect 337842 624772 337850 624794
rect 337884 624794 337940 624806
rect 337974 624794 338030 624806
rect 338064 624794 338120 624806
rect 337884 624772 337908 624794
rect 337974 624772 338008 624794
rect 338064 624772 338108 624794
rect 338154 624772 338215 624806
rect 337842 624760 337908 624772
rect 337942 624760 338008 624772
rect 338042 624760 338108 624772
rect 338142 624760 338215 624772
rect 337521 624716 338215 624760
rect 337521 624682 337580 624716
rect 337614 624694 337670 624716
rect 337642 624682 337670 624694
rect 337704 624694 337760 624716
rect 337704 624682 337708 624694
rect 337521 624660 337608 624682
rect 337642 624660 337708 624682
rect 337742 624682 337760 624694
rect 337794 624694 337850 624716
rect 337794 624682 337808 624694
rect 337742 624660 337808 624682
rect 337842 624682 337850 624694
rect 337884 624694 337940 624716
rect 337974 624694 338030 624716
rect 338064 624694 338120 624716
rect 337884 624682 337908 624694
rect 337974 624682 338008 624694
rect 338064 624682 338108 624694
rect 338154 624682 338215 624716
rect 337842 624660 337908 624682
rect 337942 624660 338008 624682
rect 338042 624660 338108 624682
rect 338142 624660 338215 624682
rect 337521 624626 338215 624660
rect 337521 624592 337580 624626
rect 337614 624594 337670 624626
rect 337642 624592 337670 624594
rect 337704 624594 337760 624626
rect 337704 624592 337708 624594
rect 337521 624560 337608 624592
rect 337642 624560 337708 624592
rect 337742 624592 337760 624594
rect 337794 624594 337850 624626
rect 337794 624592 337808 624594
rect 337742 624560 337808 624592
rect 337842 624592 337850 624594
rect 337884 624594 337940 624626
rect 337974 624594 338030 624626
rect 338064 624594 338120 624626
rect 337884 624592 337908 624594
rect 337974 624592 338008 624594
rect 338064 624592 338108 624594
rect 338154 624592 338215 624626
rect 337842 624560 337908 624592
rect 337942 624560 338008 624592
rect 338042 624560 338108 624592
rect 338142 624560 338215 624592
rect 337521 624536 338215 624560
rect 337521 624502 337580 624536
rect 337614 624502 337670 624536
rect 337704 624502 337760 624536
rect 337794 624502 337850 624536
rect 337884 624502 337940 624536
rect 337974 624502 338030 624536
rect 338064 624502 338120 624536
rect 338154 624502 338215 624536
rect 337521 624494 338215 624502
rect 337521 624460 337608 624494
rect 337642 624460 337708 624494
rect 337742 624460 337808 624494
rect 337842 624460 337908 624494
rect 337942 624460 338008 624494
rect 338042 624460 338108 624494
rect 338142 624460 338215 624494
rect 337521 624446 338215 624460
rect 337521 624412 337580 624446
rect 337614 624412 337670 624446
rect 337704 624412 337760 624446
rect 337794 624412 337850 624446
rect 337884 624412 337940 624446
rect 337974 624412 338030 624446
rect 338064 624412 338120 624446
rect 338154 624412 338215 624446
rect 337521 624394 338215 624412
rect 337521 624360 337608 624394
rect 337642 624360 337708 624394
rect 337742 624360 337808 624394
rect 337842 624360 337908 624394
rect 337942 624360 338008 624394
rect 338042 624360 338108 624394
rect 338142 624360 338215 624394
rect 337521 624356 338215 624360
rect 337521 624322 337580 624356
rect 337614 624322 337670 624356
rect 337704 624322 337760 624356
rect 337794 624322 337850 624356
rect 337884 624322 337940 624356
rect 337974 624322 338030 624356
rect 338064 624322 338120 624356
rect 338154 624322 338215 624356
rect 337521 624294 338215 624322
rect 337521 624266 337608 624294
rect 337642 624266 337708 624294
rect 337521 624232 337580 624266
rect 337642 624260 337670 624266
rect 337614 624232 337670 624260
rect 337704 624260 337708 624266
rect 337742 624266 337808 624294
rect 337742 624260 337760 624266
rect 337704 624232 337760 624260
rect 337794 624260 337808 624266
rect 337842 624266 337908 624294
rect 337942 624266 338008 624294
rect 338042 624266 338108 624294
rect 338142 624266 338215 624294
rect 337842 624260 337850 624266
rect 337794 624232 337850 624260
rect 337884 624260 337908 624266
rect 337974 624260 338008 624266
rect 338064 624260 338108 624266
rect 337884 624232 337940 624260
rect 337974 624232 338030 624260
rect 338064 624232 338120 624260
rect 338154 624232 338215 624266
rect 337521 624173 338215 624232
rect 338277 624835 338296 624869
rect 338330 624868 338694 624869
rect 338330 624835 338444 624868
rect 338277 624834 338444 624835
rect 338478 624834 338545 624868
rect 338579 624854 338694 624868
rect 338728 624854 338747 624888
rect 339565 624924 339732 624929
rect 339766 624924 339833 624958
rect 339867 624948 340074 624958
rect 340108 624948 340164 624982
rect 340198 624948 340254 624982
rect 340288 624948 340344 624982
rect 340378 624948 340434 624982
rect 340468 624948 340524 624982
rect 340558 624948 340614 624982
rect 340648 624948 340704 624982
rect 340738 624948 340794 624982
rect 340828 624958 341088 624982
rect 340828 624948 341020 624958
rect 339867 624929 341020 624948
rect 339867 624924 340035 624929
rect 339565 624888 340035 624924
rect 339565 624869 339982 624888
rect 338579 624834 338747 624854
rect 338277 624798 338747 624834
rect 338277 624779 338694 624798
rect 338277 624745 338296 624779
rect 338330 624778 338694 624779
rect 338330 624745 338444 624778
rect 338277 624744 338444 624745
rect 338478 624744 338545 624778
rect 338579 624764 338694 624778
rect 338728 624764 338747 624798
rect 338579 624744 338747 624764
rect 338277 624708 338747 624744
rect 338277 624689 338694 624708
rect 338277 624655 338296 624689
rect 338330 624688 338694 624689
rect 338330 624655 338444 624688
rect 338277 624654 338444 624655
rect 338478 624654 338545 624688
rect 338579 624674 338694 624688
rect 338728 624674 338747 624708
rect 338579 624654 338747 624674
rect 338277 624618 338747 624654
rect 338277 624599 338694 624618
rect 338277 624565 338296 624599
rect 338330 624598 338694 624599
rect 338330 624565 338444 624598
rect 338277 624564 338444 624565
rect 338478 624564 338545 624598
rect 338579 624584 338694 624598
rect 338728 624584 338747 624618
rect 338579 624564 338747 624584
rect 338277 624528 338747 624564
rect 338277 624509 338694 624528
rect 338277 624475 338296 624509
rect 338330 624508 338694 624509
rect 338330 624475 338444 624508
rect 338277 624474 338444 624475
rect 338478 624474 338545 624508
rect 338579 624494 338694 624508
rect 338728 624494 338747 624528
rect 338579 624474 338747 624494
rect 338277 624438 338747 624474
rect 338277 624419 338694 624438
rect 338277 624385 338296 624419
rect 338330 624418 338694 624419
rect 338330 624385 338444 624418
rect 338277 624384 338444 624385
rect 338478 624384 338545 624418
rect 338579 624404 338694 624418
rect 338728 624404 338747 624438
rect 338579 624384 338747 624404
rect 338277 624348 338747 624384
rect 338277 624329 338694 624348
rect 338277 624295 338296 624329
rect 338330 624328 338694 624329
rect 338330 624295 338444 624328
rect 338277 624294 338444 624295
rect 338478 624294 338545 624328
rect 338579 624314 338694 624328
rect 338728 624314 338747 624348
rect 338579 624294 338747 624314
rect 338277 624258 338747 624294
rect 338277 624239 338694 624258
rect 338277 624205 338296 624239
rect 338330 624238 338694 624239
rect 338330 624205 338444 624238
rect 338277 624204 338444 624205
rect 338478 624204 338545 624238
rect 338579 624224 338694 624238
rect 338728 624224 338747 624258
rect 338579 624204 338747 624224
rect 336988 624149 337406 624168
rect 336988 624115 337008 624149
rect 337042 624148 337406 624149
rect 337042 624115 337156 624148
rect 336988 624114 337156 624115
rect 337190 624114 337257 624148
rect 337291 624134 337406 624148
rect 337440 624134 337459 624168
rect 337291 624114 337459 624134
rect 336988 624111 337459 624114
rect 338277 624168 338747 624204
rect 338809 624806 339503 624867
rect 338809 624772 338868 624806
rect 338902 624794 338958 624806
rect 338930 624772 338958 624794
rect 338992 624794 339048 624806
rect 338992 624772 338996 624794
rect 338809 624760 338896 624772
rect 338930 624760 338996 624772
rect 339030 624772 339048 624794
rect 339082 624794 339138 624806
rect 339082 624772 339096 624794
rect 339030 624760 339096 624772
rect 339130 624772 339138 624794
rect 339172 624794 339228 624806
rect 339262 624794 339318 624806
rect 339352 624794 339408 624806
rect 339172 624772 339196 624794
rect 339262 624772 339296 624794
rect 339352 624772 339396 624794
rect 339442 624772 339503 624806
rect 339130 624760 339196 624772
rect 339230 624760 339296 624772
rect 339330 624760 339396 624772
rect 339430 624760 339503 624772
rect 338809 624716 339503 624760
rect 338809 624682 338868 624716
rect 338902 624694 338958 624716
rect 338930 624682 338958 624694
rect 338992 624694 339048 624716
rect 338992 624682 338996 624694
rect 338809 624660 338896 624682
rect 338930 624660 338996 624682
rect 339030 624682 339048 624694
rect 339082 624694 339138 624716
rect 339082 624682 339096 624694
rect 339030 624660 339096 624682
rect 339130 624682 339138 624694
rect 339172 624694 339228 624716
rect 339262 624694 339318 624716
rect 339352 624694 339408 624716
rect 339172 624682 339196 624694
rect 339262 624682 339296 624694
rect 339352 624682 339396 624694
rect 339442 624682 339503 624716
rect 339130 624660 339196 624682
rect 339230 624660 339296 624682
rect 339330 624660 339396 624682
rect 339430 624660 339503 624682
rect 338809 624626 339503 624660
rect 338809 624592 338868 624626
rect 338902 624594 338958 624626
rect 338930 624592 338958 624594
rect 338992 624594 339048 624626
rect 338992 624592 338996 624594
rect 338809 624560 338896 624592
rect 338930 624560 338996 624592
rect 339030 624592 339048 624594
rect 339082 624594 339138 624626
rect 339082 624592 339096 624594
rect 339030 624560 339096 624592
rect 339130 624592 339138 624594
rect 339172 624594 339228 624626
rect 339262 624594 339318 624626
rect 339352 624594 339408 624626
rect 339172 624592 339196 624594
rect 339262 624592 339296 624594
rect 339352 624592 339396 624594
rect 339442 624592 339503 624626
rect 339130 624560 339196 624592
rect 339230 624560 339296 624592
rect 339330 624560 339396 624592
rect 339430 624560 339503 624592
rect 338809 624536 339503 624560
rect 338809 624502 338868 624536
rect 338902 624502 338958 624536
rect 338992 624502 339048 624536
rect 339082 624502 339138 624536
rect 339172 624502 339228 624536
rect 339262 624502 339318 624536
rect 339352 624502 339408 624536
rect 339442 624502 339503 624536
rect 338809 624494 339503 624502
rect 338809 624460 338896 624494
rect 338930 624460 338996 624494
rect 339030 624460 339096 624494
rect 339130 624460 339196 624494
rect 339230 624460 339296 624494
rect 339330 624460 339396 624494
rect 339430 624460 339503 624494
rect 338809 624446 339503 624460
rect 338809 624412 338868 624446
rect 338902 624412 338958 624446
rect 338992 624412 339048 624446
rect 339082 624412 339138 624446
rect 339172 624412 339228 624446
rect 339262 624412 339318 624446
rect 339352 624412 339408 624446
rect 339442 624412 339503 624446
rect 338809 624394 339503 624412
rect 338809 624360 338896 624394
rect 338930 624360 338996 624394
rect 339030 624360 339096 624394
rect 339130 624360 339196 624394
rect 339230 624360 339296 624394
rect 339330 624360 339396 624394
rect 339430 624360 339503 624394
rect 338809 624356 339503 624360
rect 338809 624322 338868 624356
rect 338902 624322 338958 624356
rect 338992 624322 339048 624356
rect 339082 624322 339138 624356
rect 339172 624322 339228 624356
rect 339262 624322 339318 624356
rect 339352 624322 339408 624356
rect 339442 624322 339503 624356
rect 338809 624294 339503 624322
rect 338809 624266 338896 624294
rect 338930 624266 338996 624294
rect 338809 624232 338868 624266
rect 338930 624260 338958 624266
rect 338902 624232 338958 624260
rect 338992 624260 338996 624266
rect 339030 624266 339096 624294
rect 339030 624260 339048 624266
rect 338992 624232 339048 624260
rect 339082 624260 339096 624266
rect 339130 624266 339196 624294
rect 339230 624266 339296 624294
rect 339330 624266 339396 624294
rect 339430 624266 339503 624294
rect 339130 624260 339138 624266
rect 339082 624232 339138 624260
rect 339172 624260 339196 624266
rect 339262 624260 339296 624266
rect 339352 624260 339396 624266
rect 339172 624232 339228 624260
rect 339262 624232 339318 624260
rect 339352 624232 339408 624260
rect 339442 624232 339503 624266
rect 338809 624173 339503 624232
rect 339565 624835 339584 624869
rect 339618 624868 339982 624869
rect 339618 624835 339732 624868
rect 339565 624834 339732 624835
rect 339766 624834 339833 624868
rect 339867 624854 339982 624868
rect 340016 624854 340035 624888
rect 340853 624924 341020 624929
rect 341054 624924 341088 624958
rect 340853 624869 341088 624924
rect 339867 624834 340035 624854
rect 339565 624798 340035 624834
rect 339565 624779 339982 624798
rect 339565 624745 339584 624779
rect 339618 624778 339982 624779
rect 339618 624745 339732 624778
rect 339565 624744 339732 624745
rect 339766 624744 339833 624778
rect 339867 624764 339982 624778
rect 340016 624764 340035 624798
rect 339867 624744 340035 624764
rect 339565 624708 340035 624744
rect 339565 624689 339982 624708
rect 339565 624655 339584 624689
rect 339618 624688 339982 624689
rect 339618 624655 339732 624688
rect 339565 624654 339732 624655
rect 339766 624654 339833 624688
rect 339867 624674 339982 624688
rect 340016 624674 340035 624708
rect 339867 624654 340035 624674
rect 339565 624618 340035 624654
rect 339565 624599 339982 624618
rect 339565 624565 339584 624599
rect 339618 624598 339982 624599
rect 339618 624565 339732 624598
rect 339565 624564 339732 624565
rect 339766 624564 339833 624598
rect 339867 624584 339982 624598
rect 340016 624584 340035 624618
rect 339867 624564 340035 624584
rect 339565 624528 340035 624564
rect 339565 624509 339982 624528
rect 339565 624475 339584 624509
rect 339618 624508 339982 624509
rect 339618 624475 339732 624508
rect 339565 624474 339732 624475
rect 339766 624474 339833 624508
rect 339867 624494 339982 624508
rect 340016 624494 340035 624528
rect 339867 624474 340035 624494
rect 339565 624438 340035 624474
rect 339565 624419 339982 624438
rect 339565 624385 339584 624419
rect 339618 624418 339982 624419
rect 339618 624385 339732 624418
rect 339565 624384 339732 624385
rect 339766 624384 339833 624418
rect 339867 624404 339982 624418
rect 340016 624404 340035 624438
rect 339867 624384 340035 624404
rect 339565 624348 340035 624384
rect 339565 624329 339982 624348
rect 339565 624295 339584 624329
rect 339618 624328 339982 624329
rect 339618 624295 339732 624328
rect 339565 624294 339732 624295
rect 339766 624294 339833 624328
rect 339867 624314 339982 624328
rect 340016 624314 340035 624348
rect 339867 624294 340035 624314
rect 339565 624258 340035 624294
rect 339565 624239 339982 624258
rect 339565 624205 339584 624239
rect 339618 624238 339982 624239
rect 339618 624205 339732 624238
rect 339565 624204 339732 624205
rect 339766 624204 339833 624238
rect 339867 624224 339982 624238
rect 340016 624224 340035 624258
rect 339867 624204 340035 624224
rect 338277 624149 338694 624168
rect 338277 624115 338296 624149
rect 338330 624148 338694 624149
rect 338330 624115 338444 624148
rect 338277 624114 338444 624115
rect 338478 624114 338545 624148
rect 338579 624134 338694 624148
rect 338728 624134 338747 624168
rect 338579 624114 338747 624134
rect 338277 624111 338747 624114
rect 339565 624168 340035 624204
rect 340097 624806 340791 624867
rect 340097 624772 340156 624806
rect 340190 624794 340246 624806
rect 340218 624772 340246 624794
rect 340280 624794 340336 624806
rect 340280 624772 340284 624794
rect 340097 624760 340184 624772
rect 340218 624760 340284 624772
rect 340318 624772 340336 624794
rect 340370 624794 340426 624806
rect 340370 624772 340384 624794
rect 340318 624760 340384 624772
rect 340418 624772 340426 624794
rect 340460 624794 340516 624806
rect 340550 624794 340606 624806
rect 340640 624794 340696 624806
rect 340460 624772 340484 624794
rect 340550 624772 340584 624794
rect 340640 624772 340684 624794
rect 340730 624772 340791 624806
rect 340418 624760 340484 624772
rect 340518 624760 340584 624772
rect 340618 624760 340684 624772
rect 340718 624760 340791 624772
rect 340097 624716 340791 624760
rect 340097 624682 340156 624716
rect 340190 624694 340246 624716
rect 340218 624682 340246 624694
rect 340280 624694 340336 624716
rect 340280 624682 340284 624694
rect 340097 624660 340184 624682
rect 340218 624660 340284 624682
rect 340318 624682 340336 624694
rect 340370 624694 340426 624716
rect 340370 624682 340384 624694
rect 340318 624660 340384 624682
rect 340418 624682 340426 624694
rect 340460 624694 340516 624716
rect 340550 624694 340606 624716
rect 340640 624694 340696 624716
rect 340460 624682 340484 624694
rect 340550 624682 340584 624694
rect 340640 624682 340684 624694
rect 340730 624682 340791 624716
rect 340418 624660 340484 624682
rect 340518 624660 340584 624682
rect 340618 624660 340684 624682
rect 340718 624660 340791 624682
rect 340097 624626 340791 624660
rect 340097 624592 340156 624626
rect 340190 624594 340246 624626
rect 340218 624592 340246 624594
rect 340280 624594 340336 624626
rect 340280 624592 340284 624594
rect 340097 624560 340184 624592
rect 340218 624560 340284 624592
rect 340318 624592 340336 624594
rect 340370 624594 340426 624626
rect 340370 624592 340384 624594
rect 340318 624560 340384 624592
rect 340418 624592 340426 624594
rect 340460 624594 340516 624626
rect 340550 624594 340606 624626
rect 340640 624594 340696 624626
rect 340460 624592 340484 624594
rect 340550 624592 340584 624594
rect 340640 624592 340684 624594
rect 340730 624592 340791 624626
rect 340418 624560 340484 624592
rect 340518 624560 340584 624592
rect 340618 624560 340684 624592
rect 340718 624560 340791 624592
rect 340097 624536 340791 624560
rect 340097 624502 340156 624536
rect 340190 624502 340246 624536
rect 340280 624502 340336 624536
rect 340370 624502 340426 624536
rect 340460 624502 340516 624536
rect 340550 624502 340606 624536
rect 340640 624502 340696 624536
rect 340730 624502 340791 624536
rect 340097 624494 340791 624502
rect 340097 624460 340184 624494
rect 340218 624460 340284 624494
rect 340318 624460 340384 624494
rect 340418 624460 340484 624494
rect 340518 624460 340584 624494
rect 340618 624460 340684 624494
rect 340718 624460 340791 624494
rect 340097 624446 340791 624460
rect 340097 624412 340156 624446
rect 340190 624412 340246 624446
rect 340280 624412 340336 624446
rect 340370 624412 340426 624446
rect 340460 624412 340516 624446
rect 340550 624412 340606 624446
rect 340640 624412 340696 624446
rect 340730 624412 340791 624446
rect 340097 624394 340791 624412
rect 340097 624360 340184 624394
rect 340218 624360 340284 624394
rect 340318 624360 340384 624394
rect 340418 624360 340484 624394
rect 340518 624360 340584 624394
rect 340618 624360 340684 624394
rect 340718 624360 340791 624394
rect 340097 624356 340791 624360
rect 340097 624322 340156 624356
rect 340190 624322 340246 624356
rect 340280 624322 340336 624356
rect 340370 624322 340426 624356
rect 340460 624322 340516 624356
rect 340550 624322 340606 624356
rect 340640 624322 340696 624356
rect 340730 624322 340791 624356
rect 340097 624294 340791 624322
rect 340097 624266 340184 624294
rect 340218 624266 340284 624294
rect 340097 624232 340156 624266
rect 340218 624260 340246 624266
rect 340190 624232 340246 624260
rect 340280 624260 340284 624266
rect 340318 624266 340384 624294
rect 340318 624260 340336 624266
rect 340280 624232 340336 624260
rect 340370 624260 340384 624266
rect 340418 624266 340484 624294
rect 340518 624266 340584 624294
rect 340618 624266 340684 624294
rect 340718 624266 340791 624294
rect 340418 624260 340426 624266
rect 340370 624232 340426 624260
rect 340460 624260 340484 624266
rect 340550 624260 340584 624266
rect 340640 624260 340684 624266
rect 340460 624232 340516 624260
rect 340550 624232 340606 624260
rect 340640 624232 340696 624260
rect 340730 624232 340791 624266
rect 340097 624173 340791 624232
rect 340853 624835 340872 624869
rect 340906 624868 341088 624869
rect 340906 624835 341020 624868
rect 340853 624834 341020 624835
rect 341054 624834 341088 624868
rect 340853 624779 341088 624834
rect 340853 624745 340872 624779
rect 340906 624778 341088 624779
rect 340906 624745 341020 624778
rect 340853 624744 341020 624745
rect 341054 624744 341088 624778
rect 340853 624689 341088 624744
rect 340853 624655 340872 624689
rect 340906 624688 341088 624689
rect 340906 624655 341020 624688
rect 340853 624654 341020 624655
rect 341054 624654 341088 624688
rect 340853 624599 341088 624654
rect 340853 624565 340872 624599
rect 340906 624598 341088 624599
rect 340906 624565 341020 624598
rect 340853 624564 341020 624565
rect 341054 624564 341088 624598
rect 340853 624509 341088 624564
rect 340853 624475 340872 624509
rect 340906 624508 341088 624509
rect 340906 624475 341020 624508
rect 340853 624474 341020 624475
rect 341054 624474 341088 624508
rect 340853 624419 341088 624474
rect 340853 624385 340872 624419
rect 340906 624418 341088 624419
rect 340906 624385 341020 624418
rect 340853 624384 341020 624385
rect 341054 624384 341088 624418
rect 340853 624329 341088 624384
rect 340853 624295 340872 624329
rect 340906 624328 341088 624329
rect 340906 624295 341020 624328
rect 340853 624294 341020 624295
rect 341054 624294 341088 624328
rect 340853 624239 341088 624294
rect 340853 624205 340872 624239
rect 340906 624238 341088 624239
rect 340906 624205 341020 624238
rect 340853 624204 341020 624205
rect 341054 624204 341088 624238
rect 339565 624149 339982 624168
rect 339565 624115 339584 624149
rect 339618 624148 339982 624149
rect 339618 624115 339732 624148
rect 339565 624114 339732 624115
rect 339766 624114 339833 624148
rect 339867 624134 339982 624148
rect 340016 624134 340035 624168
rect 339867 624114 340035 624134
rect 339565 624111 340035 624114
rect 340853 624149 341088 624204
rect 340853 624115 340872 624149
rect 340906 624148 341088 624149
rect 340906 624115 341020 624148
rect 340853 624114 341020 624115
rect 341054 624114 341088 624148
rect 340853 624111 341088 624114
rect 334648 624092 341088 624111
rect 334648 624058 334888 624092
rect 334922 624058 334978 624092
rect 335012 624058 335068 624092
rect 335102 624058 335158 624092
rect 335192 624058 335248 624092
rect 335282 624058 335338 624092
rect 335372 624058 335428 624092
rect 335462 624058 335518 624092
rect 335552 624058 335608 624092
rect 335642 624058 336176 624092
rect 336210 624058 336266 624092
rect 336300 624058 336356 624092
rect 336390 624058 336446 624092
rect 336480 624058 336536 624092
rect 336570 624058 336626 624092
rect 336660 624058 336716 624092
rect 336750 624058 336806 624092
rect 336840 624058 336896 624092
rect 336930 624058 337464 624092
rect 337498 624058 337554 624092
rect 337588 624058 337644 624092
rect 337678 624058 337734 624092
rect 337768 624058 337824 624092
rect 337858 624058 337914 624092
rect 337948 624058 338004 624092
rect 338038 624058 338094 624092
rect 338128 624058 338184 624092
rect 338218 624058 338752 624092
rect 338786 624058 338842 624092
rect 338876 624058 338932 624092
rect 338966 624058 339022 624092
rect 339056 624058 339112 624092
rect 339146 624058 339202 624092
rect 339236 624058 339292 624092
rect 339326 624058 339382 624092
rect 339416 624058 339472 624092
rect 339506 624058 340040 624092
rect 340074 624058 340130 624092
rect 340164 624058 340220 624092
rect 340254 624058 340310 624092
rect 340344 624058 340400 624092
rect 340434 624058 340490 624092
rect 340524 624058 340580 624092
rect 340614 624058 340670 624092
rect 340704 624058 340760 624092
rect 340794 624058 341088 624092
rect 334648 624024 334681 624058
rect 334715 624039 335868 624058
rect 334715 624024 334888 624039
rect 334648 623975 334888 624024
rect 335688 624024 335868 624039
rect 335902 624024 335969 624058
rect 336003 624039 337156 624058
rect 336003 624024 336188 624039
rect 335688 623975 336188 624024
rect 336988 624024 337156 624039
rect 337190 624024 337257 624058
rect 337291 624039 338444 624058
rect 337291 624024 337388 624039
rect 336988 623975 337388 624024
rect 338288 624024 338444 624039
rect 338478 624024 338545 624058
rect 338579 624039 339732 624058
rect 338579 624024 338688 624039
rect 338288 623975 338688 624024
rect 339588 624024 339732 624039
rect 339766 624024 339833 624058
rect 339867 624039 341020 624058
rect 339867 624024 339988 624039
rect 339588 623975 339988 624024
rect 340888 624024 341020 624039
rect 341054 624024 341088 624058
rect 340888 623975 341088 624024
rect 334648 623968 341088 623975
rect 334648 623934 334681 623968
rect 334715 623945 335868 623968
rect 334715 623934 334782 623945
rect 334648 623911 334782 623934
rect 334816 623911 334872 623945
rect 334906 623911 334962 623945
rect 334996 623911 335052 623945
rect 335086 623911 335142 623945
rect 335176 623911 335232 623945
rect 335266 623911 335322 623945
rect 335356 623911 335412 623945
rect 335446 623911 335502 623945
rect 335536 623911 335592 623945
rect 335626 623911 335682 623945
rect 335716 623911 335772 623945
rect 335806 623934 335868 623945
rect 335902 623934 335969 623968
rect 336003 623945 337156 623968
rect 336003 623934 336070 623945
rect 335806 623911 336070 623934
rect 336104 623911 336160 623945
rect 336194 623911 336250 623945
rect 336284 623911 336340 623945
rect 336374 623911 336430 623945
rect 336464 623911 336520 623945
rect 336554 623911 336610 623945
rect 336644 623911 336700 623945
rect 336734 623911 336790 623945
rect 336824 623911 336880 623945
rect 336914 623911 336970 623945
rect 337004 623911 337060 623945
rect 337094 623934 337156 623945
rect 337190 623934 337257 623968
rect 337291 623945 338444 623968
rect 337291 623934 337358 623945
rect 337094 623911 337358 623934
rect 337392 623911 337448 623945
rect 337482 623911 337538 623945
rect 337572 623911 337628 623945
rect 337662 623911 337718 623945
rect 337752 623911 337808 623945
rect 337842 623911 337898 623945
rect 337932 623911 337988 623945
rect 338022 623911 338078 623945
rect 338112 623911 338168 623945
rect 338202 623911 338258 623945
rect 338292 623911 338348 623945
rect 338382 623934 338444 623945
rect 338478 623934 338545 623968
rect 338579 623945 339732 623968
rect 338579 623934 338646 623945
rect 338382 623911 338646 623934
rect 338680 623911 338736 623945
rect 338770 623911 338826 623945
rect 338860 623911 338916 623945
rect 338950 623911 339006 623945
rect 339040 623911 339096 623945
rect 339130 623911 339186 623945
rect 339220 623911 339276 623945
rect 339310 623911 339366 623945
rect 339400 623911 339456 623945
rect 339490 623911 339546 623945
rect 339580 623911 339636 623945
rect 339670 623934 339732 623945
rect 339766 623934 339833 623968
rect 339867 623945 341020 623968
rect 339867 623934 339934 623945
rect 339670 623911 339934 623934
rect 339968 623911 340024 623945
rect 340058 623911 340114 623945
rect 340148 623911 340204 623945
rect 340238 623911 340294 623945
rect 340328 623911 340384 623945
rect 340418 623911 340474 623945
rect 340508 623911 340564 623945
rect 340598 623911 340654 623945
rect 340688 623911 340744 623945
rect 340778 623911 340834 623945
rect 340868 623911 340924 623945
rect 340958 623934 341020 623945
rect 341054 623934 341088 623968
rect 340958 623911 341088 623934
rect 334648 623844 341088 623911
rect 334648 623810 334782 623844
rect 334816 623810 334872 623844
rect 334906 623810 334962 623844
rect 334996 623810 335052 623844
rect 335086 623810 335142 623844
rect 335176 623810 335232 623844
rect 335266 623810 335322 623844
rect 335356 623810 335412 623844
rect 335446 623810 335502 623844
rect 335536 623810 335592 623844
rect 335626 623810 335682 623844
rect 335716 623810 335772 623844
rect 335806 623810 336070 623844
rect 336104 623810 336160 623844
rect 336194 623810 336250 623844
rect 336284 623810 336340 623844
rect 336374 623810 336430 623844
rect 336464 623810 336520 623844
rect 336554 623810 336610 623844
rect 336644 623810 336700 623844
rect 336734 623810 336790 623844
rect 336824 623810 336880 623844
rect 336914 623810 336970 623844
rect 337004 623810 337060 623844
rect 337094 623810 337358 623844
rect 337392 623810 337448 623844
rect 337482 623810 337538 623844
rect 337572 623810 337628 623844
rect 337662 623810 337718 623844
rect 337752 623810 337808 623844
rect 337842 623810 337898 623844
rect 337932 623810 337988 623844
rect 338022 623810 338078 623844
rect 338112 623810 338168 623844
rect 338202 623810 338258 623844
rect 338292 623810 338348 623844
rect 338382 623810 338646 623844
rect 338680 623810 338736 623844
rect 338770 623810 338826 623844
rect 338860 623810 338916 623844
rect 338950 623810 339006 623844
rect 339040 623810 339096 623844
rect 339130 623810 339186 623844
rect 339220 623810 339276 623844
rect 339310 623810 339366 623844
rect 339400 623810 339456 623844
rect 339490 623810 339546 623844
rect 339580 623810 339636 623844
rect 339670 623810 339934 623844
rect 339968 623810 340024 623844
rect 340058 623810 340114 623844
rect 340148 623810 340204 623844
rect 340238 623810 340294 623844
rect 340328 623810 340384 623844
rect 340418 623810 340474 623844
rect 340508 623810 340564 623844
rect 340598 623810 340654 623844
rect 340688 623810 340744 623844
rect 340778 623810 340834 623844
rect 340868 623810 340924 623844
rect 340958 623810 341088 623844
rect 334648 623777 341088 623810
rect 334648 623760 334888 623777
rect 334648 623726 334681 623760
rect 334715 623726 334888 623760
rect 334648 623713 334888 623726
rect 335688 623760 336188 623777
rect 335688 623726 335868 623760
rect 335902 623726 335969 623760
rect 336003 623726 336188 623760
rect 335688 623713 336188 623726
rect 336988 623760 337388 623777
rect 336988 623726 337156 623760
rect 337190 623726 337257 623760
rect 337291 623726 337388 623760
rect 336988 623713 337388 623726
rect 338288 623760 338688 623777
rect 338288 623726 338444 623760
rect 338478 623726 338545 623760
rect 338579 623726 338688 623760
rect 338288 623713 338688 623726
rect 339588 623760 339988 623777
rect 339588 623726 339732 623760
rect 339766 623726 339833 623760
rect 339867 623726 339988 623760
rect 339588 623713 339988 623726
rect 340888 623760 341088 623777
rect 340888 623726 341020 623760
rect 341054 623726 341088 623760
rect 340888 623713 341088 623726
rect 334648 623694 341088 623713
rect 334648 623670 334922 623694
rect 334648 623636 334681 623670
rect 334715 623660 334922 623670
rect 334956 623660 335012 623694
rect 335046 623660 335102 623694
rect 335136 623660 335192 623694
rect 335226 623660 335282 623694
rect 335316 623660 335372 623694
rect 335406 623660 335462 623694
rect 335496 623660 335552 623694
rect 335586 623660 335642 623694
rect 335676 623670 336210 623694
rect 335676 623660 335868 623670
rect 334715 623641 335868 623660
rect 334715 623636 334888 623641
rect 334648 623600 334888 623636
rect 334648 623580 334830 623600
rect 334648 623546 334681 623580
rect 334715 623566 334830 623580
rect 334864 623566 334888 623600
rect 335688 623636 335868 623641
rect 335902 623636 335969 623670
rect 336003 623660 336210 623670
rect 336244 623660 336300 623694
rect 336334 623660 336390 623694
rect 336424 623660 336480 623694
rect 336514 623660 336570 623694
rect 336604 623660 336660 623694
rect 336694 623660 336750 623694
rect 336784 623660 336840 623694
rect 336874 623660 336930 623694
rect 336964 623670 337498 623694
rect 336964 623660 337156 623670
rect 336003 623641 337156 623660
rect 336003 623636 336188 623641
rect 335688 623600 336188 623636
rect 335688 623581 336118 623600
rect 334715 623546 334888 623566
rect 334648 623510 334888 623546
rect 334648 623490 334830 623510
rect 334648 623456 334681 623490
rect 334715 623476 334830 623490
rect 334864 623476 334888 623510
rect 334715 623456 334888 623476
rect 334648 623420 334888 623456
rect 334648 623400 334830 623420
rect 334648 623366 334681 623400
rect 334715 623386 334830 623400
rect 334864 623386 334888 623420
rect 334715 623366 334888 623386
rect 334648 623330 334888 623366
rect 334648 623310 334830 623330
rect 334648 623276 334681 623310
rect 334715 623296 334830 623310
rect 334864 623296 334888 623330
rect 334715 623276 334888 623296
rect 334648 623240 334888 623276
rect 334648 623220 334830 623240
rect 334648 623186 334681 623220
rect 334715 623206 334830 623220
rect 334864 623206 334888 623240
rect 334715 623186 334888 623206
rect 334648 623150 334888 623186
rect 334648 623130 334830 623150
rect 334648 623096 334681 623130
rect 334715 623116 334830 623130
rect 334864 623116 334888 623150
rect 334715 623096 334888 623116
rect 334648 623060 334888 623096
rect 334648 623040 334830 623060
rect 334648 623006 334681 623040
rect 334715 623026 334830 623040
rect 334864 623026 334888 623060
rect 334715 623006 334888 623026
rect 334648 622970 334888 623006
rect 334648 622950 334830 622970
rect 334648 622916 334681 622950
rect 334715 622936 334830 622950
rect 334864 622936 334888 622970
rect 334715 622916 334888 622936
rect 334648 622880 334888 622916
rect 334945 623518 335639 623579
rect 334945 623484 335004 623518
rect 335038 623506 335094 623518
rect 335066 623484 335094 623506
rect 335128 623506 335184 623518
rect 335128 623484 335132 623506
rect 334945 623472 335032 623484
rect 335066 623472 335132 623484
rect 335166 623484 335184 623506
rect 335218 623506 335274 623518
rect 335218 623484 335232 623506
rect 335166 623472 335232 623484
rect 335266 623484 335274 623506
rect 335308 623506 335364 623518
rect 335398 623506 335454 623518
rect 335488 623506 335544 623518
rect 335308 623484 335332 623506
rect 335398 623484 335432 623506
rect 335488 623484 335532 623506
rect 335578 623484 335639 623518
rect 335266 623472 335332 623484
rect 335366 623472 335432 623484
rect 335466 623472 335532 623484
rect 335566 623472 335639 623484
rect 334945 623428 335639 623472
rect 334945 623394 335004 623428
rect 335038 623406 335094 623428
rect 335066 623394 335094 623406
rect 335128 623406 335184 623428
rect 335128 623394 335132 623406
rect 334945 623372 335032 623394
rect 335066 623372 335132 623394
rect 335166 623394 335184 623406
rect 335218 623406 335274 623428
rect 335218 623394 335232 623406
rect 335166 623372 335232 623394
rect 335266 623394 335274 623406
rect 335308 623406 335364 623428
rect 335398 623406 335454 623428
rect 335488 623406 335544 623428
rect 335308 623394 335332 623406
rect 335398 623394 335432 623406
rect 335488 623394 335532 623406
rect 335578 623394 335639 623428
rect 335266 623372 335332 623394
rect 335366 623372 335432 623394
rect 335466 623372 335532 623394
rect 335566 623372 335639 623394
rect 334945 623338 335639 623372
rect 334945 623304 335004 623338
rect 335038 623306 335094 623338
rect 335066 623304 335094 623306
rect 335128 623306 335184 623338
rect 335128 623304 335132 623306
rect 334945 623272 335032 623304
rect 335066 623272 335132 623304
rect 335166 623304 335184 623306
rect 335218 623306 335274 623338
rect 335218 623304 335232 623306
rect 335166 623272 335232 623304
rect 335266 623304 335274 623306
rect 335308 623306 335364 623338
rect 335398 623306 335454 623338
rect 335488 623306 335544 623338
rect 335308 623304 335332 623306
rect 335398 623304 335432 623306
rect 335488 623304 335532 623306
rect 335578 623304 335639 623338
rect 335266 623272 335332 623304
rect 335366 623272 335432 623304
rect 335466 623272 335532 623304
rect 335566 623272 335639 623304
rect 334945 623248 335639 623272
rect 334945 623214 335004 623248
rect 335038 623214 335094 623248
rect 335128 623214 335184 623248
rect 335218 623214 335274 623248
rect 335308 623214 335364 623248
rect 335398 623214 335454 623248
rect 335488 623214 335544 623248
rect 335578 623214 335639 623248
rect 334945 623206 335639 623214
rect 334945 623172 335032 623206
rect 335066 623172 335132 623206
rect 335166 623172 335232 623206
rect 335266 623172 335332 623206
rect 335366 623172 335432 623206
rect 335466 623172 335532 623206
rect 335566 623172 335639 623206
rect 334945 623158 335639 623172
rect 334945 623124 335004 623158
rect 335038 623124 335094 623158
rect 335128 623124 335184 623158
rect 335218 623124 335274 623158
rect 335308 623124 335364 623158
rect 335398 623124 335454 623158
rect 335488 623124 335544 623158
rect 335578 623124 335639 623158
rect 334945 623106 335639 623124
rect 334945 623072 335032 623106
rect 335066 623072 335132 623106
rect 335166 623072 335232 623106
rect 335266 623072 335332 623106
rect 335366 623072 335432 623106
rect 335466 623072 335532 623106
rect 335566 623072 335639 623106
rect 334945 623068 335639 623072
rect 334945 623034 335004 623068
rect 335038 623034 335094 623068
rect 335128 623034 335184 623068
rect 335218 623034 335274 623068
rect 335308 623034 335364 623068
rect 335398 623034 335454 623068
rect 335488 623034 335544 623068
rect 335578 623034 335639 623068
rect 334945 623006 335639 623034
rect 334945 622978 335032 623006
rect 335066 622978 335132 623006
rect 334945 622944 335004 622978
rect 335066 622972 335094 622978
rect 335038 622944 335094 622972
rect 335128 622972 335132 622978
rect 335166 622978 335232 623006
rect 335166 622972 335184 622978
rect 335128 622944 335184 622972
rect 335218 622972 335232 622978
rect 335266 622978 335332 623006
rect 335366 622978 335432 623006
rect 335466 622978 335532 623006
rect 335566 622978 335639 623006
rect 335266 622972 335274 622978
rect 335218 622944 335274 622972
rect 335308 622972 335332 622978
rect 335398 622972 335432 622978
rect 335488 622972 335532 622978
rect 335308 622944 335364 622972
rect 335398 622944 335454 622972
rect 335488 622944 335544 622972
rect 335578 622944 335639 622978
rect 334945 622885 335639 622944
rect 335688 623547 335720 623581
rect 335754 623580 336118 623581
rect 335754 623547 335868 623580
rect 335688 623546 335868 623547
rect 335902 623546 335969 623580
rect 336003 623566 336118 623580
rect 336152 623566 336188 623600
rect 336988 623636 337156 623641
rect 337190 623636 337257 623670
rect 337291 623660 337498 623670
rect 337532 623660 337588 623694
rect 337622 623660 337678 623694
rect 337712 623660 337768 623694
rect 337802 623660 337858 623694
rect 337892 623660 337948 623694
rect 337982 623660 338038 623694
rect 338072 623660 338128 623694
rect 338162 623660 338218 623694
rect 338252 623670 338786 623694
rect 338252 623660 338444 623670
rect 337291 623641 338444 623660
rect 337291 623636 337459 623641
rect 336988 623600 337459 623636
rect 336988 623581 337406 623600
rect 336003 623546 336188 623566
rect 335688 623510 336188 623546
rect 335688 623491 336118 623510
rect 335688 623457 335720 623491
rect 335754 623490 336118 623491
rect 335754 623457 335868 623490
rect 335688 623456 335868 623457
rect 335902 623456 335969 623490
rect 336003 623476 336118 623490
rect 336152 623476 336188 623510
rect 336003 623456 336188 623476
rect 335688 623420 336188 623456
rect 335688 623401 336118 623420
rect 335688 623367 335720 623401
rect 335754 623400 336118 623401
rect 335754 623367 335868 623400
rect 335688 623366 335868 623367
rect 335902 623366 335969 623400
rect 336003 623386 336118 623400
rect 336152 623386 336188 623420
rect 336003 623366 336188 623386
rect 335688 623330 336188 623366
rect 335688 623311 336118 623330
rect 335688 623277 335720 623311
rect 335754 623310 336118 623311
rect 335754 623277 335868 623310
rect 335688 623276 335868 623277
rect 335902 623276 335969 623310
rect 336003 623296 336118 623310
rect 336152 623296 336188 623330
rect 336003 623276 336188 623296
rect 335688 623240 336188 623276
rect 335688 623221 336118 623240
rect 335688 623187 335720 623221
rect 335754 623220 336118 623221
rect 335754 623187 335868 623220
rect 335688 623186 335868 623187
rect 335902 623186 335969 623220
rect 336003 623206 336118 623220
rect 336152 623206 336188 623240
rect 336003 623186 336188 623206
rect 335688 623150 336188 623186
rect 335688 623131 336118 623150
rect 335688 623097 335720 623131
rect 335754 623130 336118 623131
rect 335754 623097 335868 623130
rect 335688 623096 335868 623097
rect 335902 623096 335969 623130
rect 336003 623116 336118 623130
rect 336152 623116 336188 623150
rect 336003 623096 336188 623116
rect 335688 623060 336188 623096
rect 335688 623041 336118 623060
rect 335688 623007 335720 623041
rect 335754 623040 336118 623041
rect 335754 623007 335868 623040
rect 335688 623006 335868 623007
rect 335902 623006 335969 623040
rect 336003 623026 336118 623040
rect 336152 623026 336188 623060
rect 336003 623006 336188 623026
rect 335688 622970 336188 623006
rect 335688 622951 336118 622970
rect 335688 622917 335720 622951
rect 335754 622950 336118 622951
rect 335754 622917 335868 622950
rect 335688 622916 335868 622917
rect 335902 622916 335969 622950
rect 336003 622936 336118 622950
rect 336152 622936 336188 622970
rect 336003 622916 336188 622936
rect 334648 622860 334830 622880
rect 334648 622826 334681 622860
rect 334715 622846 334830 622860
rect 334864 622846 334888 622880
rect 334715 622826 334888 622846
rect 334648 622823 334888 622826
rect 335688 622880 336188 622916
rect 336233 623518 336927 623579
rect 336233 623484 336292 623518
rect 336326 623506 336382 623518
rect 336354 623484 336382 623506
rect 336416 623506 336472 623518
rect 336416 623484 336420 623506
rect 336233 623472 336320 623484
rect 336354 623472 336420 623484
rect 336454 623484 336472 623506
rect 336506 623506 336562 623518
rect 336506 623484 336520 623506
rect 336454 623472 336520 623484
rect 336554 623484 336562 623506
rect 336596 623506 336652 623518
rect 336686 623506 336742 623518
rect 336776 623506 336832 623518
rect 336596 623484 336620 623506
rect 336686 623484 336720 623506
rect 336776 623484 336820 623506
rect 336866 623484 336927 623518
rect 336554 623472 336620 623484
rect 336654 623472 336720 623484
rect 336754 623472 336820 623484
rect 336854 623472 336927 623484
rect 336233 623428 336927 623472
rect 336233 623394 336292 623428
rect 336326 623406 336382 623428
rect 336354 623394 336382 623406
rect 336416 623406 336472 623428
rect 336416 623394 336420 623406
rect 336233 623372 336320 623394
rect 336354 623372 336420 623394
rect 336454 623394 336472 623406
rect 336506 623406 336562 623428
rect 336506 623394 336520 623406
rect 336454 623372 336520 623394
rect 336554 623394 336562 623406
rect 336596 623406 336652 623428
rect 336686 623406 336742 623428
rect 336776 623406 336832 623428
rect 336596 623394 336620 623406
rect 336686 623394 336720 623406
rect 336776 623394 336820 623406
rect 336866 623394 336927 623428
rect 336554 623372 336620 623394
rect 336654 623372 336720 623394
rect 336754 623372 336820 623394
rect 336854 623372 336927 623394
rect 336233 623338 336927 623372
rect 336233 623304 336292 623338
rect 336326 623306 336382 623338
rect 336354 623304 336382 623306
rect 336416 623306 336472 623338
rect 336416 623304 336420 623306
rect 336233 623272 336320 623304
rect 336354 623272 336420 623304
rect 336454 623304 336472 623306
rect 336506 623306 336562 623338
rect 336506 623304 336520 623306
rect 336454 623272 336520 623304
rect 336554 623304 336562 623306
rect 336596 623306 336652 623338
rect 336686 623306 336742 623338
rect 336776 623306 336832 623338
rect 336596 623304 336620 623306
rect 336686 623304 336720 623306
rect 336776 623304 336820 623306
rect 336866 623304 336927 623338
rect 336554 623272 336620 623304
rect 336654 623272 336720 623304
rect 336754 623272 336820 623304
rect 336854 623272 336927 623304
rect 336233 623248 336927 623272
rect 336233 623214 336292 623248
rect 336326 623214 336382 623248
rect 336416 623214 336472 623248
rect 336506 623214 336562 623248
rect 336596 623214 336652 623248
rect 336686 623214 336742 623248
rect 336776 623214 336832 623248
rect 336866 623214 336927 623248
rect 336233 623206 336927 623214
rect 336233 623172 336320 623206
rect 336354 623172 336420 623206
rect 336454 623172 336520 623206
rect 336554 623172 336620 623206
rect 336654 623172 336720 623206
rect 336754 623172 336820 623206
rect 336854 623172 336927 623206
rect 336233 623158 336927 623172
rect 336233 623124 336292 623158
rect 336326 623124 336382 623158
rect 336416 623124 336472 623158
rect 336506 623124 336562 623158
rect 336596 623124 336652 623158
rect 336686 623124 336742 623158
rect 336776 623124 336832 623158
rect 336866 623124 336927 623158
rect 336233 623106 336927 623124
rect 336233 623072 336320 623106
rect 336354 623072 336420 623106
rect 336454 623072 336520 623106
rect 336554 623072 336620 623106
rect 336654 623072 336720 623106
rect 336754 623072 336820 623106
rect 336854 623072 336927 623106
rect 336233 623068 336927 623072
rect 336233 623034 336292 623068
rect 336326 623034 336382 623068
rect 336416 623034 336472 623068
rect 336506 623034 336562 623068
rect 336596 623034 336652 623068
rect 336686 623034 336742 623068
rect 336776 623034 336832 623068
rect 336866 623034 336927 623068
rect 336233 623006 336927 623034
rect 336233 622978 336320 623006
rect 336354 622978 336420 623006
rect 336233 622944 336292 622978
rect 336354 622972 336382 622978
rect 336326 622944 336382 622972
rect 336416 622972 336420 622978
rect 336454 622978 336520 623006
rect 336454 622972 336472 622978
rect 336416 622944 336472 622972
rect 336506 622972 336520 622978
rect 336554 622978 336620 623006
rect 336654 622978 336720 623006
rect 336754 622978 336820 623006
rect 336854 622978 336927 623006
rect 336554 622972 336562 622978
rect 336506 622944 336562 622972
rect 336596 622972 336620 622978
rect 336686 622972 336720 622978
rect 336776 622972 336820 622978
rect 336596 622944 336652 622972
rect 336686 622944 336742 622972
rect 336776 622944 336832 622972
rect 336866 622944 336927 622978
rect 336233 622885 336927 622944
rect 336988 623547 337008 623581
rect 337042 623580 337406 623581
rect 337042 623547 337156 623580
rect 336988 623546 337156 623547
rect 337190 623546 337257 623580
rect 337291 623566 337406 623580
rect 337440 623566 337459 623600
rect 338277 623636 338444 623641
rect 338478 623636 338545 623670
rect 338579 623660 338786 623670
rect 338820 623660 338876 623694
rect 338910 623660 338966 623694
rect 339000 623660 339056 623694
rect 339090 623660 339146 623694
rect 339180 623660 339236 623694
rect 339270 623660 339326 623694
rect 339360 623660 339416 623694
rect 339450 623660 339506 623694
rect 339540 623670 340074 623694
rect 339540 623660 339732 623670
rect 338579 623641 339732 623660
rect 338579 623636 338747 623641
rect 338277 623600 338747 623636
rect 338277 623581 338694 623600
rect 337291 623546 337459 623566
rect 336988 623510 337459 623546
rect 336988 623491 337406 623510
rect 336988 623457 337008 623491
rect 337042 623490 337406 623491
rect 337042 623457 337156 623490
rect 336988 623456 337156 623457
rect 337190 623456 337257 623490
rect 337291 623476 337406 623490
rect 337440 623476 337459 623510
rect 337291 623456 337459 623476
rect 336988 623420 337459 623456
rect 336988 623401 337406 623420
rect 336988 623367 337008 623401
rect 337042 623400 337406 623401
rect 337042 623367 337156 623400
rect 336988 623366 337156 623367
rect 337190 623366 337257 623400
rect 337291 623386 337406 623400
rect 337440 623386 337459 623420
rect 337291 623366 337459 623386
rect 336988 623330 337459 623366
rect 336988 623311 337406 623330
rect 336988 623277 337008 623311
rect 337042 623310 337406 623311
rect 337042 623277 337156 623310
rect 336988 623276 337156 623277
rect 337190 623276 337257 623310
rect 337291 623296 337406 623310
rect 337440 623296 337459 623330
rect 337291 623276 337459 623296
rect 336988 623240 337459 623276
rect 336988 623221 337406 623240
rect 336988 623187 337008 623221
rect 337042 623220 337406 623221
rect 337042 623187 337156 623220
rect 336988 623186 337156 623187
rect 337190 623186 337257 623220
rect 337291 623206 337406 623220
rect 337440 623206 337459 623240
rect 337291 623186 337459 623206
rect 336988 623150 337459 623186
rect 336988 623131 337406 623150
rect 336988 623097 337008 623131
rect 337042 623130 337406 623131
rect 337042 623097 337156 623130
rect 336988 623096 337156 623097
rect 337190 623096 337257 623130
rect 337291 623116 337406 623130
rect 337440 623116 337459 623150
rect 337291 623096 337459 623116
rect 336988 623060 337459 623096
rect 336988 623041 337406 623060
rect 336988 623007 337008 623041
rect 337042 623040 337406 623041
rect 337042 623007 337156 623040
rect 336988 623006 337156 623007
rect 337190 623006 337257 623040
rect 337291 623026 337406 623040
rect 337440 623026 337459 623060
rect 337291 623006 337459 623026
rect 336988 622970 337459 623006
rect 336988 622951 337406 622970
rect 336988 622917 337008 622951
rect 337042 622950 337406 622951
rect 337042 622917 337156 622950
rect 336988 622916 337156 622917
rect 337190 622916 337257 622950
rect 337291 622936 337406 622950
rect 337440 622936 337459 622970
rect 337291 622916 337459 622936
rect 335688 622861 336118 622880
rect 335688 622827 335720 622861
rect 335754 622860 336118 622861
rect 335754 622827 335868 622860
rect 335688 622826 335868 622827
rect 335902 622826 335969 622860
rect 336003 622846 336118 622860
rect 336152 622846 336188 622880
rect 336003 622826 336188 622846
rect 335688 622823 336188 622826
rect 336988 622880 337459 622916
rect 337521 623518 338215 623579
rect 337521 623484 337580 623518
rect 337614 623506 337670 623518
rect 337642 623484 337670 623506
rect 337704 623506 337760 623518
rect 337704 623484 337708 623506
rect 337521 623472 337608 623484
rect 337642 623472 337708 623484
rect 337742 623484 337760 623506
rect 337794 623506 337850 623518
rect 337794 623484 337808 623506
rect 337742 623472 337808 623484
rect 337842 623484 337850 623506
rect 337884 623506 337940 623518
rect 337974 623506 338030 623518
rect 338064 623506 338120 623518
rect 337884 623484 337908 623506
rect 337974 623484 338008 623506
rect 338064 623484 338108 623506
rect 338154 623484 338215 623518
rect 337842 623472 337908 623484
rect 337942 623472 338008 623484
rect 338042 623472 338108 623484
rect 338142 623472 338215 623484
rect 337521 623428 338215 623472
rect 337521 623394 337580 623428
rect 337614 623406 337670 623428
rect 337642 623394 337670 623406
rect 337704 623406 337760 623428
rect 337704 623394 337708 623406
rect 337521 623372 337608 623394
rect 337642 623372 337708 623394
rect 337742 623394 337760 623406
rect 337794 623406 337850 623428
rect 337794 623394 337808 623406
rect 337742 623372 337808 623394
rect 337842 623394 337850 623406
rect 337884 623406 337940 623428
rect 337974 623406 338030 623428
rect 338064 623406 338120 623428
rect 337884 623394 337908 623406
rect 337974 623394 338008 623406
rect 338064 623394 338108 623406
rect 338154 623394 338215 623428
rect 337842 623372 337908 623394
rect 337942 623372 338008 623394
rect 338042 623372 338108 623394
rect 338142 623372 338215 623394
rect 337521 623338 338215 623372
rect 337521 623304 337580 623338
rect 337614 623306 337670 623338
rect 337642 623304 337670 623306
rect 337704 623306 337760 623338
rect 337704 623304 337708 623306
rect 337521 623272 337608 623304
rect 337642 623272 337708 623304
rect 337742 623304 337760 623306
rect 337794 623306 337850 623338
rect 337794 623304 337808 623306
rect 337742 623272 337808 623304
rect 337842 623304 337850 623306
rect 337884 623306 337940 623338
rect 337974 623306 338030 623338
rect 338064 623306 338120 623338
rect 337884 623304 337908 623306
rect 337974 623304 338008 623306
rect 338064 623304 338108 623306
rect 338154 623304 338215 623338
rect 337842 623272 337908 623304
rect 337942 623272 338008 623304
rect 338042 623272 338108 623304
rect 338142 623272 338215 623304
rect 337521 623248 338215 623272
rect 337521 623214 337580 623248
rect 337614 623214 337670 623248
rect 337704 623214 337760 623248
rect 337794 623214 337850 623248
rect 337884 623214 337940 623248
rect 337974 623214 338030 623248
rect 338064 623214 338120 623248
rect 338154 623214 338215 623248
rect 337521 623206 338215 623214
rect 337521 623172 337608 623206
rect 337642 623172 337708 623206
rect 337742 623172 337808 623206
rect 337842 623172 337908 623206
rect 337942 623172 338008 623206
rect 338042 623172 338108 623206
rect 338142 623172 338215 623206
rect 337521 623158 338215 623172
rect 337521 623124 337580 623158
rect 337614 623124 337670 623158
rect 337704 623124 337760 623158
rect 337794 623124 337850 623158
rect 337884 623124 337940 623158
rect 337974 623124 338030 623158
rect 338064 623124 338120 623158
rect 338154 623124 338215 623158
rect 337521 623106 338215 623124
rect 337521 623072 337608 623106
rect 337642 623072 337708 623106
rect 337742 623072 337808 623106
rect 337842 623072 337908 623106
rect 337942 623072 338008 623106
rect 338042 623072 338108 623106
rect 338142 623072 338215 623106
rect 337521 623068 338215 623072
rect 337521 623034 337580 623068
rect 337614 623034 337670 623068
rect 337704 623034 337760 623068
rect 337794 623034 337850 623068
rect 337884 623034 337940 623068
rect 337974 623034 338030 623068
rect 338064 623034 338120 623068
rect 338154 623034 338215 623068
rect 337521 623006 338215 623034
rect 337521 622978 337608 623006
rect 337642 622978 337708 623006
rect 337521 622944 337580 622978
rect 337642 622972 337670 622978
rect 337614 622944 337670 622972
rect 337704 622972 337708 622978
rect 337742 622978 337808 623006
rect 337742 622972 337760 622978
rect 337704 622944 337760 622972
rect 337794 622972 337808 622978
rect 337842 622978 337908 623006
rect 337942 622978 338008 623006
rect 338042 622978 338108 623006
rect 338142 622978 338215 623006
rect 337842 622972 337850 622978
rect 337794 622944 337850 622972
rect 337884 622972 337908 622978
rect 337974 622972 338008 622978
rect 338064 622972 338108 622978
rect 337884 622944 337940 622972
rect 337974 622944 338030 622972
rect 338064 622944 338120 622972
rect 338154 622944 338215 622978
rect 337521 622885 338215 622944
rect 338277 623547 338296 623581
rect 338330 623580 338694 623581
rect 338330 623547 338444 623580
rect 338277 623546 338444 623547
rect 338478 623546 338545 623580
rect 338579 623566 338694 623580
rect 338728 623566 338747 623600
rect 339565 623636 339732 623641
rect 339766 623636 339833 623670
rect 339867 623660 340074 623670
rect 340108 623660 340164 623694
rect 340198 623660 340254 623694
rect 340288 623660 340344 623694
rect 340378 623660 340434 623694
rect 340468 623660 340524 623694
rect 340558 623660 340614 623694
rect 340648 623660 340704 623694
rect 340738 623660 340794 623694
rect 340828 623670 341088 623694
rect 340828 623660 341020 623670
rect 339867 623641 341020 623660
rect 339867 623636 340035 623641
rect 339565 623600 340035 623636
rect 339565 623581 339982 623600
rect 338579 623546 338747 623566
rect 338277 623510 338747 623546
rect 338277 623491 338694 623510
rect 338277 623457 338296 623491
rect 338330 623490 338694 623491
rect 338330 623457 338444 623490
rect 338277 623456 338444 623457
rect 338478 623456 338545 623490
rect 338579 623476 338694 623490
rect 338728 623476 338747 623510
rect 338579 623456 338747 623476
rect 338277 623420 338747 623456
rect 338277 623401 338694 623420
rect 338277 623367 338296 623401
rect 338330 623400 338694 623401
rect 338330 623367 338444 623400
rect 338277 623366 338444 623367
rect 338478 623366 338545 623400
rect 338579 623386 338694 623400
rect 338728 623386 338747 623420
rect 338579 623366 338747 623386
rect 338277 623330 338747 623366
rect 338277 623311 338694 623330
rect 338277 623277 338296 623311
rect 338330 623310 338694 623311
rect 338330 623277 338444 623310
rect 338277 623276 338444 623277
rect 338478 623276 338545 623310
rect 338579 623296 338694 623310
rect 338728 623296 338747 623330
rect 338579 623276 338747 623296
rect 338277 623240 338747 623276
rect 338277 623221 338694 623240
rect 338277 623187 338296 623221
rect 338330 623220 338694 623221
rect 338330 623187 338444 623220
rect 338277 623186 338444 623187
rect 338478 623186 338545 623220
rect 338579 623206 338694 623220
rect 338728 623206 338747 623240
rect 338579 623186 338747 623206
rect 338277 623150 338747 623186
rect 338277 623131 338694 623150
rect 338277 623097 338296 623131
rect 338330 623130 338694 623131
rect 338330 623097 338444 623130
rect 338277 623096 338444 623097
rect 338478 623096 338545 623130
rect 338579 623116 338694 623130
rect 338728 623116 338747 623150
rect 338579 623096 338747 623116
rect 338277 623060 338747 623096
rect 338277 623041 338694 623060
rect 338277 623007 338296 623041
rect 338330 623040 338694 623041
rect 338330 623007 338444 623040
rect 338277 623006 338444 623007
rect 338478 623006 338545 623040
rect 338579 623026 338694 623040
rect 338728 623026 338747 623060
rect 338579 623006 338747 623026
rect 338277 622970 338747 623006
rect 338277 622951 338694 622970
rect 338277 622917 338296 622951
rect 338330 622950 338694 622951
rect 338330 622917 338444 622950
rect 338277 622916 338444 622917
rect 338478 622916 338545 622950
rect 338579 622936 338694 622950
rect 338728 622936 338747 622970
rect 338579 622916 338747 622936
rect 336988 622861 337406 622880
rect 336988 622827 337008 622861
rect 337042 622860 337406 622861
rect 337042 622827 337156 622860
rect 336988 622826 337156 622827
rect 337190 622826 337257 622860
rect 337291 622846 337406 622860
rect 337440 622846 337459 622880
rect 337291 622826 337459 622846
rect 336988 622823 337459 622826
rect 338277 622880 338747 622916
rect 338809 623518 339503 623579
rect 338809 623484 338868 623518
rect 338902 623506 338958 623518
rect 338930 623484 338958 623506
rect 338992 623506 339048 623518
rect 338992 623484 338996 623506
rect 338809 623472 338896 623484
rect 338930 623472 338996 623484
rect 339030 623484 339048 623506
rect 339082 623506 339138 623518
rect 339082 623484 339096 623506
rect 339030 623472 339096 623484
rect 339130 623484 339138 623506
rect 339172 623506 339228 623518
rect 339262 623506 339318 623518
rect 339352 623506 339408 623518
rect 339172 623484 339196 623506
rect 339262 623484 339296 623506
rect 339352 623484 339396 623506
rect 339442 623484 339503 623518
rect 339130 623472 339196 623484
rect 339230 623472 339296 623484
rect 339330 623472 339396 623484
rect 339430 623472 339503 623484
rect 338809 623428 339503 623472
rect 338809 623394 338868 623428
rect 338902 623406 338958 623428
rect 338930 623394 338958 623406
rect 338992 623406 339048 623428
rect 338992 623394 338996 623406
rect 338809 623372 338896 623394
rect 338930 623372 338996 623394
rect 339030 623394 339048 623406
rect 339082 623406 339138 623428
rect 339082 623394 339096 623406
rect 339030 623372 339096 623394
rect 339130 623394 339138 623406
rect 339172 623406 339228 623428
rect 339262 623406 339318 623428
rect 339352 623406 339408 623428
rect 339172 623394 339196 623406
rect 339262 623394 339296 623406
rect 339352 623394 339396 623406
rect 339442 623394 339503 623428
rect 339130 623372 339196 623394
rect 339230 623372 339296 623394
rect 339330 623372 339396 623394
rect 339430 623372 339503 623394
rect 338809 623338 339503 623372
rect 338809 623304 338868 623338
rect 338902 623306 338958 623338
rect 338930 623304 338958 623306
rect 338992 623306 339048 623338
rect 338992 623304 338996 623306
rect 338809 623272 338896 623304
rect 338930 623272 338996 623304
rect 339030 623304 339048 623306
rect 339082 623306 339138 623338
rect 339082 623304 339096 623306
rect 339030 623272 339096 623304
rect 339130 623304 339138 623306
rect 339172 623306 339228 623338
rect 339262 623306 339318 623338
rect 339352 623306 339408 623338
rect 339172 623304 339196 623306
rect 339262 623304 339296 623306
rect 339352 623304 339396 623306
rect 339442 623304 339503 623338
rect 339130 623272 339196 623304
rect 339230 623272 339296 623304
rect 339330 623272 339396 623304
rect 339430 623272 339503 623304
rect 338809 623248 339503 623272
rect 338809 623214 338868 623248
rect 338902 623214 338958 623248
rect 338992 623214 339048 623248
rect 339082 623214 339138 623248
rect 339172 623214 339228 623248
rect 339262 623214 339318 623248
rect 339352 623214 339408 623248
rect 339442 623214 339503 623248
rect 338809 623206 339503 623214
rect 338809 623172 338896 623206
rect 338930 623172 338996 623206
rect 339030 623172 339096 623206
rect 339130 623172 339196 623206
rect 339230 623172 339296 623206
rect 339330 623172 339396 623206
rect 339430 623172 339503 623206
rect 338809 623158 339503 623172
rect 338809 623124 338868 623158
rect 338902 623124 338958 623158
rect 338992 623124 339048 623158
rect 339082 623124 339138 623158
rect 339172 623124 339228 623158
rect 339262 623124 339318 623158
rect 339352 623124 339408 623158
rect 339442 623124 339503 623158
rect 338809 623106 339503 623124
rect 338809 623072 338896 623106
rect 338930 623072 338996 623106
rect 339030 623072 339096 623106
rect 339130 623072 339196 623106
rect 339230 623072 339296 623106
rect 339330 623072 339396 623106
rect 339430 623072 339503 623106
rect 338809 623068 339503 623072
rect 338809 623034 338868 623068
rect 338902 623034 338958 623068
rect 338992 623034 339048 623068
rect 339082 623034 339138 623068
rect 339172 623034 339228 623068
rect 339262 623034 339318 623068
rect 339352 623034 339408 623068
rect 339442 623034 339503 623068
rect 338809 623006 339503 623034
rect 338809 622978 338896 623006
rect 338930 622978 338996 623006
rect 338809 622944 338868 622978
rect 338930 622972 338958 622978
rect 338902 622944 338958 622972
rect 338992 622972 338996 622978
rect 339030 622978 339096 623006
rect 339030 622972 339048 622978
rect 338992 622944 339048 622972
rect 339082 622972 339096 622978
rect 339130 622978 339196 623006
rect 339230 622978 339296 623006
rect 339330 622978 339396 623006
rect 339430 622978 339503 623006
rect 339130 622972 339138 622978
rect 339082 622944 339138 622972
rect 339172 622972 339196 622978
rect 339262 622972 339296 622978
rect 339352 622972 339396 622978
rect 339172 622944 339228 622972
rect 339262 622944 339318 622972
rect 339352 622944 339408 622972
rect 339442 622944 339503 622978
rect 338809 622885 339503 622944
rect 339565 623547 339584 623581
rect 339618 623580 339982 623581
rect 339618 623547 339732 623580
rect 339565 623546 339732 623547
rect 339766 623546 339833 623580
rect 339867 623566 339982 623580
rect 340016 623566 340035 623600
rect 340853 623636 341020 623641
rect 341054 623636 341088 623670
rect 340853 623581 341088 623636
rect 339867 623546 340035 623566
rect 339565 623510 340035 623546
rect 339565 623491 339982 623510
rect 339565 623457 339584 623491
rect 339618 623490 339982 623491
rect 339618 623457 339732 623490
rect 339565 623456 339732 623457
rect 339766 623456 339833 623490
rect 339867 623476 339982 623490
rect 340016 623476 340035 623510
rect 339867 623456 340035 623476
rect 339565 623420 340035 623456
rect 339565 623401 339982 623420
rect 339565 623367 339584 623401
rect 339618 623400 339982 623401
rect 339618 623367 339732 623400
rect 339565 623366 339732 623367
rect 339766 623366 339833 623400
rect 339867 623386 339982 623400
rect 340016 623386 340035 623420
rect 339867 623366 340035 623386
rect 339565 623330 340035 623366
rect 339565 623311 339982 623330
rect 339565 623277 339584 623311
rect 339618 623310 339982 623311
rect 339618 623277 339732 623310
rect 339565 623276 339732 623277
rect 339766 623276 339833 623310
rect 339867 623296 339982 623310
rect 340016 623296 340035 623330
rect 339867 623276 340035 623296
rect 339565 623240 340035 623276
rect 339565 623221 339982 623240
rect 339565 623187 339584 623221
rect 339618 623220 339982 623221
rect 339618 623187 339732 623220
rect 339565 623186 339732 623187
rect 339766 623186 339833 623220
rect 339867 623206 339982 623220
rect 340016 623206 340035 623240
rect 339867 623186 340035 623206
rect 339565 623150 340035 623186
rect 339565 623131 339982 623150
rect 339565 623097 339584 623131
rect 339618 623130 339982 623131
rect 339618 623097 339732 623130
rect 339565 623096 339732 623097
rect 339766 623096 339833 623130
rect 339867 623116 339982 623130
rect 340016 623116 340035 623150
rect 339867 623096 340035 623116
rect 339565 623060 340035 623096
rect 339565 623041 339982 623060
rect 339565 623007 339584 623041
rect 339618 623040 339982 623041
rect 339618 623007 339732 623040
rect 339565 623006 339732 623007
rect 339766 623006 339833 623040
rect 339867 623026 339982 623040
rect 340016 623026 340035 623060
rect 339867 623006 340035 623026
rect 339565 622970 340035 623006
rect 339565 622951 339982 622970
rect 339565 622917 339584 622951
rect 339618 622950 339982 622951
rect 339618 622917 339732 622950
rect 339565 622916 339732 622917
rect 339766 622916 339833 622950
rect 339867 622936 339982 622950
rect 340016 622936 340035 622970
rect 339867 622916 340035 622936
rect 338277 622861 338694 622880
rect 338277 622827 338296 622861
rect 338330 622860 338694 622861
rect 338330 622827 338444 622860
rect 338277 622826 338444 622827
rect 338478 622826 338545 622860
rect 338579 622846 338694 622860
rect 338728 622846 338747 622880
rect 338579 622826 338747 622846
rect 338277 622823 338747 622826
rect 339565 622880 340035 622916
rect 340097 623518 340791 623579
rect 340097 623484 340156 623518
rect 340190 623506 340246 623518
rect 340218 623484 340246 623506
rect 340280 623506 340336 623518
rect 340280 623484 340284 623506
rect 340097 623472 340184 623484
rect 340218 623472 340284 623484
rect 340318 623484 340336 623506
rect 340370 623506 340426 623518
rect 340370 623484 340384 623506
rect 340318 623472 340384 623484
rect 340418 623484 340426 623506
rect 340460 623506 340516 623518
rect 340550 623506 340606 623518
rect 340640 623506 340696 623518
rect 340460 623484 340484 623506
rect 340550 623484 340584 623506
rect 340640 623484 340684 623506
rect 340730 623484 340791 623518
rect 340418 623472 340484 623484
rect 340518 623472 340584 623484
rect 340618 623472 340684 623484
rect 340718 623472 340791 623484
rect 340097 623428 340791 623472
rect 340097 623394 340156 623428
rect 340190 623406 340246 623428
rect 340218 623394 340246 623406
rect 340280 623406 340336 623428
rect 340280 623394 340284 623406
rect 340097 623372 340184 623394
rect 340218 623372 340284 623394
rect 340318 623394 340336 623406
rect 340370 623406 340426 623428
rect 340370 623394 340384 623406
rect 340318 623372 340384 623394
rect 340418 623394 340426 623406
rect 340460 623406 340516 623428
rect 340550 623406 340606 623428
rect 340640 623406 340696 623428
rect 340460 623394 340484 623406
rect 340550 623394 340584 623406
rect 340640 623394 340684 623406
rect 340730 623394 340791 623428
rect 340418 623372 340484 623394
rect 340518 623372 340584 623394
rect 340618 623372 340684 623394
rect 340718 623372 340791 623394
rect 340097 623338 340791 623372
rect 340097 623304 340156 623338
rect 340190 623306 340246 623338
rect 340218 623304 340246 623306
rect 340280 623306 340336 623338
rect 340280 623304 340284 623306
rect 340097 623272 340184 623304
rect 340218 623272 340284 623304
rect 340318 623304 340336 623306
rect 340370 623306 340426 623338
rect 340370 623304 340384 623306
rect 340318 623272 340384 623304
rect 340418 623304 340426 623306
rect 340460 623306 340516 623338
rect 340550 623306 340606 623338
rect 340640 623306 340696 623338
rect 340460 623304 340484 623306
rect 340550 623304 340584 623306
rect 340640 623304 340684 623306
rect 340730 623304 340791 623338
rect 340418 623272 340484 623304
rect 340518 623272 340584 623304
rect 340618 623272 340684 623304
rect 340718 623272 340791 623304
rect 340097 623248 340791 623272
rect 340097 623214 340156 623248
rect 340190 623214 340246 623248
rect 340280 623214 340336 623248
rect 340370 623214 340426 623248
rect 340460 623214 340516 623248
rect 340550 623214 340606 623248
rect 340640 623214 340696 623248
rect 340730 623214 340791 623248
rect 340097 623206 340791 623214
rect 340097 623172 340184 623206
rect 340218 623172 340284 623206
rect 340318 623172 340384 623206
rect 340418 623172 340484 623206
rect 340518 623172 340584 623206
rect 340618 623172 340684 623206
rect 340718 623172 340791 623206
rect 340097 623158 340791 623172
rect 340097 623124 340156 623158
rect 340190 623124 340246 623158
rect 340280 623124 340336 623158
rect 340370 623124 340426 623158
rect 340460 623124 340516 623158
rect 340550 623124 340606 623158
rect 340640 623124 340696 623158
rect 340730 623124 340791 623158
rect 340097 623106 340791 623124
rect 340097 623072 340184 623106
rect 340218 623072 340284 623106
rect 340318 623072 340384 623106
rect 340418 623072 340484 623106
rect 340518 623072 340584 623106
rect 340618 623072 340684 623106
rect 340718 623072 340791 623106
rect 340097 623068 340791 623072
rect 340097 623034 340156 623068
rect 340190 623034 340246 623068
rect 340280 623034 340336 623068
rect 340370 623034 340426 623068
rect 340460 623034 340516 623068
rect 340550 623034 340606 623068
rect 340640 623034 340696 623068
rect 340730 623034 340791 623068
rect 340097 623006 340791 623034
rect 340097 622978 340184 623006
rect 340218 622978 340284 623006
rect 340097 622944 340156 622978
rect 340218 622972 340246 622978
rect 340190 622944 340246 622972
rect 340280 622972 340284 622978
rect 340318 622978 340384 623006
rect 340318 622972 340336 622978
rect 340280 622944 340336 622972
rect 340370 622972 340384 622978
rect 340418 622978 340484 623006
rect 340518 622978 340584 623006
rect 340618 622978 340684 623006
rect 340718 622978 340791 623006
rect 340418 622972 340426 622978
rect 340370 622944 340426 622972
rect 340460 622972 340484 622978
rect 340550 622972 340584 622978
rect 340640 622972 340684 622978
rect 340460 622944 340516 622972
rect 340550 622944 340606 622972
rect 340640 622944 340696 622972
rect 340730 622944 340791 622978
rect 340097 622885 340791 622944
rect 340853 623547 340872 623581
rect 340906 623580 341088 623581
rect 340906 623547 341020 623580
rect 340853 623546 341020 623547
rect 341054 623546 341088 623580
rect 340853 623491 341088 623546
rect 340853 623457 340872 623491
rect 340906 623490 341088 623491
rect 340906 623457 341020 623490
rect 340853 623456 341020 623457
rect 341054 623456 341088 623490
rect 340853 623401 341088 623456
rect 340853 623367 340872 623401
rect 340906 623400 341088 623401
rect 340906 623367 341020 623400
rect 340853 623366 341020 623367
rect 341054 623366 341088 623400
rect 340853 623311 341088 623366
rect 340853 623277 340872 623311
rect 340906 623310 341088 623311
rect 340906 623277 341020 623310
rect 340853 623276 341020 623277
rect 341054 623276 341088 623310
rect 340853 623221 341088 623276
rect 340853 623187 340872 623221
rect 340906 623220 341088 623221
rect 340906 623187 341020 623220
rect 340853 623186 341020 623187
rect 341054 623186 341088 623220
rect 340853 623131 341088 623186
rect 340853 623097 340872 623131
rect 340906 623130 341088 623131
rect 340906 623097 341020 623130
rect 340853 623096 341020 623097
rect 341054 623096 341088 623130
rect 340853 623041 341088 623096
rect 340853 623007 340872 623041
rect 340906 623040 341088 623041
rect 340906 623007 341020 623040
rect 340853 623006 341020 623007
rect 341054 623006 341088 623040
rect 340853 622951 341088 623006
rect 340853 622917 340872 622951
rect 340906 622950 341088 622951
rect 340906 622917 341020 622950
rect 340853 622916 341020 622917
rect 341054 622916 341088 622950
rect 339565 622861 339982 622880
rect 339565 622827 339584 622861
rect 339618 622860 339982 622861
rect 339618 622827 339732 622860
rect 339565 622826 339732 622827
rect 339766 622826 339833 622860
rect 339867 622846 339982 622860
rect 340016 622846 340035 622880
rect 339867 622826 340035 622846
rect 339565 622823 340035 622826
rect 340853 622861 341088 622916
rect 340853 622827 340872 622861
rect 340906 622860 341088 622861
rect 340906 622827 341020 622860
rect 340853 622826 341020 622827
rect 341054 622826 341088 622860
rect 340853 622823 341088 622826
rect 334648 622804 341088 622823
rect 334648 622770 334888 622804
rect 334922 622770 334978 622804
rect 335012 622770 335068 622804
rect 335102 622770 335158 622804
rect 335192 622770 335248 622804
rect 335282 622770 335338 622804
rect 335372 622770 335428 622804
rect 335462 622770 335518 622804
rect 335552 622770 335608 622804
rect 335642 622770 336176 622804
rect 336210 622770 336266 622804
rect 336300 622770 336356 622804
rect 336390 622770 336446 622804
rect 336480 622770 336536 622804
rect 336570 622770 336626 622804
rect 336660 622770 336716 622804
rect 336750 622770 336806 622804
rect 336840 622770 336896 622804
rect 336930 622770 337464 622804
rect 337498 622770 337554 622804
rect 337588 622770 337644 622804
rect 337678 622770 337734 622804
rect 337768 622770 337824 622804
rect 337858 622770 337914 622804
rect 337948 622770 338004 622804
rect 338038 622770 338094 622804
rect 338128 622770 338184 622804
rect 338218 622770 338752 622804
rect 338786 622770 338842 622804
rect 338876 622770 338932 622804
rect 338966 622770 339022 622804
rect 339056 622770 339112 622804
rect 339146 622770 339202 622804
rect 339236 622770 339292 622804
rect 339326 622770 339382 622804
rect 339416 622770 339472 622804
rect 339506 622770 340040 622804
rect 340074 622770 340130 622804
rect 340164 622770 340220 622804
rect 340254 622770 340310 622804
rect 340344 622770 340400 622804
rect 340434 622770 340490 622804
rect 340524 622770 340580 622804
rect 340614 622770 340670 622804
rect 340704 622770 340760 622804
rect 340794 622770 341088 622804
rect 334648 622736 334681 622770
rect 334715 622751 335868 622770
rect 334715 622736 334888 622751
rect 334648 622687 334888 622736
rect 335688 622736 335868 622751
rect 335902 622736 335969 622770
rect 336003 622751 337156 622770
rect 336003 622736 336188 622751
rect 335688 622687 336188 622736
rect 336988 622736 337156 622751
rect 337190 622736 337257 622770
rect 337291 622751 338444 622770
rect 337291 622736 337388 622751
rect 336988 622687 337388 622736
rect 338288 622736 338444 622751
rect 338478 622736 338545 622770
rect 338579 622751 339732 622770
rect 338579 622736 338688 622751
rect 338288 622687 338688 622736
rect 339588 622736 339732 622751
rect 339766 622736 339833 622770
rect 339867 622751 341020 622770
rect 339867 622736 339988 622751
rect 339588 622687 339988 622736
rect 340888 622736 341020 622751
rect 341054 622736 341088 622770
rect 340888 622687 341088 622736
rect 334648 622680 341088 622687
rect 334648 622646 334681 622680
rect 334715 622657 335868 622680
rect 334715 622646 334782 622657
rect 334648 622623 334782 622646
rect 334816 622623 334872 622657
rect 334906 622623 334962 622657
rect 334996 622623 335052 622657
rect 335086 622623 335142 622657
rect 335176 622623 335232 622657
rect 335266 622623 335322 622657
rect 335356 622623 335412 622657
rect 335446 622623 335502 622657
rect 335536 622623 335592 622657
rect 335626 622623 335682 622657
rect 335716 622623 335772 622657
rect 335806 622646 335868 622657
rect 335902 622646 335969 622680
rect 336003 622657 337156 622680
rect 336003 622646 336070 622657
rect 335806 622623 336070 622646
rect 336104 622623 336160 622657
rect 336194 622623 336250 622657
rect 336284 622623 336340 622657
rect 336374 622623 336430 622657
rect 336464 622623 336520 622657
rect 336554 622623 336610 622657
rect 336644 622623 336700 622657
rect 336734 622623 336790 622657
rect 336824 622623 336880 622657
rect 336914 622623 336970 622657
rect 337004 622623 337060 622657
rect 337094 622646 337156 622657
rect 337190 622646 337257 622680
rect 337291 622657 338444 622680
rect 337291 622646 337358 622657
rect 337094 622623 337358 622646
rect 337392 622623 337448 622657
rect 337482 622623 337538 622657
rect 337572 622623 337628 622657
rect 337662 622623 337718 622657
rect 337752 622623 337808 622657
rect 337842 622623 337898 622657
rect 337932 622623 337988 622657
rect 338022 622623 338078 622657
rect 338112 622623 338168 622657
rect 338202 622623 338258 622657
rect 338292 622623 338348 622657
rect 338382 622646 338444 622657
rect 338478 622646 338545 622680
rect 338579 622657 339732 622680
rect 338579 622646 338646 622657
rect 338382 622623 338646 622646
rect 338680 622623 338736 622657
rect 338770 622623 338826 622657
rect 338860 622623 338916 622657
rect 338950 622623 339006 622657
rect 339040 622623 339096 622657
rect 339130 622623 339186 622657
rect 339220 622623 339276 622657
rect 339310 622623 339366 622657
rect 339400 622623 339456 622657
rect 339490 622623 339546 622657
rect 339580 622623 339636 622657
rect 339670 622646 339732 622657
rect 339766 622646 339833 622680
rect 339867 622657 341020 622680
rect 339867 622646 339934 622657
rect 339670 622623 339934 622646
rect 339968 622623 340024 622657
rect 340058 622623 340114 622657
rect 340148 622623 340204 622657
rect 340238 622623 340294 622657
rect 340328 622623 340384 622657
rect 340418 622623 340474 622657
rect 340508 622623 340564 622657
rect 340598 622623 340654 622657
rect 340688 622623 340744 622657
rect 340778 622623 340834 622657
rect 340868 622623 340924 622657
rect 340958 622646 341020 622657
rect 341054 622646 341088 622680
rect 340958 622623 341088 622646
rect 334648 622556 341088 622623
rect 334648 622522 334782 622556
rect 334816 622522 334872 622556
rect 334906 622522 334962 622556
rect 334996 622522 335052 622556
rect 335086 622522 335142 622556
rect 335176 622522 335232 622556
rect 335266 622522 335322 622556
rect 335356 622522 335412 622556
rect 335446 622522 335502 622556
rect 335536 622522 335592 622556
rect 335626 622522 335682 622556
rect 335716 622522 335772 622556
rect 335806 622522 336070 622556
rect 336104 622522 336160 622556
rect 336194 622522 336250 622556
rect 336284 622522 336340 622556
rect 336374 622522 336430 622556
rect 336464 622522 336520 622556
rect 336554 622522 336610 622556
rect 336644 622522 336700 622556
rect 336734 622522 336790 622556
rect 336824 622522 336880 622556
rect 336914 622522 336970 622556
rect 337004 622522 337060 622556
rect 337094 622522 337358 622556
rect 337392 622522 337448 622556
rect 337482 622522 337538 622556
rect 337572 622522 337628 622556
rect 337662 622522 337718 622556
rect 337752 622522 337808 622556
rect 337842 622522 337898 622556
rect 337932 622522 337988 622556
rect 338022 622522 338078 622556
rect 338112 622522 338168 622556
rect 338202 622522 338258 622556
rect 338292 622522 338348 622556
rect 338382 622522 338646 622556
rect 338680 622522 338736 622556
rect 338770 622522 338826 622556
rect 338860 622522 338916 622556
rect 338950 622522 339006 622556
rect 339040 622522 339096 622556
rect 339130 622522 339186 622556
rect 339220 622522 339276 622556
rect 339310 622522 339366 622556
rect 339400 622522 339456 622556
rect 339490 622522 339546 622556
rect 339580 622522 339636 622556
rect 339670 622522 339934 622556
rect 339968 622522 340024 622556
rect 340058 622522 340114 622556
rect 340148 622522 340204 622556
rect 340238 622522 340294 622556
rect 340328 622522 340384 622556
rect 340418 622522 340474 622556
rect 340508 622522 340564 622556
rect 340598 622522 340654 622556
rect 340688 622522 340744 622556
rect 340778 622522 340834 622556
rect 340868 622522 340924 622556
rect 340958 622522 341088 622556
rect 334648 622489 341088 622522
rect 334648 622472 334888 622489
rect 334648 622438 334681 622472
rect 334715 622438 334888 622472
rect 334648 622425 334888 622438
rect 335688 622472 336188 622489
rect 335688 622438 335868 622472
rect 335902 622438 335969 622472
rect 336003 622438 336188 622472
rect 335688 622425 336188 622438
rect 336988 622472 337388 622489
rect 336988 622438 337156 622472
rect 337190 622438 337257 622472
rect 337291 622438 337388 622472
rect 336988 622425 337388 622438
rect 338288 622472 338688 622489
rect 338288 622438 338444 622472
rect 338478 622438 338545 622472
rect 338579 622438 338688 622472
rect 338288 622425 338688 622438
rect 339588 622472 339988 622489
rect 339588 622438 339732 622472
rect 339766 622438 339833 622472
rect 339867 622438 339988 622472
rect 339588 622425 339988 622438
rect 340888 622472 341088 622489
rect 340888 622438 341020 622472
rect 341054 622438 341088 622472
rect 340888 622425 341088 622438
rect 334648 622406 341088 622425
rect 334648 622382 334922 622406
rect 334648 622348 334681 622382
rect 334715 622372 334922 622382
rect 334956 622372 335012 622406
rect 335046 622372 335102 622406
rect 335136 622372 335192 622406
rect 335226 622372 335282 622406
rect 335316 622372 335372 622406
rect 335406 622372 335462 622406
rect 335496 622372 335552 622406
rect 335586 622372 335642 622406
rect 335676 622382 336210 622406
rect 335676 622372 335868 622382
rect 334715 622353 335868 622372
rect 334715 622348 334888 622353
rect 334648 622312 334888 622348
rect 334648 622292 334830 622312
rect 334648 622258 334681 622292
rect 334715 622278 334830 622292
rect 334864 622278 334888 622312
rect 335688 622348 335868 622353
rect 335902 622348 335969 622382
rect 336003 622372 336210 622382
rect 336244 622372 336300 622406
rect 336334 622372 336390 622406
rect 336424 622372 336480 622406
rect 336514 622372 336570 622406
rect 336604 622372 336660 622406
rect 336694 622372 336750 622406
rect 336784 622372 336840 622406
rect 336874 622372 336930 622406
rect 336964 622382 337498 622406
rect 336964 622372 337156 622382
rect 336003 622353 337156 622372
rect 336003 622348 336188 622353
rect 335688 622312 336188 622348
rect 335688 622293 336118 622312
rect 334715 622258 334888 622278
rect 334648 622222 334888 622258
rect 334648 622202 334830 622222
rect 334648 622168 334681 622202
rect 334715 622188 334830 622202
rect 334864 622188 334888 622222
rect 334715 622168 334888 622188
rect 334648 622132 334888 622168
rect 334648 622112 334830 622132
rect 334648 622078 334681 622112
rect 334715 622098 334830 622112
rect 334864 622098 334888 622132
rect 334715 622078 334888 622098
rect 334648 622042 334888 622078
rect 334648 622022 334830 622042
rect 334648 621988 334681 622022
rect 334715 622008 334830 622022
rect 334864 622008 334888 622042
rect 334715 621988 334888 622008
rect 334648 621952 334888 621988
rect 334648 621932 334830 621952
rect 334648 621898 334681 621932
rect 334715 621918 334830 621932
rect 334864 621918 334888 621952
rect 334715 621898 334888 621918
rect 334648 621862 334888 621898
rect 334648 621842 334830 621862
rect 334648 621808 334681 621842
rect 334715 621828 334830 621842
rect 334864 621828 334888 621862
rect 334715 621808 334888 621828
rect 334648 621772 334888 621808
rect 334648 621752 334830 621772
rect 334648 621718 334681 621752
rect 334715 621738 334830 621752
rect 334864 621738 334888 621772
rect 334715 621718 334888 621738
rect 334648 621682 334888 621718
rect 334648 621662 334830 621682
rect 334648 621628 334681 621662
rect 334715 621648 334830 621662
rect 334864 621648 334888 621682
rect 334715 621628 334888 621648
rect 334648 621592 334888 621628
rect 334945 622230 335639 622291
rect 334945 622196 335004 622230
rect 335038 622218 335094 622230
rect 335066 622196 335094 622218
rect 335128 622218 335184 622230
rect 335128 622196 335132 622218
rect 334945 622184 335032 622196
rect 335066 622184 335132 622196
rect 335166 622196 335184 622218
rect 335218 622218 335274 622230
rect 335218 622196 335232 622218
rect 335166 622184 335232 622196
rect 335266 622196 335274 622218
rect 335308 622218 335364 622230
rect 335398 622218 335454 622230
rect 335488 622218 335544 622230
rect 335308 622196 335332 622218
rect 335398 622196 335432 622218
rect 335488 622196 335532 622218
rect 335578 622196 335639 622230
rect 335266 622184 335332 622196
rect 335366 622184 335432 622196
rect 335466 622184 335532 622196
rect 335566 622184 335639 622196
rect 334945 622140 335639 622184
rect 334945 622106 335004 622140
rect 335038 622118 335094 622140
rect 335066 622106 335094 622118
rect 335128 622118 335184 622140
rect 335128 622106 335132 622118
rect 334945 622084 335032 622106
rect 335066 622084 335132 622106
rect 335166 622106 335184 622118
rect 335218 622118 335274 622140
rect 335218 622106 335232 622118
rect 335166 622084 335232 622106
rect 335266 622106 335274 622118
rect 335308 622118 335364 622140
rect 335398 622118 335454 622140
rect 335488 622118 335544 622140
rect 335308 622106 335332 622118
rect 335398 622106 335432 622118
rect 335488 622106 335532 622118
rect 335578 622106 335639 622140
rect 335266 622084 335332 622106
rect 335366 622084 335432 622106
rect 335466 622084 335532 622106
rect 335566 622084 335639 622106
rect 334945 622050 335639 622084
rect 334945 622016 335004 622050
rect 335038 622018 335094 622050
rect 335066 622016 335094 622018
rect 335128 622018 335184 622050
rect 335128 622016 335132 622018
rect 334945 621984 335032 622016
rect 335066 621984 335132 622016
rect 335166 622016 335184 622018
rect 335218 622018 335274 622050
rect 335218 622016 335232 622018
rect 335166 621984 335232 622016
rect 335266 622016 335274 622018
rect 335308 622018 335364 622050
rect 335398 622018 335454 622050
rect 335488 622018 335544 622050
rect 335308 622016 335332 622018
rect 335398 622016 335432 622018
rect 335488 622016 335532 622018
rect 335578 622016 335639 622050
rect 335266 621984 335332 622016
rect 335366 621984 335432 622016
rect 335466 621984 335532 622016
rect 335566 621984 335639 622016
rect 334945 621960 335639 621984
rect 334945 621926 335004 621960
rect 335038 621926 335094 621960
rect 335128 621926 335184 621960
rect 335218 621926 335274 621960
rect 335308 621926 335364 621960
rect 335398 621926 335454 621960
rect 335488 621926 335544 621960
rect 335578 621926 335639 621960
rect 334945 621918 335639 621926
rect 334945 621884 335032 621918
rect 335066 621884 335132 621918
rect 335166 621884 335232 621918
rect 335266 621884 335332 621918
rect 335366 621884 335432 621918
rect 335466 621884 335532 621918
rect 335566 621884 335639 621918
rect 334945 621870 335639 621884
rect 334945 621836 335004 621870
rect 335038 621836 335094 621870
rect 335128 621836 335184 621870
rect 335218 621836 335274 621870
rect 335308 621836 335364 621870
rect 335398 621836 335454 621870
rect 335488 621836 335544 621870
rect 335578 621836 335639 621870
rect 334945 621818 335639 621836
rect 334945 621784 335032 621818
rect 335066 621784 335132 621818
rect 335166 621784 335232 621818
rect 335266 621784 335332 621818
rect 335366 621784 335432 621818
rect 335466 621784 335532 621818
rect 335566 621784 335639 621818
rect 334945 621780 335639 621784
rect 334945 621746 335004 621780
rect 335038 621746 335094 621780
rect 335128 621746 335184 621780
rect 335218 621746 335274 621780
rect 335308 621746 335364 621780
rect 335398 621746 335454 621780
rect 335488 621746 335544 621780
rect 335578 621746 335639 621780
rect 334945 621718 335639 621746
rect 334945 621690 335032 621718
rect 335066 621690 335132 621718
rect 334945 621656 335004 621690
rect 335066 621684 335094 621690
rect 335038 621656 335094 621684
rect 335128 621684 335132 621690
rect 335166 621690 335232 621718
rect 335166 621684 335184 621690
rect 335128 621656 335184 621684
rect 335218 621684 335232 621690
rect 335266 621690 335332 621718
rect 335366 621690 335432 621718
rect 335466 621690 335532 621718
rect 335566 621690 335639 621718
rect 335266 621684 335274 621690
rect 335218 621656 335274 621684
rect 335308 621684 335332 621690
rect 335398 621684 335432 621690
rect 335488 621684 335532 621690
rect 335308 621656 335364 621684
rect 335398 621656 335454 621684
rect 335488 621656 335544 621684
rect 335578 621656 335639 621690
rect 334945 621597 335639 621656
rect 335688 622259 335720 622293
rect 335754 622292 336118 622293
rect 335754 622259 335868 622292
rect 335688 622258 335868 622259
rect 335902 622258 335969 622292
rect 336003 622278 336118 622292
rect 336152 622278 336188 622312
rect 336988 622348 337156 622353
rect 337190 622348 337257 622382
rect 337291 622372 337498 622382
rect 337532 622372 337588 622406
rect 337622 622372 337678 622406
rect 337712 622372 337768 622406
rect 337802 622372 337858 622406
rect 337892 622372 337948 622406
rect 337982 622372 338038 622406
rect 338072 622372 338128 622406
rect 338162 622372 338218 622406
rect 338252 622382 338786 622406
rect 338252 622372 338444 622382
rect 337291 622353 338444 622372
rect 337291 622348 337459 622353
rect 336988 622312 337459 622348
rect 336988 622293 337406 622312
rect 336003 622258 336188 622278
rect 335688 622222 336188 622258
rect 335688 622203 336118 622222
rect 335688 622169 335720 622203
rect 335754 622202 336118 622203
rect 335754 622169 335868 622202
rect 335688 622168 335868 622169
rect 335902 622168 335969 622202
rect 336003 622188 336118 622202
rect 336152 622188 336188 622222
rect 336003 622168 336188 622188
rect 335688 622132 336188 622168
rect 335688 622113 336118 622132
rect 335688 622079 335720 622113
rect 335754 622112 336118 622113
rect 335754 622079 335868 622112
rect 335688 622078 335868 622079
rect 335902 622078 335969 622112
rect 336003 622098 336118 622112
rect 336152 622098 336188 622132
rect 336003 622078 336188 622098
rect 335688 622042 336188 622078
rect 335688 622023 336118 622042
rect 335688 621989 335720 622023
rect 335754 622022 336118 622023
rect 335754 621989 335868 622022
rect 335688 621988 335868 621989
rect 335902 621988 335969 622022
rect 336003 622008 336118 622022
rect 336152 622008 336188 622042
rect 336003 621988 336188 622008
rect 335688 621952 336188 621988
rect 335688 621933 336118 621952
rect 335688 621899 335720 621933
rect 335754 621932 336118 621933
rect 335754 621899 335868 621932
rect 335688 621898 335868 621899
rect 335902 621898 335969 621932
rect 336003 621918 336118 621932
rect 336152 621918 336188 621952
rect 336003 621898 336188 621918
rect 335688 621862 336188 621898
rect 335688 621843 336118 621862
rect 335688 621809 335720 621843
rect 335754 621842 336118 621843
rect 335754 621809 335868 621842
rect 335688 621808 335868 621809
rect 335902 621808 335969 621842
rect 336003 621828 336118 621842
rect 336152 621828 336188 621862
rect 336003 621808 336188 621828
rect 335688 621772 336188 621808
rect 335688 621753 336118 621772
rect 335688 621719 335720 621753
rect 335754 621752 336118 621753
rect 335754 621719 335868 621752
rect 335688 621718 335868 621719
rect 335902 621718 335969 621752
rect 336003 621738 336118 621752
rect 336152 621738 336188 621772
rect 336003 621718 336188 621738
rect 335688 621682 336188 621718
rect 335688 621663 336118 621682
rect 335688 621629 335720 621663
rect 335754 621662 336118 621663
rect 335754 621629 335868 621662
rect 335688 621628 335868 621629
rect 335902 621628 335969 621662
rect 336003 621648 336118 621662
rect 336152 621648 336188 621682
rect 336003 621628 336188 621648
rect 334648 621572 334830 621592
rect 334648 621538 334681 621572
rect 334715 621558 334830 621572
rect 334864 621558 334888 621592
rect 334715 621538 334888 621558
rect 334648 621535 334888 621538
rect 335688 621592 336188 621628
rect 336233 622230 336927 622291
rect 336233 622196 336292 622230
rect 336326 622218 336382 622230
rect 336354 622196 336382 622218
rect 336416 622218 336472 622230
rect 336416 622196 336420 622218
rect 336233 622184 336320 622196
rect 336354 622184 336420 622196
rect 336454 622196 336472 622218
rect 336506 622218 336562 622230
rect 336506 622196 336520 622218
rect 336454 622184 336520 622196
rect 336554 622196 336562 622218
rect 336596 622218 336652 622230
rect 336686 622218 336742 622230
rect 336776 622218 336832 622230
rect 336596 622196 336620 622218
rect 336686 622196 336720 622218
rect 336776 622196 336820 622218
rect 336866 622196 336927 622230
rect 336554 622184 336620 622196
rect 336654 622184 336720 622196
rect 336754 622184 336820 622196
rect 336854 622184 336927 622196
rect 336233 622140 336927 622184
rect 336233 622106 336292 622140
rect 336326 622118 336382 622140
rect 336354 622106 336382 622118
rect 336416 622118 336472 622140
rect 336416 622106 336420 622118
rect 336233 622084 336320 622106
rect 336354 622084 336420 622106
rect 336454 622106 336472 622118
rect 336506 622118 336562 622140
rect 336506 622106 336520 622118
rect 336454 622084 336520 622106
rect 336554 622106 336562 622118
rect 336596 622118 336652 622140
rect 336686 622118 336742 622140
rect 336776 622118 336832 622140
rect 336596 622106 336620 622118
rect 336686 622106 336720 622118
rect 336776 622106 336820 622118
rect 336866 622106 336927 622140
rect 336554 622084 336620 622106
rect 336654 622084 336720 622106
rect 336754 622084 336820 622106
rect 336854 622084 336927 622106
rect 336233 622050 336927 622084
rect 336233 622016 336292 622050
rect 336326 622018 336382 622050
rect 336354 622016 336382 622018
rect 336416 622018 336472 622050
rect 336416 622016 336420 622018
rect 336233 621984 336320 622016
rect 336354 621984 336420 622016
rect 336454 622016 336472 622018
rect 336506 622018 336562 622050
rect 336506 622016 336520 622018
rect 336454 621984 336520 622016
rect 336554 622016 336562 622018
rect 336596 622018 336652 622050
rect 336686 622018 336742 622050
rect 336776 622018 336832 622050
rect 336596 622016 336620 622018
rect 336686 622016 336720 622018
rect 336776 622016 336820 622018
rect 336866 622016 336927 622050
rect 336554 621984 336620 622016
rect 336654 621984 336720 622016
rect 336754 621984 336820 622016
rect 336854 621984 336927 622016
rect 336233 621960 336927 621984
rect 336233 621926 336292 621960
rect 336326 621926 336382 621960
rect 336416 621926 336472 621960
rect 336506 621926 336562 621960
rect 336596 621926 336652 621960
rect 336686 621926 336742 621960
rect 336776 621926 336832 621960
rect 336866 621926 336927 621960
rect 336233 621918 336927 621926
rect 336233 621884 336320 621918
rect 336354 621884 336420 621918
rect 336454 621884 336520 621918
rect 336554 621884 336620 621918
rect 336654 621884 336720 621918
rect 336754 621884 336820 621918
rect 336854 621884 336927 621918
rect 336233 621870 336927 621884
rect 336233 621836 336292 621870
rect 336326 621836 336382 621870
rect 336416 621836 336472 621870
rect 336506 621836 336562 621870
rect 336596 621836 336652 621870
rect 336686 621836 336742 621870
rect 336776 621836 336832 621870
rect 336866 621836 336927 621870
rect 336233 621818 336927 621836
rect 336233 621784 336320 621818
rect 336354 621784 336420 621818
rect 336454 621784 336520 621818
rect 336554 621784 336620 621818
rect 336654 621784 336720 621818
rect 336754 621784 336820 621818
rect 336854 621784 336927 621818
rect 336233 621780 336927 621784
rect 336233 621746 336292 621780
rect 336326 621746 336382 621780
rect 336416 621746 336472 621780
rect 336506 621746 336562 621780
rect 336596 621746 336652 621780
rect 336686 621746 336742 621780
rect 336776 621746 336832 621780
rect 336866 621746 336927 621780
rect 336233 621718 336927 621746
rect 336233 621690 336320 621718
rect 336354 621690 336420 621718
rect 336233 621656 336292 621690
rect 336354 621684 336382 621690
rect 336326 621656 336382 621684
rect 336416 621684 336420 621690
rect 336454 621690 336520 621718
rect 336454 621684 336472 621690
rect 336416 621656 336472 621684
rect 336506 621684 336520 621690
rect 336554 621690 336620 621718
rect 336654 621690 336720 621718
rect 336754 621690 336820 621718
rect 336854 621690 336927 621718
rect 336554 621684 336562 621690
rect 336506 621656 336562 621684
rect 336596 621684 336620 621690
rect 336686 621684 336720 621690
rect 336776 621684 336820 621690
rect 336596 621656 336652 621684
rect 336686 621656 336742 621684
rect 336776 621656 336832 621684
rect 336866 621656 336927 621690
rect 336233 621597 336927 621656
rect 336988 622259 337008 622293
rect 337042 622292 337406 622293
rect 337042 622259 337156 622292
rect 336988 622258 337156 622259
rect 337190 622258 337257 622292
rect 337291 622278 337406 622292
rect 337440 622278 337459 622312
rect 338277 622348 338444 622353
rect 338478 622348 338545 622382
rect 338579 622372 338786 622382
rect 338820 622372 338876 622406
rect 338910 622372 338966 622406
rect 339000 622372 339056 622406
rect 339090 622372 339146 622406
rect 339180 622372 339236 622406
rect 339270 622372 339326 622406
rect 339360 622372 339416 622406
rect 339450 622372 339506 622406
rect 339540 622382 340074 622406
rect 339540 622372 339732 622382
rect 338579 622353 339732 622372
rect 338579 622348 338747 622353
rect 338277 622312 338747 622348
rect 338277 622293 338694 622312
rect 337291 622258 337459 622278
rect 336988 622222 337459 622258
rect 336988 622203 337406 622222
rect 336988 622169 337008 622203
rect 337042 622202 337406 622203
rect 337042 622169 337156 622202
rect 336988 622168 337156 622169
rect 337190 622168 337257 622202
rect 337291 622188 337406 622202
rect 337440 622188 337459 622222
rect 337291 622168 337459 622188
rect 336988 622132 337459 622168
rect 336988 622113 337406 622132
rect 336988 622079 337008 622113
rect 337042 622112 337406 622113
rect 337042 622079 337156 622112
rect 336988 622078 337156 622079
rect 337190 622078 337257 622112
rect 337291 622098 337406 622112
rect 337440 622098 337459 622132
rect 337291 622078 337459 622098
rect 336988 622042 337459 622078
rect 336988 622023 337406 622042
rect 336988 621989 337008 622023
rect 337042 622022 337406 622023
rect 337042 621989 337156 622022
rect 336988 621988 337156 621989
rect 337190 621988 337257 622022
rect 337291 622008 337406 622022
rect 337440 622008 337459 622042
rect 337291 621988 337459 622008
rect 336988 621952 337459 621988
rect 336988 621933 337406 621952
rect 336988 621899 337008 621933
rect 337042 621932 337406 621933
rect 337042 621899 337156 621932
rect 336988 621898 337156 621899
rect 337190 621898 337257 621932
rect 337291 621918 337406 621932
rect 337440 621918 337459 621952
rect 337291 621898 337459 621918
rect 336988 621862 337459 621898
rect 336988 621843 337406 621862
rect 336988 621809 337008 621843
rect 337042 621842 337406 621843
rect 337042 621809 337156 621842
rect 336988 621808 337156 621809
rect 337190 621808 337257 621842
rect 337291 621828 337406 621842
rect 337440 621828 337459 621862
rect 337291 621808 337459 621828
rect 336988 621772 337459 621808
rect 336988 621753 337406 621772
rect 336988 621719 337008 621753
rect 337042 621752 337406 621753
rect 337042 621719 337156 621752
rect 336988 621718 337156 621719
rect 337190 621718 337257 621752
rect 337291 621738 337406 621752
rect 337440 621738 337459 621772
rect 337291 621718 337459 621738
rect 336988 621682 337459 621718
rect 336988 621663 337406 621682
rect 336988 621629 337008 621663
rect 337042 621662 337406 621663
rect 337042 621629 337156 621662
rect 336988 621628 337156 621629
rect 337190 621628 337257 621662
rect 337291 621648 337406 621662
rect 337440 621648 337459 621682
rect 337291 621628 337459 621648
rect 335688 621573 336118 621592
rect 335688 621539 335720 621573
rect 335754 621572 336118 621573
rect 335754 621539 335868 621572
rect 335688 621538 335868 621539
rect 335902 621538 335969 621572
rect 336003 621558 336118 621572
rect 336152 621558 336188 621592
rect 336003 621538 336188 621558
rect 335688 621535 336188 621538
rect 336988 621592 337459 621628
rect 337521 622230 338215 622291
rect 337521 622196 337580 622230
rect 337614 622218 337670 622230
rect 337642 622196 337670 622218
rect 337704 622218 337760 622230
rect 337704 622196 337708 622218
rect 337521 622184 337608 622196
rect 337642 622184 337708 622196
rect 337742 622196 337760 622218
rect 337794 622218 337850 622230
rect 337794 622196 337808 622218
rect 337742 622184 337808 622196
rect 337842 622196 337850 622218
rect 337884 622218 337940 622230
rect 337974 622218 338030 622230
rect 338064 622218 338120 622230
rect 337884 622196 337908 622218
rect 337974 622196 338008 622218
rect 338064 622196 338108 622218
rect 338154 622196 338215 622230
rect 337842 622184 337908 622196
rect 337942 622184 338008 622196
rect 338042 622184 338108 622196
rect 338142 622184 338215 622196
rect 337521 622140 338215 622184
rect 337521 622106 337580 622140
rect 337614 622118 337670 622140
rect 337642 622106 337670 622118
rect 337704 622118 337760 622140
rect 337704 622106 337708 622118
rect 337521 622084 337608 622106
rect 337642 622084 337708 622106
rect 337742 622106 337760 622118
rect 337794 622118 337850 622140
rect 337794 622106 337808 622118
rect 337742 622084 337808 622106
rect 337842 622106 337850 622118
rect 337884 622118 337940 622140
rect 337974 622118 338030 622140
rect 338064 622118 338120 622140
rect 337884 622106 337908 622118
rect 337974 622106 338008 622118
rect 338064 622106 338108 622118
rect 338154 622106 338215 622140
rect 337842 622084 337908 622106
rect 337942 622084 338008 622106
rect 338042 622084 338108 622106
rect 338142 622084 338215 622106
rect 337521 622050 338215 622084
rect 337521 622016 337580 622050
rect 337614 622018 337670 622050
rect 337642 622016 337670 622018
rect 337704 622018 337760 622050
rect 337704 622016 337708 622018
rect 337521 621984 337608 622016
rect 337642 621984 337708 622016
rect 337742 622016 337760 622018
rect 337794 622018 337850 622050
rect 337794 622016 337808 622018
rect 337742 621984 337808 622016
rect 337842 622016 337850 622018
rect 337884 622018 337940 622050
rect 337974 622018 338030 622050
rect 338064 622018 338120 622050
rect 337884 622016 337908 622018
rect 337974 622016 338008 622018
rect 338064 622016 338108 622018
rect 338154 622016 338215 622050
rect 337842 621984 337908 622016
rect 337942 621984 338008 622016
rect 338042 621984 338108 622016
rect 338142 621984 338215 622016
rect 337521 621960 338215 621984
rect 337521 621926 337580 621960
rect 337614 621926 337670 621960
rect 337704 621926 337760 621960
rect 337794 621926 337850 621960
rect 337884 621926 337940 621960
rect 337974 621926 338030 621960
rect 338064 621926 338120 621960
rect 338154 621926 338215 621960
rect 337521 621918 338215 621926
rect 337521 621884 337608 621918
rect 337642 621884 337708 621918
rect 337742 621884 337808 621918
rect 337842 621884 337908 621918
rect 337942 621884 338008 621918
rect 338042 621884 338108 621918
rect 338142 621884 338215 621918
rect 337521 621870 338215 621884
rect 337521 621836 337580 621870
rect 337614 621836 337670 621870
rect 337704 621836 337760 621870
rect 337794 621836 337850 621870
rect 337884 621836 337940 621870
rect 337974 621836 338030 621870
rect 338064 621836 338120 621870
rect 338154 621836 338215 621870
rect 337521 621818 338215 621836
rect 337521 621784 337608 621818
rect 337642 621784 337708 621818
rect 337742 621784 337808 621818
rect 337842 621784 337908 621818
rect 337942 621784 338008 621818
rect 338042 621784 338108 621818
rect 338142 621784 338215 621818
rect 337521 621780 338215 621784
rect 337521 621746 337580 621780
rect 337614 621746 337670 621780
rect 337704 621746 337760 621780
rect 337794 621746 337850 621780
rect 337884 621746 337940 621780
rect 337974 621746 338030 621780
rect 338064 621746 338120 621780
rect 338154 621746 338215 621780
rect 337521 621718 338215 621746
rect 337521 621690 337608 621718
rect 337642 621690 337708 621718
rect 337521 621656 337580 621690
rect 337642 621684 337670 621690
rect 337614 621656 337670 621684
rect 337704 621684 337708 621690
rect 337742 621690 337808 621718
rect 337742 621684 337760 621690
rect 337704 621656 337760 621684
rect 337794 621684 337808 621690
rect 337842 621690 337908 621718
rect 337942 621690 338008 621718
rect 338042 621690 338108 621718
rect 338142 621690 338215 621718
rect 337842 621684 337850 621690
rect 337794 621656 337850 621684
rect 337884 621684 337908 621690
rect 337974 621684 338008 621690
rect 338064 621684 338108 621690
rect 337884 621656 337940 621684
rect 337974 621656 338030 621684
rect 338064 621656 338120 621684
rect 338154 621656 338215 621690
rect 337521 621597 338215 621656
rect 338277 622259 338296 622293
rect 338330 622292 338694 622293
rect 338330 622259 338444 622292
rect 338277 622258 338444 622259
rect 338478 622258 338545 622292
rect 338579 622278 338694 622292
rect 338728 622278 338747 622312
rect 339565 622348 339732 622353
rect 339766 622348 339833 622382
rect 339867 622372 340074 622382
rect 340108 622372 340164 622406
rect 340198 622372 340254 622406
rect 340288 622372 340344 622406
rect 340378 622372 340434 622406
rect 340468 622372 340524 622406
rect 340558 622372 340614 622406
rect 340648 622372 340704 622406
rect 340738 622372 340794 622406
rect 340828 622382 341088 622406
rect 340828 622372 341020 622382
rect 339867 622353 341020 622372
rect 339867 622348 340035 622353
rect 339565 622312 340035 622348
rect 339565 622293 339982 622312
rect 338579 622258 338747 622278
rect 338277 622222 338747 622258
rect 338277 622203 338694 622222
rect 338277 622169 338296 622203
rect 338330 622202 338694 622203
rect 338330 622169 338444 622202
rect 338277 622168 338444 622169
rect 338478 622168 338545 622202
rect 338579 622188 338694 622202
rect 338728 622188 338747 622222
rect 338579 622168 338747 622188
rect 338277 622132 338747 622168
rect 338277 622113 338694 622132
rect 338277 622079 338296 622113
rect 338330 622112 338694 622113
rect 338330 622079 338444 622112
rect 338277 622078 338444 622079
rect 338478 622078 338545 622112
rect 338579 622098 338694 622112
rect 338728 622098 338747 622132
rect 338579 622078 338747 622098
rect 338277 622042 338747 622078
rect 338277 622023 338694 622042
rect 338277 621989 338296 622023
rect 338330 622022 338694 622023
rect 338330 621989 338444 622022
rect 338277 621988 338444 621989
rect 338478 621988 338545 622022
rect 338579 622008 338694 622022
rect 338728 622008 338747 622042
rect 338579 621988 338747 622008
rect 338277 621952 338747 621988
rect 338277 621933 338694 621952
rect 338277 621899 338296 621933
rect 338330 621932 338694 621933
rect 338330 621899 338444 621932
rect 338277 621898 338444 621899
rect 338478 621898 338545 621932
rect 338579 621918 338694 621932
rect 338728 621918 338747 621952
rect 338579 621898 338747 621918
rect 338277 621862 338747 621898
rect 338277 621843 338694 621862
rect 338277 621809 338296 621843
rect 338330 621842 338694 621843
rect 338330 621809 338444 621842
rect 338277 621808 338444 621809
rect 338478 621808 338545 621842
rect 338579 621828 338694 621842
rect 338728 621828 338747 621862
rect 338579 621808 338747 621828
rect 338277 621772 338747 621808
rect 338277 621753 338694 621772
rect 338277 621719 338296 621753
rect 338330 621752 338694 621753
rect 338330 621719 338444 621752
rect 338277 621718 338444 621719
rect 338478 621718 338545 621752
rect 338579 621738 338694 621752
rect 338728 621738 338747 621772
rect 338579 621718 338747 621738
rect 338277 621682 338747 621718
rect 338277 621663 338694 621682
rect 338277 621629 338296 621663
rect 338330 621662 338694 621663
rect 338330 621629 338444 621662
rect 338277 621628 338444 621629
rect 338478 621628 338545 621662
rect 338579 621648 338694 621662
rect 338728 621648 338747 621682
rect 338579 621628 338747 621648
rect 336988 621573 337406 621592
rect 336988 621539 337008 621573
rect 337042 621572 337406 621573
rect 337042 621539 337156 621572
rect 336988 621538 337156 621539
rect 337190 621538 337257 621572
rect 337291 621558 337406 621572
rect 337440 621558 337459 621592
rect 337291 621538 337459 621558
rect 336988 621535 337459 621538
rect 338277 621592 338747 621628
rect 338809 622230 339503 622291
rect 338809 622196 338868 622230
rect 338902 622218 338958 622230
rect 338930 622196 338958 622218
rect 338992 622218 339048 622230
rect 338992 622196 338996 622218
rect 338809 622184 338896 622196
rect 338930 622184 338996 622196
rect 339030 622196 339048 622218
rect 339082 622218 339138 622230
rect 339082 622196 339096 622218
rect 339030 622184 339096 622196
rect 339130 622196 339138 622218
rect 339172 622218 339228 622230
rect 339262 622218 339318 622230
rect 339352 622218 339408 622230
rect 339172 622196 339196 622218
rect 339262 622196 339296 622218
rect 339352 622196 339396 622218
rect 339442 622196 339503 622230
rect 339130 622184 339196 622196
rect 339230 622184 339296 622196
rect 339330 622184 339396 622196
rect 339430 622184 339503 622196
rect 338809 622140 339503 622184
rect 338809 622106 338868 622140
rect 338902 622118 338958 622140
rect 338930 622106 338958 622118
rect 338992 622118 339048 622140
rect 338992 622106 338996 622118
rect 338809 622084 338896 622106
rect 338930 622084 338996 622106
rect 339030 622106 339048 622118
rect 339082 622118 339138 622140
rect 339082 622106 339096 622118
rect 339030 622084 339096 622106
rect 339130 622106 339138 622118
rect 339172 622118 339228 622140
rect 339262 622118 339318 622140
rect 339352 622118 339408 622140
rect 339172 622106 339196 622118
rect 339262 622106 339296 622118
rect 339352 622106 339396 622118
rect 339442 622106 339503 622140
rect 339130 622084 339196 622106
rect 339230 622084 339296 622106
rect 339330 622084 339396 622106
rect 339430 622084 339503 622106
rect 338809 622050 339503 622084
rect 338809 622016 338868 622050
rect 338902 622018 338958 622050
rect 338930 622016 338958 622018
rect 338992 622018 339048 622050
rect 338992 622016 338996 622018
rect 338809 621984 338896 622016
rect 338930 621984 338996 622016
rect 339030 622016 339048 622018
rect 339082 622018 339138 622050
rect 339082 622016 339096 622018
rect 339030 621984 339096 622016
rect 339130 622016 339138 622018
rect 339172 622018 339228 622050
rect 339262 622018 339318 622050
rect 339352 622018 339408 622050
rect 339172 622016 339196 622018
rect 339262 622016 339296 622018
rect 339352 622016 339396 622018
rect 339442 622016 339503 622050
rect 339130 621984 339196 622016
rect 339230 621984 339296 622016
rect 339330 621984 339396 622016
rect 339430 621984 339503 622016
rect 338809 621960 339503 621984
rect 338809 621926 338868 621960
rect 338902 621926 338958 621960
rect 338992 621926 339048 621960
rect 339082 621926 339138 621960
rect 339172 621926 339228 621960
rect 339262 621926 339318 621960
rect 339352 621926 339408 621960
rect 339442 621926 339503 621960
rect 338809 621918 339503 621926
rect 338809 621884 338896 621918
rect 338930 621884 338996 621918
rect 339030 621884 339096 621918
rect 339130 621884 339196 621918
rect 339230 621884 339296 621918
rect 339330 621884 339396 621918
rect 339430 621884 339503 621918
rect 338809 621870 339503 621884
rect 338809 621836 338868 621870
rect 338902 621836 338958 621870
rect 338992 621836 339048 621870
rect 339082 621836 339138 621870
rect 339172 621836 339228 621870
rect 339262 621836 339318 621870
rect 339352 621836 339408 621870
rect 339442 621836 339503 621870
rect 338809 621818 339503 621836
rect 338809 621784 338896 621818
rect 338930 621784 338996 621818
rect 339030 621784 339096 621818
rect 339130 621784 339196 621818
rect 339230 621784 339296 621818
rect 339330 621784 339396 621818
rect 339430 621784 339503 621818
rect 338809 621780 339503 621784
rect 338809 621746 338868 621780
rect 338902 621746 338958 621780
rect 338992 621746 339048 621780
rect 339082 621746 339138 621780
rect 339172 621746 339228 621780
rect 339262 621746 339318 621780
rect 339352 621746 339408 621780
rect 339442 621746 339503 621780
rect 338809 621718 339503 621746
rect 338809 621690 338896 621718
rect 338930 621690 338996 621718
rect 338809 621656 338868 621690
rect 338930 621684 338958 621690
rect 338902 621656 338958 621684
rect 338992 621684 338996 621690
rect 339030 621690 339096 621718
rect 339030 621684 339048 621690
rect 338992 621656 339048 621684
rect 339082 621684 339096 621690
rect 339130 621690 339196 621718
rect 339230 621690 339296 621718
rect 339330 621690 339396 621718
rect 339430 621690 339503 621718
rect 339130 621684 339138 621690
rect 339082 621656 339138 621684
rect 339172 621684 339196 621690
rect 339262 621684 339296 621690
rect 339352 621684 339396 621690
rect 339172 621656 339228 621684
rect 339262 621656 339318 621684
rect 339352 621656 339408 621684
rect 339442 621656 339503 621690
rect 338809 621597 339503 621656
rect 339565 622259 339584 622293
rect 339618 622292 339982 622293
rect 339618 622259 339732 622292
rect 339565 622258 339732 622259
rect 339766 622258 339833 622292
rect 339867 622278 339982 622292
rect 340016 622278 340035 622312
rect 340853 622348 341020 622353
rect 341054 622348 341088 622382
rect 340853 622293 341088 622348
rect 339867 622258 340035 622278
rect 339565 622222 340035 622258
rect 339565 622203 339982 622222
rect 339565 622169 339584 622203
rect 339618 622202 339982 622203
rect 339618 622169 339732 622202
rect 339565 622168 339732 622169
rect 339766 622168 339833 622202
rect 339867 622188 339982 622202
rect 340016 622188 340035 622222
rect 339867 622168 340035 622188
rect 339565 622132 340035 622168
rect 339565 622113 339982 622132
rect 339565 622079 339584 622113
rect 339618 622112 339982 622113
rect 339618 622079 339732 622112
rect 339565 622078 339732 622079
rect 339766 622078 339833 622112
rect 339867 622098 339982 622112
rect 340016 622098 340035 622132
rect 339867 622078 340035 622098
rect 339565 622042 340035 622078
rect 339565 622023 339982 622042
rect 339565 621989 339584 622023
rect 339618 622022 339982 622023
rect 339618 621989 339732 622022
rect 339565 621988 339732 621989
rect 339766 621988 339833 622022
rect 339867 622008 339982 622022
rect 340016 622008 340035 622042
rect 339867 621988 340035 622008
rect 339565 621952 340035 621988
rect 339565 621933 339982 621952
rect 339565 621899 339584 621933
rect 339618 621932 339982 621933
rect 339618 621899 339732 621932
rect 339565 621898 339732 621899
rect 339766 621898 339833 621932
rect 339867 621918 339982 621932
rect 340016 621918 340035 621952
rect 339867 621898 340035 621918
rect 339565 621862 340035 621898
rect 339565 621843 339982 621862
rect 339565 621809 339584 621843
rect 339618 621842 339982 621843
rect 339618 621809 339732 621842
rect 339565 621808 339732 621809
rect 339766 621808 339833 621842
rect 339867 621828 339982 621842
rect 340016 621828 340035 621862
rect 339867 621808 340035 621828
rect 339565 621772 340035 621808
rect 339565 621753 339982 621772
rect 339565 621719 339584 621753
rect 339618 621752 339982 621753
rect 339618 621719 339732 621752
rect 339565 621718 339732 621719
rect 339766 621718 339833 621752
rect 339867 621738 339982 621752
rect 340016 621738 340035 621772
rect 339867 621718 340035 621738
rect 339565 621682 340035 621718
rect 339565 621663 339982 621682
rect 339565 621629 339584 621663
rect 339618 621662 339982 621663
rect 339618 621629 339732 621662
rect 339565 621628 339732 621629
rect 339766 621628 339833 621662
rect 339867 621648 339982 621662
rect 340016 621648 340035 621682
rect 339867 621628 340035 621648
rect 338277 621573 338694 621592
rect 338277 621539 338296 621573
rect 338330 621572 338694 621573
rect 338330 621539 338444 621572
rect 338277 621538 338444 621539
rect 338478 621538 338545 621572
rect 338579 621558 338694 621572
rect 338728 621558 338747 621592
rect 338579 621538 338747 621558
rect 338277 621535 338747 621538
rect 339565 621592 340035 621628
rect 340097 622230 340791 622291
rect 340097 622196 340156 622230
rect 340190 622218 340246 622230
rect 340218 622196 340246 622218
rect 340280 622218 340336 622230
rect 340280 622196 340284 622218
rect 340097 622184 340184 622196
rect 340218 622184 340284 622196
rect 340318 622196 340336 622218
rect 340370 622218 340426 622230
rect 340370 622196 340384 622218
rect 340318 622184 340384 622196
rect 340418 622196 340426 622218
rect 340460 622218 340516 622230
rect 340550 622218 340606 622230
rect 340640 622218 340696 622230
rect 340460 622196 340484 622218
rect 340550 622196 340584 622218
rect 340640 622196 340684 622218
rect 340730 622196 340791 622230
rect 340418 622184 340484 622196
rect 340518 622184 340584 622196
rect 340618 622184 340684 622196
rect 340718 622184 340791 622196
rect 340097 622140 340791 622184
rect 340097 622106 340156 622140
rect 340190 622118 340246 622140
rect 340218 622106 340246 622118
rect 340280 622118 340336 622140
rect 340280 622106 340284 622118
rect 340097 622084 340184 622106
rect 340218 622084 340284 622106
rect 340318 622106 340336 622118
rect 340370 622118 340426 622140
rect 340370 622106 340384 622118
rect 340318 622084 340384 622106
rect 340418 622106 340426 622118
rect 340460 622118 340516 622140
rect 340550 622118 340606 622140
rect 340640 622118 340696 622140
rect 340460 622106 340484 622118
rect 340550 622106 340584 622118
rect 340640 622106 340684 622118
rect 340730 622106 340791 622140
rect 340418 622084 340484 622106
rect 340518 622084 340584 622106
rect 340618 622084 340684 622106
rect 340718 622084 340791 622106
rect 340097 622050 340791 622084
rect 340097 622016 340156 622050
rect 340190 622018 340246 622050
rect 340218 622016 340246 622018
rect 340280 622018 340336 622050
rect 340280 622016 340284 622018
rect 340097 621984 340184 622016
rect 340218 621984 340284 622016
rect 340318 622016 340336 622018
rect 340370 622018 340426 622050
rect 340370 622016 340384 622018
rect 340318 621984 340384 622016
rect 340418 622016 340426 622018
rect 340460 622018 340516 622050
rect 340550 622018 340606 622050
rect 340640 622018 340696 622050
rect 340460 622016 340484 622018
rect 340550 622016 340584 622018
rect 340640 622016 340684 622018
rect 340730 622016 340791 622050
rect 340418 621984 340484 622016
rect 340518 621984 340584 622016
rect 340618 621984 340684 622016
rect 340718 621984 340791 622016
rect 340097 621960 340791 621984
rect 340097 621926 340156 621960
rect 340190 621926 340246 621960
rect 340280 621926 340336 621960
rect 340370 621926 340426 621960
rect 340460 621926 340516 621960
rect 340550 621926 340606 621960
rect 340640 621926 340696 621960
rect 340730 621926 340791 621960
rect 340097 621918 340791 621926
rect 340097 621884 340184 621918
rect 340218 621884 340284 621918
rect 340318 621884 340384 621918
rect 340418 621884 340484 621918
rect 340518 621884 340584 621918
rect 340618 621884 340684 621918
rect 340718 621884 340791 621918
rect 340097 621870 340791 621884
rect 340097 621836 340156 621870
rect 340190 621836 340246 621870
rect 340280 621836 340336 621870
rect 340370 621836 340426 621870
rect 340460 621836 340516 621870
rect 340550 621836 340606 621870
rect 340640 621836 340696 621870
rect 340730 621836 340791 621870
rect 340097 621818 340791 621836
rect 340097 621784 340184 621818
rect 340218 621784 340284 621818
rect 340318 621784 340384 621818
rect 340418 621784 340484 621818
rect 340518 621784 340584 621818
rect 340618 621784 340684 621818
rect 340718 621784 340791 621818
rect 340097 621780 340791 621784
rect 340097 621746 340156 621780
rect 340190 621746 340246 621780
rect 340280 621746 340336 621780
rect 340370 621746 340426 621780
rect 340460 621746 340516 621780
rect 340550 621746 340606 621780
rect 340640 621746 340696 621780
rect 340730 621746 340791 621780
rect 340097 621718 340791 621746
rect 340097 621690 340184 621718
rect 340218 621690 340284 621718
rect 340097 621656 340156 621690
rect 340218 621684 340246 621690
rect 340190 621656 340246 621684
rect 340280 621684 340284 621690
rect 340318 621690 340384 621718
rect 340318 621684 340336 621690
rect 340280 621656 340336 621684
rect 340370 621684 340384 621690
rect 340418 621690 340484 621718
rect 340518 621690 340584 621718
rect 340618 621690 340684 621718
rect 340718 621690 340791 621718
rect 340418 621684 340426 621690
rect 340370 621656 340426 621684
rect 340460 621684 340484 621690
rect 340550 621684 340584 621690
rect 340640 621684 340684 621690
rect 340460 621656 340516 621684
rect 340550 621656 340606 621684
rect 340640 621656 340696 621684
rect 340730 621656 340791 621690
rect 340097 621597 340791 621656
rect 340853 622259 340872 622293
rect 340906 622292 341088 622293
rect 340906 622259 341020 622292
rect 340853 622258 341020 622259
rect 341054 622258 341088 622292
rect 340853 622203 341088 622258
rect 340853 622169 340872 622203
rect 340906 622202 341088 622203
rect 340906 622169 341020 622202
rect 340853 622168 341020 622169
rect 341054 622168 341088 622202
rect 340853 622113 341088 622168
rect 340853 622079 340872 622113
rect 340906 622112 341088 622113
rect 340906 622079 341020 622112
rect 340853 622078 341020 622079
rect 341054 622078 341088 622112
rect 340853 622023 341088 622078
rect 340853 621989 340872 622023
rect 340906 622022 341088 622023
rect 340906 621989 341020 622022
rect 340853 621988 341020 621989
rect 341054 621988 341088 622022
rect 340853 621933 341088 621988
rect 340853 621899 340872 621933
rect 340906 621932 341088 621933
rect 340906 621899 341020 621932
rect 340853 621898 341020 621899
rect 341054 621898 341088 621932
rect 340853 621843 341088 621898
rect 340853 621809 340872 621843
rect 340906 621842 341088 621843
rect 340906 621809 341020 621842
rect 340853 621808 341020 621809
rect 341054 621808 341088 621842
rect 340853 621753 341088 621808
rect 340853 621719 340872 621753
rect 340906 621752 341088 621753
rect 340906 621719 341020 621752
rect 340853 621718 341020 621719
rect 341054 621718 341088 621752
rect 340853 621663 341088 621718
rect 340853 621629 340872 621663
rect 340906 621662 341088 621663
rect 340906 621629 341020 621662
rect 340853 621628 341020 621629
rect 341054 621628 341088 621662
rect 339565 621573 339982 621592
rect 339565 621539 339584 621573
rect 339618 621572 339982 621573
rect 339618 621539 339732 621572
rect 339565 621538 339732 621539
rect 339766 621538 339833 621572
rect 339867 621558 339982 621572
rect 340016 621558 340035 621592
rect 339867 621538 340035 621558
rect 339565 621535 340035 621538
rect 340853 621573 341088 621628
rect 340853 621539 340872 621573
rect 340906 621572 341088 621573
rect 340906 621539 341020 621572
rect 340853 621538 341020 621539
rect 341054 621538 341088 621572
rect 340853 621535 341088 621538
rect 334648 621516 341088 621535
rect 334648 621482 334888 621516
rect 334922 621482 334978 621516
rect 335012 621482 335068 621516
rect 335102 621482 335158 621516
rect 335192 621482 335248 621516
rect 335282 621482 335338 621516
rect 335372 621482 335428 621516
rect 335462 621482 335518 621516
rect 335552 621482 335608 621516
rect 335642 621482 336176 621516
rect 336210 621482 336266 621516
rect 336300 621482 336356 621516
rect 336390 621482 336446 621516
rect 336480 621482 336536 621516
rect 336570 621482 336626 621516
rect 336660 621482 336716 621516
rect 336750 621482 336806 621516
rect 336840 621482 336896 621516
rect 336930 621482 337464 621516
rect 337498 621482 337554 621516
rect 337588 621482 337644 621516
rect 337678 621482 337734 621516
rect 337768 621482 337824 621516
rect 337858 621482 337914 621516
rect 337948 621482 338004 621516
rect 338038 621482 338094 621516
rect 338128 621482 338184 621516
rect 338218 621482 338752 621516
rect 338786 621482 338842 621516
rect 338876 621482 338932 621516
rect 338966 621482 339022 621516
rect 339056 621482 339112 621516
rect 339146 621482 339202 621516
rect 339236 621482 339292 621516
rect 339326 621482 339382 621516
rect 339416 621482 339472 621516
rect 339506 621482 340040 621516
rect 340074 621482 340130 621516
rect 340164 621482 340220 621516
rect 340254 621482 340310 621516
rect 340344 621482 340400 621516
rect 340434 621482 340490 621516
rect 340524 621482 340580 621516
rect 340614 621482 340670 621516
rect 340704 621482 340760 621516
rect 340794 621482 341088 621516
rect 334648 621448 334681 621482
rect 334715 621463 335868 621482
rect 334715 621448 334888 621463
rect 334648 621399 334888 621448
rect 335688 621448 335868 621463
rect 335902 621448 335969 621482
rect 336003 621463 337156 621482
rect 336003 621448 336188 621463
rect 335688 621399 336188 621448
rect 336988 621448 337156 621463
rect 337190 621448 337257 621482
rect 337291 621463 338444 621482
rect 337291 621448 337388 621463
rect 336988 621399 337388 621448
rect 338288 621448 338444 621463
rect 338478 621448 338545 621482
rect 338579 621463 339732 621482
rect 338579 621448 338688 621463
rect 338288 621399 338688 621448
rect 339588 621448 339732 621463
rect 339766 621448 339833 621482
rect 339867 621463 341020 621482
rect 339867 621448 339988 621463
rect 339588 621399 339988 621448
rect 340888 621448 341020 621463
rect 341054 621448 341088 621482
rect 340888 621399 341088 621448
rect 334648 621392 341088 621399
rect 334648 621358 334681 621392
rect 334715 621369 335868 621392
rect 334715 621358 334782 621369
rect 334648 621335 334782 621358
rect 334816 621335 334872 621369
rect 334906 621335 334962 621369
rect 334996 621335 335052 621369
rect 335086 621335 335142 621369
rect 335176 621335 335232 621369
rect 335266 621335 335322 621369
rect 335356 621335 335412 621369
rect 335446 621335 335502 621369
rect 335536 621335 335592 621369
rect 335626 621335 335682 621369
rect 335716 621335 335772 621369
rect 335806 621358 335868 621369
rect 335902 621358 335969 621392
rect 336003 621369 337156 621392
rect 336003 621358 336070 621369
rect 335806 621335 336070 621358
rect 336104 621335 336160 621369
rect 336194 621335 336250 621369
rect 336284 621335 336340 621369
rect 336374 621335 336430 621369
rect 336464 621335 336520 621369
rect 336554 621335 336610 621369
rect 336644 621335 336700 621369
rect 336734 621335 336790 621369
rect 336824 621335 336880 621369
rect 336914 621335 336970 621369
rect 337004 621335 337060 621369
rect 337094 621358 337156 621369
rect 337190 621358 337257 621392
rect 337291 621369 338444 621392
rect 337291 621358 337358 621369
rect 337094 621335 337358 621358
rect 337392 621335 337448 621369
rect 337482 621335 337538 621369
rect 337572 621335 337628 621369
rect 337662 621335 337718 621369
rect 337752 621335 337808 621369
rect 337842 621335 337898 621369
rect 337932 621335 337988 621369
rect 338022 621335 338078 621369
rect 338112 621335 338168 621369
rect 338202 621335 338258 621369
rect 338292 621335 338348 621369
rect 338382 621358 338444 621369
rect 338478 621358 338545 621392
rect 338579 621369 339732 621392
rect 338579 621358 338646 621369
rect 338382 621335 338646 621358
rect 338680 621335 338736 621369
rect 338770 621335 338826 621369
rect 338860 621335 338916 621369
rect 338950 621335 339006 621369
rect 339040 621335 339096 621369
rect 339130 621335 339186 621369
rect 339220 621335 339276 621369
rect 339310 621335 339366 621369
rect 339400 621335 339456 621369
rect 339490 621335 339546 621369
rect 339580 621335 339636 621369
rect 339670 621358 339732 621369
rect 339766 621358 339833 621392
rect 339867 621369 341020 621392
rect 339867 621358 339934 621369
rect 339670 621335 339934 621358
rect 339968 621335 340024 621369
rect 340058 621335 340114 621369
rect 340148 621335 340204 621369
rect 340238 621335 340294 621369
rect 340328 621335 340384 621369
rect 340418 621335 340474 621369
rect 340508 621335 340564 621369
rect 340598 621335 340654 621369
rect 340688 621335 340744 621369
rect 340778 621335 340834 621369
rect 340868 621335 340924 621369
rect 340958 621358 341020 621369
rect 341054 621358 341088 621392
rect 340958 621335 341088 621358
rect 334648 621268 341088 621335
rect 334648 621234 334782 621268
rect 334816 621234 334872 621268
rect 334906 621234 334962 621268
rect 334996 621234 335052 621268
rect 335086 621234 335142 621268
rect 335176 621234 335232 621268
rect 335266 621234 335322 621268
rect 335356 621234 335412 621268
rect 335446 621234 335502 621268
rect 335536 621234 335592 621268
rect 335626 621234 335682 621268
rect 335716 621234 335772 621268
rect 335806 621234 336070 621268
rect 336104 621234 336160 621268
rect 336194 621234 336250 621268
rect 336284 621234 336340 621268
rect 336374 621234 336430 621268
rect 336464 621234 336520 621268
rect 336554 621234 336610 621268
rect 336644 621234 336700 621268
rect 336734 621234 336790 621268
rect 336824 621234 336880 621268
rect 336914 621234 336970 621268
rect 337004 621234 337060 621268
rect 337094 621234 337358 621268
rect 337392 621234 337448 621268
rect 337482 621234 337538 621268
rect 337572 621234 337628 621268
rect 337662 621234 337718 621268
rect 337752 621234 337808 621268
rect 337842 621234 337898 621268
rect 337932 621234 337988 621268
rect 338022 621234 338078 621268
rect 338112 621234 338168 621268
rect 338202 621234 338258 621268
rect 338292 621234 338348 621268
rect 338382 621234 338646 621268
rect 338680 621234 338736 621268
rect 338770 621234 338826 621268
rect 338860 621234 338916 621268
rect 338950 621234 339006 621268
rect 339040 621234 339096 621268
rect 339130 621234 339186 621268
rect 339220 621234 339276 621268
rect 339310 621234 339366 621268
rect 339400 621234 339456 621268
rect 339490 621234 339546 621268
rect 339580 621234 339636 621268
rect 339670 621234 339934 621268
rect 339968 621234 340024 621268
rect 340058 621234 340114 621268
rect 340148 621234 340204 621268
rect 340238 621234 340294 621268
rect 340328 621234 340384 621268
rect 340418 621234 340474 621268
rect 340508 621234 340564 621268
rect 340598 621234 340654 621268
rect 340688 621234 340744 621268
rect 340778 621234 340834 621268
rect 340868 621234 340924 621268
rect 340958 621234 341088 621268
rect 334648 621201 341088 621234
rect 334648 621184 334888 621201
rect 334648 621150 334681 621184
rect 334715 621150 334888 621184
rect 334648 621137 334888 621150
rect 335688 621184 336188 621201
rect 335688 621150 335868 621184
rect 335902 621150 335969 621184
rect 336003 621150 336188 621184
rect 335688 621137 336188 621150
rect 336988 621184 337388 621201
rect 336988 621150 337156 621184
rect 337190 621150 337257 621184
rect 337291 621150 337388 621184
rect 336988 621137 337388 621150
rect 338288 621184 338688 621201
rect 338288 621150 338444 621184
rect 338478 621150 338545 621184
rect 338579 621150 338688 621184
rect 338288 621137 338688 621150
rect 339588 621184 339988 621201
rect 339588 621150 339732 621184
rect 339766 621150 339833 621184
rect 339867 621150 339988 621184
rect 339588 621137 339988 621150
rect 340888 621184 341088 621201
rect 340888 621150 341020 621184
rect 341054 621150 341088 621184
rect 340888 621137 341088 621150
rect 334648 621118 341088 621137
rect 334648 621094 334922 621118
rect 334648 621060 334681 621094
rect 334715 621084 334922 621094
rect 334956 621084 335012 621118
rect 335046 621084 335102 621118
rect 335136 621084 335192 621118
rect 335226 621084 335282 621118
rect 335316 621084 335372 621118
rect 335406 621084 335462 621118
rect 335496 621084 335552 621118
rect 335586 621084 335642 621118
rect 335676 621094 336210 621118
rect 335676 621084 335868 621094
rect 334715 621065 335868 621084
rect 334715 621060 334888 621065
rect 334648 621024 334888 621060
rect 334648 621004 334830 621024
rect 334648 620970 334681 621004
rect 334715 620990 334830 621004
rect 334864 620990 334888 621024
rect 335688 621060 335868 621065
rect 335902 621060 335969 621094
rect 336003 621084 336210 621094
rect 336244 621084 336300 621118
rect 336334 621084 336390 621118
rect 336424 621084 336480 621118
rect 336514 621084 336570 621118
rect 336604 621084 336660 621118
rect 336694 621084 336750 621118
rect 336784 621084 336840 621118
rect 336874 621084 336930 621118
rect 336964 621094 337498 621118
rect 336964 621084 337156 621094
rect 336003 621065 337156 621084
rect 336003 621060 336188 621065
rect 335688 621024 336188 621060
rect 335688 621005 336118 621024
rect 334715 620970 334888 620990
rect 334648 620934 334888 620970
rect 334648 620914 334830 620934
rect 334648 620880 334681 620914
rect 334715 620900 334830 620914
rect 334864 620900 334888 620934
rect 334715 620880 334888 620900
rect 334648 620844 334888 620880
rect 334648 620824 334830 620844
rect 334648 620790 334681 620824
rect 334715 620810 334830 620824
rect 334864 620810 334888 620844
rect 334715 620790 334888 620810
rect 334648 620754 334888 620790
rect 334648 620734 334830 620754
rect 334648 620700 334681 620734
rect 334715 620720 334830 620734
rect 334864 620720 334888 620754
rect 334715 620700 334888 620720
rect 334648 620664 334888 620700
rect 334648 620644 334830 620664
rect 334648 620610 334681 620644
rect 334715 620630 334830 620644
rect 334864 620630 334888 620664
rect 334715 620610 334888 620630
rect 334648 620574 334888 620610
rect 334648 620554 334830 620574
rect 334648 620520 334681 620554
rect 334715 620540 334830 620554
rect 334864 620540 334888 620574
rect 334715 620520 334888 620540
rect 334648 620484 334888 620520
rect 334648 620464 334830 620484
rect 334648 620430 334681 620464
rect 334715 620450 334830 620464
rect 334864 620450 334888 620484
rect 334715 620430 334888 620450
rect 334648 620394 334888 620430
rect 334648 620374 334830 620394
rect 334648 620340 334681 620374
rect 334715 620360 334830 620374
rect 334864 620360 334888 620394
rect 334715 620340 334888 620360
rect 334648 620304 334888 620340
rect 334945 620942 335639 621003
rect 334945 620908 335004 620942
rect 335038 620930 335094 620942
rect 335066 620908 335094 620930
rect 335128 620930 335184 620942
rect 335128 620908 335132 620930
rect 334945 620896 335032 620908
rect 335066 620896 335132 620908
rect 335166 620908 335184 620930
rect 335218 620930 335274 620942
rect 335218 620908 335232 620930
rect 335166 620896 335232 620908
rect 335266 620908 335274 620930
rect 335308 620930 335364 620942
rect 335398 620930 335454 620942
rect 335488 620930 335544 620942
rect 335308 620908 335332 620930
rect 335398 620908 335432 620930
rect 335488 620908 335532 620930
rect 335578 620908 335639 620942
rect 335266 620896 335332 620908
rect 335366 620896 335432 620908
rect 335466 620896 335532 620908
rect 335566 620896 335639 620908
rect 334945 620852 335639 620896
rect 334945 620818 335004 620852
rect 335038 620830 335094 620852
rect 335066 620818 335094 620830
rect 335128 620830 335184 620852
rect 335128 620818 335132 620830
rect 334945 620796 335032 620818
rect 335066 620796 335132 620818
rect 335166 620818 335184 620830
rect 335218 620830 335274 620852
rect 335218 620818 335232 620830
rect 335166 620796 335232 620818
rect 335266 620818 335274 620830
rect 335308 620830 335364 620852
rect 335398 620830 335454 620852
rect 335488 620830 335544 620852
rect 335308 620818 335332 620830
rect 335398 620818 335432 620830
rect 335488 620818 335532 620830
rect 335578 620818 335639 620852
rect 335266 620796 335332 620818
rect 335366 620796 335432 620818
rect 335466 620796 335532 620818
rect 335566 620796 335639 620818
rect 334945 620762 335639 620796
rect 334945 620728 335004 620762
rect 335038 620730 335094 620762
rect 335066 620728 335094 620730
rect 335128 620730 335184 620762
rect 335128 620728 335132 620730
rect 334945 620696 335032 620728
rect 335066 620696 335132 620728
rect 335166 620728 335184 620730
rect 335218 620730 335274 620762
rect 335218 620728 335232 620730
rect 335166 620696 335232 620728
rect 335266 620728 335274 620730
rect 335308 620730 335364 620762
rect 335398 620730 335454 620762
rect 335488 620730 335544 620762
rect 335308 620728 335332 620730
rect 335398 620728 335432 620730
rect 335488 620728 335532 620730
rect 335578 620728 335639 620762
rect 335266 620696 335332 620728
rect 335366 620696 335432 620728
rect 335466 620696 335532 620728
rect 335566 620696 335639 620728
rect 334945 620672 335639 620696
rect 334945 620638 335004 620672
rect 335038 620638 335094 620672
rect 335128 620638 335184 620672
rect 335218 620638 335274 620672
rect 335308 620638 335364 620672
rect 335398 620638 335454 620672
rect 335488 620638 335544 620672
rect 335578 620638 335639 620672
rect 334945 620630 335639 620638
rect 334945 620596 335032 620630
rect 335066 620596 335132 620630
rect 335166 620596 335232 620630
rect 335266 620596 335332 620630
rect 335366 620596 335432 620630
rect 335466 620596 335532 620630
rect 335566 620596 335639 620630
rect 334945 620582 335639 620596
rect 334945 620548 335004 620582
rect 335038 620548 335094 620582
rect 335128 620548 335184 620582
rect 335218 620548 335274 620582
rect 335308 620548 335364 620582
rect 335398 620548 335454 620582
rect 335488 620548 335544 620582
rect 335578 620548 335639 620582
rect 334945 620530 335639 620548
rect 334945 620496 335032 620530
rect 335066 620496 335132 620530
rect 335166 620496 335232 620530
rect 335266 620496 335332 620530
rect 335366 620496 335432 620530
rect 335466 620496 335532 620530
rect 335566 620496 335639 620530
rect 334945 620492 335639 620496
rect 334945 620458 335004 620492
rect 335038 620458 335094 620492
rect 335128 620458 335184 620492
rect 335218 620458 335274 620492
rect 335308 620458 335364 620492
rect 335398 620458 335454 620492
rect 335488 620458 335544 620492
rect 335578 620458 335639 620492
rect 334945 620430 335639 620458
rect 334945 620402 335032 620430
rect 335066 620402 335132 620430
rect 334945 620368 335004 620402
rect 335066 620396 335094 620402
rect 335038 620368 335094 620396
rect 335128 620396 335132 620402
rect 335166 620402 335232 620430
rect 335166 620396 335184 620402
rect 335128 620368 335184 620396
rect 335218 620396 335232 620402
rect 335266 620402 335332 620430
rect 335366 620402 335432 620430
rect 335466 620402 335532 620430
rect 335566 620402 335639 620430
rect 335266 620396 335274 620402
rect 335218 620368 335274 620396
rect 335308 620396 335332 620402
rect 335398 620396 335432 620402
rect 335488 620396 335532 620402
rect 335308 620368 335364 620396
rect 335398 620368 335454 620396
rect 335488 620368 335544 620396
rect 335578 620368 335639 620402
rect 334945 620309 335639 620368
rect 335688 620971 335720 621005
rect 335754 621004 336118 621005
rect 335754 620971 335868 621004
rect 335688 620970 335868 620971
rect 335902 620970 335969 621004
rect 336003 620990 336118 621004
rect 336152 620990 336188 621024
rect 336988 621060 337156 621065
rect 337190 621060 337257 621094
rect 337291 621084 337498 621094
rect 337532 621084 337588 621118
rect 337622 621084 337678 621118
rect 337712 621084 337768 621118
rect 337802 621084 337858 621118
rect 337892 621084 337948 621118
rect 337982 621084 338038 621118
rect 338072 621084 338128 621118
rect 338162 621084 338218 621118
rect 338252 621094 338786 621118
rect 338252 621084 338444 621094
rect 337291 621065 338444 621084
rect 337291 621060 337459 621065
rect 336988 621024 337459 621060
rect 336988 621005 337406 621024
rect 336003 620970 336188 620990
rect 335688 620934 336188 620970
rect 335688 620915 336118 620934
rect 335688 620881 335720 620915
rect 335754 620914 336118 620915
rect 335754 620881 335868 620914
rect 335688 620880 335868 620881
rect 335902 620880 335969 620914
rect 336003 620900 336118 620914
rect 336152 620900 336188 620934
rect 336003 620880 336188 620900
rect 335688 620844 336188 620880
rect 335688 620825 336118 620844
rect 335688 620791 335720 620825
rect 335754 620824 336118 620825
rect 335754 620791 335868 620824
rect 335688 620790 335868 620791
rect 335902 620790 335969 620824
rect 336003 620810 336118 620824
rect 336152 620810 336188 620844
rect 336003 620790 336188 620810
rect 335688 620754 336188 620790
rect 335688 620735 336118 620754
rect 335688 620701 335720 620735
rect 335754 620734 336118 620735
rect 335754 620701 335868 620734
rect 335688 620700 335868 620701
rect 335902 620700 335969 620734
rect 336003 620720 336118 620734
rect 336152 620720 336188 620754
rect 336003 620700 336188 620720
rect 335688 620664 336188 620700
rect 335688 620645 336118 620664
rect 335688 620611 335720 620645
rect 335754 620644 336118 620645
rect 335754 620611 335868 620644
rect 335688 620610 335868 620611
rect 335902 620610 335969 620644
rect 336003 620630 336118 620644
rect 336152 620630 336188 620664
rect 336003 620610 336188 620630
rect 335688 620574 336188 620610
rect 335688 620555 336118 620574
rect 335688 620521 335720 620555
rect 335754 620554 336118 620555
rect 335754 620521 335868 620554
rect 335688 620520 335868 620521
rect 335902 620520 335969 620554
rect 336003 620540 336118 620554
rect 336152 620540 336188 620574
rect 336003 620520 336188 620540
rect 335688 620484 336188 620520
rect 335688 620465 336118 620484
rect 335688 620431 335720 620465
rect 335754 620464 336118 620465
rect 335754 620431 335868 620464
rect 335688 620430 335868 620431
rect 335902 620430 335969 620464
rect 336003 620450 336118 620464
rect 336152 620450 336188 620484
rect 336003 620430 336188 620450
rect 335688 620394 336188 620430
rect 335688 620375 336118 620394
rect 335688 620341 335720 620375
rect 335754 620374 336118 620375
rect 335754 620341 335868 620374
rect 335688 620340 335868 620341
rect 335902 620340 335969 620374
rect 336003 620360 336118 620374
rect 336152 620360 336188 620394
rect 336003 620340 336188 620360
rect 334648 620284 334830 620304
rect 334648 620250 334681 620284
rect 334715 620270 334830 620284
rect 334864 620270 334888 620304
rect 334715 620250 334888 620270
rect 334648 620247 334888 620250
rect 335688 620304 336188 620340
rect 336233 620942 336927 621003
rect 336233 620908 336292 620942
rect 336326 620930 336382 620942
rect 336354 620908 336382 620930
rect 336416 620930 336472 620942
rect 336416 620908 336420 620930
rect 336233 620896 336320 620908
rect 336354 620896 336420 620908
rect 336454 620908 336472 620930
rect 336506 620930 336562 620942
rect 336506 620908 336520 620930
rect 336454 620896 336520 620908
rect 336554 620908 336562 620930
rect 336596 620930 336652 620942
rect 336686 620930 336742 620942
rect 336776 620930 336832 620942
rect 336596 620908 336620 620930
rect 336686 620908 336720 620930
rect 336776 620908 336820 620930
rect 336866 620908 336927 620942
rect 336554 620896 336620 620908
rect 336654 620896 336720 620908
rect 336754 620896 336820 620908
rect 336854 620896 336927 620908
rect 336233 620852 336927 620896
rect 336233 620818 336292 620852
rect 336326 620830 336382 620852
rect 336354 620818 336382 620830
rect 336416 620830 336472 620852
rect 336416 620818 336420 620830
rect 336233 620796 336320 620818
rect 336354 620796 336420 620818
rect 336454 620818 336472 620830
rect 336506 620830 336562 620852
rect 336506 620818 336520 620830
rect 336454 620796 336520 620818
rect 336554 620818 336562 620830
rect 336596 620830 336652 620852
rect 336686 620830 336742 620852
rect 336776 620830 336832 620852
rect 336596 620818 336620 620830
rect 336686 620818 336720 620830
rect 336776 620818 336820 620830
rect 336866 620818 336927 620852
rect 336554 620796 336620 620818
rect 336654 620796 336720 620818
rect 336754 620796 336820 620818
rect 336854 620796 336927 620818
rect 336233 620762 336927 620796
rect 336233 620728 336292 620762
rect 336326 620730 336382 620762
rect 336354 620728 336382 620730
rect 336416 620730 336472 620762
rect 336416 620728 336420 620730
rect 336233 620696 336320 620728
rect 336354 620696 336420 620728
rect 336454 620728 336472 620730
rect 336506 620730 336562 620762
rect 336506 620728 336520 620730
rect 336454 620696 336520 620728
rect 336554 620728 336562 620730
rect 336596 620730 336652 620762
rect 336686 620730 336742 620762
rect 336776 620730 336832 620762
rect 336596 620728 336620 620730
rect 336686 620728 336720 620730
rect 336776 620728 336820 620730
rect 336866 620728 336927 620762
rect 336554 620696 336620 620728
rect 336654 620696 336720 620728
rect 336754 620696 336820 620728
rect 336854 620696 336927 620728
rect 336233 620672 336927 620696
rect 336233 620638 336292 620672
rect 336326 620638 336382 620672
rect 336416 620638 336472 620672
rect 336506 620638 336562 620672
rect 336596 620638 336652 620672
rect 336686 620638 336742 620672
rect 336776 620638 336832 620672
rect 336866 620638 336927 620672
rect 336233 620630 336927 620638
rect 336233 620596 336320 620630
rect 336354 620596 336420 620630
rect 336454 620596 336520 620630
rect 336554 620596 336620 620630
rect 336654 620596 336720 620630
rect 336754 620596 336820 620630
rect 336854 620596 336927 620630
rect 336233 620582 336927 620596
rect 336233 620548 336292 620582
rect 336326 620548 336382 620582
rect 336416 620548 336472 620582
rect 336506 620548 336562 620582
rect 336596 620548 336652 620582
rect 336686 620548 336742 620582
rect 336776 620548 336832 620582
rect 336866 620548 336927 620582
rect 336233 620530 336927 620548
rect 336233 620496 336320 620530
rect 336354 620496 336420 620530
rect 336454 620496 336520 620530
rect 336554 620496 336620 620530
rect 336654 620496 336720 620530
rect 336754 620496 336820 620530
rect 336854 620496 336927 620530
rect 336233 620492 336927 620496
rect 336233 620458 336292 620492
rect 336326 620458 336382 620492
rect 336416 620458 336472 620492
rect 336506 620458 336562 620492
rect 336596 620458 336652 620492
rect 336686 620458 336742 620492
rect 336776 620458 336832 620492
rect 336866 620458 336927 620492
rect 336233 620430 336927 620458
rect 336233 620402 336320 620430
rect 336354 620402 336420 620430
rect 336233 620368 336292 620402
rect 336354 620396 336382 620402
rect 336326 620368 336382 620396
rect 336416 620396 336420 620402
rect 336454 620402 336520 620430
rect 336454 620396 336472 620402
rect 336416 620368 336472 620396
rect 336506 620396 336520 620402
rect 336554 620402 336620 620430
rect 336654 620402 336720 620430
rect 336754 620402 336820 620430
rect 336854 620402 336927 620430
rect 336554 620396 336562 620402
rect 336506 620368 336562 620396
rect 336596 620396 336620 620402
rect 336686 620396 336720 620402
rect 336776 620396 336820 620402
rect 336596 620368 336652 620396
rect 336686 620368 336742 620396
rect 336776 620368 336832 620396
rect 336866 620368 336927 620402
rect 336233 620309 336927 620368
rect 336988 620971 337008 621005
rect 337042 621004 337406 621005
rect 337042 620971 337156 621004
rect 336988 620970 337156 620971
rect 337190 620970 337257 621004
rect 337291 620990 337406 621004
rect 337440 620990 337459 621024
rect 338277 621060 338444 621065
rect 338478 621060 338545 621094
rect 338579 621084 338786 621094
rect 338820 621084 338876 621118
rect 338910 621084 338966 621118
rect 339000 621084 339056 621118
rect 339090 621084 339146 621118
rect 339180 621084 339236 621118
rect 339270 621084 339326 621118
rect 339360 621084 339416 621118
rect 339450 621084 339506 621118
rect 339540 621094 340074 621118
rect 339540 621084 339732 621094
rect 338579 621065 339732 621084
rect 338579 621060 338747 621065
rect 338277 621024 338747 621060
rect 338277 621005 338694 621024
rect 337291 620970 337459 620990
rect 336988 620934 337459 620970
rect 336988 620915 337406 620934
rect 336988 620881 337008 620915
rect 337042 620914 337406 620915
rect 337042 620881 337156 620914
rect 336988 620880 337156 620881
rect 337190 620880 337257 620914
rect 337291 620900 337406 620914
rect 337440 620900 337459 620934
rect 337291 620880 337459 620900
rect 336988 620844 337459 620880
rect 336988 620825 337406 620844
rect 336988 620791 337008 620825
rect 337042 620824 337406 620825
rect 337042 620791 337156 620824
rect 336988 620790 337156 620791
rect 337190 620790 337257 620824
rect 337291 620810 337406 620824
rect 337440 620810 337459 620844
rect 337291 620790 337459 620810
rect 336988 620754 337459 620790
rect 336988 620735 337406 620754
rect 336988 620701 337008 620735
rect 337042 620734 337406 620735
rect 337042 620701 337156 620734
rect 336988 620700 337156 620701
rect 337190 620700 337257 620734
rect 337291 620720 337406 620734
rect 337440 620720 337459 620754
rect 337291 620700 337459 620720
rect 336988 620664 337459 620700
rect 336988 620645 337406 620664
rect 336988 620611 337008 620645
rect 337042 620644 337406 620645
rect 337042 620611 337156 620644
rect 336988 620610 337156 620611
rect 337190 620610 337257 620644
rect 337291 620630 337406 620644
rect 337440 620630 337459 620664
rect 337291 620610 337459 620630
rect 336988 620574 337459 620610
rect 336988 620555 337406 620574
rect 336988 620521 337008 620555
rect 337042 620554 337406 620555
rect 337042 620521 337156 620554
rect 336988 620520 337156 620521
rect 337190 620520 337257 620554
rect 337291 620540 337406 620554
rect 337440 620540 337459 620574
rect 337291 620520 337459 620540
rect 336988 620484 337459 620520
rect 336988 620465 337406 620484
rect 336988 620431 337008 620465
rect 337042 620464 337406 620465
rect 337042 620431 337156 620464
rect 336988 620430 337156 620431
rect 337190 620430 337257 620464
rect 337291 620450 337406 620464
rect 337440 620450 337459 620484
rect 337291 620430 337459 620450
rect 336988 620394 337459 620430
rect 336988 620375 337406 620394
rect 336988 620341 337008 620375
rect 337042 620374 337406 620375
rect 337042 620341 337156 620374
rect 336988 620340 337156 620341
rect 337190 620340 337257 620374
rect 337291 620360 337406 620374
rect 337440 620360 337459 620394
rect 337291 620340 337459 620360
rect 335688 620285 336118 620304
rect 335688 620251 335720 620285
rect 335754 620284 336118 620285
rect 335754 620251 335868 620284
rect 335688 620250 335868 620251
rect 335902 620250 335969 620284
rect 336003 620270 336118 620284
rect 336152 620270 336188 620304
rect 336003 620250 336188 620270
rect 335688 620247 336188 620250
rect 336988 620304 337459 620340
rect 337521 620942 338215 621003
rect 337521 620908 337580 620942
rect 337614 620930 337670 620942
rect 337642 620908 337670 620930
rect 337704 620930 337760 620942
rect 337704 620908 337708 620930
rect 337521 620896 337608 620908
rect 337642 620896 337708 620908
rect 337742 620908 337760 620930
rect 337794 620930 337850 620942
rect 337794 620908 337808 620930
rect 337742 620896 337808 620908
rect 337842 620908 337850 620930
rect 337884 620930 337940 620942
rect 337974 620930 338030 620942
rect 338064 620930 338120 620942
rect 337884 620908 337908 620930
rect 337974 620908 338008 620930
rect 338064 620908 338108 620930
rect 338154 620908 338215 620942
rect 337842 620896 337908 620908
rect 337942 620896 338008 620908
rect 338042 620896 338108 620908
rect 338142 620896 338215 620908
rect 337521 620852 338215 620896
rect 337521 620818 337580 620852
rect 337614 620830 337670 620852
rect 337642 620818 337670 620830
rect 337704 620830 337760 620852
rect 337704 620818 337708 620830
rect 337521 620796 337608 620818
rect 337642 620796 337708 620818
rect 337742 620818 337760 620830
rect 337794 620830 337850 620852
rect 337794 620818 337808 620830
rect 337742 620796 337808 620818
rect 337842 620818 337850 620830
rect 337884 620830 337940 620852
rect 337974 620830 338030 620852
rect 338064 620830 338120 620852
rect 337884 620818 337908 620830
rect 337974 620818 338008 620830
rect 338064 620818 338108 620830
rect 338154 620818 338215 620852
rect 337842 620796 337908 620818
rect 337942 620796 338008 620818
rect 338042 620796 338108 620818
rect 338142 620796 338215 620818
rect 337521 620762 338215 620796
rect 337521 620728 337580 620762
rect 337614 620730 337670 620762
rect 337642 620728 337670 620730
rect 337704 620730 337760 620762
rect 337704 620728 337708 620730
rect 337521 620696 337608 620728
rect 337642 620696 337708 620728
rect 337742 620728 337760 620730
rect 337794 620730 337850 620762
rect 337794 620728 337808 620730
rect 337742 620696 337808 620728
rect 337842 620728 337850 620730
rect 337884 620730 337940 620762
rect 337974 620730 338030 620762
rect 338064 620730 338120 620762
rect 337884 620728 337908 620730
rect 337974 620728 338008 620730
rect 338064 620728 338108 620730
rect 338154 620728 338215 620762
rect 337842 620696 337908 620728
rect 337942 620696 338008 620728
rect 338042 620696 338108 620728
rect 338142 620696 338215 620728
rect 337521 620672 338215 620696
rect 337521 620638 337580 620672
rect 337614 620638 337670 620672
rect 337704 620638 337760 620672
rect 337794 620638 337850 620672
rect 337884 620638 337940 620672
rect 337974 620638 338030 620672
rect 338064 620638 338120 620672
rect 338154 620638 338215 620672
rect 337521 620630 338215 620638
rect 337521 620596 337608 620630
rect 337642 620596 337708 620630
rect 337742 620596 337808 620630
rect 337842 620596 337908 620630
rect 337942 620596 338008 620630
rect 338042 620596 338108 620630
rect 338142 620596 338215 620630
rect 337521 620582 338215 620596
rect 337521 620548 337580 620582
rect 337614 620548 337670 620582
rect 337704 620548 337760 620582
rect 337794 620548 337850 620582
rect 337884 620548 337940 620582
rect 337974 620548 338030 620582
rect 338064 620548 338120 620582
rect 338154 620548 338215 620582
rect 337521 620530 338215 620548
rect 337521 620496 337608 620530
rect 337642 620496 337708 620530
rect 337742 620496 337808 620530
rect 337842 620496 337908 620530
rect 337942 620496 338008 620530
rect 338042 620496 338108 620530
rect 338142 620496 338215 620530
rect 337521 620492 338215 620496
rect 337521 620458 337580 620492
rect 337614 620458 337670 620492
rect 337704 620458 337760 620492
rect 337794 620458 337850 620492
rect 337884 620458 337940 620492
rect 337974 620458 338030 620492
rect 338064 620458 338120 620492
rect 338154 620458 338215 620492
rect 337521 620430 338215 620458
rect 337521 620402 337608 620430
rect 337642 620402 337708 620430
rect 337521 620368 337580 620402
rect 337642 620396 337670 620402
rect 337614 620368 337670 620396
rect 337704 620396 337708 620402
rect 337742 620402 337808 620430
rect 337742 620396 337760 620402
rect 337704 620368 337760 620396
rect 337794 620396 337808 620402
rect 337842 620402 337908 620430
rect 337942 620402 338008 620430
rect 338042 620402 338108 620430
rect 338142 620402 338215 620430
rect 337842 620396 337850 620402
rect 337794 620368 337850 620396
rect 337884 620396 337908 620402
rect 337974 620396 338008 620402
rect 338064 620396 338108 620402
rect 337884 620368 337940 620396
rect 337974 620368 338030 620396
rect 338064 620368 338120 620396
rect 338154 620368 338215 620402
rect 337521 620309 338215 620368
rect 338277 620971 338296 621005
rect 338330 621004 338694 621005
rect 338330 620971 338444 621004
rect 338277 620970 338444 620971
rect 338478 620970 338545 621004
rect 338579 620990 338694 621004
rect 338728 620990 338747 621024
rect 339565 621060 339732 621065
rect 339766 621060 339833 621094
rect 339867 621084 340074 621094
rect 340108 621084 340164 621118
rect 340198 621084 340254 621118
rect 340288 621084 340344 621118
rect 340378 621084 340434 621118
rect 340468 621084 340524 621118
rect 340558 621084 340614 621118
rect 340648 621084 340704 621118
rect 340738 621084 340794 621118
rect 340828 621094 341088 621118
rect 340828 621084 341020 621094
rect 339867 621065 341020 621084
rect 339867 621060 340035 621065
rect 339565 621024 340035 621060
rect 339565 621005 339982 621024
rect 338579 620970 338747 620990
rect 338277 620934 338747 620970
rect 338277 620915 338694 620934
rect 338277 620881 338296 620915
rect 338330 620914 338694 620915
rect 338330 620881 338444 620914
rect 338277 620880 338444 620881
rect 338478 620880 338545 620914
rect 338579 620900 338694 620914
rect 338728 620900 338747 620934
rect 338579 620880 338747 620900
rect 338277 620844 338747 620880
rect 338277 620825 338694 620844
rect 338277 620791 338296 620825
rect 338330 620824 338694 620825
rect 338330 620791 338444 620824
rect 338277 620790 338444 620791
rect 338478 620790 338545 620824
rect 338579 620810 338694 620824
rect 338728 620810 338747 620844
rect 338579 620790 338747 620810
rect 338277 620754 338747 620790
rect 338277 620735 338694 620754
rect 338277 620701 338296 620735
rect 338330 620734 338694 620735
rect 338330 620701 338444 620734
rect 338277 620700 338444 620701
rect 338478 620700 338545 620734
rect 338579 620720 338694 620734
rect 338728 620720 338747 620754
rect 338579 620700 338747 620720
rect 338277 620664 338747 620700
rect 338277 620645 338694 620664
rect 338277 620611 338296 620645
rect 338330 620644 338694 620645
rect 338330 620611 338444 620644
rect 338277 620610 338444 620611
rect 338478 620610 338545 620644
rect 338579 620630 338694 620644
rect 338728 620630 338747 620664
rect 338579 620610 338747 620630
rect 338277 620574 338747 620610
rect 338277 620555 338694 620574
rect 338277 620521 338296 620555
rect 338330 620554 338694 620555
rect 338330 620521 338444 620554
rect 338277 620520 338444 620521
rect 338478 620520 338545 620554
rect 338579 620540 338694 620554
rect 338728 620540 338747 620574
rect 338579 620520 338747 620540
rect 338277 620484 338747 620520
rect 338277 620465 338694 620484
rect 338277 620431 338296 620465
rect 338330 620464 338694 620465
rect 338330 620431 338444 620464
rect 338277 620430 338444 620431
rect 338478 620430 338545 620464
rect 338579 620450 338694 620464
rect 338728 620450 338747 620484
rect 338579 620430 338747 620450
rect 338277 620394 338747 620430
rect 338277 620375 338694 620394
rect 338277 620341 338296 620375
rect 338330 620374 338694 620375
rect 338330 620341 338444 620374
rect 338277 620340 338444 620341
rect 338478 620340 338545 620374
rect 338579 620360 338694 620374
rect 338728 620360 338747 620394
rect 338579 620340 338747 620360
rect 336988 620285 337406 620304
rect 336988 620251 337008 620285
rect 337042 620284 337406 620285
rect 337042 620251 337156 620284
rect 336988 620250 337156 620251
rect 337190 620250 337257 620284
rect 337291 620270 337406 620284
rect 337440 620270 337459 620304
rect 337291 620250 337459 620270
rect 336988 620247 337459 620250
rect 338277 620304 338747 620340
rect 338809 620942 339503 621003
rect 338809 620908 338868 620942
rect 338902 620930 338958 620942
rect 338930 620908 338958 620930
rect 338992 620930 339048 620942
rect 338992 620908 338996 620930
rect 338809 620896 338896 620908
rect 338930 620896 338996 620908
rect 339030 620908 339048 620930
rect 339082 620930 339138 620942
rect 339082 620908 339096 620930
rect 339030 620896 339096 620908
rect 339130 620908 339138 620930
rect 339172 620930 339228 620942
rect 339262 620930 339318 620942
rect 339352 620930 339408 620942
rect 339172 620908 339196 620930
rect 339262 620908 339296 620930
rect 339352 620908 339396 620930
rect 339442 620908 339503 620942
rect 339130 620896 339196 620908
rect 339230 620896 339296 620908
rect 339330 620896 339396 620908
rect 339430 620896 339503 620908
rect 338809 620852 339503 620896
rect 338809 620818 338868 620852
rect 338902 620830 338958 620852
rect 338930 620818 338958 620830
rect 338992 620830 339048 620852
rect 338992 620818 338996 620830
rect 338809 620796 338896 620818
rect 338930 620796 338996 620818
rect 339030 620818 339048 620830
rect 339082 620830 339138 620852
rect 339082 620818 339096 620830
rect 339030 620796 339096 620818
rect 339130 620818 339138 620830
rect 339172 620830 339228 620852
rect 339262 620830 339318 620852
rect 339352 620830 339408 620852
rect 339172 620818 339196 620830
rect 339262 620818 339296 620830
rect 339352 620818 339396 620830
rect 339442 620818 339503 620852
rect 339130 620796 339196 620818
rect 339230 620796 339296 620818
rect 339330 620796 339396 620818
rect 339430 620796 339503 620818
rect 338809 620762 339503 620796
rect 338809 620728 338868 620762
rect 338902 620730 338958 620762
rect 338930 620728 338958 620730
rect 338992 620730 339048 620762
rect 338992 620728 338996 620730
rect 338809 620696 338896 620728
rect 338930 620696 338996 620728
rect 339030 620728 339048 620730
rect 339082 620730 339138 620762
rect 339082 620728 339096 620730
rect 339030 620696 339096 620728
rect 339130 620728 339138 620730
rect 339172 620730 339228 620762
rect 339262 620730 339318 620762
rect 339352 620730 339408 620762
rect 339172 620728 339196 620730
rect 339262 620728 339296 620730
rect 339352 620728 339396 620730
rect 339442 620728 339503 620762
rect 339130 620696 339196 620728
rect 339230 620696 339296 620728
rect 339330 620696 339396 620728
rect 339430 620696 339503 620728
rect 338809 620672 339503 620696
rect 338809 620638 338868 620672
rect 338902 620638 338958 620672
rect 338992 620638 339048 620672
rect 339082 620638 339138 620672
rect 339172 620638 339228 620672
rect 339262 620638 339318 620672
rect 339352 620638 339408 620672
rect 339442 620638 339503 620672
rect 338809 620630 339503 620638
rect 338809 620596 338896 620630
rect 338930 620596 338996 620630
rect 339030 620596 339096 620630
rect 339130 620596 339196 620630
rect 339230 620596 339296 620630
rect 339330 620596 339396 620630
rect 339430 620596 339503 620630
rect 338809 620582 339503 620596
rect 338809 620548 338868 620582
rect 338902 620548 338958 620582
rect 338992 620548 339048 620582
rect 339082 620548 339138 620582
rect 339172 620548 339228 620582
rect 339262 620548 339318 620582
rect 339352 620548 339408 620582
rect 339442 620548 339503 620582
rect 338809 620530 339503 620548
rect 338809 620496 338896 620530
rect 338930 620496 338996 620530
rect 339030 620496 339096 620530
rect 339130 620496 339196 620530
rect 339230 620496 339296 620530
rect 339330 620496 339396 620530
rect 339430 620496 339503 620530
rect 338809 620492 339503 620496
rect 338809 620458 338868 620492
rect 338902 620458 338958 620492
rect 338992 620458 339048 620492
rect 339082 620458 339138 620492
rect 339172 620458 339228 620492
rect 339262 620458 339318 620492
rect 339352 620458 339408 620492
rect 339442 620458 339503 620492
rect 338809 620430 339503 620458
rect 338809 620402 338896 620430
rect 338930 620402 338996 620430
rect 338809 620368 338868 620402
rect 338930 620396 338958 620402
rect 338902 620368 338958 620396
rect 338992 620396 338996 620402
rect 339030 620402 339096 620430
rect 339030 620396 339048 620402
rect 338992 620368 339048 620396
rect 339082 620396 339096 620402
rect 339130 620402 339196 620430
rect 339230 620402 339296 620430
rect 339330 620402 339396 620430
rect 339430 620402 339503 620430
rect 339130 620396 339138 620402
rect 339082 620368 339138 620396
rect 339172 620396 339196 620402
rect 339262 620396 339296 620402
rect 339352 620396 339396 620402
rect 339172 620368 339228 620396
rect 339262 620368 339318 620396
rect 339352 620368 339408 620396
rect 339442 620368 339503 620402
rect 338809 620309 339503 620368
rect 339565 620971 339584 621005
rect 339618 621004 339982 621005
rect 339618 620971 339732 621004
rect 339565 620970 339732 620971
rect 339766 620970 339833 621004
rect 339867 620990 339982 621004
rect 340016 620990 340035 621024
rect 340853 621060 341020 621065
rect 341054 621060 341088 621094
rect 340853 621005 341088 621060
rect 339867 620970 340035 620990
rect 339565 620934 340035 620970
rect 339565 620915 339982 620934
rect 339565 620881 339584 620915
rect 339618 620914 339982 620915
rect 339618 620881 339732 620914
rect 339565 620880 339732 620881
rect 339766 620880 339833 620914
rect 339867 620900 339982 620914
rect 340016 620900 340035 620934
rect 339867 620880 340035 620900
rect 339565 620844 340035 620880
rect 339565 620825 339982 620844
rect 339565 620791 339584 620825
rect 339618 620824 339982 620825
rect 339618 620791 339732 620824
rect 339565 620790 339732 620791
rect 339766 620790 339833 620824
rect 339867 620810 339982 620824
rect 340016 620810 340035 620844
rect 339867 620790 340035 620810
rect 339565 620754 340035 620790
rect 339565 620735 339982 620754
rect 339565 620701 339584 620735
rect 339618 620734 339982 620735
rect 339618 620701 339732 620734
rect 339565 620700 339732 620701
rect 339766 620700 339833 620734
rect 339867 620720 339982 620734
rect 340016 620720 340035 620754
rect 339867 620700 340035 620720
rect 339565 620664 340035 620700
rect 339565 620645 339982 620664
rect 339565 620611 339584 620645
rect 339618 620644 339982 620645
rect 339618 620611 339732 620644
rect 339565 620610 339732 620611
rect 339766 620610 339833 620644
rect 339867 620630 339982 620644
rect 340016 620630 340035 620664
rect 339867 620610 340035 620630
rect 339565 620574 340035 620610
rect 339565 620555 339982 620574
rect 339565 620521 339584 620555
rect 339618 620554 339982 620555
rect 339618 620521 339732 620554
rect 339565 620520 339732 620521
rect 339766 620520 339833 620554
rect 339867 620540 339982 620554
rect 340016 620540 340035 620574
rect 339867 620520 340035 620540
rect 339565 620484 340035 620520
rect 339565 620465 339982 620484
rect 339565 620431 339584 620465
rect 339618 620464 339982 620465
rect 339618 620431 339732 620464
rect 339565 620430 339732 620431
rect 339766 620430 339833 620464
rect 339867 620450 339982 620464
rect 340016 620450 340035 620484
rect 339867 620430 340035 620450
rect 339565 620394 340035 620430
rect 339565 620375 339982 620394
rect 339565 620341 339584 620375
rect 339618 620374 339982 620375
rect 339618 620341 339732 620374
rect 339565 620340 339732 620341
rect 339766 620340 339833 620374
rect 339867 620360 339982 620374
rect 340016 620360 340035 620394
rect 339867 620340 340035 620360
rect 338277 620285 338694 620304
rect 338277 620251 338296 620285
rect 338330 620284 338694 620285
rect 338330 620251 338444 620284
rect 338277 620250 338444 620251
rect 338478 620250 338545 620284
rect 338579 620270 338694 620284
rect 338728 620270 338747 620304
rect 338579 620250 338747 620270
rect 338277 620247 338747 620250
rect 339565 620304 340035 620340
rect 340097 620942 340791 621003
rect 340097 620908 340156 620942
rect 340190 620930 340246 620942
rect 340218 620908 340246 620930
rect 340280 620930 340336 620942
rect 340280 620908 340284 620930
rect 340097 620896 340184 620908
rect 340218 620896 340284 620908
rect 340318 620908 340336 620930
rect 340370 620930 340426 620942
rect 340370 620908 340384 620930
rect 340318 620896 340384 620908
rect 340418 620908 340426 620930
rect 340460 620930 340516 620942
rect 340550 620930 340606 620942
rect 340640 620930 340696 620942
rect 340460 620908 340484 620930
rect 340550 620908 340584 620930
rect 340640 620908 340684 620930
rect 340730 620908 340791 620942
rect 340418 620896 340484 620908
rect 340518 620896 340584 620908
rect 340618 620896 340684 620908
rect 340718 620896 340791 620908
rect 340097 620852 340791 620896
rect 340097 620818 340156 620852
rect 340190 620830 340246 620852
rect 340218 620818 340246 620830
rect 340280 620830 340336 620852
rect 340280 620818 340284 620830
rect 340097 620796 340184 620818
rect 340218 620796 340284 620818
rect 340318 620818 340336 620830
rect 340370 620830 340426 620852
rect 340370 620818 340384 620830
rect 340318 620796 340384 620818
rect 340418 620818 340426 620830
rect 340460 620830 340516 620852
rect 340550 620830 340606 620852
rect 340640 620830 340696 620852
rect 340460 620818 340484 620830
rect 340550 620818 340584 620830
rect 340640 620818 340684 620830
rect 340730 620818 340791 620852
rect 340418 620796 340484 620818
rect 340518 620796 340584 620818
rect 340618 620796 340684 620818
rect 340718 620796 340791 620818
rect 340097 620762 340791 620796
rect 340097 620728 340156 620762
rect 340190 620730 340246 620762
rect 340218 620728 340246 620730
rect 340280 620730 340336 620762
rect 340280 620728 340284 620730
rect 340097 620696 340184 620728
rect 340218 620696 340284 620728
rect 340318 620728 340336 620730
rect 340370 620730 340426 620762
rect 340370 620728 340384 620730
rect 340318 620696 340384 620728
rect 340418 620728 340426 620730
rect 340460 620730 340516 620762
rect 340550 620730 340606 620762
rect 340640 620730 340696 620762
rect 340460 620728 340484 620730
rect 340550 620728 340584 620730
rect 340640 620728 340684 620730
rect 340730 620728 340791 620762
rect 340418 620696 340484 620728
rect 340518 620696 340584 620728
rect 340618 620696 340684 620728
rect 340718 620696 340791 620728
rect 340097 620672 340791 620696
rect 340097 620638 340156 620672
rect 340190 620638 340246 620672
rect 340280 620638 340336 620672
rect 340370 620638 340426 620672
rect 340460 620638 340516 620672
rect 340550 620638 340606 620672
rect 340640 620638 340696 620672
rect 340730 620638 340791 620672
rect 340097 620630 340791 620638
rect 340097 620596 340184 620630
rect 340218 620596 340284 620630
rect 340318 620596 340384 620630
rect 340418 620596 340484 620630
rect 340518 620596 340584 620630
rect 340618 620596 340684 620630
rect 340718 620596 340791 620630
rect 340097 620582 340791 620596
rect 340097 620548 340156 620582
rect 340190 620548 340246 620582
rect 340280 620548 340336 620582
rect 340370 620548 340426 620582
rect 340460 620548 340516 620582
rect 340550 620548 340606 620582
rect 340640 620548 340696 620582
rect 340730 620548 340791 620582
rect 340097 620530 340791 620548
rect 340097 620496 340184 620530
rect 340218 620496 340284 620530
rect 340318 620496 340384 620530
rect 340418 620496 340484 620530
rect 340518 620496 340584 620530
rect 340618 620496 340684 620530
rect 340718 620496 340791 620530
rect 340097 620492 340791 620496
rect 340097 620458 340156 620492
rect 340190 620458 340246 620492
rect 340280 620458 340336 620492
rect 340370 620458 340426 620492
rect 340460 620458 340516 620492
rect 340550 620458 340606 620492
rect 340640 620458 340696 620492
rect 340730 620458 340791 620492
rect 340097 620430 340791 620458
rect 340097 620402 340184 620430
rect 340218 620402 340284 620430
rect 340097 620368 340156 620402
rect 340218 620396 340246 620402
rect 340190 620368 340246 620396
rect 340280 620396 340284 620402
rect 340318 620402 340384 620430
rect 340318 620396 340336 620402
rect 340280 620368 340336 620396
rect 340370 620396 340384 620402
rect 340418 620402 340484 620430
rect 340518 620402 340584 620430
rect 340618 620402 340684 620430
rect 340718 620402 340791 620430
rect 340418 620396 340426 620402
rect 340370 620368 340426 620396
rect 340460 620396 340484 620402
rect 340550 620396 340584 620402
rect 340640 620396 340684 620402
rect 340460 620368 340516 620396
rect 340550 620368 340606 620396
rect 340640 620368 340696 620396
rect 340730 620368 340791 620402
rect 340097 620309 340791 620368
rect 340853 620971 340872 621005
rect 340906 621004 341088 621005
rect 340906 620971 341020 621004
rect 340853 620970 341020 620971
rect 341054 620970 341088 621004
rect 340853 620915 341088 620970
rect 340853 620881 340872 620915
rect 340906 620914 341088 620915
rect 340906 620881 341020 620914
rect 340853 620880 341020 620881
rect 341054 620880 341088 620914
rect 340853 620825 341088 620880
rect 340853 620791 340872 620825
rect 340906 620824 341088 620825
rect 340906 620791 341020 620824
rect 340853 620790 341020 620791
rect 341054 620790 341088 620824
rect 340853 620735 341088 620790
rect 340853 620701 340872 620735
rect 340906 620734 341088 620735
rect 340906 620701 341020 620734
rect 340853 620700 341020 620701
rect 341054 620700 341088 620734
rect 340853 620645 341088 620700
rect 340853 620611 340872 620645
rect 340906 620644 341088 620645
rect 340906 620611 341020 620644
rect 340853 620610 341020 620611
rect 341054 620610 341088 620644
rect 340853 620555 341088 620610
rect 340853 620521 340872 620555
rect 340906 620554 341088 620555
rect 340906 620521 341020 620554
rect 340853 620520 341020 620521
rect 341054 620520 341088 620554
rect 340853 620465 341088 620520
rect 340853 620431 340872 620465
rect 340906 620464 341088 620465
rect 340906 620431 341020 620464
rect 340853 620430 341020 620431
rect 341054 620430 341088 620464
rect 340853 620375 341088 620430
rect 340853 620341 340872 620375
rect 340906 620374 341088 620375
rect 340906 620341 341020 620374
rect 340853 620340 341020 620341
rect 341054 620340 341088 620374
rect 339565 620285 339982 620304
rect 339565 620251 339584 620285
rect 339618 620284 339982 620285
rect 339618 620251 339732 620284
rect 339565 620250 339732 620251
rect 339766 620250 339833 620284
rect 339867 620270 339982 620284
rect 340016 620270 340035 620304
rect 339867 620250 340035 620270
rect 339565 620247 340035 620250
rect 340853 620285 341088 620340
rect 340853 620251 340872 620285
rect 340906 620284 341088 620285
rect 340906 620251 341020 620284
rect 340853 620250 341020 620251
rect 341054 620250 341088 620284
rect 340853 620247 341088 620250
rect 334648 620228 341088 620247
rect 334648 620194 334888 620228
rect 334922 620194 334978 620228
rect 335012 620194 335068 620228
rect 335102 620194 335158 620228
rect 335192 620194 335248 620228
rect 335282 620194 335338 620228
rect 335372 620194 335428 620228
rect 335462 620194 335518 620228
rect 335552 620194 335608 620228
rect 335642 620194 336176 620228
rect 336210 620194 336266 620228
rect 336300 620194 336356 620228
rect 336390 620194 336446 620228
rect 336480 620194 336536 620228
rect 336570 620194 336626 620228
rect 336660 620194 336716 620228
rect 336750 620194 336806 620228
rect 336840 620194 336896 620228
rect 336930 620194 337464 620228
rect 337498 620194 337554 620228
rect 337588 620194 337644 620228
rect 337678 620194 337734 620228
rect 337768 620194 337824 620228
rect 337858 620194 337914 620228
rect 337948 620194 338004 620228
rect 338038 620194 338094 620228
rect 338128 620194 338184 620228
rect 338218 620194 338752 620228
rect 338786 620194 338842 620228
rect 338876 620194 338932 620228
rect 338966 620194 339022 620228
rect 339056 620194 339112 620228
rect 339146 620194 339202 620228
rect 339236 620194 339292 620228
rect 339326 620194 339382 620228
rect 339416 620194 339472 620228
rect 339506 620194 340040 620228
rect 340074 620194 340130 620228
rect 340164 620194 340220 620228
rect 340254 620194 340310 620228
rect 340344 620194 340400 620228
rect 340434 620194 340490 620228
rect 340524 620194 340580 620228
rect 340614 620194 340670 620228
rect 340704 620194 340760 620228
rect 340794 620194 341088 620228
rect 334648 620160 334681 620194
rect 334715 620175 335868 620194
rect 334715 620160 334888 620175
rect 334648 620111 334888 620160
rect 335688 620160 335868 620175
rect 335902 620160 335969 620194
rect 336003 620175 337156 620194
rect 336003 620160 336188 620175
rect 335688 620111 336188 620160
rect 336988 620160 337156 620175
rect 337190 620160 337257 620194
rect 337291 620175 338444 620194
rect 337291 620160 337388 620175
rect 336988 620111 337388 620160
rect 338288 620160 338444 620175
rect 338478 620160 338545 620194
rect 338579 620175 339732 620194
rect 338579 620160 338688 620175
rect 338288 620111 338688 620160
rect 339588 620160 339732 620175
rect 339766 620160 339833 620194
rect 339867 620175 341020 620194
rect 339867 620160 339988 620175
rect 339588 620111 339988 620160
rect 340888 620160 341020 620175
rect 341054 620160 341088 620194
rect 340888 620111 341088 620160
rect 334648 620104 341088 620111
rect 334648 620070 334681 620104
rect 334715 620081 335868 620104
rect 334715 620070 334782 620081
rect 334648 620047 334782 620070
rect 334816 620047 334872 620081
rect 334906 620047 334962 620081
rect 334996 620047 335052 620081
rect 335086 620047 335142 620081
rect 335176 620047 335232 620081
rect 335266 620047 335322 620081
rect 335356 620047 335412 620081
rect 335446 620047 335502 620081
rect 335536 620047 335592 620081
rect 335626 620047 335682 620081
rect 335716 620047 335772 620081
rect 335806 620070 335868 620081
rect 335902 620070 335969 620104
rect 336003 620081 337156 620104
rect 336003 620070 336070 620081
rect 335806 620047 336070 620070
rect 336104 620047 336160 620081
rect 336194 620047 336250 620081
rect 336284 620047 336340 620081
rect 336374 620047 336430 620081
rect 336464 620047 336520 620081
rect 336554 620047 336610 620081
rect 336644 620047 336700 620081
rect 336734 620047 336790 620081
rect 336824 620047 336880 620081
rect 336914 620047 336970 620081
rect 337004 620047 337060 620081
rect 337094 620070 337156 620081
rect 337190 620070 337257 620104
rect 337291 620081 338444 620104
rect 337291 620070 337358 620081
rect 337094 620047 337358 620070
rect 337392 620047 337448 620081
rect 337482 620047 337538 620081
rect 337572 620047 337628 620081
rect 337662 620047 337718 620081
rect 337752 620047 337808 620081
rect 337842 620047 337898 620081
rect 337932 620047 337988 620081
rect 338022 620047 338078 620081
rect 338112 620047 338168 620081
rect 338202 620047 338258 620081
rect 338292 620047 338348 620081
rect 338382 620070 338444 620081
rect 338478 620070 338545 620104
rect 338579 620081 339732 620104
rect 338579 620070 338646 620081
rect 338382 620047 338646 620070
rect 338680 620047 338736 620081
rect 338770 620047 338826 620081
rect 338860 620047 338916 620081
rect 338950 620047 339006 620081
rect 339040 620047 339096 620081
rect 339130 620047 339186 620081
rect 339220 620047 339276 620081
rect 339310 620047 339366 620081
rect 339400 620047 339456 620081
rect 339490 620047 339546 620081
rect 339580 620047 339636 620081
rect 339670 620070 339732 620081
rect 339766 620070 339833 620104
rect 339867 620081 341020 620104
rect 339867 620070 339934 620081
rect 339670 620047 339934 620070
rect 339968 620047 340024 620081
rect 340058 620047 340114 620081
rect 340148 620047 340204 620081
rect 340238 620047 340294 620081
rect 340328 620047 340384 620081
rect 340418 620047 340474 620081
rect 340508 620047 340564 620081
rect 340598 620047 340654 620081
rect 340688 620047 340744 620081
rect 340778 620047 340834 620081
rect 340868 620047 340924 620081
rect 340958 620070 341020 620081
rect 341054 620070 341088 620104
rect 340958 620047 341088 620070
rect 334648 619980 341088 620047
rect 334648 619946 334782 619980
rect 334816 619946 334872 619980
rect 334906 619946 334962 619980
rect 334996 619946 335052 619980
rect 335086 619946 335142 619980
rect 335176 619946 335232 619980
rect 335266 619946 335322 619980
rect 335356 619946 335412 619980
rect 335446 619946 335502 619980
rect 335536 619946 335592 619980
rect 335626 619946 335682 619980
rect 335716 619946 335772 619980
rect 335806 619946 336070 619980
rect 336104 619946 336160 619980
rect 336194 619946 336250 619980
rect 336284 619946 336340 619980
rect 336374 619946 336430 619980
rect 336464 619946 336520 619980
rect 336554 619946 336610 619980
rect 336644 619946 336700 619980
rect 336734 619946 336790 619980
rect 336824 619946 336880 619980
rect 336914 619946 336970 619980
rect 337004 619946 337060 619980
rect 337094 619946 337358 619980
rect 337392 619946 337448 619980
rect 337482 619946 337538 619980
rect 337572 619946 337628 619980
rect 337662 619946 337718 619980
rect 337752 619946 337808 619980
rect 337842 619946 337898 619980
rect 337932 619946 337988 619980
rect 338022 619946 338078 619980
rect 338112 619946 338168 619980
rect 338202 619946 338258 619980
rect 338292 619946 338348 619980
rect 338382 619946 338646 619980
rect 338680 619946 338736 619980
rect 338770 619946 338826 619980
rect 338860 619946 338916 619980
rect 338950 619946 339006 619980
rect 339040 619946 339096 619980
rect 339130 619946 339186 619980
rect 339220 619946 339276 619980
rect 339310 619946 339366 619980
rect 339400 619946 339456 619980
rect 339490 619946 339546 619980
rect 339580 619946 339636 619980
rect 339670 619946 339934 619980
rect 339968 619946 340024 619980
rect 340058 619946 340114 619980
rect 340148 619946 340204 619980
rect 340238 619946 340294 619980
rect 340328 619946 340384 619980
rect 340418 619946 340474 619980
rect 340508 619946 340564 619980
rect 340598 619946 340654 619980
rect 340688 619946 340744 619980
rect 340778 619946 340834 619980
rect 340868 619946 340924 619980
rect 340958 619946 341088 619980
rect 334648 619913 341088 619946
rect 334648 619896 334888 619913
rect 334648 619862 334681 619896
rect 334715 619862 334888 619896
rect 334648 619849 334888 619862
rect 335688 619896 336188 619913
rect 335688 619862 335868 619896
rect 335902 619862 335969 619896
rect 336003 619862 336188 619896
rect 335688 619849 336188 619862
rect 336988 619896 337388 619913
rect 336988 619862 337156 619896
rect 337190 619862 337257 619896
rect 337291 619862 337388 619896
rect 336988 619849 337388 619862
rect 338288 619896 338688 619913
rect 338288 619862 338444 619896
rect 338478 619862 338545 619896
rect 338579 619862 338688 619896
rect 338288 619849 338688 619862
rect 339588 619896 339988 619913
rect 339588 619862 339732 619896
rect 339766 619862 339833 619896
rect 339867 619862 339988 619896
rect 339588 619849 339988 619862
rect 340888 619896 341088 619913
rect 340888 619862 341020 619896
rect 341054 619862 341088 619896
rect 340888 619849 341088 619862
rect 334648 619830 341088 619849
rect 334648 619806 334922 619830
rect 334648 619772 334681 619806
rect 334715 619796 334922 619806
rect 334956 619796 335012 619830
rect 335046 619796 335102 619830
rect 335136 619796 335192 619830
rect 335226 619796 335282 619830
rect 335316 619796 335372 619830
rect 335406 619796 335462 619830
rect 335496 619796 335552 619830
rect 335586 619796 335642 619830
rect 335676 619806 336210 619830
rect 335676 619796 335868 619806
rect 334715 619777 335868 619796
rect 334715 619772 334888 619777
rect 334648 619736 334888 619772
rect 334648 619716 334830 619736
rect 334648 619682 334681 619716
rect 334715 619702 334830 619716
rect 334864 619702 334888 619736
rect 335688 619772 335868 619777
rect 335902 619772 335969 619806
rect 336003 619796 336210 619806
rect 336244 619796 336300 619830
rect 336334 619796 336390 619830
rect 336424 619796 336480 619830
rect 336514 619796 336570 619830
rect 336604 619796 336660 619830
rect 336694 619796 336750 619830
rect 336784 619796 336840 619830
rect 336874 619796 336930 619830
rect 336964 619806 337498 619830
rect 336964 619796 337156 619806
rect 336003 619777 337156 619796
rect 336003 619772 336188 619777
rect 335688 619736 336188 619772
rect 335688 619717 336118 619736
rect 334715 619682 334888 619702
rect 334648 619646 334888 619682
rect 334648 619626 334830 619646
rect 334648 619592 334681 619626
rect 334715 619612 334830 619626
rect 334864 619612 334888 619646
rect 334715 619592 334888 619612
rect 334648 619556 334888 619592
rect 334648 619536 334830 619556
rect 334648 619502 334681 619536
rect 334715 619522 334830 619536
rect 334864 619522 334888 619556
rect 334715 619502 334888 619522
rect 334648 619466 334888 619502
rect 334648 619446 334830 619466
rect 334648 619412 334681 619446
rect 334715 619432 334830 619446
rect 334864 619432 334888 619466
rect 334715 619412 334888 619432
rect 334648 619376 334888 619412
rect 334648 619356 334830 619376
rect 334648 619322 334681 619356
rect 334715 619342 334830 619356
rect 334864 619342 334888 619376
rect 334715 619322 334888 619342
rect 334648 619286 334888 619322
rect 334648 619266 334830 619286
rect 334648 619232 334681 619266
rect 334715 619252 334830 619266
rect 334864 619252 334888 619286
rect 334715 619232 334888 619252
rect 334648 619196 334888 619232
rect 334648 619176 334830 619196
rect 334648 619142 334681 619176
rect 334715 619162 334830 619176
rect 334864 619162 334888 619196
rect 334715 619142 334888 619162
rect 334648 619106 334888 619142
rect 334648 619086 334830 619106
rect 334648 619052 334681 619086
rect 334715 619072 334830 619086
rect 334864 619072 334888 619106
rect 334715 619052 334888 619072
rect 334648 619016 334888 619052
rect 334945 619654 335639 619715
rect 334945 619620 335004 619654
rect 335038 619642 335094 619654
rect 335066 619620 335094 619642
rect 335128 619642 335184 619654
rect 335128 619620 335132 619642
rect 334945 619608 335032 619620
rect 335066 619608 335132 619620
rect 335166 619620 335184 619642
rect 335218 619642 335274 619654
rect 335218 619620 335232 619642
rect 335166 619608 335232 619620
rect 335266 619620 335274 619642
rect 335308 619642 335364 619654
rect 335398 619642 335454 619654
rect 335488 619642 335544 619654
rect 335308 619620 335332 619642
rect 335398 619620 335432 619642
rect 335488 619620 335532 619642
rect 335578 619620 335639 619654
rect 335266 619608 335332 619620
rect 335366 619608 335432 619620
rect 335466 619608 335532 619620
rect 335566 619608 335639 619620
rect 334945 619564 335639 619608
rect 334945 619530 335004 619564
rect 335038 619542 335094 619564
rect 335066 619530 335094 619542
rect 335128 619542 335184 619564
rect 335128 619530 335132 619542
rect 334945 619508 335032 619530
rect 335066 619508 335132 619530
rect 335166 619530 335184 619542
rect 335218 619542 335274 619564
rect 335218 619530 335232 619542
rect 335166 619508 335232 619530
rect 335266 619530 335274 619542
rect 335308 619542 335364 619564
rect 335398 619542 335454 619564
rect 335488 619542 335544 619564
rect 335308 619530 335332 619542
rect 335398 619530 335432 619542
rect 335488 619530 335532 619542
rect 335578 619530 335639 619564
rect 335266 619508 335332 619530
rect 335366 619508 335432 619530
rect 335466 619508 335532 619530
rect 335566 619508 335639 619530
rect 334945 619474 335639 619508
rect 334945 619440 335004 619474
rect 335038 619442 335094 619474
rect 335066 619440 335094 619442
rect 335128 619442 335184 619474
rect 335128 619440 335132 619442
rect 334945 619408 335032 619440
rect 335066 619408 335132 619440
rect 335166 619440 335184 619442
rect 335218 619442 335274 619474
rect 335218 619440 335232 619442
rect 335166 619408 335232 619440
rect 335266 619440 335274 619442
rect 335308 619442 335364 619474
rect 335398 619442 335454 619474
rect 335488 619442 335544 619474
rect 335308 619440 335332 619442
rect 335398 619440 335432 619442
rect 335488 619440 335532 619442
rect 335578 619440 335639 619474
rect 335266 619408 335332 619440
rect 335366 619408 335432 619440
rect 335466 619408 335532 619440
rect 335566 619408 335639 619440
rect 334945 619384 335639 619408
rect 334945 619350 335004 619384
rect 335038 619350 335094 619384
rect 335128 619350 335184 619384
rect 335218 619350 335274 619384
rect 335308 619350 335364 619384
rect 335398 619350 335454 619384
rect 335488 619350 335544 619384
rect 335578 619350 335639 619384
rect 334945 619342 335639 619350
rect 334945 619308 335032 619342
rect 335066 619308 335132 619342
rect 335166 619308 335232 619342
rect 335266 619308 335332 619342
rect 335366 619308 335432 619342
rect 335466 619308 335532 619342
rect 335566 619308 335639 619342
rect 334945 619294 335639 619308
rect 334945 619260 335004 619294
rect 335038 619260 335094 619294
rect 335128 619260 335184 619294
rect 335218 619260 335274 619294
rect 335308 619260 335364 619294
rect 335398 619260 335454 619294
rect 335488 619260 335544 619294
rect 335578 619260 335639 619294
rect 334945 619242 335639 619260
rect 334945 619208 335032 619242
rect 335066 619208 335132 619242
rect 335166 619208 335232 619242
rect 335266 619208 335332 619242
rect 335366 619208 335432 619242
rect 335466 619208 335532 619242
rect 335566 619208 335639 619242
rect 334945 619204 335639 619208
rect 334945 619170 335004 619204
rect 335038 619170 335094 619204
rect 335128 619170 335184 619204
rect 335218 619170 335274 619204
rect 335308 619170 335364 619204
rect 335398 619170 335454 619204
rect 335488 619170 335544 619204
rect 335578 619170 335639 619204
rect 334945 619142 335639 619170
rect 334945 619114 335032 619142
rect 335066 619114 335132 619142
rect 334945 619080 335004 619114
rect 335066 619108 335094 619114
rect 335038 619080 335094 619108
rect 335128 619108 335132 619114
rect 335166 619114 335232 619142
rect 335166 619108 335184 619114
rect 335128 619080 335184 619108
rect 335218 619108 335232 619114
rect 335266 619114 335332 619142
rect 335366 619114 335432 619142
rect 335466 619114 335532 619142
rect 335566 619114 335639 619142
rect 335266 619108 335274 619114
rect 335218 619080 335274 619108
rect 335308 619108 335332 619114
rect 335398 619108 335432 619114
rect 335488 619108 335532 619114
rect 335308 619080 335364 619108
rect 335398 619080 335454 619108
rect 335488 619080 335544 619108
rect 335578 619080 335639 619114
rect 334945 619021 335639 619080
rect 335688 619683 335720 619717
rect 335754 619716 336118 619717
rect 335754 619683 335868 619716
rect 335688 619682 335868 619683
rect 335902 619682 335969 619716
rect 336003 619702 336118 619716
rect 336152 619702 336188 619736
rect 336988 619772 337156 619777
rect 337190 619772 337257 619806
rect 337291 619796 337498 619806
rect 337532 619796 337588 619830
rect 337622 619796 337678 619830
rect 337712 619796 337768 619830
rect 337802 619796 337858 619830
rect 337892 619796 337948 619830
rect 337982 619796 338038 619830
rect 338072 619796 338128 619830
rect 338162 619796 338218 619830
rect 338252 619806 338786 619830
rect 338252 619796 338444 619806
rect 337291 619777 338444 619796
rect 337291 619772 337459 619777
rect 336988 619736 337459 619772
rect 336988 619717 337406 619736
rect 336003 619682 336188 619702
rect 335688 619646 336188 619682
rect 335688 619627 336118 619646
rect 335688 619593 335720 619627
rect 335754 619626 336118 619627
rect 335754 619593 335868 619626
rect 335688 619592 335868 619593
rect 335902 619592 335969 619626
rect 336003 619612 336118 619626
rect 336152 619612 336188 619646
rect 336003 619592 336188 619612
rect 335688 619556 336188 619592
rect 335688 619537 336118 619556
rect 335688 619503 335720 619537
rect 335754 619536 336118 619537
rect 335754 619503 335868 619536
rect 335688 619502 335868 619503
rect 335902 619502 335969 619536
rect 336003 619522 336118 619536
rect 336152 619522 336188 619556
rect 336003 619502 336188 619522
rect 335688 619466 336188 619502
rect 335688 619447 336118 619466
rect 335688 619413 335720 619447
rect 335754 619446 336118 619447
rect 335754 619413 335868 619446
rect 335688 619412 335868 619413
rect 335902 619412 335969 619446
rect 336003 619432 336118 619446
rect 336152 619432 336188 619466
rect 336003 619412 336188 619432
rect 335688 619376 336188 619412
rect 335688 619357 336118 619376
rect 335688 619323 335720 619357
rect 335754 619356 336118 619357
rect 335754 619323 335868 619356
rect 335688 619322 335868 619323
rect 335902 619322 335969 619356
rect 336003 619342 336118 619356
rect 336152 619342 336188 619376
rect 336003 619322 336188 619342
rect 335688 619286 336188 619322
rect 335688 619267 336118 619286
rect 335688 619233 335720 619267
rect 335754 619266 336118 619267
rect 335754 619233 335868 619266
rect 335688 619232 335868 619233
rect 335902 619232 335969 619266
rect 336003 619252 336118 619266
rect 336152 619252 336188 619286
rect 336003 619232 336188 619252
rect 335688 619196 336188 619232
rect 335688 619177 336118 619196
rect 335688 619143 335720 619177
rect 335754 619176 336118 619177
rect 335754 619143 335868 619176
rect 335688 619142 335868 619143
rect 335902 619142 335969 619176
rect 336003 619162 336118 619176
rect 336152 619162 336188 619196
rect 336003 619142 336188 619162
rect 335688 619106 336188 619142
rect 335688 619087 336118 619106
rect 335688 619053 335720 619087
rect 335754 619086 336118 619087
rect 335754 619053 335868 619086
rect 335688 619052 335868 619053
rect 335902 619052 335969 619086
rect 336003 619072 336118 619086
rect 336152 619072 336188 619106
rect 336003 619052 336188 619072
rect 334648 618996 334830 619016
rect 334648 618962 334681 618996
rect 334715 618982 334830 618996
rect 334864 618982 334888 619016
rect 334715 618962 334888 618982
rect 334648 618959 334888 618962
rect 335688 619016 336188 619052
rect 336233 619654 336927 619715
rect 336233 619620 336292 619654
rect 336326 619642 336382 619654
rect 336354 619620 336382 619642
rect 336416 619642 336472 619654
rect 336416 619620 336420 619642
rect 336233 619608 336320 619620
rect 336354 619608 336420 619620
rect 336454 619620 336472 619642
rect 336506 619642 336562 619654
rect 336506 619620 336520 619642
rect 336454 619608 336520 619620
rect 336554 619620 336562 619642
rect 336596 619642 336652 619654
rect 336686 619642 336742 619654
rect 336776 619642 336832 619654
rect 336596 619620 336620 619642
rect 336686 619620 336720 619642
rect 336776 619620 336820 619642
rect 336866 619620 336927 619654
rect 336554 619608 336620 619620
rect 336654 619608 336720 619620
rect 336754 619608 336820 619620
rect 336854 619608 336927 619620
rect 336233 619564 336927 619608
rect 336233 619530 336292 619564
rect 336326 619542 336382 619564
rect 336354 619530 336382 619542
rect 336416 619542 336472 619564
rect 336416 619530 336420 619542
rect 336233 619508 336320 619530
rect 336354 619508 336420 619530
rect 336454 619530 336472 619542
rect 336506 619542 336562 619564
rect 336506 619530 336520 619542
rect 336454 619508 336520 619530
rect 336554 619530 336562 619542
rect 336596 619542 336652 619564
rect 336686 619542 336742 619564
rect 336776 619542 336832 619564
rect 336596 619530 336620 619542
rect 336686 619530 336720 619542
rect 336776 619530 336820 619542
rect 336866 619530 336927 619564
rect 336554 619508 336620 619530
rect 336654 619508 336720 619530
rect 336754 619508 336820 619530
rect 336854 619508 336927 619530
rect 336233 619474 336927 619508
rect 336233 619440 336292 619474
rect 336326 619442 336382 619474
rect 336354 619440 336382 619442
rect 336416 619442 336472 619474
rect 336416 619440 336420 619442
rect 336233 619408 336320 619440
rect 336354 619408 336420 619440
rect 336454 619440 336472 619442
rect 336506 619442 336562 619474
rect 336506 619440 336520 619442
rect 336454 619408 336520 619440
rect 336554 619440 336562 619442
rect 336596 619442 336652 619474
rect 336686 619442 336742 619474
rect 336776 619442 336832 619474
rect 336596 619440 336620 619442
rect 336686 619440 336720 619442
rect 336776 619440 336820 619442
rect 336866 619440 336927 619474
rect 336554 619408 336620 619440
rect 336654 619408 336720 619440
rect 336754 619408 336820 619440
rect 336854 619408 336927 619440
rect 336233 619384 336927 619408
rect 336233 619350 336292 619384
rect 336326 619350 336382 619384
rect 336416 619350 336472 619384
rect 336506 619350 336562 619384
rect 336596 619350 336652 619384
rect 336686 619350 336742 619384
rect 336776 619350 336832 619384
rect 336866 619350 336927 619384
rect 336233 619342 336927 619350
rect 336233 619308 336320 619342
rect 336354 619308 336420 619342
rect 336454 619308 336520 619342
rect 336554 619308 336620 619342
rect 336654 619308 336720 619342
rect 336754 619308 336820 619342
rect 336854 619308 336927 619342
rect 336233 619294 336927 619308
rect 336233 619260 336292 619294
rect 336326 619260 336382 619294
rect 336416 619260 336472 619294
rect 336506 619260 336562 619294
rect 336596 619260 336652 619294
rect 336686 619260 336742 619294
rect 336776 619260 336832 619294
rect 336866 619260 336927 619294
rect 336233 619242 336927 619260
rect 336233 619208 336320 619242
rect 336354 619208 336420 619242
rect 336454 619208 336520 619242
rect 336554 619208 336620 619242
rect 336654 619208 336720 619242
rect 336754 619208 336820 619242
rect 336854 619208 336927 619242
rect 336233 619204 336927 619208
rect 336233 619170 336292 619204
rect 336326 619170 336382 619204
rect 336416 619170 336472 619204
rect 336506 619170 336562 619204
rect 336596 619170 336652 619204
rect 336686 619170 336742 619204
rect 336776 619170 336832 619204
rect 336866 619170 336927 619204
rect 336233 619142 336927 619170
rect 336233 619114 336320 619142
rect 336354 619114 336420 619142
rect 336233 619080 336292 619114
rect 336354 619108 336382 619114
rect 336326 619080 336382 619108
rect 336416 619108 336420 619114
rect 336454 619114 336520 619142
rect 336454 619108 336472 619114
rect 336416 619080 336472 619108
rect 336506 619108 336520 619114
rect 336554 619114 336620 619142
rect 336654 619114 336720 619142
rect 336754 619114 336820 619142
rect 336854 619114 336927 619142
rect 336554 619108 336562 619114
rect 336506 619080 336562 619108
rect 336596 619108 336620 619114
rect 336686 619108 336720 619114
rect 336776 619108 336820 619114
rect 336596 619080 336652 619108
rect 336686 619080 336742 619108
rect 336776 619080 336832 619108
rect 336866 619080 336927 619114
rect 336233 619021 336927 619080
rect 336988 619683 337008 619717
rect 337042 619716 337406 619717
rect 337042 619683 337156 619716
rect 336988 619682 337156 619683
rect 337190 619682 337257 619716
rect 337291 619702 337406 619716
rect 337440 619702 337459 619736
rect 338277 619772 338444 619777
rect 338478 619772 338545 619806
rect 338579 619796 338786 619806
rect 338820 619796 338876 619830
rect 338910 619796 338966 619830
rect 339000 619796 339056 619830
rect 339090 619796 339146 619830
rect 339180 619796 339236 619830
rect 339270 619796 339326 619830
rect 339360 619796 339416 619830
rect 339450 619796 339506 619830
rect 339540 619806 340074 619830
rect 339540 619796 339732 619806
rect 338579 619777 339732 619796
rect 338579 619772 338747 619777
rect 338277 619736 338747 619772
rect 338277 619717 338694 619736
rect 337291 619682 337459 619702
rect 336988 619646 337459 619682
rect 336988 619627 337406 619646
rect 336988 619593 337008 619627
rect 337042 619626 337406 619627
rect 337042 619593 337156 619626
rect 336988 619592 337156 619593
rect 337190 619592 337257 619626
rect 337291 619612 337406 619626
rect 337440 619612 337459 619646
rect 337291 619592 337459 619612
rect 336988 619556 337459 619592
rect 336988 619537 337406 619556
rect 336988 619503 337008 619537
rect 337042 619536 337406 619537
rect 337042 619503 337156 619536
rect 336988 619502 337156 619503
rect 337190 619502 337257 619536
rect 337291 619522 337406 619536
rect 337440 619522 337459 619556
rect 337291 619502 337459 619522
rect 336988 619466 337459 619502
rect 336988 619447 337406 619466
rect 336988 619413 337008 619447
rect 337042 619446 337406 619447
rect 337042 619413 337156 619446
rect 336988 619412 337156 619413
rect 337190 619412 337257 619446
rect 337291 619432 337406 619446
rect 337440 619432 337459 619466
rect 337291 619412 337459 619432
rect 336988 619376 337459 619412
rect 336988 619357 337406 619376
rect 336988 619323 337008 619357
rect 337042 619356 337406 619357
rect 337042 619323 337156 619356
rect 336988 619322 337156 619323
rect 337190 619322 337257 619356
rect 337291 619342 337406 619356
rect 337440 619342 337459 619376
rect 337291 619322 337459 619342
rect 336988 619286 337459 619322
rect 336988 619267 337406 619286
rect 336988 619233 337008 619267
rect 337042 619266 337406 619267
rect 337042 619233 337156 619266
rect 336988 619232 337156 619233
rect 337190 619232 337257 619266
rect 337291 619252 337406 619266
rect 337440 619252 337459 619286
rect 337291 619232 337459 619252
rect 336988 619196 337459 619232
rect 336988 619177 337406 619196
rect 336988 619143 337008 619177
rect 337042 619176 337406 619177
rect 337042 619143 337156 619176
rect 336988 619142 337156 619143
rect 337190 619142 337257 619176
rect 337291 619162 337406 619176
rect 337440 619162 337459 619196
rect 337291 619142 337459 619162
rect 336988 619106 337459 619142
rect 336988 619087 337406 619106
rect 336988 619053 337008 619087
rect 337042 619086 337406 619087
rect 337042 619053 337156 619086
rect 336988 619052 337156 619053
rect 337190 619052 337257 619086
rect 337291 619072 337406 619086
rect 337440 619072 337459 619106
rect 337291 619052 337459 619072
rect 335688 618997 336118 619016
rect 335688 618963 335720 618997
rect 335754 618996 336118 618997
rect 335754 618963 335868 618996
rect 335688 618962 335868 618963
rect 335902 618962 335969 618996
rect 336003 618982 336118 618996
rect 336152 618982 336188 619016
rect 336003 618962 336188 618982
rect 335688 618959 336188 618962
rect 336988 619016 337459 619052
rect 337521 619654 338215 619715
rect 337521 619620 337580 619654
rect 337614 619642 337670 619654
rect 337642 619620 337670 619642
rect 337704 619642 337760 619654
rect 337704 619620 337708 619642
rect 337521 619608 337608 619620
rect 337642 619608 337708 619620
rect 337742 619620 337760 619642
rect 337794 619642 337850 619654
rect 337794 619620 337808 619642
rect 337742 619608 337808 619620
rect 337842 619620 337850 619642
rect 337884 619642 337940 619654
rect 337974 619642 338030 619654
rect 338064 619642 338120 619654
rect 337884 619620 337908 619642
rect 337974 619620 338008 619642
rect 338064 619620 338108 619642
rect 338154 619620 338215 619654
rect 337842 619608 337908 619620
rect 337942 619608 338008 619620
rect 338042 619608 338108 619620
rect 338142 619608 338215 619620
rect 337521 619564 338215 619608
rect 337521 619530 337580 619564
rect 337614 619542 337670 619564
rect 337642 619530 337670 619542
rect 337704 619542 337760 619564
rect 337704 619530 337708 619542
rect 337521 619508 337608 619530
rect 337642 619508 337708 619530
rect 337742 619530 337760 619542
rect 337794 619542 337850 619564
rect 337794 619530 337808 619542
rect 337742 619508 337808 619530
rect 337842 619530 337850 619542
rect 337884 619542 337940 619564
rect 337974 619542 338030 619564
rect 338064 619542 338120 619564
rect 337884 619530 337908 619542
rect 337974 619530 338008 619542
rect 338064 619530 338108 619542
rect 338154 619530 338215 619564
rect 337842 619508 337908 619530
rect 337942 619508 338008 619530
rect 338042 619508 338108 619530
rect 338142 619508 338215 619530
rect 337521 619474 338215 619508
rect 337521 619440 337580 619474
rect 337614 619442 337670 619474
rect 337642 619440 337670 619442
rect 337704 619442 337760 619474
rect 337704 619440 337708 619442
rect 337521 619408 337608 619440
rect 337642 619408 337708 619440
rect 337742 619440 337760 619442
rect 337794 619442 337850 619474
rect 337794 619440 337808 619442
rect 337742 619408 337808 619440
rect 337842 619440 337850 619442
rect 337884 619442 337940 619474
rect 337974 619442 338030 619474
rect 338064 619442 338120 619474
rect 337884 619440 337908 619442
rect 337974 619440 338008 619442
rect 338064 619440 338108 619442
rect 338154 619440 338215 619474
rect 337842 619408 337908 619440
rect 337942 619408 338008 619440
rect 338042 619408 338108 619440
rect 338142 619408 338215 619440
rect 337521 619384 338215 619408
rect 337521 619350 337580 619384
rect 337614 619350 337670 619384
rect 337704 619350 337760 619384
rect 337794 619350 337850 619384
rect 337884 619350 337940 619384
rect 337974 619350 338030 619384
rect 338064 619350 338120 619384
rect 338154 619350 338215 619384
rect 337521 619342 338215 619350
rect 337521 619308 337608 619342
rect 337642 619308 337708 619342
rect 337742 619308 337808 619342
rect 337842 619308 337908 619342
rect 337942 619308 338008 619342
rect 338042 619308 338108 619342
rect 338142 619308 338215 619342
rect 337521 619294 338215 619308
rect 337521 619260 337580 619294
rect 337614 619260 337670 619294
rect 337704 619260 337760 619294
rect 337794 619260 337850 619294
rect 337884 619260 337940 619294
rect 337974 619260 338030 619294
rect 338064 619260 338120 619294
rect 338154 619260 338215 619294
rect 337521 619242 338215 619260
rect 337521 619208 337608 619242
rect 337642 619208 337708 619242
rect 337742 619208 337808 619242
rect 337842 619208 337908 619242
rect 337942 619208 338008 619242
rect 338042 619208 338108 619242
rect 338142 619208 338215 619242
rect 337521 619204 338215 619208
rect 337521 619170 337580 619204
rect 337614 619170 337670 619204
rect 337704 619170 337760 619204
rect 337794 619170 337850 619204
rect 337884 619170 337940 619204
rect 337974 619170 338030 619204
rect 338064 619170 338120 619204
rect 338154 619170 338215 619204
rect 337521 619142 338215 619170
rect 337521 619114 337608 619142
rect 337642 619114 337708 619142
rect 337521 619080 337580 619114
rect 337642 619108 337670 619114
rect 337614 619080 337670 619108
rect 337704 619108 337708 619114
rect 337742 619114 337808 619142
rect 337742 619108 337760 619114
rect 337704 619080 337760 619108
rect 337794 619108 337808 619114
rect 337842 619114 337908 619142
rect 337942 619114 338008 619142
rect 338042 619114 338108 619142
rect 338142 619114 338215 619142
rect 337842 619108 337850 619114
rect 337794 619080 337850 619108
rect 337884 619108 337908 619114
rect 337974 619108 338008 619114
rect 338064 619108 338108 619114
rect 337884 619080 337940 619108
rect 337974 619080 338030 619108
rect 338064 619080 338120 619108
rect 338154 619080 338215 619114
rect 337521 619021 338215 619080
rect 338277 619683 338296 619717
rect 338330 619716 338694 619717
rect 338330 619683 338444 619716
rect 338277 619682 338444 619683
rect 338478 619682 338545 619716
rect 338579 619702 338694 619716
rect 338728 619702 338747 619736
rect 339565 619772 339732 619777
rect 339766 619772 339833 619806
rect 339867 619796 340074 619806
rect 340108 619796 340164 619830
rect 340198 619796 340254 619830
rect 340288 619796 340344 619830
rect 340378 619796 340434 619830
rect 340468 619796 340524 619830
rect 340558 619796 340614 619830
rect 340648 619796 340704 619830
rect 340738 619796 340794 619830
rect 340828 619806 341088 619830
rect 340828 619796 341020 619806
rect 339867 619777 341020 619796
rect 339867 619772 340035 619777
rect 339565 619736 340035 619772
rect 339565 619717 339982 619736
rect 338579 619682 338747 619702
rect 338277 619646 338747 619682
rect 338277 619627 338694 619646
rect 338277 619593 338296 619627
rect 338330 619626 338694 619627
rect 338330 619593 338444 619626
rect 338277 619592 338444 619593
rect 338478 619592 338545 619626
rect 338579 619612 338694 619626
rect 338728 619612 338747 619646
rect 338579 619592 338747 619612
rect 338277 619556 338747 619592
rect 338277 619537 338694 619556
rect 338277 619503 338296 619537
rect 338330 619536 338694 619537
rect 338330 619503 338444 619536
rect 338277 619502 338444 619503
rect 338478 619502 338545 619536
rect 338579 619522 338694 619536
rect 338728 619522 338747 619556
rect 338579 619502 338747 619522
rect 338277 619466 338747 619502
rect 338277 619447 338694 619466
rect 338277 619413 338296 619447
rect 338330 619446 338694 619447
rect 338330 619413 338444 619446
rect 338277 619412 338444 619413
rect 338478 619412 338545 619446
rect 338579 619432 338694 619446
rect 338728 619432 338747 619466
rect 338579 619412 338747 619432
rect 338277 619376 338747 619412
rect 338277 619357 338694 619376
rect 338277 619323 338296 619357
rect 338330 619356 338694 619357
rect 338330 619323 338444 619356
rect 338277 619322 338444 619323
rect 338478 619322 338545 619356
rect 338579 619342 338694 619356
rect 338728 619342 338747 619376
rect 338579 619322 338747 619342
rect 338277 619286 338747 619322
rect 338277 619267 338694 619286
rect 338277 619233 338296 619267
rect 338330 619266 338694 619267
rect 338330 619233 338444 619266
rect 338277 619232 338444 619233
rect 338478 619232 338545 619266
rect 338579 619252 338694 619266
rect 338728 619252 338747 619286
rect 338579 619232 338747 619252
rect 338277 619196 338747 619232
rect 338277 619177 338694 619196
rect 338277 619143 338296 619177
rect 338330 619176 338694 619177
rect 338330 619143 338444 619176
rect 338277 619142 338444 619143
rect 338478 619142 338545 619176
rect 338579 619162 338694 619176
rect 338728 619162 338747 619196
rect 338579 619142 338747 619162
rect 338277 619106 338747 619142
rect 338277 619087 338694 619106
rect 338277 619053 338296 619087
rect 338330 619086 338694 619087
rect 338330 619053 338444 619086
rect 338277 619052 338444 619053
rect 338478 619052 338545 619086
rect 338579 619072 338694 619086
rect 338728 619072 338747 619106
rect 338579 619052 338747 619072
rect 336988 618997 337406 619016
rect 336988 618963 337008 618997
rect 337042 618996 337406 618997
rect 337042 618963 337156 618996
rect 336988 618962 337156 618963
rect 337190 618962 337257 618996
rect 337291 618982 337406 618996
rect 337440 618982 337459 619016
rect 337291 618962 337459 618982
rect 336988 618959 337459 618962
rect 338277 619016 338747 619052
rect 338809 619654 339503 619715
rect 338809 619620 338868 619654
rect 338902 619642 338958 619654
rect 338930 619620 338958 619642
rect 338992 619642 339048 619654
rect 338992 619620 338996 619642
rect 338809 619608 338896 619620
rect 338930 619608 338996 619620
rect 339030 619620 339048 619642
rect 339082 619642 339138 619654
rect 339082 619620 339096 619642
rect 339030 619608 339096 619620
rect 339130 619620 339138 619642
rect 339172 619642 339228 619654
rect 339262 619642 339318 619654
rect 339352 619642 339408 619654
rect 339172 619620 339196 619642
rect 339262 619620 339296 619642
rect 339352 619620 339396 619642
rect 339442 619620 339503 619654
rect 339130 619608 339196 619620
rect 339230 619608 339296 619620
rect 339330 619608 339396 619620
rect 339430 619608 339503 619620
rect 338809 619564 339503 619608
rect 338809 619530 338868 619564
rect 338902 619542 338958 619564
rect 338930 619530 338958 619542
rect 338992 619542 339048 619564
rect 338992 619530 338996 619542
rect 338809 619508 338896 619530
rect 338930 619508 338996 619530
rect 339030 619530 339048 619542
rect 339082 619542 339138 619564
rect 339082 619530 339096 619542
rect 339030 619508 339096 619530
rect 339130 619530 339138 619542
rect 339172 619542 339228 619564
rect 339262 619542 339318 619564
rect 339352 619542 339408 619564
rect 339172 619530 339196 619542
rect 339262 619530 339296 619542
rect 339352 619530 339396 619542
rect 339442 619530 339503 619564
rect 339130 619508 339196 619530
rect 339230 619508 339296 619530
rect 339330 619508 339396 619530
rect 339430 619508 339503 619530
rect 338809 619474 339503 619508
rect 338809 619440 338868 619474
rect 338902 619442 338958 619474
rect 338930 619440 338958 619442
rect 338992 619442 339048 619474
rect 338992 619440 338996 619442
rect 338809 619408 338896 619440
rect 338930 619408 338996 619440
rect 339030 619440 339048 619442
rect 339082 619442 339138 619474
rect 339082 619440 339096 619442
rect 339030 619408 339096 619440
rect 339130 619440 339138 619442
rect 339172 619442 339228 619474
rect 339262 619442 339318 619474
rect 339352 619442 339408 619474
rect 339172 619440 339196 619442
rect 339262 619440 339296 619442
rect 339352 619440 339396 619442
rect 339442 619440 339503 619474
rect 339130 619408 339196 619440
rect 339230 619408 339296 619440
rect 339330 619408 339396 619440
rect 339430 619408 339503 619440
rect 338809 619384 339503 619408
rect 338809 619350 338868 619384
rect 338902 619350 338958 619384
rect 338992 619350 339048 619384
rect 339082 619350 339138 619384
rect 339172 619350 339228 619384
rect 339262 619350 339318 619384
rect 339352 619350 339408 619384
rect 339442 619350 339503 619384
rect 338809 619342 339503 619350
rect 338809 619308 338896 619342
rect 338930 619308 338996 619342
rect 339030 619308 339096 619342
rect 339130 619308 339196 619342
rect 339230 619308 339296 619342
rect 339330 619308 339396 619342
rect 339430 619308 339503 619342
rect 338809 619294 339503 619308
rect 338809 619260 338868 619294
rect 338902 619260 338958 619294
rect 338992 619260 339048 619294
rect 339082 619260 339138 619294
rect 339172 619260 339228 619294
rect 339262 619260 339318 619294
rect 339352 619260 339408 619294
rect 339442 619260 339503 619294
rect 338809 619242 339503 619260
rect 338809 619208 338896 619242
rect 338930 619208 338996 619242
rect 339030 619208 339096 619242
rect 339130 619208 339196 619242
rect 339230 619208 339296 619242
rect 339330 619208 339396 619242
rect 339430 619208 339503 619242
rect 338809 619204 339503 619208
rect 338809 619170 338868 619204
rect 338902 619170 338958 619204
rect 338992 619170 339048 619204
rect 339082 619170 339138 619204
rect 339172 619170 339228 619204
rect 339262 619170 339318 619204
rect 339352 619170 339408 619204
rect 339442 619170 339503 619204
rect 338809 619142 339503 619170
rect 338809 619114 338896 619142
rect 338930 619114 338996 619142
rect 338809 619080 338868 619114
rect 338930 619108 338958 619114
rect 338902 619080 338958 619108
rect 338992 619108 338996 619114
rect 339030 619114 339096 619142
rect 339030 619108 339048 619114
rect 338992 619080 339048 619108
rect 339082 619108 339096 619114
rect 339130 619114 339196 619142
rect 339230 619114 339296 619142
rect 339330 619114 339396 619142
rect 339430 619114 339503 619142
rect 339130 619108 339138 619114
rect 339082 619080 339138 619108
rect 339172 619108 339196 619114
rect 339262 619108 339296 619114
rect 339352 619108 339396 619114
rect 339172 619080 339228 619108
rect 339262 619080 339318 619108
rect 339352 619080 339408 619108
rect 339442 619080 339503 619114
rect 338809 619021 339503 619080
rect 339565 619683 339584 619717
rect 339618 619716 339982 619717
rect 339618 619683 339732 619716
rect 339565 619682 339732 619683
rect 339766 619682 339833 619716
rect 339867 619702 339982 619716
rect 340016 619702 340035 619736
rect 340853 619772 341020 619777
rect 341054 619772 341088 619806
rect 340853 619717 341088 619772
rect 339867 619682 340035 619702
rect 339565 619646 340035 619682
rect 339565 619627 339982 619646
rect 339565 619593 339584 619627
rect 339618 619626 339982 619627
rect 339618 619593 339732 619626
rect 339565 619592 339732 619593
rect 339766 619592 339833 619626
rect 339867 619612 339982 619626
rect 340016 619612 340035 619646
rect 339867 619592 340035 619612
rect 339565 619556 340035 619592
rect 339565 619537 339982 619556
rect 339565 619503 339584 619537
rect 339618 619536 339982 619537
rect 339618 619503 339732 619536
rect 339565 619502 339732 619503
rect 339766 619502 339833 619536
rect 339867 619522 339982 619536
rect 340016 619522 340035 619556
rect 339867 619502 340035 619522
rect 339565 619466 340035 619502
rect 339565 619447 339982 619466
rect 339565 619413 339584 619447
rect 339618 619446 339982 619447
rect 339618 619413 339732 619446
rect 339565 619412 339732 619413
rect 339766 619412 339833 619446
rect 339867 619432 339982 619446
rect 340016 619432 340035 619466
rect 339867 619412 340035 619432
rect 339565 619376 340035 619412
rect 339565 619357 339982 619376
rect 339565 619323 339584 619357
rect 339618 619356 339982 619357
rect 339618 619323 339732 619356
rect 339565 619322 339732 619323
rect 339766 619322 339833 619356
rect 339867 619342 339982 619356
rect 340016 619342 340035 619376
rect 339867 619322 340035 619342
rect 339565 619286 340035 619322
rect 339565 619267 339982 619286
rect 339565 619233 339584 619267
rect 339618 619266 339982 619267
rect 339618 619233 339732 619266
rect 339565 619232 339732 619233
rect 339766 619232 339833 619266
rect 339867 619252 339982 619266
rect 340016 619252 340035 619286
rect 339867 619232 340035 619252
rect 339565 619196 340035 619232
rect 339565 619177 339982 619196
rect 339565 619143 339584 619177
rect 339618 619176 339982 619177
rect 339618 619143 339732 619176
rect 339565 619142 339732 619143
rect 339766 619142 339833 619176
rect 339867 619162 339982 619176
rect 340016 619162 340035 619196
rect 339867 619142 340035 619162
rect 339565 619106 340035 619142
rect 339565 619087 339982 619106
rect 339565 619053 339584 619087
rect 339618 619086 339982 619087
rect 339618 619053 339732 619086
rect 339565 619052 339732 619053
rect 339766 619052 339833 619086
rect 339867 619072 339982 619086
rect 340016 619072 340035 619106
rect 339867 619052 340035 619072
rect 338277 618997 338694 619016
rect 338277 618963 338296 618997
rect 338330 618996 338694 618997
rect 338330 618963 338444 618996
rect 338277 618962 338444 618963
rect 338478 618962 338545 618996
rect 338579 618982 338694 618996
rect 338728 618982 338747 619016
rect 338579 618962 338747 618982
rect 338277 618959 338747 618962
rect 339565 619016 340035 619052
rect 340097 619654 340791 619715
rect 340097 619620 340156 619654
rect 340190 619642 340246 619654
rect 340218 619620 340246 619642
rect 340280 619642 340336 619654
rect 340280 619620 340284 619642
rect 340097 619608 340184 619620
rect 340218 619608 340284 619620
rect 340318 619620 340336 619642
rect 340370 619642 340426 619654
rect 340370 619620 340384 619642
rect 340318 619608 340384 619620
rect 340418 619620 340426 619642
rect 340460 619642 340516 619654
rect 340550 619642 340606 619654
rect 340640 619642 340696 619654
rect 340460 619620 340484 619642
rect 340550 619620 340584 619642
rect 340640 619620 340684 619642
rect 340730 619620 340791 619654
rect 340418 619608 340484 619620
rect 340518 619608 340584 619620
rect 340618 619608 340684 619620
rect 340718 619608 340791 619620
rect 340097 619564 340791 619608
rect 340097 619530 340156 619564
rect 340190 619542 340246 619564
rect 340218 619530 340246 619542
rect 340280 619542 340336 619564
rect 340280 619530 340284 619542
rect 340097 619508 340184 619530
rect 340218 619508 340284 619530
rect 340318 619530 340336 619542
rect 340370 619542 340426 619564
rect 340370 619530 340384 619542
rect 340318 619508 340384 619530
rect 340418 619530 340426 619542
rect 340460 619542 340516 619564
rect 340550 619542 340606 619564
rect 340640 619542 340696 619564
rect 340460 619530 340484 619542
rect 340550 619530 340584 619542
rect 340640 619530 340684 619542
rect 340730 619530 340791 619564
rect 340418 619508 340484 619530
rect 340518 619508 340584 619530
rect 340618 619508 340684 619530
rect 340718 619508 340791 619530
rect 340097 619474 340791 619508
rect 340097 619440 340156 619474
rect 340190 619442 340246 619474
rect 340218 619440 340246 619442
rect 340280 619442 340336 619474
rect 340280 619440 340284 619442
rect 340097 619408 340184 619440
rect 340218 619408 340284 619440
rect 340318 619440 340336 619442
rect 340370 619442 340426 619474
rect 340370 619440 340384 619442
rect 340318 619408 340384 619440
rect 340418 619440 340426 619442
rect 340460 619442 340516 619474
rect 340550 619442 340606 619474
rect 340640 619442 340696 619474
rect 340460 619440 340484 619442
rect 340550 619440 340584 619442
rect 340640 619440 340684 619442
rect 340730 619440 340791 619474
rect 340418 619408 340484 619440
rect 340518 619408 340584 619440
rect 340618 619408 340684 619440
rect 340718 619408 340791 619440
rect 340097 619384 340791 619408
rect 340097 619350 340156 619384
rect 340190 619350 340246 619384
rect 340280 619350 340336 619384
rect 340370 619350 340426 619384
rect 340460 619350 340516 619384
rect 340550 619350 340606 619384
rect 340640 619350 340696 619384
rect 340730 619350 340791 619384
rect 340097 619342 340791 619350
rect 340097 619308 340184 619342
rect 340218 619308 340284 619342
rect 340318 619308 340384 619342
rect 340418 619308 340484 619342
rect 340518 619308 340584 619342
rect 340618 619308 340684 619342
rect 340718 619308 340791 619342
rect 340097 619294 340791 619308
rect 340097 619260 340156 619294
rect 340190 619260 340246 619294
rect 340280 619260 340336 619294
rect 340370 619260 340426 619294
rect 340460 619260 340516 619294
rect 340550 619260 340606 619294
rect 340640 619260 340696 619294
rect 340730 619260 340791 619294
rect 340097 619242 340791 619260
rect 340097 619208 340184 619242
rect 340218 619208 340284 619242
rect 340318 619208 340384 619242
rect 340418 619208 340484 619242
rect 340518 619208 340584 619242
rect 340618 619208 340684 619242
rect 340718 619208 340791 619242
rect 340097 619204 340791 619208
rect 340097 619170 340156 619204
rect 340190 619170 340246 619204
rect 340280 619170 340336 619204
rect 340370 619170 340426 619204
rect 340460 619170 340516 619204
rect 340550 619170 340606 619204
rect 340640 619170 340696 619204
rect 340730 619170 340791 619204
rect 340097 619142 340791 619170
rect 340097 619114 340184 619142
rect 340218 619114 340284 619142
rect 340097 619080 340156 619114
rect 340218 619108 340246 619114
rect 340190 619080 340246 619108
rect 340280 619108 340284 619114
rect 340318 619114 340384 619142
rect 340318 619108 340336 619114
rect 340280 619080 340336 619108
rect 340370 619108 340384 619114
rect 340418 619114 340484 619142
rect 340518 619114 340584 619142
rect 340618 619114 340684 619142
rect 340718 619114 340791 619142
rect 340418 619108 340426 619114
rect 340370 619080 340426 619108
rect 340460 619108 340484 619114
rect 340550 619108 340584 619114
rect 340640 619108 340684 619114
rect 340460 619080 340516 619108
rect 340550 619080 340606 619108
rect 340640 619080 340696 619108
rect 340730 619080 340791 619114
rect 340097 619021 340791 619080
rect 340853 619683 340872 619717
rect 340906 619716 341088 619717
rect 340906 619683 341020 619716
rect 340853 619682 341020 619683
rect 341054 619682 341088 619716
rect 340853 619627 341088 619682
rect 340853 619593 340872 619627
rect 340906 619626 341088 619627
rect 340906 619593 341020 619626
rect 340853 619592 341020 619593
rect 341054 619592 341088 619626
rect 340853 619537 341088 619592
rect 340853 619503 340872 619537
rect 340906 619536 341088 619537
rect 340906 619503 341020 619536
rect 340853 619502 341020 619503
rect 341054 619502 341088 619536
rect 340853 619447 341088 619502
rect 340853 619413 340872 619447
rect 340906 619446 341088 619447
rect 340906 619413 341020 619446
rect 340853 619412 341020 619413
rect 341054 619412 341088 619446
rect 340853 619357 341088 619412
rect 340853 619323 340872 619357
rect 340906 619356 341088 619357
rect 340906 619323 341020 619356
rect 340853 619322 341020 619323
rect 341054 619322 341088 619356
rect 340853 619267 341088 619322
rect 340853 619233 340872 619267
rect 340906 619266 341088 619267
rect 340906 619233 341020 619266
rect 340853 619232 341020 619233
rect 341054 619232 341088 619266
rect 340853 619177 341088 619232
rect 340853 619143 340872 619177
rect 340906 619176 341088 619177
rect 340906 619143 341020 619176
rect 340853 619142 341020 619143
rect 341054 619142 341088 619176
rect 340853 619087 341088 619142
rect 340853 619053 340872 619087
rect 340906 619086 341088 619087
rect 340906 619053 341020 619086
rect 340853 619052 341020 619053
rect 341054 619052 341088 619086
rect 339565 618997 339982 619016
rect 339565 618963 339584 618997
rect 339618 618996 339982 618997
rect 339618 618963 339732 618996
rect 339565 618962 339732 618963
rect 339766 618962 339833 618996
rect 339867 618982 339982 618996
rect 340016 618982 340035 619016
rect 339867 618962 340035 618982
rect 339565 618959 340035 618962
rect 340853 618997 341088 619052
rect 340853 618963 340872 618997
rect 340906 618996 341088 618997
rect 340906 618963 341020 618996
rect 340853 618962 341020 618963
rect 341054 618962 341088 618996
rect 340853 618959 341088 618962
rect 334648 618940 341088 618959
rect 334648 618906 334888 618940
rect 334922 618906 334978 618940
rect 335012 618906 335068 618940
rect 335102 618906 335158 618940
rect 335192 618906 335248 618940
rect 335282 618906 335338 618940
rect 335372 618906 335428 618940
rect 335462 618906 335518 618940
rect 335552 618906 335608 618940
rect 335642 618906 336176 618940
rect 336210 618906 336266 618940
rect 336300 618906 336356 618940
rect 336390 618906 336446 618940
rect 336480 618906 336536 618940
rect 336570 618906 336626 618940
rect 336660 618906 336716 618940
rect 336750 618906 336806 618940
rect 336840 618906 336896 618940
rect 336930 618906 337464 618940
rect 337498 618906 337554 618940
rect 337588 618906 337644 618940
rect 337678 618906 337734 618940
rect 337768 618906 337824 618940
rect 337858 618906 337914 618940
rect 337948 618906 338004 618940
rect 338038 618906 338094 618940
rect 338128 618906 338184 618940
rect 338218 618906 338752 618940
rect 338786 618906 338842 618940
rect 338876 618906 338932 618940
rect 338966 618906 339022 618940
rect 339056 618906 339112 618940
rect 339146 618906 339202 618940
rect 339236 618906 339292 618940
rect 339326 618906 339382 618940
rect 339416 618906 339472 618940
rect 339506 618906 340040 618940
rect 340074 618906 340130 618940
rect 340164 618906 340220 618940
rect 340254 618906 340310 618940
rect 340344 618906 340400 618940
rect 340434 618906 340490 618940
rect 340524 618906 340580 618940
rect 340614 618906 340670 618940
rect 340704 618906 340760 618940
rect 340794 618906 341088 618940
rect 334648 618872 334681 618906
rect 334715 618887 335868 618906
rect 334715 618872 334888 618887
rect 334648 618823 334888 618872
rect 335688 618872 335868 618887
rect 335902 618872 335969 618906
rect 336003 618887 337156 618906
rect 336003 618872 336188 618887
rect 335688 618823 336188 618872
rect 336988 618872 337156 618887
rect 337190 618872 337257 618906
rect 337291 618887 338444 618906
rect 337291 618872 337388 618887
rect 336988 618823 337388 618872
rect 338288 618872 338444 618887
rect 338478 618872 338545 618906
rect 338579 618887 339732 618906
rect 338579 618872 338688 618887
rect 338288 618823 338688 618872
rect 339588 618872 339732 618887
rect 339766 618872 339833 618906
rect 339867 618887 341020 618906
rect 339867 618872 339988 618887
rect 339588 618823 339988 618872
rect 340888 618872 341020 618887
rect 341054 618872 341088 618906
rect 340888 618823 341088 618872
rect 334648 618816 341088 618823
rect 334648 618782 334681 618816
rect 334715 618793 335868 618816
rect 334715 618782 334782 618793
rect 334648 618759 334782 618782
rect 334816 618759 334872 618793
rect 334906 618759 334962 618793
rect 334996 618759 335052 618793
rect 335086 618759 335142 618793
rect 335176 618759 335232 618793
rect 335266 618759 335322 618793
rect 335356 618759 335412 618793
rect 335446 618759 335502 618793
rect 335536 618759 335592 618793
rect 335626 618759 335682 618793
rect 335716 618759 335772 618793
rect 335806 618782 335868 618793
rect 335902 618782 335969 618816
rect 336003 618793 337156 618816
rect 336003 618782 336070 618793
rect 335806 618759 336070 618782
rect 336104 618759 336160 618793
rect 336194 618759 336250 618793
rect 336284 618759 336340 618793
rect 336374 618759 336430 618793
rect 336464 618759 336520 618793
rect 336554 618759 336610 618793
rect 336644 618759 336700 618793
rect 336734 618759 336790 618793
rect 336824 618759 336880 618793
rect 336914 618759 336970 618793
rect 337004 618759 337060 618793
rect 337094 618782 337156 618793
rect 337190 618782 337257 618816
rect 337291 618793 338444 618816
rect 337291 618782 337358 618793
rect 337094 618759 337358 618782
rect 337392 618759 337448 618793
rect 337482 618759 337538 618793
rect 337572 618759 337628 618793
rect 337662 618759 337718 618793
rect 337752 618759 337808 618793
rect 337842 618759 337898 618793
rect 337932 618759 337988 618793
rect 338022 618759 338078 618793
rect 338112 618759 338168 618793
rect 338202 618759 338258 618793
rect 338292 618759 338348 618793
rect 338382 618782 338444 618793
rect 338478 618782 338545 618816
rect 338579 618793 339732 618816
rect 338579 618782 338646 618793
rect 338382 618759 338646 618782
rect 338680 618759 338736 618793
rect 338770 618759 338826 618793
rect 338860 618759 338916 618793
rect 338950 618759 339006 618793
rect 339040 618759 339096 618793
rect 339130 618759 339186 618793
rect 339220 618759 339276 618793
rect 339310 618759 339366 618793
rect 339400 618759 339456 618793
rect 339490 618759 339546 618793
rect 339580 618759 339636 618793
rect 339670 618782 339732 618793
rect 339766 618782 339833 618816
rect 339867 618793 341020 618816
rect 339867 618782 339934 618793
rect 339670 618759 339934 618782
rect 339968 618759 340024 618793
rect 340058 618759 340114 618793
rect 340148 618759 340204 618793
rect 340238 618759 340294 618793
rect 340328 618759 340384 618793
rect 340418 618759 340474 618793
rect 340508 618759 340564 618793
rect 340598 618759 340654 618793
rect 340688 618759 340744 618793
rect 340778 618759 340834 618793
rect 340868 618759 340924 618793
rect 340958 618782 341020 618793
rect 341054 618782 341088 618816
rect 340958 618759 341088 618782
rect 334648 618692 341088 618759
rect 334648 618658 334782 618692
rect 334816 618658 334872 618692
rect 334906 618658 334962 618692
rect 334996 618658 335052 618692
rect 335086 618658 335142 618692
rect 335176 618658 335232 618692
rect 335266 618658 335322 618692
rect 335356 618658 335412 618692
rect 335446 618658 335502 618692
rect 335536 618658 335592 618692
rect 335626 618658 335682 618692
rect 335716 618658 335772 618692
rect 335806 618658 336070 618692
rect 336104 618658 336160 618692
rect 336194 618658 336250 618692
rect 336284 618658 336340 618692
rect 336374 618658 336430 618692
rect 336464 618658 336520 618692
rect 336554 618658 336610 618692
rect 336644 618658 336700 618692
rect 336734 618658 336790 618692
rect 336824 618658 336880 618692
rect 336914 618658 336970 618692
rect 337004 618658 337060 618692
rect 337094 618658 337358 618692
rect 337392 618658 337448 618692
rect 337482 618658 337538 618692
rect 337572 618658 337628 618692
rect 337662 618658 337718 618692
rect 337752 618658 337808 618692
rect 337842 618658 337898 618692
rect 337932 618658 337988 618692
rect 338022 618658 338078 618692
rect 338112 618658 338168 618692
rect 338202 618658 338258 618692
rect 338292 618658 338348 618692
rect 338382 618658 338646 618692
rect 338680 618658 338736 618692
rect 338770 618658 338826 618692
rect 338860 618658 338916 618692
rect 338950 618658 339006 618692
rect 339040 618658 339096 618692
rect 339130 618658 339186 618692
rect 339220 618658 339276 618692
rect 339310 618658 339366 618692
rect 339400 618658 339456 618692
rect 339490 618658 339546 618692
rect 339580 618658 339636 618692
rect 339670 618658 339934 618692
rect 339968 618658 340024 618692
rect 340058 618658 340114 618692
rect 340148 618658 340204 618692
rect 340238 618658 340294 618692
rect 340328 618658 340384 618692
rect 340418 618658 340474 618692
rect 340508 618658 340564 618692
rect 340598 618658 340654 618692
rect 340688 618658 340744 618692
rect 340778 618658 340834 618692
rect 340868 618658 340924 618692
rect 340958 618658 341088 618692
rect 334648 618625 341088 618658
rect 334648 618608 334888 618625
rect 334648 618574 334681 618608
rect 334715 618574 334888 618608
rect 334648 618561 334888 618574
rect 335688 618608 336188 618625
rect 335688 618574 335868 618608
rect 335902 618574 335969 618608
rect 336003 618574 336188 618608
rect 335688 618561 336188 618574
rect 336988 618608 337388 618625
rect 336988 618574 337156 618608
rect 337190 618574 337257 618608
rect 337291 618574 337388 618608
rect 336988 618561 337388 618574
rect 338288 618608 338688 618625
rect 338288 618574 338444 618608
rect 338478 618574 338545 618608
rect 338579 618574 338688 618608
rect 338288 618561 338688 618574
rect 339588 618608 339988 618625
rect 339588 618574 339732 618608
rect 339766 618574 339833 618608
rect 339867 618574 339988 618608
rect 339588 618561 339988 618574
rect 340888 618608 341088 618625
rect 340888 618574 341020 618608
rect 341054 618574 341088 618608
rect 340888 618561 341088 618574
rect 334648 618542 341088 618561
rect 334648 618518 334922 618542
rect 334648 618484 334681 618518
rect 334715 618508 334922 618518
rect 334956 618508 335012 618542
rect 335046 618508 335102 618542
rect 335136 618508 335192 618542
rect 335226 618508 335282 618542
rect 335316 618508 335372 618542
rect 335406 618508 335462 618542
rect 335496 618508 335552 618542
rect 335586 618508 335642 618542
rect 335676 618518 336210 618542
rect 335676 618508 335868 618518
rect 334715 618489 335868 618508
rect 334715 618484 334888 618489
rect 334648 618448 334888 618484
rect 334648 618428 334830 618448
rect 334648 618394 334681 618428
rect 334715 618414 334830 618428
rect 334864 618414 334888 618448
rect 335688 618484 335868 618489
rect 335902 618484 335969 618518
rect 336003 618508 336210 618518
rect 336244 618508 336300 618542
rect 336334 618508 336390 618542
rect 336424 618508 336480 618542
rect 336514 618508 336570 618542
rect 336604 618508 336660 618542
rect 336694 618508 336750 618542
rect 336784 618508 336840 618542
rect 336874 618508 336930 618542
rect 336964 618518 337498 618542
rect 336964 618508 337156 618518
rect 336003 618489 337156 618508
rect 336003 618484 336188 618489
rect 335688 618448 336188 618484
rect 335688 618429 336118 618448
rect 334715 618394 334888 618414
rect 334648 618358 334888 618394
rect 334648 618338 334830 618358
rect 334648 618304 334681 618338
rect 334715 618324 334830 618338
rect 334864 618324 334888 618358
rect 334715 618304 334888 618324
rect 334648 618268 334888 618304
rect 334648 618248 334830 618268
rect 334648 618214 334681 618248
rect 334715 618234 334830 618248
rect 334864 618234 334888 618268
rect 334715 618214 334888 618234
rect 334648 618178 334888 618214
rect 334648 618158 334830 618178
rect 334648 618124 334681 618158
rect 334715 618144 334830 618158
rect 334864 618144 334888 618178
rect 334715 618124 334888 618144
rect 334648 618088 334888 618124
rect 334648 618068 334830 618088
rect 334648 618034 334681 618068
rect 334715 618054 334830 618068
rect 334864 618054 334888 618088
rect 334715 618034 334888 618054
rect 334648 617998 334888 618034
rect 334648 617978 334830 617998
rect 334648 617944 334681 617978
rect 334715 617964 334830 617978
rect 334864 617964 334888 617998
rect 334715 617944 334888 617964
rect 334648 617908 334888 617944
rect 334648 617888 334830 617908
rect 334648 617854 334681 617888
rect 334715 617874 334830 617888
rect 334864 617874 334888 617908
rect 334715 617854 334888 617874
rect 334648 617818 334888 617854
rect 334648 617798 334830 617818
rect 334648 617764 334681 617798
rect 334715 617784 334830 617798
rect 334864 617784 334888 617818
rect 334715 617764 334888 617784
rect 334648 617728 334888 617764
rect 334945 618366 335639 618427
rect 334945 618332 335004 618366
rect 335038 618354 335094 618366
rect 335066 618332 335094 618354
rect 335128 618354 335184 618366
rect 335128 618332 335132 618354
rect 334945 618320 335032 618332
rect 335066 618320 335132 618332
rect 335166 618332 335184 618354
rect 335218 618354 335274 618366
rect 335218 618332 335232 618354
rect 335166 618320 335232 618332
rect 335266 618332 335274 618354
rect 335308 618354 335364 618366
rect 335398 618354 335454 618366
rect 335488 618354 335544 618366
rect 335308 618332 335332 618354
rect 335398 618332 335432 618354
rect 335488 618332 335532 618354
rect 335578 618332 335639 618366
rect 335266 618320 335332 618332
rect 335366 618320 335432 618332
rect 335466 618320 335532 618332
rect 335566 618320 335639 618332
rect 334945 618276 335639 618320
rect 334945 618242 335004 618276
rect 335038 618254 335094 618276
rect 335066 618242 335094 618254
rect 335128 618254 335184 618276
rect 335128 618242 335132 618254
rect 334945 618220 335032 618242
rect 335066 618220 335132 618242
rect 335166 618242 335184 618254
rect 335218 618254 335274 618276
rect 335218 618242 335232 618254
rect 335166 618220 335232 618242
rect 335266 618242 335274 618254
rect 335308 618254 335364 618276
rect 335398 618254 335454 618276
rect 335488 618254 335544 618276
rect 335308 618242 335332 618254
rect 335398 618242 335432 618254
rect 335488 618242 335532 618254
rect 335578 618242 335639 618276
rect 335266 618220 335332 618242
rect 335366 618220 335432 618242
rect 335466 618220 335532 618242
rect 335566 618220 335639 618242
rect 334945 618186 335639 618220
rect 334945 618152 335004 618186
rect 335038 618154 335094 618186
rect 335066 618152 335094 618154
rect 335128 618154 335184 618186
rect 335128 618152 335132 618154
rect 334945 618120 335032 618152
rect 335066 618120 335132 618152
rect 335166 618152 335184 618154
rect 335218 618154 335274 618186
rect 335218 618152 335232 618154
rect 335166 618120 335232 618152
rect 335266 618152 335274 618154
rect 335308 618154 335364 618186
rect 335398 618154 335454 618186
rect 335488 618154 335544 618186
rect 335308 618152 335332 618154
rect 335398 618152 335432 618154
rect 335488 618152 335532 618154
rect 335578 618152 335639 618186
rect 335266 618120 335332 618152
rect 335366 618120 335432 618152
rect 335466 618120 335532 618152
rect 335566 618120 335639 618152
rect 334945 618096 335639 618120
rect 334945 618062 335004 618096
rect 335038 618062 335094 618096
rect 335128 618062 335184 618096
rect 335218 618062 335274 618096
rect 335308 618062 335364 618096
rect 335398 618062 335454 618096
rect 335488 618062 335544 618096
rect 335578 618062 335639 618096
rect 334945 618054 335639 618062
rect 334945 618020 335032 618054
rect 335066 618020 335132 618054
rect 335166 618020 335232 618054
rect 335266 618020 335332 618054
rect 335366 618020 335432 618054
rect 335466 618020 335532 618054
rect 335566 618020 335639 618054
rect 334945 618006 335639 618020
rect 334945 617972 335004 618006
rect 335038 617972 335094 618006
rect 335128 617972 335184 618006
rect 335218 617972 335274 618006
rect 335308 617972 335364 618006
rect 335398 617972 335454 618006
rect 335488 617972 335544 618006
rect 335578 617972 335639 618006
rect 334945 617954 335639 617972
rect 334945 617920 335032 617954
rect 335066 617920 335132 617954
rect 335166 617920 335232 617954
rect 335266 617920 335332 617954
rect 335366 617920 335432 617954
rect 335466 617920 335532 617954
rect 335566 617920 335639 617954
rect 334945 617916 335639 617920
rect 334945 617882 335004 617916
rect 335038 617882 335094 617916
rect 335128 617882 335184 617916
rect 335218 617882 335274 617916
rect 335308 617882 335364 617916
rect 335398 617882 335454 617916
rect 335488 617882 335544 617916
rect 335578 617882 335639 617916
rect 334945 617854 335639 617882
rect 334945 617826 335032 617854
rect 335066 617826 335132 617854
rect 334945 617792 335004 617826
rect 335066 617820 335094 617826
rect 335038 617792 335094 617820
rect 335128 617820 335132 617826
rect 335166 617826 335232 617854
rect 335166 617820 335184 617826
rect 335128 617792 335184 617820
rect 335218 617820 335232 617826
rect 335266 617826 335332 617854
rect 335366 617826 335432 617854
rect 335466 617826 335532 617854
rect 335566 617826 335639 617854
rect 335266 617820 335274 617826
rect 335218 617792 335274 617820
rect 335308 617820 335332 617826
rect 335398 617820 335432 617826
rect 335488 617820 335532 617826
rect 335308 617792 335364 617820
rect 335398 617792 335454 617820
rect 335488 617792 335544 617820
rect 335578 617792 335639 617826
rect 334945 617733 335639 617792
rect 335688 618395 335720 618429
rect 335754 618428 336118 618429
rect 335754 618395 335868 618428
rect 335688 618394 335868 618395
rect 335902 618394 335969 618428
rect 336003 618414 336118 618428
rect 336152 618414 336188 618448
rect 336988 618484 337156 618489
rect 337190 618484 337257 618518
rect 337291 618508 337498 618518
rect 337532 618508 337588 618542
rect 337622 618508 337678 618542
rect 337712 618508 337768 618542
rect 337802 618508 337858 618542
rect 337892 618508 337948 618542
rect 337982 618508 338038 618542
rect 338072 618508 338128 618542
rect 338162 618508 338218 618542
rect 338252 618518 338786 618542
rect 338252 618508 338444 618518
rect 337291 618489 338444 618508
rect 337291 618484 337459 618489
rect 336988 618448 337459 618484
rect 336988 618429 337406 618448
rect 336003 618394 336188 618414
rect 335688 618358 336188 618394
rect 335688 618339 336118 618358
rect 335688 618305 335720 618339
rect 335754 618338 336118 618339
rect 335754 618305 335868 618338
rect 335688 618304 335868 618305
rect 335902 618304 335969 618338
rect 336003 618324 336118 618338
rect 336152 618324 336188 618358
rect 336003 618304 336188 618324
rect 335688 618268 336188 618304
rect 335688 618249 336118 618268
rect 335688 618215 335720 618249
rect 335754 618248 336118 618249
rect 335754 618215 335868 618248
rect 335688 618214 335868 618215
rect 335902 618214 335969 618248
rect 336003 618234 336118 618248
rect 336152 618234 336188 618268
rect 336003 618214 336188 618234
rect 335688 618178 336188 618214
rect 335688 618159 336118 618178
rect 335688 618125 335720 618159
rect 335754 618158 336118 618159
rect 335754 618125 335868 618158
rect 335688 618124 335868 618125
rect 335902 618124 335969 618158
rect 336003 618144 336118 618158
rect 336152 618144 336188 618178
rect 336003 618124 336188 618144
rect 335688 618088 336188 618124
rect 335688 618069 336118 618088
rect 335688 618035 335720 618069
rect 335754 618068 336118 618069
rect 335754 618035 335868 618068
rect 335688 618034 335868 618035
rect 335902 618034 335969 618068
rect 336003 618054 336118 618068
rect 336152 618054 336188 618088
rect 336003 618034 336188 618054
rect 335688 617998 336188 618034
rect 335688 617979 336118 617998
rect 335688 617945 335720 617979
rect 335754 617978 336118 617979
rect 335754 617945 335868 617978
rect 335688 617944 335868 617945
rect 335902 617944 335969 617978
rect 336003 617964 336118 617978
rect 336152 617964 336188 617998
rect 336003 617944 336188 617964
rect 335688 617908 336188 617944
rect 335688 617889 336118 617908
rect 335688 617855 335720 617889
rect 335754 617888 336118 617889
rect 335754 617855 335868 617888
rect 335688 617854 335868 617855
rect 335902 617854 335969 617888
rect 336003 617874 336118 617888
rect 336152 617874 336188 617908
rect 336003 617854 336188 617874
rect 335688 617818 336188 617854
rect 335688 617799 336118 617818
rect 335688 617765 335720 617799
rect 335754 617798 336118 617799
rect 335754 617765 335868 617798
rect 335688 617764 335868 617765
rect 335902 617764 335969 617798
rect 336003 617784 336118 617798
rect 336152 617784 336188 617818
rect 336003 617764 336188 617784
rect 334648 617708 334830 617728
rect 334648 617674 334681 617708
rect 334715 617694 334830 617708
rect 334864 617694 334888 617728
rect 334715 617674 334888 617694
rect 334648 617671 334888 617674
rect 335688 617728 336188 617764
rect 336233 618366 336927 618427
rect 336233 618332 336292 618366
rect 336326 618354 336382 618366
rect 336354 618332 336382 618354
rect 336416 618354 336472 618366
rect 336416 618332 336420 618354
rect 336233 618320 336320 618332
rect 336354 618320 336420 618332
rect 336454 618332 336472 618354
rect 336506 618354 336562 618366
rect 336506 618332 336520 618354
rect 336454 618320 336520 618332
rect 336554 618332 336562 618354
rect 336596 618354 336652 618366
rect 336686 618354 336742 618366
rect 336776 618354 336832 618366
rect 336596 618332 336620 618354
rect 336686 618332 336720 618354
rect 336776 618332 336820 618354
rect 336866 618332 336927 618366
rect 336554 618320 336620 618332
rect 336654 618320 336720 618332
rect 336754 618320 336820 618332
rect 336854 618320 336927 618332
rect 336233 618276 336927 618320
rect 336233 618242 336292 618276
rect 336326 618254 336382 618276
rect 336354 618242 336382 618254
rect 336416 618254 336472 618276
rect 336416 618242 336420 618254
rect 336233 618220 336320 618242
rect 336354 618220 336420 618242
rect 336454 618242 336472 618254
rect 336506 618254 336562 618276
rect 336506 618242 336520 618254
rect 336454 618220 336520 618242
rect 336554 618242 336562 618254
rect 336596 618254 336652 618276
rect 336686 618254 336742 618276
rect 336776 618254 336832 618276
rect 336596 618242 336620 618254
rect 336686 618242 336720 618254
rect 336776 618242 336820 618254
rect 336866 618242 336927 618276
rect 336554 618220 336620 618242
rect 336654 618220 336720 618242
rect 336754 618220 336820 618242
rect 336854 618220 336927 618242
rect 336233 618186 336927 618220
rect 336233 618152 336292 618186
rect 336326 618154 336382 618186
rect 336354 618152 336382 618154
rect 336416 618154 336472 618186
rect 336416 618152 336420 618154
rect 336233 618120 336320 618152
rect 336354 618120 336420 618152
rect 336454 618152 336472 618154
rect 336506 618154 336562 618186
rect 336506 618152 336520 618154
rect 336454 618120 336520 618152
rect 336554 618152 336562 618154
rect 336596 618154 336652 618186
rect 336686 618154 336742 618186
rect 336776 618154 336832 618186
rect 336596 618152 336620 618154
rect 336686 618152 336720 618154
rect 336776 618152 336820 618154
rect 336866 618152 336927 618186
rect 336554 618120 336620 618152
rect 336654 618120 336720 618152
rect 336754 618120 336820 618152
rect 336854 618120 336927 618152
rect 336233 618096 336927 618120
rect 336233 618062 336292 618096
rect 336326 618062 336382 618096
rect 336416 618062 336472 618096
rect 336506 618062 336562 618096
rect 336596 618062 336652 618096
rect 336686 618062 336742 618096
rect 336776 618062 336832 618096
rect 336866 618062 336927 618096
rect 336233 618054 336927 618062
rect 336233 618020 336320 618054
rect 336354 618020 336420 618054
rect 336454 618020 336520 618054
rect 336554 618020 336620 618054
rect 336654 618020 336720 618054
rect 336754 618020 336820 618054
rect 336854 618020 336927 618054
rect 336233 618006 336927 618020
rect 336233 617972 336292 618006
rect 336326 617972 336382 618006
rect 336416 617972 336472 618006
rect 336506 617972 336562 618006
rect 336596 617972 336652 618006
rect 336686 617972 336742 618006
rect 336776 617972 336832 618006
rect 336866 617972 336927 618006
rect 336233 617954 336927 617972
rect 336233 617920 336320 617954
rect 336354 617920 336420 617954
rect 336454 617920 336520 617954
rect 336554 617920 336620 617954
rect 336654 617920 336720 617954
rect 336754 617920 336820 617954
rect 336854 617920 336927 617954
rect 336233 617916 336927 617920
rect 336233 617882 336292 617916
rect 336326 617882 336382 617916
rect 336416 617882 336472 617916
rect 336506 617882 336562 617916
rect 336596 617882 336652 617916
rect 336686 617882 336742 617916
rect 336776 617882 336832 617916
rect 336866 617882 336927 617916
rect 336233 617854 336927 617882
rect 336233 617826 336320 617854
rect 336354 617826 336420 617854
rect 336233 617792 336292 617826
rect 336354 617820 336382 617826
rect 336326 617792 336382 617820
rect 336416 617820 336420 617826
rect 336454 617826 336520 617854
rect 336454 617820 336472 617826
rect 336416 617792 336472 617820
rect 336506 617820 336520 617826
rect 336554 617826 336620 617854
rect 336654 617826 336720 617854
rect 336754 617826 336820 617854
rect 336854 617826 336927 617854
rect 336554 617820 336562 617826
rect 336506 617792 336562 617820
rect 336596 617820 336620 617826
rect 336686 617820 336720 617826
rect 336776 617820 336820 617826
rect 336596 617792 336652 617820
rect 336686 617792 336742 617820
rect 336776 617792 336832 617820
rect 336866 617792 336927 617826
rect 336233 617733 336927 617792
rect 336988 618395 337008 618429
rect 337042 618428 337406 618429
rect 337042 618395 337156 618428
rect 336988 618394 337156 618395
rect 337190 618394 337257 618428
rect 337291 618414 337406 618428
rect 337440 618414 337459 618448
rect 338277 618484 338444 618489
rect 338478 618484 338545 618518
rect 338579 618508 338786 618518
rect 338820 618508 338876 618542
rect 338910 618508 338966 618542
rect 339000 618508 339056 618542
rect 339090 618508 339146 618542
rect 339180 618508 339236 618542
rect 339270 618508 339326 618542
rect 339360 618508 339416 618542
rect 339450 618508 339506 618542
rect 339540 618518 340074 618542
rect 339540 618508 339732 618518
rect 338579 618489 339732 618508
rect 338579 618484 338747 618489
rect 338277 618448 338747 618484
rect 338277 618429 338694 618448
rect 337291 618394 337459 618414
rect 336988 618358 337459 618394
rect 336988 618339 337406 618358
rect 336988 618305 337008 618339
rect 337042 618338 337406 618339
rect 337042 618305 337156 618338
rect 336988 618304 337156 618305
rect 337190 618304 337257 618338
rect 337291 618324 337406 618338
rect 337440 618324 337459 618358
rect 337291 618304 337459 618324
rect 336988 618268 337459 618304
rect 336988 618249 337406 618268
rect 336988 618215 337008 618249
rect 337042 618248 337406 618249
rect 337042 618215 337156 618248
rect 336988 618214 337156 618215
rect 337190 618214 337257 618248
rect 337291 618234 337406 618248
rect 337440 618234 337459 618268
rect 337291 618214 337459 618234
rect 336988 618178 337459 618214
rect 336988 618159 337406 618178
rect 336988 618125 337008 618159
rect 337042 618158 337406 618159
rect 337042 618125 337156 618158
rect 336988 618124 337156 618125
rect 337190 618124 337257 618158
rect 337291 618144 337406 618158
rect 337440 618144 337459 618178
rect 337291 618124 337459 618144
rect 336988 618088 337459 618124
rect 336988 618069 337406 618088
rect 336988 618035 337008 618069
rect 337042 618068 337406 618069
rect 337042 618035 337156 618068
rect 336988 618034 337156 618035
rect 337190 618034 337257 618068
rect 337291 618054 337406 618068
rect 337440 618054 337459 618088
rect 337291 618034 337459 618054
rect 336988 617998 337459 618034
rect 336988 617979 337406 617998
rect 336988 617945 337008 617979
rect 337042 617978 337406 617979
rect 337042 617945 337156 617978
rect 336988 617944 337156 617945
rect 337190 617944 337257 617978
rect 337291 617964 337406 617978
rect 337440 617964 337459 617998
rect 337291 617944 337459 617964
rect 336988 617908 337459 617944
rect 336988 617889 337406 617908
rect 336988 617855 337008 617889
rect 337042 617888 337406 617889
rect 337042 617855 337156 617888
rect 336988 617854 337156 617855
rect 337190 617854 337257 617888
rect 337291 617874 337406 617888
rect 337440 617874 337459 617908
rect 337291 617854 337459 617874
rect 336988 617818 337459 617854
rect 336988 617799 337406 617818
rect 336988 617765 337008 617799
rect 337042 617798 337406 617799
rect 337042 617765 337156 617798
rect 336988 617764 337156 617765
rect 337190 617764 337257 617798
rect 337291 617784 337406 617798
rect 337440 617784 337459 617818
rect 337291 617764 337459 617784
rect 335688 617709 336118 617728
rect 335688 617675 335720 617709
rect 335754 617708 336118 617709
rect 335754 617675 335868 617708
rect 335688 617674 335868 617675
rect 335902 617674 335969 617708
rect 336003 617694 336118 617708
rect 336152 617694 336188 617728
rect 336003 617674 336188 617694
rect 335688 617671 336188 617674
rect 336988 617728 337459 617764
rect 337521 618366 338215 618427
rect 337521 618332 337580 618366
rect 337614 618354 337670 618366
rect 337642 618332 337670 618354
rect 337704 618354 337760 618366
rect 337704 618332 337708 618354
rect 337521 618320 337608 618332
rect 337642 618320 337708 618332
rect 337742 618332 337760 618354
rect 337794 618354 337850 618366
rect 337794 618332 337808 618354
rect 337742 618320 337808 618332
rect 337842 618332 337850 618354
rect 337884 618354 337940 618366
rect 337974 618354 338030 618366
rect 338064 618354 338120 618366
rect 337884 618332 337908 618354
rect 337974 618332 338008 618354
rect 338064 618332 338108 618354
rect 338154 618332 338215 618366
rect 337842 618320 337908 618332
rect 337942 618320 338008 618332
rect 338042 618320 338108 618332
rect 338142 618320 338215 618332
rect 337521 618276 338215 618320
rect 337521 618242 337580 618276
rect 337614 618254 337670 618276
rect 337642 618242 337670 618254
rect 337704 618254 337760 618276
rect 337704 618242 337708 618254
rect 337521 618220 337608 618242
rect 337642 618220 337708 618242
rect 337742 618242 337760 618254
rect 337794 618254 337850 618276
rect 337794 618242 337808 618254
rect 337742 618220 337808 618242
rect 337842 618242 337850 618254
rect 337884 618254 337940 618276
rect 337974 618254 338030 618276
rect 338064 618254 338120 618276
rect 337884 618242 337908 618254
rect 337974 618242 338008 618254
rect 338064 618242 338108 618254
rect 338154 618242 338215 618276
rect 337842 618220 337908 618242
rect 337942 618220 338008 618242
rect 338042 618220 338108 618242
rect 338142 618220 338215 618242
rect 337521 618186 338215 618220
rect 337521 618152 337580 618186
rect 337614 618154 337670 618186
rect 337642 618152 337670 618154
rect 337704 618154 337760 618186
rect 337704 618152 337708 618154
rect 337521 618120 337608 618152
rect 337642 618120 337708 618152
rect 337742 618152 337760 618154
rect 337794 618154 337850 618186
rect 337794 618152 337808 618154
rect 337742 618120 337808 618152
rect 337842 618152 337850 618154
rect 337884 618154 337940 618186
rect 337974 618154 338030 618186
rect 338064 618154 338120 618186
rect 337884 618152 337908 618154
rect 337974 618152 338008 618154
rect 338064 618152 338108 618154
rect 338154 618152 338215 618186
rect 337842 618120 337908 618152
rect 337942 618120 338008 618152
rect 338042 618120 338108 618152
rect 338142 618120 338215 618152
rect 337521 618096 338215 618120
rect 337521 618062 337580 618096
rect 337614 618062 337670 618096
rect 337704 618062 337760 618096
rect 337794 618062 337850 618096
rect 337884 618062 337940 618096
rect 337974 618062 338030 618096
rect 338064 618062 338120 618096
rect 338154 618062 338215 618096
rect 337521 618054 338215 618062
rect 337521 618020 337608 618054
rect 337642 618020 337708 618054
rect 337742 618020 337808 618054
rect 337842 618020 337908 618054
rect 337942 618020 338008 618054
rect 338042 618020 338108 618054
rect 338142 618020 338215 618054
rect 337521 618006 338215 618020
rect 337521 617972 337580 618006
rect 337614 617972 337670 618006
rect 337704 617972 337760 618006
rect 337794 617972 337850 618006
rect 337884 617972 337940 618006
rect 337974 617972 338030 618006
rect 338064 617972 338120 618006
rect 338154 617972 338215 618006
rect 337521 617954 338215 617972
rect 337521 617920 337608 617954
rect 337642 617920 337708 617954
rect 337742 617920 337808 617954
rect 337842 617920 337908 617954
rect 337942 617920 338008 617954
rect 338042 617920 338108 617954
rect 338142 617920 338215 617954
rect 337521 617916 338215 617920
rect 337521 617882 337580 617916
rect 337614 617882 337670 617916
rect 337704 617882 337760 617916
rect 337794 617882 337850 617916
rect 337884 617882 337940 617916
rect 337974 617882 338030 617916
rect 338064 617882 338120 617916
rect 338154 617882 338215 617916
rect 337521 617854 338215 617882
rect 337521 617826 337608 617854
rect 337642 617826 337708 617854
rect 337521 617792 337580 617826
rect 337642 617820 337670 617826
rect 337614 617792 337670 617820
rect 337704 617820 337708 617826
rect 337742 617826 337808 617854
rect 337742 617820 337760 617826
rect 337704 617792 337760 617820
rect 337794 617820 337808 617826
rect 337842 617826 337908 617854
rect 337942 617826 338008 617854
rect 338042 617826 338108 617854
rect 338142 617826 338215 617854
rect 337842 617820 337850 617826
rect 337794 617792 337850 617820
rect 337884 617820 337908 617826
rect 337974 617820 338008 617826
rect 338064 617820 338108 617826
rect 337884 617792 337940 617820
rect 337974 617792 338030 617820
rect 338064 617792 338120 617820
rect 338154 617792 338215 617826
rect 337521 617733 338215 617792
rect 338277 618395 338296 618429
rect 338330 618428 338694 618429
rect 338330 618395 338444 618428
rect 338277 618394 338444 618395
rect 338478 618394 338545 618428
rect 338579 618414 338694 618428
rect 338728 618414 338747 618448
rect 339565 618484 339732 618489
rect 339766 618484 339833 618518
rect 339867 618508 340074 618518
rect 340108 618508 340164 618542
rect 340198 618508 340254 618542
rect 340288 618508 340344 618542
rect 340378 618508 340434 618542
rect 340468 618508 340524 618542
rect 340558 618508 340614 618542
rect 340648 618508 340704 618542
rect 340738 618508 340794 618542
rect 340828 618518 341088 618542
rect 340828 618508 341020 618518
rect 339867 618489 341020 618508
rect 339867 618484 340035 618489
rect 339565 618448 340035 618484
rect 339565 618429 339982 618448
rect 338579 618394 338747 618414
rect 338277 618358 338747 618394
rect 338277 618339 338694 618358
rect 338277 618305 338296 618339
rect 338330 618338 338694 618339
rect 338330 618305 338444 618338
rect 338277 618304 338444 618305
rect 338478 618304 338545 618338
rect 338579 618324 338694 618338
rect 338728 618324 338747 618358
rect 338579 618304 338747 618324
rect 338277 618268 338747 618304
rect 338277 618249 338694 618268
rect 338277 618215 338296 618249
rect 338330 618248 338694 618249
rect 338330 618215 338444 618248
rect 338277 618214 338444 618215
rect 338478 618214 338545 618248
rect 338579 618234 338694 618248
rect 338728 618234 338747 618268
rect 338579 618214 338747 618234
rect 338277 618178 338747 618214
rect 338277 618159 338694 618178
rect 338277 618125 338296 618159
rect 338330 618158 338694 618159
rect 338330 618125 338444 618158
rect 338277 618124 338444 618125
rect 338478 618124 338545 618158
rect 338579 618144 338694 618158
rect 338728 618144 338747 618178
rect 338579 618124 338747 618144
rect 338277 618088 338747 618124
rect 338277 618069 338694 618088
rect 338277 618035 338296 618069
rect 338330 618068 338694 618069
rect 338330 618035 338444 618068
rect 338277 618034 338444 618035
rect 338478 618034 338545 618068
rect 338579 618054 338694 618068
rect 338728 618054 338747 618088
rect 338579 618034 338747 618054
rect 338277 617998 338747 618034
rect 338277 617979 338694 617998
rect 338277 617945 338296 617979
rect 338330 617978 338694 617979
rect 338330 617945 338444 617978
rect 338277 617944 338444 617945
rect 338478 617944 338545 617978
rect 338579 617964 338694 617978
rect 338728 617964 338747 617998
rect 338579 617944 338747 617964
rect 338277 617908 338747 617944
rect 338277 617889 338694 617908
rect 338277 617855 338296 617889
rect 338330 617888 338694 617889
rect 338330 617855 338444 617888
rect 338277 617854 338444 617855
rect 338478 617854 338545 617888
rect 338579 617874 338694 617888
rect 338728 617874 338747 617908
rect 338579 617854 338747 617874
rect 338277 617818 338747 617854
rect 338277 617799 338694 617818
rect 338277 617765 338296 617799
rect 338330 617798 338694 617799
rect 338330 617765 338444 617798
rect 338277 617764 338444 617765
rect 338478 617764 338545 617798
rect 338579 617784 338694 617798
rect 338728 617784 338747 617818
rect 338579 617764 338747 617784
rect 336988 617709 337406 617728
rect 336988 617675 337008 617709
rect 337042 617708 337406 617709
rect 337042 617675 337156 617708
rect 336988 617674 337156 617675
rect 337190 617674 337257 617708
rect 337291 617694 337406 617708
rect 337440 617694 337459 617728
rect 337291 617674 337459 617694
rect 336988 617671 337459 617674
rect 338277 617728 338747 617764
rect 338809 618366 339503 618427
rect 338809 618332 338868 618366
rect 338902 618354 338958 618366
rect 338930 618332 338958 618354
rect 338992 618354 339048 618366
rect 338992 618332 338996 618354
rect 338809 618320 338896 618332
rect 338930 618320 338996 618332
rect 339030 618332 339048 618354
rect 339082 618354 339138 618366
rect 339082 618332 339096 618354
rect 339030 618320 339096 618332
rect 339130 618332 339138 618354
rect 339172 618354 339228 618366
rect 339262 618354 339318 618366
rect 339352 618354 339408 618366
rect 339172 618332 339196 618354
rect 339262 618332 339296 618354
rect 339352 618332 339396 618354
rect 339442 618332 339503 618366
rect 339130 618320 339196 618332
rect 339230 618320 339296 618332
rect 339330 618320 339396 618332
rect 339430 618320 339503 618332
rect 338809 618276 339503 618320
rect 338809 618242 338868 618276
rect 338902 618254 338958 618276
rect 338930 618242 338958 618254
rect 338992 618254 339048 618276
rect 338992 618242 338996 618254
rect 338809 618220 338896 618242
rect 338930 618220 338996 618242
rect 339030 618242 339048 618254
rect 339082 618254 339138 618276
rect 339082 618242 339096 618254
rect 339030 618220 339096 618242
rect 339130 618242 339138 618254
rect 339172 618254 339228 618276
rect 339262 618254 339318 618276
rect 339352 618254 339408 618276
rect 339172 618242 339196 618254
rect 339262 618242 339296 618254
rect 339352 618242 339396 618254
rect 339442 618242 339503 618276
rect 339130 618220 339196 618242
rect 339230 618220 339296 618242
rect 339330 618220 339396 618242
rect 339430 618220 339503 618242
rect 338809 618186 339503 618220
rect 338809 618152 338868 618186
rect 338902 618154 338958 618186
rect 338930 618152 338958 618154
rect 338992 618154 339048 618186
rect 338992 618152 338996 618154
rect 338809 618120 338896 618152
rect 338930 618120 338996 618152
rect 339030 618152 339048 618154
rect 339082 618154 339138 618186
rect 339082 618152 339096 618154
rect 339030 618120 339096 618152
rect 339130 618152 339138 618154
rect 339172 618154 339228 618186
rect 339262 618154 339318 618186
rect 339352 618154 339408 618186
rect 339172 618152 339196 618154
rect 339262 618152 339296 618154
rect 339352 618152 339396 618154
rect 339442 618152 339503 618186
rect 339130 618120 339196 618152
rect 339230 618120 339296 618152
rect 339330 618120 339396 618152
rect 339430 618120 339503 618152
rect 338809 618096 339503 618120
rect 338809 618062 338868 618096
rect 338902 618062 338958 618096
rect 338992 618062 339048 618096
rect 339082 618062 339138 618096
rect 339172 618062 339228 618096
rect 339262 618062 339318 618096
rect 339352 618062 339408 618096
rect 339442 618062 339503 618096
rect 338809 618054 339503 618062
rect 338809 618020 338896 618054
rect 338930 618020 338996 618054
rect 339030 618020 339096 618054
rect 339130 618020 339196 618054
rect 339230 618020 339296 618054
rect 339330 618020 339396 618054
rect 339430 618020 339503 618054
rect 338809 618006 339503 618020
rect 338809 617972 338868 618006
rect 338902 617972 338958 618006
rect 338992 617972 339048 618006
rect 339082 617972 339138 618006
rect 339172 617972 339228 618006
rect 339262 617972 339318 618006
rect 339352 617972 339408 618006
rect 339442 617972 339503 618006
rect 338809 617954 339503 617972
rect 338809 617920 338896 617954
rect 338930 617920 338996 617954
rect 339030 617920 339096 617954
rect 339130 617920 339196 617954
rect 339230 617920 339296 617954
rect 339330 617920 339396 617954
rect 339430 617920 339503 617954
rect 338809 617916 339503 617920
rect 338809 617882 338868 617916
rect 338902 617882 338958 617916
rect 338992 617882 339048 617916
rect 339082 617882 339138 617916
rect 339172 617882 339228 617916
rect 339262 617882 339318 617916
rect 339352 617882 339408 617916
rect 339442 617882 339503 617916
rect 338809 617854 339503 617882
rect 338809 617826 338896 617854
rect 338930 617826 338996 617854
rect 338809 617792 338868 617826
rect 338930 617820 338958 617826
rect 338902 617792 338958 617820
rect 338992 617820 338996 617826
rect 339030 617826 339096 617854
rect 339030 617820 339048 617826
rect 338992 617792 339048 617820
rect 339082 617820 339096 617826
rect 339130 617826 339196 617854
rect 339230 617826 339296 617854
rect 339330 617826 339396 617854
rect 339430 617826 339503 617854
rect 339130 617820 339138 617826
rect 339082 617792 339138 617820
rect 339172 617820 339196 617826
rect 339262 617820 339296 617826
rect 339352 617820 339396 617826
rect 339172 617792 339228 617820
rect 339262 617792 339318 617820
rect 339352 617792 339408 617820
rect 339442 617792 339503 617826
rect 338809 617733 339503 617792
rect 339565 618395 339584 618429
rect 339618 618428 339982 618429
rect 339618 618395 339732 618428
rect 339565 618394 339732 618395
rect 339766 618394 339833 618428
rect 339867 618414 339982 618428
rect 340016 618414 340035 618448
rect 340853 618484 341020 618489
rect 341054 618484 341088 618518
rect 340853 618429 341088 618484
rect 339867 618394 340035 618414
rect 339565 618358 340035 618394
rect 339565 618339 339982 618358
rect 339565 618305 339584 618339
rect 339618 618338 339982 618339
rect 339618 618305 339732 618338
rect 339565 618304 339732 618305
rect 339766 618304 339833 618338
rect 339867 618324 339982 618338
rect 340016 618324 340035 618358
rect 339867 618304 340035 618324
rect 339565 618268 340035 618304
rect 339565 618249 339982 618268
rect 339565 618215 339584 618249
rect 339618 618248 339982 618249
rect 339618 618215 339732 618248
rect 339565 618214 339732 618215
rect 339766 618214 339833 618248
rect 339867 618234 339982 618248
rect 340016 618234 340035 618268
rect 339867 618214 340035 618234
rect 339565 618178 340035 618214
rect 339565 618159 339982 618178
rect 339565 618125 339584 618159
rect 339618 618158 339982 618159
rect 339618 618125 339732 618158
rect 339565 618124 339732 618125
rect 339766 618124 339833 618158
rect 339867 618144 339982 618158
rect 340016 618144 340035 618178
rect 339867 618124 340035 618144
rect 339565 618088 340035 618124
rect 339565 618069 339982 618088
rect 339565 618035 339584 618069
rect 339618 618068 339982 618069
rect 339618 618035 339732 618068
rect 339565 618034 339732 618035
rect 339766 618034 339833 618068
rect 339867 618054 339982 618068
rect 340016 618054 340035 618088
rect 339867 618034 340035 618054
rect 339565 617998 340035 618034
rect 339565 617979 339982 617998
rect 339565 617945 339584 617979
rect 339618 617978 339982 617979
rect 339618 617945 339732 617978
rect 339565 617944 339732 617945
rect 339766 617944 339833 617978
rect 339867 617964 339982 617978
rect 340016 617964 340035 617998
rect 339867 617944 340035 617964
rect 339565 617908 340035 617944
rect 339565 617889 339982 617908
rect 339565 617855 339584 617889
rect 339618 617888 339982 617889
rect 339618 617855 339732 617888
rect 339565 617854 339732 617855
rect 339766 617854 339833 617888
rect 339867 617874 339982 617888
rect 340016 617874 340035 617908
rect 339867 617854 340035 617874
rect 339565 617818 340035 617854
rect 339565 617799 339982 617818
rect 339565 617765 339584 617799
rect 339618 617798 339982 617799
rect 339618 617765 339732 617798
rect 339565 617764 339732 617765
rect 339766 617764 339833 617798
rect 339867 617784 339982 617798
rect 340016 617784 340035 617818
rect 339867 617764 340035 617784
rect 338277 617709 338694 617728
rect 338277 617675 338296 617709
rect 338330 617708 338694 617709
rect 338330 617675 338444 617708
rect 338277 617674 338444 617675
rect 338478 617674 338545 617708
rect 338579 617694 338694 617708
rect 338728 617694 338747 617728
rect 338579 617674 338747 617694
rect 338277 617671 338747 617674
rect 339565 617728 340035 617764
rect 340097 618366 340791 618427
rect 340097 618332 340156 618366
rect 340190 618354 340246 618366
rect 340218 618332 340246 618354
rect 340280 618354 340336 618366
rect 340280 618332 340284 618354
rect 340097 618320 340184 618332
rect 340218 618320 340284 618332
rect 340318 618332 340336 618354
rect 340370 618354 340426 618366
rect 340370 618332 340384 618354
rect 340318 618320 340384 618332
rect 340418 618332 340426 618354
rect 340460 618354 340516 618366
rect 340550 618354 340606 618366
rect 340640 618354 340696 618366
rect 340460 618332 340484 618354
rect 340550 618332 340584 618354
rect 340640 618332 340684 618354
rect 340730 618332 340791 618366
rect 340418 618320 340484 618332
rect 340518 618320 340584 618332
rect 340618 618320 340684 618332
rect 340718 618320 340791 618332
rect 340097 618276 340791 618320
rect 340097 618242 340156 618276
rect 340190 618254 340246 618276
rect 340218 618242 340246 618254
rect 340280 618254 340336 618276
rect 340280 618242 340284 618254
rect 340097 618220 340184 618242
rect 340218 618220 340284 618242
rect 340318 618242 340336 618254
rect 340370 618254 340426 618276
rect 340370 618242 340384 618254
rect 340318 618220 340384 618242
rect 340418 618242 340426 618254
rect 340460 618254 340516 618276
rect 340550 618254 340606 618276
rect 340640 618254 340696 618276
rect 340460 618242 340484 618254
rect 340550 618242 340584 618254
rect 340640 618242 340684 618254
rect 340730 618242 340791 618276
rect 340418 618220 340484 618242
rect 340518 618220 340584 618242
rect 340618 618220 340684 618242
rect 340718 618220 340791 618242
rect 340097 618186 340791 618220
rect 340097 618152 340156 618186
rect 340190 618154 340246 618186
rect 340218 618152 340246 618154
rect 340280 618154 340336 618186
rect 340280 618152 340284 618154
rect 340097 618120 340184 618152
rect 340218 618120 340284 618152
rect 340318 618152 340336 618154
rect 340370 618154 340426 618186
rect 340370 618152 340384 618154
rect 340318 618120 340384 618152
rect 340418 618152 340426 618154
rect 340460 618154 340516 618186
rect 340550 618154 340606 618186
rect 340640 618154 340696 618186
rect 340460 618152 340484 618154
rect 340550 618152 340584 618154
rect 340640 618152 340684 618154
rect 340730 618152 340791 618186
rect 340418 618120 340484 618152
rect 340518 618120 340584 618152
rect 340618 618120 340684 618152
rect 340718 618120 340791 618152
rect 340097 618096 340791 618120
rect 340097 618062 340156 618096
rect 340190 618062 340246 618096
rect 340280 618062 340336 618096
rect 340370 618062 340426 618096
rect 340460 618062 340516 618096
rect 340550 618062 340606 618096
rect 340640 618062 340696 618096
rect 340730 618062 340791 618096
rect 340097 618054 340791 618062
rect 340097 618020 340184 618054
rect 340218 618020 340284 618054
rect 340318 618020 340384 618054
rect 340418 618020 340484 618054
rect 340518 618020 340584 618054
rect 340618 618020 340684 618054
rect 340718 618020 340791 618054
rect 340097 618006 340791 618020
rect 340097 617972 340156 618006
rect 340190 617972 340246 618006
rect 340280 617972 340336 618006
rect 340370 617972 340426 618006
rect 340460 617972 340516 618006
rect 340550 617972 340606 618006
rect 340640 617972 340696 618006
rect 340730 617972 340791 618006
rect 340097 617954 340791 617972
rect 340097 617920 340184 617954
rect 340218 617920 340284 617954
rect 340318 617920 340384 617954
rect 340418 617920 340484 617954
rect 340518 617920 340584 617954
rect 340618 617920 340684 617954
rect 340718 617920 340791 617954
rect 340097 617916 340791 617920
rect 340097 617882 340156 617916
rect 340190 617882 340246 617916
rect 340280 617882 340336 617916
rect 340370 617882 340426 617916
rect 340460 617882 340516 617916
rect 340550 617882 340606 617916
rect 340640 617882 340696 617916
rect 340730 617882 340791 617916
rect 340097 617854 340791 617882
rect 340097 617826 340184 617854
rect 340218 617826 340284 617854
rect 340097 617792 340156 617826
rect 340218 617820 340246 617826
rect 340190 617792 340246 617820
rect 340280 617820 340284 617826
rect 340318 617826 340384 617854
rect 340318 617820 340336 617826
rect 340280 617792 340336 617820
rect 340370 617820 340384 617826
rect 340418 617826 340484 617854
rect 340518 617826 340584 617854
rect 340618 617826 340684 617854
rect 340718 617826 340791 617854
rect 340418 617820 340426 617826
rect 340370 617792 340426 617820
rect 340460 617820 340484 617826
rect 340550 617820 340584 617826
rect 340640 617820 340684 617826
rect 340460 617792 340516 617820
rect 340550 617792 340606 617820
rect 340640 617792 340696 617820
rect 340730 617792 340791 617826
rect 340097 617733 340791 617792
rect 340853 618395 340872 618429
rect 340906 618428 341088 618429
rect 340906 618395 341020 618428
rect 340853 618394 341020 618395
rect 341054 618394 341088 618428
rect 340853 618339 341088 618394
rect 340853 618305 340872 618339
rect 340906 618338 341088 618339
rect 340906 618305 341020 618338
rect 340853 618304 341020 618305
rect 341054 618304 341088 618338
rect 340853 618249 341088 618304
rect 340853 618215 340872 618249
rect 340906 618248 341088 618249
rect 340906 618215 341020 618248
rect 340853 618214 341020 618215
rect 341054 618214 341088 618248
rect 340853 618159 341088 618214
rect 340853 618125 340872 618159
rect 340906 618158 341088 618159
rect 340906 618125 341020 618158
rect 340853 618124 341020 618125
rect 341054 618124 341088 618158
rect 340853 618069 341088 618124
rect 340853 618035 340872 618069
rect 340906 618068 341088 618069
rect 340906 618035 341020 618068
rect 340853 618034 341020 618035
rect 341054 618034 341088 618068
rect 340853 617979 341088 618034
rect 340853 617945 340872 617979
rect 340906 617978 341088 617979
rect 340906 617945 341020 617978
rect 340853 617944 341020 617945
rect 341054 617944 341088 617978
rect 340853 617889 341088 617944
rect 340853 617855 340872 617889
rect 340906 617888 341088 617889
rect 340906 617855 341020 617888
rect 340853 617854 341020 617855
rect 341054 617854 341088 617888
rect 340853 617799 341088 617854
rect 340853 617765 340872 617799
rect 340906 617798 341088 617799
rect 340906 617765 341020 617798
rect 340853 617764 341020 617765
rect 341054 617764 341088 617798
rect 339565 617709 339982 617728
rect 339565 617675 339584 617709
rect 339618 617708 339982 617709
rect 339618 617675 339732 617708
rect 339565 617674 339732 617675
rect 339766 617674 339833 617708
rect 339867 617694 339982 617708
rect 340016 617694 340035 617728
rect 339867 617674 340035 617694
rect 339565 617671 340035 617674
rect 340853 617709 341088 617764
rect 340853 617675 340872 617709
rect 340906 617708 341088 617709
rect 340906 617675 341020 617708
rect 340853 617674 341020 617675
rect 341054 617674 341088 617708
rect 340853 617671 341088 617674
rect 334648 617652 341088 617671
rect 334648 617618 334888 617652
rect 334922 617618 334978 617652
rect 335012 617618 335068 617652
rect 335102 617618 335158 617652
rect 335192 617618 335248 617652
rect 335282 617618 335338 617652
rect 335372 617618 335428 617652
rect 335462 617618 335518 617652
rect 335552 617618 335608 617652
rect 335642 617618 336176 617652
rect 336210 617618 336266 617652
rect 336300 617618 336356 617652
rect 336390 617618 336446 617652
rect 336480 617618 336536 617652
rect 336570 617618 336626 617652
rect 336660 617618 336716 617652
rect 336750 617618 336806 617652
rect 336840 617618 336896 617652
rect 336930 617618 337464 617652
rect 337498 617618 337554 617652
rect 337588 617618 337644 617652
rect 337678 617618 337734 617652
rect 337768 617618 337824 617652
rect 337858 617618 337914 617652
rect 337948 617618 338004 617652
rect 338038 617618 338094 617652
rect 338128 617618 338184 617652
rect 338218 617618 338752 617652
rect 338786 617618 338842 617652
rect 338876 617618 338932 617652
rect 338966 617618 339022 617652
rect 339056 617618 339112 617652
rect 339146 617618 339202 617652
rect 339236 617618 339292 617652
rect 339326 617618 339382 617652
rect 339416 617618 339472 617652
rect 339506 617618 340040 617652
rect 340074 617618 340130 617652
rect 340164 617618 340220 617652
rect 340254 617618 340310 617652
rect 340344 617618 340400 617652
rect 340434 617618 340490 617652
rect 340524 617618 340580 617652
rect 340614 617618 340670 617652
rect 340704 617618 340760 617652
rect 340794 617618 341088 617652
rect 334648 617584 334681 617618
rect 334715 617599 335868 617618
rect 334715 617584 334888 617599
rect 334648 617535 334888 617584
rect 335688 617584 335868 617599
rect 335902 617584 335969 617618
rect 336003 617599 337156 617618
rect 336003 617584 336188 617599
rect 335688 617535 336188 617584
rect 336988 617584 337156 617599
rect 337190 617584 337257 617618
rect 337291 617599 338444 617618
rect 337291 617584 337388 617599
rect 336988 617535 337388 617584
rect 338288 617584 338444 617599
rect 338478 617584 338545 617618
rect 338579 617599 339732 617618
rect 338579 617584 338688 617599
rect 338288 617535 338688 617584
rect 339588 617584 339732 617599
rect 339766 617584 339833 617618
rect 339867 617599 341020 617618
rect 339867 617584 339988 617599
rect 339588 617535 339988 617584
rect 340888 617584 341020 617599
rect 341054 617584 341088 617618
rect 340888 617535 341088 617584
rect 334648 617528 341088 617535
rect 334648 617494 334681 617528
rect 334715 617505 335868 617528
rect 334715 617494 334782 617505
rect 334648 617471 334782 617494
rect 334816 617471 334872 617505
rect 334906 617471 334962 617505
rect 334996 617471 335052 617505
rect 335086 617471 335142 617505
rect 335176 617471 335232 617505
rect 335266 617471 335322 617505
rect 335356 617471 335412 617505
rect 335446 617471 335502 617505
rect 335536 617471 335592 617505
rect 335626 617471 335682 617505
rect 335716 617471 335772 617505
rect 335806 617494 335868 617505
rect 335902 617494 335969 617528
rect 336003 617505 337156 617528
rect 336003 617494 336070 617505
rect 335806 617471 336070 617494
rect 336104 617471 336160 617505
rect 336194 617471 336250 617505
rect 336284 617471 336340 617505
rect 336374 617471 336430 617505
rect 336464 617471 336520 617505
rect 336554 617471 336610 617505
rect 336644 617471 336700 617505
rect 336734 617471 336790 617505
rect 336824 617471 336880 617505
rect 336914 617471 336970 617505
rect 337004 617471 337060 617505
rect 337094 617494 337156 617505
rect 337190 617494 337257 617528
rect 337291 617505 338444 617528
rect 337291 617494 337358 617505
rect 337094 617471 337358 617494
rect 337392 617471 337448 617505
rect 337482 617471 337538 617505
rect 337572 617471 337628 617505
rect 337662 617471 337718 617505
rect 337752 617471 337808 617505
rect 337842 617471 337898 617505
rect 337932 617471 337988 617505
rect 338022 617471 338078 617505
rect 338112 617471 338168 617505
rect 338202 617471 338258 617505
rect 338292 617471 338348 617505
rect 338382 617494 338444 617505
rect 338478 617494 338545 617528
rect 338579 617505 339732 617528
rect 338579 617494 338646 617505
rect 338382 617471 338646 617494
rect 338680 617471 338736 617505
rect 338770 617471 338826 617505
rect 338860 617471 338916 617505
rect 338950 617471 339006 617505
rect 339040 617471 339096 617505
rect 339130 617471 339186 617505
rect 339220 617471 339276 617505
rect 339310 617471 339366 617505
rect 339400 617471 339456 617505
rect 339490 617471 339546 617505
rect 339580 617471 339636 617505
rect 339670 617494 339732 617505
rect 339766 617494 339833 617528
rect 339867 617505 341020 617528
rect 339867 617494 339934 617505
rect 339670 617471 339934 617494
rect 339968 617471 340024 617505
rect 340058 617471 340114 617505
rect 340148 617471 340204 617505
rect 340238 617471 340294 617505
rect 340328 617471 340384 617505
rect 340418 617471 340474 617505
rect 340508 617471 340564 617505
rect 340598 617471 340654 617505
rect 340688 617471 340744 617505
rect 340778 617471 340834 617505
rect 340868 617471 340924 617505
rect 340958 617494 341020 617505
rect 341054 617494 341088 617528
rect 340958 617471 341088 617494
rect 334648 617436 341088 617471
rect 334688 617424 334888 617436
rect 335688 617424 336188 617436
rect 340888 617424 341088 617436
rect 330070 616606 330170 616706
rect 330570 616606 330670 616706
rect 330070 616506 330670 616606
rect 297800 616456 298888 616472
rect 297800 615464 298824 616456
rect 297800 615448 298876 615464
rect 298976 615448 299100 615464
rect 299200 615448 299324 615464
rect 299424 615448 299548 615464
rect 299648 615448 299772 615464
rect 299872 615448 299996 615464
rect 300096 615448 300220 615464
rect 300320 615448 300444 615464
rect 300544 615448 300668 615464
rect 300768 615448 300892 615464
rect 300992 615448 301116 615464
rect 301216 615448 301340 615464
rect 301440 615448 301564 615464
rect 301664 615448 301788 615464
rect 301888 615448 302012 615464
rect 302112 615448 302236 615464
rect 302336 615448 302460 615464
rect 302560 615448 302684 615464
rect 302784 615448 302908 615464
rect 303008 615448 303132 615464
rect 303232 615448 303356 615464
rect 303456 615448 303580 615464
rect 303680 615448 303804 615464
rect 303904 615448 304028 615464
rect 304128 615448 304252 615464
rect 304352 615448 304476 615464
rect 304576 615448 304700 615464
rect 304800 615448 304924 615464
rect 305024 615448 305148 615464
rect 305248 615448 305372 615464
rect 305472 615448 309346 615464
rect 309446 615448 309570 615464
rect 309670 615448 309794 615464
rect 309894 615448 310018 615464
rect 310118 615448 310242 615464
rect 310342 615448 310466 615464
rect 310566 615448 310690 615464
rect 310790 615448 310914 615464
rect 311014 615448 311138 615464
rect 311238 615448 311362 615464
rect 311462 615448 311586 615464
rect 311686 615448 311810 615464
rect 311910 615448 312034 615464
rect 312134 615448 312258 615464
rect 312358 615448 312482 615464
rect 312582 615448 312706 615464
rect 312806 615448 312930 615464
rect 313030 615448 313154 615464
rect 313254 615448 313378 615464
rect 313478 615448 313602 615464
rect 313702 615448 313826 615464
rect 313926 615448 314050 615464
rect 314150 615448 314274 615464
rect 314374 615448 314498 615464
rect 314598 615448 314722 615464
rect 314822 615448 314946 615464
rect 315046 615448 315170 615464
rect 315270 615448 315394 615464
rect 315494 615448 315618 615464
rect 315718 615448 315842 615464
rect 315942 615448 335616 615464
rect 335716 615448 335840 615464
rect 335940 615448 336064 615464
rect 336164 615448 336288 615464
rect 336388 615448 336512 615464
rect 336612 615448 336736 615464
rect 336836 615448 336960 615464
rect 337060 615448 337184 615464
rect 337284 615448 337408 615464
rect 337508 615448 337632 615464
rect 337732 615448 337856 615464
rect 337956 615448 338080 615464
rect 338180 615448 338304 615464
rect 338404 615448 338528 615464
rect 338628 615448 338752 615464
rect 338852 615448 338976 615464
rect 339076 615448 339200 615464
rect 339300 615448 339424 615464
rect 339524 615448 339648 615464
rect 339748 615448 339872 615464
rect 339972 615448 340096 615464
rect 340196 615448 340320 615464
rect 340420 615448 340544 615464
rect 340644 615448 340768 615464
rect 340868 615448 340992 615464
rect 297800 614448 297848 615448
rect 341092 615424 341104 615464
rect 341092 615394 341216 615424
rect 341316 615394 341440 615424
rect 341540 615394 341664 615424
rect 341764 615394 341888 615424
rect 342096 615424 342112 640648
rect 343112 637996 343160 640648
rect 343126 637896 343160 637996
rect 343112 637772 343160 637896
rect 343126 637672 343160 637772
rect 343112 637548 343160 637672
rect 343126 637448 343160 637548
rect 343112 637324 343160 637448
rect 343126 637224 343160 637324
rect 343112 637100 343160 637224
rect 343126 637000 343160 637100
rect 343112 636876 343160 637000
rect 343126 636776 343160 636876
rect 343112 636652 343160 636776
rect 343126 636552 343160 636652
rect 343112 636428 343160 636552
rect 343126 636328 343160 636428
rect 343112 636204 343160 636328
rect 343126 636104 343160 636204
rect 343112 635980 343160 636104
rect 343126 635880 343160 635980
rect 343112 635756 343160 635880
rect 343126 635656 343160 635756
rect 343112 635532 343160 635656
rect 343126 635432 343160 635532
rect 343112 635308 343160 635432
rect 343126 635208 343160 635308
rect 343112 635084 343160 635208
rect 343126 634984 343160 635084
rect 343112 634860 343160 634984
rect 343126 634760 343160 634860
rect 343112 634636 343160 634760
rect 343126 634536 343160 634636
rect 343112 634412 343160 634536
rect 343126 634312 343160 634412
rect 343112 634188 343160 634312
rect 343126 634088 343160 634188
rect 343112 633964 343160 634088
rect 343126 633864 343160 633964
rect 343112 633740 343160 633864
rect 343126 633640 343160 633740
rect 343112 633516 343160 633640
rect 343126 633416 343160 633516
rect 343112 633292 343160 633416
rect 343126 633192 343160 633292
rect 343112 633068 343160 633192
rect 343126 632968 343160 633068
rect 343112 632844 343160 632968
rect 343126 632744 343160 632844
rect 343112 632620 343160 632744
rect 343126 632520 343160 632620
rect 343112 632396 343160 632520
rect 343126 632296 343160 632396
rect 343112 632172 343160 632296
rect 343126 632072 343160 632172
rect 343112 631948 343160 632072
rect 343126 631848 343160 631948
rect 343112 631724 343160 631848
rect 343126 631624 343160 631724
rect 343112 631500 343160 631624
rect 343126 631400 343160 631500
rect 343112 624596 343160 631400
rect 343126 624496 343160 624596
rect 343112 624372 343160 624496
rect 343126 624272 343160 624372
rect 343112 624148 343160 624272
rect 343126 624048 343160 624148
rect 343112 623924 343160 624048
rect 343126 623824 343160 623924
rect 343112 623700 343160 623824
rect 343126 623600 343160 623700
rect 343112 623476 343160 623600
rect 343126 623376 343160 623476
rect 343112 623252 343160 623376
rect 343126 623152 343160 623252
rect 343112 623028 343160 623152
rect 343126 622928 343160 623028
rect 343112 622804 343160 622928
rect 343126 622704 343160 622804
rect 343112 622580 343160 622704
rect 343126 622480 343160 622580
rect 343112 622356 343160 622480
rect 343126 622256 343160 622356
rect 343112 622132 343160 622256
rect 343126 622032 343160 622132
rect 343112 621908 343160 622032
rect 343126 621808 343160 621908
rect 343112 621684 343160 621808
rect 343126 621584 343160 621684
rect 343112 621460 343160 621584
rect 343126 621360 343160 621460
rect 343112 621236 343160 621360
rect 343126 621136 343160 621236
rect 343112 621012 343160 621136
rect 343126 620912 343160 621012
rect 343112 620788 343160 620912
rect 343126 620688 343160 620788
rect 343112 620564 343160 620688
rect 343126 620464 343160 620564
rect 343112 620340 343160 620464
rect 343126 620240 343160 620340
rect 343112 620116 343160 620240
rect 343126 620016 343160 620116
rect 343112 619892 343160 620016
rect 343126 619792 343160 619892
rect 343112 619668 343160 619792
rect 343126 619568 343160 619668
rect 343112 619444 343160 619568
rect 343126 619344 343160 619444
rect 343112 619220 343160 619344
rect 343126 619120 343160 619220
rect 343112 618996 343160 619120
rect 343126 618896 343160 618996
rect 343112 618772 343160 618896
rect 343126 618672 343160 618772
rect 343112 618548 343160 618672
rect 343126 618448 343160 618548
rect 343112 618324 343160 618448
rect 343126 618224 343160 618324
rect 343112 618100 343160 618224
rect 343126 618000 343160 618100
rect 341988 615394 342112 615424
rect 341088 615270 342112 615394
rect 341092 615170 341216 615270
rect 341316 615170 341440 615270
rect 341540 615170 341664 615270
rect 341764 615170 341888 615270
rect 341988 615170 342112 615270
rect 341088 615046 342112 615170
rect 341092 614946 341216 615046
rect 341316 614946 341440 615046
rect 341540 614946 341664 615046
rect 341764 614946 341888 615046
rect 341988 614946 342112 615046
rect 341088 614822 342112 614946
rect 341092 614722 341216 614822
rect 341316 614722 341440 614822
rect 341540 614722 341664 614822
rect 341764 614722 341888 614822
rect 341988 614722 342112 614822
rect 341088 614598 342112 614722
rect 341092 614498 341216 614598
rect 341316 614498 341440 614598
rect 341540 614498 341664 614598
rect 341764 614498 341888 614598
rect 341988 614498 342112 614598
rect 341088 614448 342112 614498
rect 297800 614432 342112 614448
rect 297800 614400 298824 614432
rect 340112 614424 342112 614432
rect 343112 614424 343160 618000
rect 340112 614400 343160 614424
<< viali >>
rect 298876 642672 298976 642694
rect 299100 642672 299200 642694
rect 299324 642672 299424 642694
rect 299548 642672 299648 642694
rect 299772 642672 299872 642694
rect 299996 642672 300096 642694
rect 300220 642672 300320 642694
rect 300444 642672 300544 642694
rect 300668 642672 300768 642694
rect 300892 642672 300992 642694
rect 301116 642672 301216 642694
rect 301340 642672 301440 642694
rect 301564 642672 301664 642694
rect 301788 642672 301888 642694
rect 302012 642672 302112 642694
rect 302236 642672 302336 642694
rect 302460 642672 302560 642694
rect 302684 642672 302784 642694
rect 302908 642672 303008 642694
rect 303132 642672 303232 642694
rect 303356 642672 303456 642694
rect 303580 642672 303680 642694
rect 303804 642672 303904 642694
rect 304028 642672 304128 642694
rect 304252 642672 304352 642694
rect 304476 642672 304576 642694
rect 304700 642672 304800 642694
rect 304924 642672 305024 642694
rect 305148 642672 305248 642694
rect 305372 642672 305472 642694
rect 309346 642672 309446 642694
rect 309570 642672 309670 642694
rect 309794 642672 309894 642694
rect 310018 642672 310118 642694
rect 310242 642672 310342 642694
rect 310466 642672 310566 642694
rect 310690 642672 310790 642694
rect 310914 642672 311014 642694
rect 311138 642672 311238 642694
rect 311362 642672 311462 642694
rect 311586 642672 311686 642694
rect 311810 642672 311910 642694
rect 312034 642672 312134 642694
rect 312258 642672 312358 642694
rect 312482 642672 312582 642694
rect 312706 642672 312806 642694
rect 312930 642672 313030 642694
rect 313154 642672 313254 642694
rect 313378 642672 313478 642694
rect 313602 642672 313702 642694
rect 313826 642672 313926 642694
rect 314050 642672 314150 642694
rect 314274 642672 314374 642694
rect 314498 642672 314598 642694
rect 314722 642672 314822 642694
rect 314946 642672 315046 642694
rect 315170 642672 315270 642694
rect 315394 642672 315494 642694
rect 315618 642672 315718 642694
rect 315842 642672 315942 642694
rect 335616 642672 335716 642714
rect 335840 642672 335940 642714
rect 336064 642672 336164 642714
rect 336288 642672 336388 642714
rect 336512 642672 336612 642714
rect 336736 642672 336836 642714
rect 336960 642672 337060 642714
rect 337184 642672 337284 642714
rect 337408 642672 337508 642714
rect 337632 642672 337732 642714
rect 337856 642672 337956 642714
rect 338080 642672 338180 642714
rect 338304 642672 338404 642714
rect 338528 642672 338628 642714
rect 338752 642672 338852 642714
rect 338976 642672 339076 642714
rect 339200 642672 339300 642714
rect 339424 642672 339524 642714
rect 339648 642672 339748 642714
rect 339872 642672 339972 642714
rect 340096 642672 340196 642714
rect 340320 642672 340420 642714
rect 340544 642672 340644 642714
rect 340768 642672 340868 642714
rect 340992 642672 341092 642714
rect 341216 642672 341316 642714
rect 341440 642672 341540 642714
rect 341664 642672 341764 642714
rect 341888 642672 341988 642714
rect 342112 642672 342212 642714
rect 298876 642594 298976 642672
rect 299100 642594 299200 642672
rect 299324 642594 299424 642672
rect 299548 642594 299648 642672
rect 299772 642594 299872 642672
rect 299996 642594 300096 642672
rect 300220 642594 300320 642672
rect 300444 642594 300544 642672
rect 300668 642594 300768 642672
rect 300892 642594 300992 642672
rect 301116 642594 301216 642672
rect 301340 642594 301440 642672
rect 301564 642594 301664 642672
rect 301788 642594 301888 642672
rect 302012 642594 302112 642672
rect 302236 642594 302336 642672
rect 302460 642594 302560 642672
rect 302684 642594 302784 642672
rect 302908 642594 303008 642672
rect 303132 642594 303232 642672
rect 303356 642594 303456 642672
rect 303580 642594 303680 642672
rect 303804 642594 303904 642672
rect 304028 642594 304128 642672
rect 304252 642594 304352 642672
rect 304476 642594 304576 642672
rect 304700 642594 304800 642672
rect 304924 642594 305024 642672
rect 305148 642594 305248 642672
rect 305372 642594 305472 642672
rect 309346 642594 309446 642672
rect 309570 642594 309670 642672
rect 309794 642594 309894 642672
rect 310018 642594 310118 642672
rect 310242 642594 310342 642672
rect 310466 642594 310566 642672
rect 310690 642594 310790 642672
rect 310914 642594 311014 642672
rect 311138 642594 311238 642672
rect 311362 642594 311462 642672
rect 311586 642594 311686 642672
rect 311810 642594 311910 642672
rect 312034 642594 312134 642672
rect 312258 642594 312358 642672
rect 312482 642594 312582 642672
rect 312706 642594 312806 642672
rect 312930 642594 313030 642672
rect 313154 642594 313254 642672
rect 313378 642594 313478 642672
rect 313602 642594 313702 642672
rect 313826 642594 313926 642672
rect 314050 642594 314150 642672
rect 314274 642594 314374 642672
rect 314498 642594 314598 642672
rect 314722 642594 314822 642672
rect 314946 642594 315046 642672
rect 315170 642594 315270 642672
rect 315394 642594 315494 642672
rect 315618 642594 315718 642672
rect 315842 642594 315942 642672
rect 335616 642614 335716 642672
rect 335840 642614 335940 642672
rect 336064 642614 336164 642672
rect 336288 642614 336388 642672
rect 336512 642614 336612 642672
rect 336736 642614 336836 642672
rect 336960 642614 337060 642672
rect 337184 642614 337284 642672
rect 337408 642614 337508 642672
rect 337632 642614 337732 642672
rect 337856 642614 337956 642672
rect 338080 642614 338180 642672
rect 338304 642614 338404 642672
rect 338528 642614 338628 642672
rect 338752 642614 338852 642672
rect 338976 642614 339076 642672
rect 339200 642614 339300 642672
rect 339424 642614 339524 642672
rect 339648 642614 339748 642672
rect 339872 642614 339972 642672
rect 340096 642614 340196 642672
rect 340320 642614 340420 642672
rect 340544 642614 340644 642672
rect 340768 642614 340868 642672
rect 340992 642614 341092 642672
rect 341216 642614 341316 642672
rect 341440 642614 341540 642672
rect 341664 642614 341764 642672
rect 341888 642614 341988 642672
rect 342112 642614 342212 642672
rect 298876 642370 298976 642470
rect 299100 642370 299200 642470
rect 299324 642370 299424 642470
rect 299548 642370 299648 642470
rect 299772 642370 299872 642470
rect 299996 642370 300096 642470
rect 300220 642370 300320 642470
rect 300444 642370 300544 642470
rect 300668 642370 300768 642470
rect 300892 642370 300992 642470
rect 301116 642370 301216 642470
rect 301340 642370 301440 642470
rect 301564 642370 301664 642470
rect 301788 642370 301888 642470
rect 302012 642370 302112 642470
rect 302236 642370 302336 642470
rect 302460 642370 302560 642470
rect 302684 642370 302784 642470
rect 302908 642370 303008 642470
rect 303132 642370 303232 642470
rect 303356 642370 303456 642470
rect 303580 642370 303680 642470
rect 303804 642370 303904 642470
rect 304028 642370 304128 642470
rect 304252 642370 304352 642470
rect 304476 642370 304576 642470
rect 304700 642370 304800 642470
rect 304924 642370 305024 642470
rect 305148 642370 305248 642470
rect 305372 642370 305472 642470
rect 309346 642370 309446 642470
rect 309570 642370 309670 642470
rect 309794 642370 309894 642470
rect 310018 642370 310118 642470
rect 310242 642370 310342 642470
rect 310466 642370 310566 642470
rect 310690 642370 310790 642470
rect 310914 642370 311014 642470
rect 311138 642370 311238 642470
rect 311362 642370 311462 642470
rect 311586 642370 311686 642470
rect 311810 642370 311910 642470
rect 312034 642370 312134 642470
rect 312258 642370 312358 642470
rect 312482 642370 312582 642470
rect 312706 642370 312806 642470
rect 312930 642370 313030 642470
rect 313154 642370 313254 642470
rect 313378 642370 313478 642470
rect 313602 642370 313702 642470
rect 313826 642370 313926 642470
rect 314050 642370 314150 642470
rect 314274 642370 314374 642470
rect 314498 642370 314598 642470
rect 314722 642370 314822 642470
rect 314946 642370 315046 642470
rect 315170 642370 315270 642470
rect 315394 642370 315494 642470
rect 315618 642370 315718 642470
rect 315842 642370 315942 642470
rect 335616 642390 335716 642490
rect 335840 642390 335940 642490
rect 336064 642390 336164 642490
rect 336288 642390 336388 642490
rect 336512 642390 336612 642490
rect 336736 642390 336836 642490
rect 336960 642390 337060 642490
rect 337184 642390 337284 642490
rect 337408 642390 337508 642490
rect 337632 642390 337732 642490
rect 337856 642390 337956 642490
rect 338080 642390 338180 642490
rect 338304 642390 338404 642490
rect 338528 642390 338628 642490
rect 338752 642390 338852 642490
rect 338976 642390 339076 642490
rect 339200 642390 339300 642490
rect 339424 642390 339524 642490
rect 339648 642390 339748 642490
rect 339872 642390 339972 642490
rect 340096 642390 340196 642490
rect 340320 642390 340420 642490
rect 340544 642390 340644 642490
rect 340768 642390 340868 642490
rect 340992 642390 341092 642490
rect 341216 642390 341316 642490
rect 341440 642390 341540 642490
rect 341664 642390 341764 642490
rect 341888 642390 341988 642490
rect 342112 642390 342212 642490
rect 298876 642146 298976 642246
rect 299100 642146 299200 642246
rect 299324 642146 299424 642246
rect 299548 642146 299648 642246
rect 299772 642146 299872 642246
rect 299996 642146 300096 642246
rect 300220 642146 300320 642246
rect 300444 642146 300544 642246
rect 300668 642146 300768 642246
rect 300892 642146 300992 642246
rect 301116 642146 301216 642246
rect 301340 642146 301440 642246
rect 301564 642146 301664 642246
rect 301788 642146 301888 642246
rect 302012 642146 302112 642246
rect 302236 642146 302336 642246
rect 302460 642146 302560 642246
rect 302684 642146 302784 642246
rect 302908 642146 303008 642246
rect 303132 642146 303232 642246
rect 303356 642146 303456 642246
rect 303580 642146 303680 642246
rect 303804 642146 303904 642246
rect 304028 642146 304128 642246
rect 304252 642146 304352 642246
rect 304476 642146 304576 642246
rect 304700 642146 304800 642246
rect 304924 642146 305024 642246
rect 305148 642146 305248 642246
rect 305372 642146 305472 642246
rect 309346 642146 309446 642246
rect 309570 642146 309670 642246
rect 309794 642146 309894 642246
rect 310018 642146 310118 642246
rect 310242 642146 310342 642246
rect 310466 642146 310566 642246
rect 310690 642146 310790 642246
rect 310914 642146 311014 642246
rect 311138 642146 311238 642246
rect 311362 642146 311462 642246
rect 311586 642146 311686 642246
rect 311810 642146 311910 642246
rect 312034 642146 312134 642246
rect 312258 642146 312358 642246
rect 312482 642146 312582 642246
rect 312706 642146 312806 642246
rect 312930 642146 313030 642246
rect 313154 642146 313254 642246
rect 313378 642146 313478 642246
rect 313602 642146 313702 642246
rect 313826 642146 313926 642246
rect 314050 642146 314150 642246
rect 314274 642146 314374 642246
rect 314498 642146 314598 642246
rect 314722 642146 314822 642246
rect 314946 642146 315046 642246
rect 315170 642146 315270 642246
rect 315394 642146 315494 642246
rect 315618 642146 315718 642246
rect 315842 642146 315942 642246
rect 335616 642166 335716 642266
rect 335840 642166 335940 642266
rect 336064 642166 336164 642266
rect 336288 642166 336388 642266
rect 336512 642166 336612 642266
rect 336736 642166 336836 642266
rect 336960 642166 337060 642266
rect 337184 642166 337284 642266
rect 337408 642166 337508 642266
rect 337632 642166 337732 642266
rect 337856 642166 337956 642266
rect 338080 642166 338180 642266
rect 338304 642166 338404 642266
rect 338528 642166 338628 642266
rect 338752 642166 338852 642266
rect 338976 642166 339076 642266
rect 339200 642166 339300 642266
rect 339424 642166 339524 642266
rect 339648 642166 339748 642266
rect 339872 642166 339972 642266
rect 340096 642166 340196 642266
rect 340320 642166 340420 642266
rect 340544 642166 340644 642266
rect 340768 642166 340868 642266
rect 340992 642166 341092 642266
rect 341216 642166 341316 642266
rect 341440 642166 341540 642266
rect 341664 642166 341764 642266
rect 341888 642166 341988 642266
rect 342112 642166 342212 642266
rect 298876 641922 298976 642022
rect 299100 641922 299200 642022
rect 299324 641922 299424 642022
rect 299548 641922 299648 642022
rect 299772 641922 299872 642022
rect 299996 641922 300096 642022
rect 300220 641922 300320 642022
rect 300444 641922 300544 642022
rect 300668 641922 300768 642022
rect 300892 641922 300992 642022
rect 301116 641922 301216 642022
rect 301340 641922 301440 642022
rect 301564 641922 301664 642022
rect 301788 641922 301888 642022
rect 302012 641922 302112 642022
rect 302236 641922 302336 642022
rect 302460 641922 302560 642022
rect 302684 641922 302784 642022
rect 302908 641922 303008 642022
rect 303132 641922 303232 642022
rect 303356 641922 303456 642022
rect 303580 641922 303680 642022
rect 303804 641922 303904 642022
rect 304028 641922 304128 642022
rect 304252 641922 304352 642022
rect 304476 641922 304576 642022
rect 304700 641922 304800 642022
rect 304924 641922 305024 642022
rect 305148 641922 305248 642022
rect 305372 641922 305472 642022
rect 309346 641922 309446 642022
rect 309570 641922 309670 642022
rect 309794 641922 309894 642022
rect 310018 641922 310118 642022
rect 310242 641922 310342 642022
rect 310466 641922 310566 642022
rect 310690 641922 310790 642022
rect 310914 641922 311014 642022
rect 311138 641922 311238 642022
rect 311362 641922 311462 642022
rect 311586 641922 311686 642022
rect 311810 641922 311910 642022
rect 312034 641922 312134 642022
rect 312258 641922 312358 642022
rect 312482 641922 312582 642022
rect 312706 641922 312806 642022
rect 312930 641922 313030 642022
rect 313154 641922 313254 642022
rect 313378 641922 313478 642022
rect 313602 641922 313702 642022
rect 313826 641922 313926 642022
rect 314050 641922 314150 642022
rect 314274 641922 314374 642022
rect 314498 641922 314598 642022
rect 314722 641922 314822 642022
rect 314946 641922 315046 642022
rect 315170 641922 315270 642022
rect 315394 641922 315494 642022
rect 315618 641922 315718 642022
rect 315842 641922 315942 642022
rect 335616 641942 335716 642042
rect 335840 641942 335940 642042
rect 336064 641942 336164 642042
rect 336288 641942 336388 642042
rect 336512 641942 336612 642042
rect 336736 641942 336836 642042
rect 336960 641942 337060 642042
rect 337184 641942 337284 642042
rect 337408 641942 337508 642042
rect 337632 641942 337732 642042
rect 337856 641942 337956 642042
rect 338080 641942 338180 642042
rect 338304 641942 338404 642042
rect 338528 641942 338628 642042
rect 338752 641942 338852 642042
rect 338976 641942 339076 642042
rect 339200 641942 339300 642042
rect 339424 641942 339524 642042
rect 339648 641942 339748 642042
rect 339872 641942 339972 642042
rect 340096 641942 340196 642042
rect 340320 641942 340420 642042
rect 340544 641942 340644 642042
rect 340768 641942 340868 642042
rect 340992 641942 341092 642042
rect 341216 641942 341316 642042
rect 341440 641942 341540 642042
rect 341664 641942 341764 642042
rect 341888 641942 341988 642042
rect 342112 641942 342212 642042
rect 298876 641698 298976 641798
rect 299100 641698 299200 641798
rect 299324 641698 299424 641798
rect 299548 641698 299648 641798
rect 299772 641698 299872 641798
rect 299996 641698 300096 641798
rect 300220 641698 300320 641798
rect 300444 641698 300544 641798
rect 300668 641698 300768 641798
rect 300892 641698 300992 641798
rect 301116 641698 301216 641798
rect 301340 641698 301440 641798
rect 301564 641698 301664 641798
rect 301788 641698 301888 641798
rect 302012 641698 302112 641798
rect 302236 641698 302336 641798
rect 302460 641698 302560 641798
rect 302684 641698 302784 641798
rect 302908 641698 303008 641798
rect 303132 641698 303232 641798
rect 303356 641698 303456 641798
rect 303580 641698 303680 641798
rect 303804 641698 303904 641798
rect 304028 641698 304128 641798
rect 304252 641698 304352 641798
rect 304476 641698 304576 641798
rect 304700 641698 304800 641798
rect 304924 641698 305024 641798
rect 305148 641698 305248 641798
rect 305372 641698 305472 641798
rect 309346 641698 309446 641798
rect 309570 641698 309670 641798
rect 309794 641698 309894 641798
rect 310018 641698 310118 641798
rect 310242 641698 310342 641798
rect 310466 641698 310566 641798
rect 310690 641698 310790 641798
rect 310914 641698 311014 641798
rect 311138 641698 311238 641798
rect 311362 641698 311462 641798
rect 311586 641698 311686 641798
rect 311810 641698 311910 641798
rect 312034 641698 312134 641798
rect 312258 641698 312358 641798
rect 312482 641698 312582 641798
rect 312706 641698 312806 641798
rect 312930 641698 313030 641798
rect 313154 641698 313254 641798
rect 313378 641698 313478 641798
rect 313602 641698 313702 641798
rect 313826 641698 313926 641798
rect 314050 641698 314150 641798
rect 314274 641698 314374 641798
rect 314498 641698 314598 641798
rect 314722 641698 314822 641798
rect 314946 641698 315046 641798
rect 315170 641698 315270 641798
rect 315394 641698 315494 641798
rect 315618 641698 315718 641798
rect 315842 641698 315942 641798
rect 335616 641718 335716 641818
rect 335840 641718 335940 641818
rect 336064 641718 336164 641818
rect 336288 641718 336388 641818
rect 336512 641718 336612 641818
rect 336736 641718 336836 641818
rect 336960 641718 337060 641818
rect 337184 641718 337284 641818
rect 337408 641718 337508 641818
rect 337632 641718 337732 641818
rect 337856 641718 337956 641818
rect 338080 641718 338180 641818
rect 338304 641718 338404 641818
rect 338528 641718 338628 641818
rect 338752 641718 338852 641818
rect 338976 641718 339076 641818
rect 339200 641718 339300 641818
rect 339424 641718 339524 641818
rect 339648 641718 339748 641818
rect 339872 641718 339972 641818
rect 340096 641718 340196 641818
rect 340320 641718 340420 641818
rect 340544 641718 340644 641818
rect 340768 641718 340868 641818
rect 340992 641718 341092 641818
rect 341216 641718 341316 641818
rect 341440 641718 341540 641818
rect 341664 641718 341764 641818
rect 341888 641718 341988 641818
rect 342112 641718 342212 641818
rect 297850 637896 297872 637996
rect 297872 637896 297950 637996
rect 298074 637896 298174 637996
rect 298298 637896 298398 637996
rect 298522 637896 298622 637996
rect 298746 637896 298846 637996
rect 297850 637672 297872 637772
rect 297872 637672 297950 637772
rect 298074 637672 298174 637772
rect 298298 637672 298398 637772
rect 298522 637672 298622 637772
rect 298746 637672 298846 637772
rect 297850 637448 297872 637548
rect 297872 637448 297950 637548
rect 298074 637448 298174 637548
rect 298298 637448 298398 637548
rect 298522 637448 298622 637548
rect 298746 637448 298846 637548
rect 297850 637224 297872 637324
rect 297872 637224 297950 637324
rect 298074 637224 298174 637324
rect 298298 637224 298398 637324
rect 298522 637224 298622 637324
rect 298746 637224 298846 637324
rect 297850 637000 297872 637100
rect 297872 637000 297950 637100
rect 298074 637000 298174 637100
rect 298298 637000 298398 637100
rect 298522 637000 298622 637100
rect 298746 637000 298846 637100
rect 297850 636776 297872 636876
rect 297872 636776 297950 636876
rect 298074 636776 298174 636876
rect 298298 636776 298398 636876
rect 298522 636776 298622 636876
rect 298746 636776 298846 636876
rect 297850 636552 297872 636652
rect 297872 636552 297950 636652
rect 298074 636552 298174 636652
rect 298298 636552 298398 636652
rect 298522 636552 298622 636652
rect 298746 636552 298846 636652
rect 297850 636328 297872 636428
rect 297872 636328 297950 636428
rect 298074 636328 298174 636428
rect 298298 636328 298398 636428
rect 298522 636328 298622 636428
rect 298746 636328 298846 636428
rect 297850 636104 297872 636204
rect 297872 636104 297950 636204
rect 298074 636104 298174 636204
rect 298298 636104 298398 636204
rect 298522 636104 298622 636204
rect 298746 636104 298846 636204
rect 297850 635880 297872 635980
rect 297872 635880 297950 635980
rect 298074 635880 298174 635980
rect 298298 635880 298398 635980
rect 298522 635880 298622 635980
rect 298746 635880 298846 635980
rect 297850 635656 297872 635756
rect 297872 635656 297950 635756
rect 298074 635656 298174 635756
rect 298298 635656 298398 635756
rect 298522 635656 298622 635756
rect 298746 635656 298846 635756
rect 297850 635432 297872 635532
rect 297872 635432 297950 635532
rect 298074 635432 298174 635532
rect 298298 635432 298398 635532
rect 298522 635432 298622 635532
rect 298746 635432 298846 635532
rect 297850 635208 297872 635308
rect 297872 635208 297950 635308
rect 298074 635208 298174 635308
rect 298298 635208 298398 635308
rect 298522 635208 298622 635308
rect 298746 635208 298846 635308
rect 297850 634984 297872 635084
rect 297872 634984 297950 635084
rect 298074 634984 298174 635084
rect 298298 634984 298398 635084
rect 298522 634984 298622 635084
rect 298746 634984 298846 635084
rect 297850 634760 297872 634860
rect 297872 634760 297950 634860
rect 298074 634760 298174 634860
rect 298298 634760 298398 634860
rect 298522 634760 298622 634860
rect 298746 634760 298846 634860
rect 297850 634536 297872 634636
rect 297872 634536 297950 634636
rect 298074 634536 298174 634636
rect 298298 634536 298398 634636
rect 298522 634536 298622 634636
rect 298746 634536 298846 634636
rect 297850 634312 297872 634412
rect 297872 634312 297950 634412
rect 298074 634312 298174 634412
rect 298298 634312 298398 634412
rect 298522 634312 298622 634412
rect 298746 634312 298846 634412
rect 297850 634088 297872 634188
rect 297872 634088 297950 634188
rect 298074 634088 298174 634188
rect 298298 634088 298398 634188
rect 298522 634088 298622 634188
rect 298746 634088 298846 634188
rect 297850 633864 297872 633964
rect 297872 633864 297950 633964
rect 298074 633864 298174 633964
rect 298298 633864 298398 633964
rect 298522 633864 298622 633964
rect 298746 633864 298846 633964
rect 297850 633640 297872 633740
rect 297872 633640 297950 633740
rect 298074 633640 298174 633740
rect 298298 633640 298398 633740
rect 298522 633640 298622 633740
rect 298746 633640 298846 633740
rect 297850 633416 297872 633516
rect 297872 633416 297950 633516
rect 298074 633416 298174 633516
rect 298298 633416 298398 633516
rect 298522 633416 298622 633516
rect 298746 633416 298846 633516
rect 297850 633192 297872 633292
rect 297872 633192 297950 633292
rect 298074 633192 298174 633292
rect 298298 633192 298398 633292
rect 298522 633192 298622 633292
rect 298746 633192 298846 633292
rect 297850 632968 297872 633068
rect 297872 632968 297950 633068
rect 298074 632968 298174 633068
rect 298298 632968 298398 633068
rect 298522 632968 298622 633068
rect 298746 632968 298846 633068
rect 297850 632744 297872 632844
rect 297872 632744 297950 632844
rect 298074 632744 298174 632844
rect 298298 632744 298398 632844
rect 298522 632744 298622 632844
rect 298746 632744 298846 632844
rect 297850 632520 297872 632620
rect 297872 632520 297950 632620
rect 298074 632520 298174 632620
rect 298298 632520 298398 632620
rect 298522 632520 298622 632620
rect 298746 632520 298846 632620
rect 297850 632296 297872 632396
rect 297872 632296 297950 632396
rect 298074 632296 298174 632396
rect 298298 632296 298398 632396
rect 298522 632296 298622 632396
rect 298746 632296 298846 632396
rect 297850 632072 297872 632172
rect 297872 632072 297950 632172
rect 298074 632072 298174 632172
rect 298298 632072 298398 632172
rect 298522 632072 298622 632172
rect 298746 632072 298846 632172
rect 297850 631848 297872 631948
rect 297872 631848 297950 631948
rect 298074 631848 298174 631948
rect 298298 631848 298398 631948
rect 298522 631848 298622 631948
rect 298746 631848 298846 631948
rect 297850 631624 297872 631724
rect 297872 631624 297950 631724
rect 298074 631624 298174 631724
rect 298298 631624 298398 631724
rect 298522 631624 298622 631724
rect 298746 631624 298846 631724
rect 297850 631400 297872 631500
rect 297872 631400 297950 631500
rect 298074 631400 298174 631500
rect 298298 631400 298398 631500
rect 298522 631400 298622 631500
rect 298746 631400 298846 631500
rect 297850 624496 297872 624596
rect 297872 624496 297950 624596
rect 298074 624496 298174 624596
rect 298298 624496 298398 624596
rect 298522 624496 298622 624596
rect 298746 624496 298846 624596
rect 297850 624272 297872 624372
rect 297872 624272 297950 624372
rect 298074 624272 298174 624372
rect 298298 624272 298398 624372
rect 298522 624272 298622 624372
rect 298746 624272 298846 624372
rect 297850 624048 297872 624148
rect 297872 624048 297950 624148
rect 298074 624048 298174 624148
rect 298298 624048 298398 624148
rect 298522 624048 298622 624148
rect 298746 624048 298846 624148
rect 297850 623824 297872 623924
rect 297872 623824 297950 623924
rect 298074 623824 298174 623924
rect 298298 623824 298398 623924
rect 298522 623824 298622 623924
rect 298746 623824 298846 623924
rect 297850 623600 297872 623700
rect 297872 623600 297950 623700
rect 298074 623600 298174 623700
rect 298298 623600 298398 623700
rect 298522 623600 298622 623700
rect 298746 623600 298846 623700
rect 297850 623376 297872 623476
rect 297872 623376 297950 623476
rect 298074 623376 298174 623476
rect 298298 623376 298398 623476
rect 298522 623376 298622 623476
rect 298746 623376 298846 623476
rect 297850 623152 297872 623252
rect 297872 623152 297950 623252
rect 298074 623152 298174 623252
rect 298298 623152 298398 623252
rect 298522 623152 298622 623252
rect 298746 623152 298846 623252
rect 297850 622928 297872 623028
rect 297872 622928 297950 623028
rect 298074 622928 298174 623028
rect 298298 622928 298398 623028
rect 298522 622928 298622 623028
rect 298746 622928 298846 623028
rect 297850 622704 297872 622804
rect 297872 622704 297950 622804
rect 298074 622704 298174 622804
rect 298298 622704 298398 622804
rect 298522 622704 298622 622804
rect 298746 622704 298846 622804
rect 297850 622480 297872 622580
rect 297872 622480 297950 622580
rect 298074 622480 298174 622580
rect 298298 622480 298398 622580
rect 298522 622480 298622 622580
rect 298746 622480 298846 622580
rect 297850 622256 297872 622356
rect 297872 622256 297950 622356
rect 298074 622256 298174 622356
rect 298298 622256 298398 622356
rect 298522 622256 298622 622356
rect 298746 622256 298846 622356
rect 297850 622032 297872 622132
rect 297872 622032 297950 622132
rect 298074 622032 298174 622132
rect 298298 622032 298398 622132
rect 298522 622032 298622 622132
rect 298746 622032 298846 622132
rect 297850 621808 297872 621908
rect 297872 621808 297950 621908
rect 298074 621808 298174 621908
rect 298298 621808 298398 621908
rect 298522 621808 298622 621908
rect 298746 621808 298846 621908
rect 297850 621584 297872 621684
rect 297872 621584 297950 621684
rect 298074 621584 298174 621684
rect 298298 621584 298398 621684
rect 298522 621584 298622 621684
rect 298746 621584 298846 621684
rect 297850 621360 297872 621460
rect 297872 621360 297950 621460
rect 298074 621360 298174 621460
rect 298298 621360 298398 621460
rect 298522 621360 298622 621460
rect 298746 621360 298846 621460
rect 297850 621136 297872 621236
rect 297872 621136 297950 621236
rect 298074 621136 298174 621236
rect 298298 621136 298398 621236
rect 298522 621136 298622 621236
rect 298746 621136 298846 621236
rect 297850 620912 297872 621012
rect 297872 620912 297950 621012
rect 298074 620912 298174 621012
rect 298298 620912 298398 621012
rect 298522 620912 298622 621012
rect 298746 620912 298846 621012
rect 297850 620688 297872 620788
rect 297872 620688 297950 620788
rect 298074 620688 298174 620788
rect 298298 620688 298398 620788
rect 298522 620688 298622 620788
rect 298746 620688 298846 620788
rect 297850 620464 297872 620564
rect 297872 620464 297950 620564
rect 298074 620464 298174 620564
rect 298298 620464 298398 620564
rect 298522 620464 298622 620564
rect 298746 620464 298846 620564
rect 297850 620240 297872 620340
rect 297872 620240 297950 620340
rect 298074 620240 298174 620340
rect 298298 620240 298398 620340
rect 298522 620240 298622 620340
rect 298746 620240 298846 620340
rect 297850 620016 297872 620116
rect 297872 620016 297950 620116
rect 298074 620016 298174 620116
rect 298298 620016 298398 620116
rect 298522 620016 298622 620116
rect 298746 620016 298846 620116
rect 297850 619792 297872 619892
rect 297872 619792 297950 619892
rect 298074 619792 298174 619892
rect 298298 619792 298398 619892
rect 298522 619792 298622 619892
rect 298746 619792 298846 619892
rect 297850 619568 297872 619668
rect 297872 619568 297950 619668
rect 298074 619568 298174 619668
rect 298298 619568 298398 619668
rect 298522 619568 298622 619668
rect 298746 619568 298846 619668
rect 297850 619344 297872 619444
rect 297872 619344 297950 619444
rect 298074 619344 298174 619444
rect 298298 619344 298398 619444
rect 298522 619344 298622 619444
rect 298746 619344 298846 619444
rect 297850 619120 297872 619220
rect 297872 619120 297950 619220
rect 298074 619120 298174 619220
rect 298298 619120 298398 619220
rect 298522 619120 298622 619220
rect 298746 619120 298846 619220
rect 297850 618896 297872 618996
rect 297872 618896 297950 618996
rect 298074 618896 298174 618996
rect 298298 618896 298398 618996
rect 298522 618896 298622 618996
rect 298746 618896 298846 618996
rect 297850 618672 297872 618772
rect 297872 618672 297950 618772
rect 298074 618672 298174 618772
rect 298298 618672 298398 618772
rect 298522 618672 298622 618772
rect 298746 618672 298846 618772
rect 297850 618448 297872 618548
rect 297872 618448 297950 618548
rect 298074 618448 298174 618548
rect 298298 618448 298398 618548
rect 298522 618448 298622 618548
rect 298746 618448 298846 618548
rect 297850 618224 297872 618324
rect 297872 618224 297950 618324
rect 298074 618224 298174 618324
rect 298298 618224 298398 618324
rect 298522 618224 298622 618324
rect 298746 618224 298846 618324
rect 297850 618000 297872 618100
rect 297872 618000 297950 618100
rect 298074 618000 298174 618100
rect 298298 618000 298398 618100
rect 298522 618000 298622 618100
rect 298746 618000 298846 618100
rect 300672 640542 311888 640558
rect 300672 639776 300688 640542
rect 300688 639776 311872 640542
rect 311872 639776 311888 640542
rect 300672 639760 311888 639776
rect 316560 637085 317098 637482
rect 317378 637085 317916 637482
rect 318196 637085 318734 637482
rect 319014 637085 319552 637482
rect 321468 637023 322006 637420
rect 322286 637023 322824 637420
rect 323104 637023 323642 637420
rect 323922 637023 324460 637420
rect 324740 637023 325278 637420
rect 325558 637023 326096 637420
rect 326376 637023 326914 637420
rect 327194 637023 327732 637420
rect 328012 637023 328550 637420
rect 328830 637023 329368 637420
rect 329648 637023 330186 637420
rect 330466 637023 331004 637420
rect 331284 637023 331822 637420
rect 332102 637023 332640 637420
rect 332920 637023 333458 637420
rect 333738 637023 334276 637420
rect 334556 637023 335094 637420
rect 313288 635699 313826 636096
rect 314106 635699 314644 636096
rect 314924 635699 315462 636096
rect 313288 631944 313826 632341
rect 314106 631944 314644 632341
rect 314924 631944 315462 632341
rect 315744 631674 316238 632740
rect 316560 632354 317098 632751
rect 317378 632354 317916 632751
rect 318196 632354 318734 632751
rect 319014 632354 319552 632751
rect 320696 631686 321208 632738
rect 321468 630288 322006 630685
rect 322286 630287 322824 630685
rect 323104 630288 323642 630685
rect 323922 630288 324460 630685
rect 324740 630287 325278 630685
rect 325558 630288 326096 630685
rect 326376 630288 326914 630685
rect 327194 630287 327732 630685
rect 328012 630288 328550 630685
rect 328830 630288 329368 630685
rect 329648 630288 330186 630685
rect 330466 630287 331004 630685
rect 331284 630288 331822 630685
rect 332102 630288 332640 630685
rect 332920 630288 333458 630685
rect 333738 630288 334276 630685
rect 334556 630288 335094 630685
rect 335032 627348 335038 627370
rect 335038 627348 335066 627370
rect 335032 627336 335066 627348
rect 335132 627336 335166 627370
rect 335232 627336 335266 627370
rect 335332 627348 335364 627370
rect 335364 627348 335366 627370
rect 335432 627348 335454 627370
rect 335454 627348 335466 627370
rect 335532 627348 335544 627370
rect 335544 627348 335566 627370
rect 335332 627336 335366 627348
rect 335432 627336 335466 627348
rect 335532 627336 335566 627348
rect 335032 627258 335038 627270
rect 335038 627258 335066 627270
rect 335032 627236 335066 627258
rect 335132 627236 335166 627270
rect 335232 627236 335266 627270
rect 335332 627258 335364 627270
rect 335364 627258 335366 627270
rect 335432 627258 335454 627270
rect 335454 627258 335466 627270
rect 335532 627258 335544 627270
rect 335544 627258 335566 627270
rect 335332 627236 335366 627258
rect 335432 627236 335466 627258
rect 335532 627236 335566 627258
rect 335032 627168 335038 627170
rect 335038 627168 335066 627170
rect 335032 627136 335066 627168
rect 335132 627136 335166 627170
rect 335232 627136 335266 627170
rect 335332 627168 335364 627170
rect 335364 627168 335366 627170
rect 335432 627168 335454 627170
rect 335454 627168 335466 627170
rect 335532 627168 335544 627170
rect 335544 627168 335566 627170
rect 335332 627136 335366 627168
rect 335432 627136 335466 627168
rect 335532 627136 335566 627168
rect 335032 627036 335066 627070
rect 335132 627036 335166 627070
rect 335232 627036 335266 627070
rect 335332 627036 335366 627070
rect 335432 627036 335466 627070
rect 335532 627036 335566 627070
rect 335032 626936 335066 626970
rect 335132 626936 335166 626970
rect 335232 626936 335266 626970
rect 335332 626936 335366 626970
rect 335432 626936 335466 626970
rect 335532 626936 335566 626970
rect 335032 626842 335066 626870
rect 335032 626836 335038 626842
rect 335038 626836 335066 626842
rect 335132 626836 335166 626870
rect 335232 626836 335266 626870
rect 335332 626842 335366 626870
rect 335432 626842 335466 626870
rect 335532 626842 335566 626870
rect 335332 626836 335364 626842
rect 335364 626836 335366 626842
rect 335432 626836 335454 626842
rect 335454 626836 335466 626842
rect 335532 626836 335544 626842
rect 335544 626836 335566 626842
rect 336320 627348 336326 627370
rect 336326 627348 336354 627370
rect 336320 627336 336354 627348
rect 336420 627336 336454 627370
rect 336520 627336 336554 627370
rect 336620 627348 336652 627370
rect 336652 627348 336654 627370
rect 336720 627348 336742 627370
rect 336742 627348 336754 627370
rect 336820 627348 336832 627370
rect 336832 627348 336854 627370
rect 336620 627336 336654 627348
rect 336720 627336 336754 627348
rect 336820 627336 336854 627348
rect 336320 627258 336326 627270
rect 336326 627258 336354 627270
rect 336320 627236 336354 627258
rect 336420 627236 336454 627270
rect 336520 627236 336554 627270
rect 336620 627258 336652 627270
rect 336652 627258 336654 627270
rect 336720 627258 336742 627270
rect 336742 627258 336754 627270
rect 336820 627258 336832 627270
rect 336832 627258 336854 627270
rect 336620 627236 336654 627258
rect 336720 627236 336754 627258
rect 336820 627236 336854 627258
rect 336320 627168 336326 627170
rect 336326 627168 336354 627170
rect 336320 627136 336354 627168
rect 336420 627136 336454 627170
rect 336520 627136 336554 627170
rect 336620 627168 336652 627170
rect 336652 627168 336654 627170
rect 336720 627168 336742 627170
rect 336742 627168 336754 627170
rect 336820 627168 336832 627170
rect 336832 627168 336854 627170
rect 336620 627136 336654 627168
rect 336720 627136 336754 627168
rect 336820 627136 336854 627168
rect 336320 627036 336354 627070
rect 336420 627036 336454 627070
rect 336520 627036 336554 627070
rect 336620 627036 336654 627070
rect 336720 627036 336754 627070
rect 336820 627036 336854 627070
rect 336320 626936 336354 626970
rect 336420 626936 336454 626970
rect 336520 626936 336554 626970
rect 336620 626936 336654 626970
rect 336720 626936 336754 626970
rect 336820 626936 336854 626970
rect 336320 626842 336354 626870
rect 336320 626836 336326 626842
rect 336326 626836 336354 626842
rect 336420 626836 336454 626870
rect 336520 626836 336554 626870
rect 336620 626842 336654 626870
rect 336720 626842 336754 626870
rect 336820 626842 336854 626870
rect 336620 626836 336652 626842
rect 336652 626836 336654 626842
rect 336720 626836 336742 626842
rect 336742 626836 336754 626842
rect 336820 626836 336832 626842
rect 336832 626836 336854 626842
rect 337608 627348 337614 627370
rect 337614 627348 337642 627370
rect 337608 627336 337642 627348
rect 337708 627336 337742 627370
rect 337808 627336 337842 627370
rect 337908 627348 337940 627370
rect 337940 627348 337942 627370
rect 338008 627348 338030 627370
rect 338030 627348 338042 627370
rect 338108 627348 338120 627370
rect 338120 627348 338142 627370
rect 337908 627336 337942 627348
rect 338008 627336 338042 627348
rect 338108 627336 338142 627348
rect 337608 627258 337614 627270
rect 337614 627258 337642 627270
rect 337608 627236 337642 627258
rect 337708 627236 337742 627270
rect 337808 627236 337842 627270
rect 337908 627258 337940 627270
rect 337940 627258 337942 627270
rect 338008 627258 338030 627270
rect 338030 627258 338042 627270
rect 338108 627258 338120 627270
rect 338120 627258 338142 627270
rect 337908 627236 337942 627258
rect 338008 627236 338042 627258
rect 338108 627236 338142 627258
rect 337608 627168 337614 627170
rect 337614 627168 337642 627170
rect 337608 627136 337642 627168
rect 337708 627136 337742 627170
rect 337808 627136 337842 627170
rect 337908 627168 337940 627170
rect 337940 627168 337942 627170
rect 338008 627168 338030 627170
rect 338030 627168 338042 627170
rect 338108 627168 338120 627170
rect 338120 627168 338142 627170
rect 337908 627136 337942 627168
rect 338008 627136 338042 627168
rect 338108 627136 338142 627168
rect 337608 627036 337642 627070
rect 337708 627036 337742 627070
rect 337808 627036 337842 627070
rect 337908 627036 337942 627070
rect 338008 627036 338042 627070
rect 338108 627036 338142 627070
rect 337608 626936 337642 626970
rect 337708 626936 337742 626970
rect 337808 626936 337842 626970
rect 337908 626936 337942 626970
rect 338008 626936 338042 626970
rect 338108 626936 338142 626970
rect 337608 626842 337642 626870
rect 337608 626836 337614 626842
rect 337614 626836 337642 626842
rect 337708 626836 337742 626870
rect 337808 626836 337842 626870
rect 337908 626842 337942 626870
rect 338008 626842 338042 626870
rect 338108 626842 338142 626870
rect 337908 626836 337940 626842
rect 337940 626836 337942 626842
rect 338008 626836 338030 626842
rect 338030 626836 338042 626842
rect 338108 626836 338120 626842
rect 338120 626836 338142 626842
rect 338896 627348 338902 627370
rect 338902 627348 338930 627370
rect 338896 627336 338930 627348
rect 338996 627336 339030 627370
rect 339096 627336 339130 627370
rect 339196 627348 339228 627370
rect 339228 627348 339230 627370
rect 339296 627348 339318 627370
rect 339318 627348 339330 627370
rect 339396 627348 339408 627370
rect 339408 627348 339430 627370
rect 339196 627336 339230 627348
rect 339296 627336 339330 627348
rect 339396 627336 339430 627348
rect 338896 627258 338902 627270
rect 338902 627258 338930 627270
rect 338896 627236 338930 627258
rect 338996 627236 339030 627270
rect 339096 627236 339130 627270
rect 339196 627258 339228 627270
rect 339228 627258 339230 627270
rect 339296 627258 339318 627270
rect 339318 627258 339330 627270
rect 339396 627258 339408 627270
rect 339408 627258 339430 627270
rect 339196 627236 339230 627258
rect 339296 627236 339330 627258
rect 339396 627236 339430 627258
rect 338896 627168 338902 627170
rect 338902 627168 338930 627170
rect 338896 627136 338930 627168
rect 338996 627136 339030 627170
rect 339096 627136 339130 627170
rect 339196 627168 339228 627170
rect 339228 627168 339230 627170
rect 339296 627168 339318 627170
rect 339318 627168 339330 627170
rect 339396 627168 339408 627170
rect 339408 627168 339430 627170
rect 339196 627136 339230 627168
rect 339296 627136 339330 627168
rect 339396 627136 339430 627168
rect 338896 627036 338930 627070
rect 338996 627036 339030 627070
rect 339096 627036 339130 627070
rect 339196 627036 339230 627070
rect 339296 627036 339330 627070
rect 339396 627036 339430 627070
rect 338896 626936 338930 626970
rect 338996 626936 339030 626970
rect 339096 626936 339130 626970
rect 339196 626936 339230 626970
rect 339296 626936 339330 626970
rect 339396 626936 339430 626970
rect 338896 626842 338930 626870
rect 338896 626836 338902 626842
rect 338902 626836 338930 626842
rect 338996 626836 339030 626870
rect 339096 626836 339130 626870
rect 339196 626842 339230 626870
rect 339296 626842 339330 626870
rect 339396 626842 339430 626870
rect 339196 626836 339228 626842
rect 339228 626836 339230 626842
rect 339296 626836 339318 626842
rect 339318 626836 339330 626842
rect 339396 626836 339408 626842
rect 339408 626836 339430 626842
rect 340184 627348 340190 627370
rect 340190 627348 340218 627370
rect 340184 627336 340218 627348
rect 340284 627336 340318 627370
rect 340384 627336 340418 627370
rect 340484 627348 340516 627370
rect 340516 627348 340518 627370
rect 340584 627348 340606 627370
rect 340606 627348 340618 627370
rect 340684 627348 340696 627370
rect 340696 627348 340718 627370
rect 340484 627336 340518 627348
rect 340584 627336 340618 627348
rect 340684 627336 340718 627348
rect 340184 627258 340190 627270
rect 340190 627258 340218 627270
rect 340184 627236 340218 627258
rect 340284 627236 340318 627270
rect 340384 627236 340418 627270
rect 340484 627258 340516 627270
rect 340516 627258 340518 627270
rect 340584 627258 340606 627270
rect 340606 627258 340618 627270
rect 340684 627258 340696 627270
rect 340696 627258 340718 627270
rect 340484 627236 340518 627258
rect 340584 627236 340618 627258
rect 340684 627236 340718 627258
rect 340184 627168 340190 627170
rect 340190 627168 340218 627170
rect 340184 627136 340218 627168
rect 340284 627136 340318 627170
rect 340384 627136 340418 627170
rect 340484 627168 340516 627170
rect 340516 627168 340518 627170
rect 340584 627168 340606 627170
rect 340606 627168 340618 627170
rect 340684 627168 340696 627170
rect 340696 627168 340718 627170
rect 340484 627136 340518 627168
rect 340584 627136 340618 627168
rect 340684 627136 340718 627168
rect 340184 627036 340218 627070
rect 340284 627036 340318 627070
rect 340384 627036 340418 627070
rect 340484 627036 340518 627070
rect 340584 627036 340618 627070
rect 340684 627036 340718 627070
rect 340184 626936 340218 626970
rect 340284 626936 340318 626970
rect 340384 626936 340418 626970
rect 340484 626936 340518 626970
rect 340584 626936 340618 626970
rect 340684 626936 340718 626970
rect 340184 626842 340218 626870
rect 340184 626836 340190 626842
rect 340190 626836 340218 626842
rect 340284 626836 340318 626870
rect 340384 626836 340418 626870
rect 340484 626842 340518 626870
rect 340584 626842 340618 626870
rect 340684 626842 340718 626870
rect 340484 626836 340516 626842
rect 340516 626836 340518 626842
rect 340584 626836 340606 626842
rect 340606 626836 340618 626842
rect 340684 626836 340696 626842
rect 340696 626836 340718 626842
rect 335032 626060 335038 626082
rect 335038 626060 335066 626082
rect 335032 626048 335066 626060
rect 335132 626048 335166 626082
rect 335232 626048 335266 626082
rect 335332 626060 335364 626082
rect 335364 626060 335366 626082
rect 335432 626060 335454 626082
rect 335454 626060 335466 626082
rect 335532 626060 335544 626082
rect 335544 626060 335566 626082
rect 335332 626048 335366 626060
rect 335432 626048 335466 626060
rect 335532 626048 335566 626060
rect 335032 625970 335038 625982
rect 335038 625970 335066 625982
rect 335032 625948 335066 625970
rect 335132 625948 335166 625982
rect 335232 625948 335266 625982
rect 335332 625970 335364 625982
rect 335364 625970 335366 625982
rect 335432 625970 335454 625982
rect 335454 625970 335466 625982
rect 335532 625970 335544 625982
rect 335544 625970 335566 625982
rect 335332 625948 335366 625970
rect 335432 625948 335466 625970
rect 335532 625948 335566 625970
rect 335032 625880 335038 625882
rect 335038 625880 335066 625882
rect 335032 625848 335066 625880
rect 335132 625848 335166 625882
rect 335232 625848 335266 625882
rect 335332 625880 335364 625882
rect 335364 625880 335366 625882
rect 335432 625880 335454 625882
rect 335454 625880 335466 625882
rect 335532 625880 335544 625882
rect 335544 625880 335566 625882
rect 335332 625848 335366 625880
rect 335432 625848 335466 625880
rect 335532 625848 335566 625880
rect 335032 625748 335066 625782
rect 335132 625748 335166 625782
rect 335232 625748 335266 625782
rect 335332 625748 335366 625782
rect 335432 625748 335466 625782
rect 335532 625748 335566 625782
rect 335032 625648 335066 625682
rect 335132 625648 335166 625682
rect 335232 625648 335266 625682
rect 335332 625648 335366 625682
rect 335432 625648 335466 625682
rect 335532 625648 335566 625682
rect 335032 625554 335066 625582
rect 335032 625548 335038 625554
rect 335038 625548 335066 625554
rect 335132 625548 335166 625582
rect 335232 625548 335266 625582
rect 335332 625554 335366 625582
rect 335432 625554 335466 625582
rect 335532 625554 335566 625582
rect 335332 625548 335364 625554
rect 335364 625548 335366 625554
rect 335432 625548 335454 625554
rect 335454 625548 335466 625554
rect 335532 625548 335544 625554
rect 335544 625548 335566 625554
rect 336320 626060 336326 626082
rect 336326 626060 336354 626082
rect 336320 626048 336354 626060
rect 336420 626048 336454 626082
rect 336520 626048 336554 626082
rect 336620 626060 336652 626082
rect 336652 626060 336654 626082
rect 336720 626060 336742 626082
rect 336742 626060 336754 626082
rect 336820 626060 336832 626082
rect 336832 626060 336854 626082
rect 336620 626048 336654 626060
rect 336720 626048 336754 626060
rect 336820 626048 336854 626060
rect 336320 625970 336326 625982
rect 336326 625970 336354 625982
rect 336320 625948 336354 625970
rect 336420 625948 336454 625982
rect 336520 625948 336554 625982
rect 336620 625970 336652 625982
rect 336652 625970 336654 625982
rect 336720 625970 336742 625982
rect 336742 625970 336754 625982
rect 336820 625970 336832 625982
rect 336832 625970 336854 625982
rect 336620 625948 336654 625970
rect 336720 625948 336754 625970
rect 336820 625948 336854 625970
rect 336320 625880 336326 625882
rect 336326 625880 336354 625882
rect 336320 625848 336354 625880
rect 336420 625848 336454 625882
rect 336520 625848 336554 625882
rect 336620 625880 336652 625882
rect 336652 625880 336654 625882
rect 336720 625880 336742 625882
rect 336742 625880 336754 625882
rect 336820 625880 336832 625882
rect 336832 625880 336854 625882
rect 336620 625848 336654 625880
rect 336720 625848 336754 625880
rect 336820 625848 336854 625880
rect 336320 625748 336354 625782
rect 336420 625748 336454 625782
rect 336520 625748 336554 625782
rect 336620 625748 336654 625782
rect 336720 625748 336754 625782
rect 336820 625748 336854 625782
rect 336320 625648 336354 625682
rect 336420 625648 336454 625682
rect 336520 625648 336554 625682
rect 336620 625648 336654 625682
rect 336720 625648 336754 625682
rect 336820 625648 336854 625682
rect 336320 625554 336354 625582
rect 336320 625548 336326 625554
rect 336326 625548 336354 625554
rect 336420 625548 336454 625582
rect 336520 625548 336554 625582
rect 336620 625554 336654 625582
rect 336720 625554 336754 625582
rect 336820 625554 336854 625582
rect 336620 625548 336652 625554
rect 336652 625548 336654 625554
rect 336720 625548 336742 625554
rect 336742 625548 336754 625554
rect 336820 625548 336832 625554
rect 336832 625548 336854 625554
rect 337608 626060 337614 626082
rect 337614 626060 337642 626082
rect 337608 626048 337642 626060
rect 337708 626048 337742 626082
rect 337808 626048 337842 626082
rect 337908 626060 337940 626082
rect 337940 626060 337942 626082
rect 338008 626060 338030 626082
rect 338030 626060 338042 626082
rect 338108 626060 338120 626082
rect 338120 626060 338142 626082
rect 337908 626048 337942 626060
rect 338008 626048 338042 626060
rect 338108 626048 338142 626060
rect 337608 625970 337614 625982
rect 337614 625970 337642 625982
rect 337608 625948 337642 625970
rect 337708 625948 337742 625982
rect 337808 625948 337842 625982
rect 337908 625970 337940 625982
rect 337940 625970 337942 625982
rect 338008 625970 338030 625982
rect 338030 625970 338042 625982
rect 338108 625970 338120 625982
rect 338120 625970 338142 625982
rect 337908 625948 337942 625970
rect 338008 625948 338042 625970
rect 338108 625948 338142 625970
rect 337608 625880 337614 625882
rect 337614 625880 337642 625882
rect 337608 625848 337642 625880
rect 337708 625848 337742 625882
rect 337808 625848 337842 625882
rect 337908 625880 337940 625882
rect 337940 625880 337942 625882
rect 338008 625880 338030 625882
rect 338030 625880 338042 625882
rect 338108 625880 338120 625882
rect 338120 625880 338142 625882
rect 337908 625848 337942 625880
rect 338008 625848 338042 625880
rect 338108 625848 338142 625880
rect 337608 625748 337642 625782
rect 337708 625748 337742 625782
rect 337808 625748 337842 625782
rect 337908 625748 337942 625782
rect 338008 625748 338042 625782
rect 338108 625748 338142 625782
rect 337608 625648 337642 625682
rect 337708 625648 337742 625682
rect 337808 625648 337842 625682
rect 337908 625648 337942 625682
rect 338008 625648 338042 625682
rect 338108 625648 338142 625682
rect 337608 625554 337642 625582
rect 337608 625548 337614 625554
rect 337614 625548 337642 625554
rect 337708 625548 337742 625582
rect 337808 625548 337842 625582
rect 337908 625554 337942 625582
rect 338008 625554 338042 625582
rect 338108 625554 338142 625582
rect 337908 625548 337940 625554
rect 337940 625548 337942 625554
rect 338008 625548 338030 625554
rect 338030 625548 338042 625554
rect 338108 625548 338120 625554
rect 338120 625548 338142 625554
rect 338896 626060 338902 626082
rect 338902 626060 338930 626082
rect 338896 626048 338930 626060
rect 338996 626048 339030 626082
rect 339096 626048 339130 626082
rect 339196 626060 339228 626082
rect 339228 626060 339230 626082
rect 339296 626060 339318 626082
rect 339318 626060 339330 626082
rect 339396 626060 339408 626082
rect 339408 626060 339430 626082
rect 339196 626048 339230 626060
rect 339296 626048 339330 626060
rect 339396 626048 339430 626060
rect 338896 625970 338902 625982
rect 338902 625970 338930 625982
rect 338896 625948 338930 625970
rect 338996 625948 339030 625982
rect 339096 625948 339130 625982
rect 339196 625970 339228 625982
rect 339228 625970 339230 625982
rect 339296 625970 339318 625982
rect 339318 625970 339330 625982
rect 339396 625970 339408 625982
rect 339408 625970 339430 625982
rect 339196 625948 339230 625970
rect 339296 625948 339330 625970
rect 339396 625948 339430 625970
rect 338896 625880 338902 625882
rect 338902 625880 338930 625882
rect 338896 625848 338930 625880
rect 338996 625848 339030 625882
rect 339096 625848 339130 625882
rect 339196 625880 339228 625882
rect 339228 625880 339230 625882
rect 339296 625880 339318 625882
rect 339318 625880 339330 625882
rect 339396 625880 339408 625882
rect 339408 625880 339430 625882
rect 339196 625848 339230 625880
rect 339296 625848 339330 625880
rect 339396 625848 339430 625880
rect 338896 625748 338930 625782
rect 338996 625748 339030 625782
rect 339096 625748 339130 625782
rect 339196 625748 339230 625782
rect 339296 625748 339330 625782
rect 339396 625748 339430 625782
rect 338896 625648 338930 625682
rect 338996 625648 339030 625682
rect 339096 625648 339130 625682
rect 339196 625648 339230 625682
rect 339296 625648 339330 625682
rect 339396 625648 339430 625682
rect 338896 625554 338930 625582
rect 338896 625548 338902 625554
rect 338902 625548 338930 625554
rect 338996 625548 339030 625582
rect 339096 625548 339130 625582
rect 339196 625554 339230 625582
rect 339296 625554 339330 625582
rect 339396 625554 339430 625582
rect 339196 625548 339228 625554
rect 339228 625548 339230 625554
rect 339296 625548 339318 625554
rect 339318 625548 339330 625554
rect 339396 625548 339408 625554
rect 339408 625548 339430 625554
rect 340184 626060 340190 626082
rect 340190 626060 340218 626082
rect 340184 626048 340218 626060
rect 340284 626048 340318 626082
rect 340384 626048 340418 626082
rect 340484 626060 340516 626082
rect 340516 626060 340518 626082
rect 340584 626060 340606 626082
rect 340606 626060 340618 626082
rect 340684 626060 340696 626082
rect 340696 626060 340718 626082
rect 340484 626048 340518 626060
rect 340584 626048 340618 626060
rect 340684 626048 340718 626060
rect 340184 625970 340190 625982
rect 340190 625970 340218 625982
rect 340184 625948 340218 625970
rect 340284 625948 340318 625982
rect 340384 625948 340418 625982
rect 340484 625970 340516 625982
rect 340516 625970 340518 625982
rect 340584 625970 340606 625982
rect 340606 625970 340618 625982
rect 340684 625970 340696 625982
rect 340696 625970 340718 625982
rect 340484 625948 340518 625970
rect 340584 625948 340618 625970
rect 340684 625948 340718 625970
rect 340184 625880 340190 625882
rect 340190 625880 340218 625882
rect 340184 625848 340218 625880
rect 340284 625848 340318 625882
rect 340384 625848 340418 625882
rect 340484 625880 340516 625882
rect 340516 625880 340518 625882
rect 340584 625880 340606 625882
rect 340606 625880 340618 625882
rect 340684 625880 340696 625882
rect 340696 625880 340718 625882
rect 340484 625848 340518 625880
rect 340584 625848 340618 625880
rect 340684 625848 340718 625880
rect 340184 625748 340218 625782
rect 340284 625748 340318 625782
rect 340384 625748 340418 625782
rect 340484 625748 340518 625782
rect 340584 625748 340618 625782
rect 340684 625748 340718 625782
rect 340184 625648 340218 625682
rect 340284 625648 340318 625682
rect 340384 625648 340418 625682
rect 340484 625648 340518 625682
rect 340584 625648 340618 625682
rect 340684 625648 340718 625682
rect 340184 625554 340218 625582
rect 340184 625548 340190 625554
rect 340190 625548 340218 625554
rect 340284 625548 340318 625582
rect 340384 625548 340418 625582
rect 340484 625554 340518 625582
rect 340584 625554 340618 625582
rect 340684 625554 340718 625582
rect 340484 625548 340516 625554
rect 340516 625548 340518 625554
rect 340584 625548 340606 625554
rect 340606 625548 340618 625554
rect 340684 625548 340696 625554
rect 340696 625548 340718 625554
rect 304316 624888 310780 624894
rect 304316 624556 304322 624888
rect 304322 624556 310774 624888
rect 310774 624556 310780 624888
rect 304316 624550 310780 624556
rect 305040 624324 310416 624358
rect 304956 624020 304990 624204
rect 305040 623866 310416 623900
rect 305476 622198 305660 622232
rect 306048 622198 306232 622232
rect 306620 622198 306804 622232
rect 307192 622198 307376 622232
rect 307764 622198 307948 622232
rect 308336 622198 308520 622232
rect 308908 622198 309092 622232
rect 309480 622198 309664 622232
rect 301298 621174 301350 621226
rect 302214 621174 302266 621226
rect 300546 621076 300730 621110
rect 301004 621076 301188 621110
rect 301462 621076 301646 621110
rect 301920 621076 302104 621110
rect 302378 621076 302562 621110
rect 302836 621076 303020 621110
rect 300392 620650 300426 621026
rect 300850 620650 300884 621026
rect 301308 620650 301342 621026
rect 301766 620650 301800 621026
rect 302224 620650 302258 621026
rect 302682 620650 302716 621026
rect 303140 620650 303174 621026
rect 304770 620550 304870 622148
rect 305322 620372 305356 622148
rect 305780 620372 305814 622148
rect 305894 620372 305928 622148
rect 306352 620372 306386 622148
rect 306466 620372 306500 622148
rect 306924 620372 306958 622148
rect 307038 620372 307072 622148
rect 307496 620372 307530 622148
rect 307610 620372 307644 622148
rect 308068 620372 308102 622148
rect 308182 620372 308216 622148
rect 308640 620372 308674 622148
rect 308754 620372 308788 622148
rect 309212 620372 309246 622148
rect 309326 620372 309360 622148
rect 309784 620372 309818 622148
rect 310270 620550 310370 622148
rect 303750 619795 303934 619829
rect 304322 619795 304506 619829
rect 304894 619795 305078 619829
rect 305466 619795 305650 619829
rect 306038 619795 306222 619829
rect 306610 619795 306794 619829
rect 307182 619795 307366 619829
rect 307754 619795 307938 619829
rect 308326 619795 308510 619829
rect 308898 619795 309082 619829
rect 309470 619795 309654 619829
rect 310042 619795 310226 619829
rect 310614 619795 310798 619829
rect 311186 619795 311370 619829
rect 302954 617306 303054 619648
rect 303596 617180 303630 619736
rect 304054 617180 304088 619736
rect 304168 617180 304202 619736
rect 304626 617180 304660 619736
rect 304740 617180 304774 619736
rect 305198 617180 305232 619736
rect 305312 617180 305346 619736
rect 305770 617180 305804 619736
rect 305884 617180 305918 619736
rect 306342 617180 306376 619736
rect 306456 617180 306490 619736
rect 306914 617180 306948 619736
rect 307028 617180 307062 619736
rect 307486 617180 307520 619736
rect 307600 617180 307634 619736
rect 308058 617180 308092 619736
rect 308172 617180 308206 619736
rect 308630 617180 308664 619736
rect 308744 617180 308778 619736
rect 309202 617180 309236 619736
rect 309316 617180 309350 619736
rect 309774 617180 309808 619736
rect 309888 617180 309922 619736
rect 310346 617180 310380 619736
rect 310460 617180 310494 619736
rect 310918 617180 310952 619736
rect 311032 617180 311066 619736
rect 311490 617180 311524 619736
rect 312082 617306 312182 619648
rect 306536 616702 308878 616802
rect 313404 617218 313438 624934
rect 313862 617218 313896 624934
rect 314320 617218 314354 624934
rect 314778 617218 314812 624934
rect 315236 617218 315270 624934
rect 315694 617218 315728 624934
rect 316152 617218 316186 624934
rect 316610 617218 316644 624934
rect 317068 617218 317102 624934
rect 317526 617218 317560 624934
rect 317984 617218 318018 624934
rect 318442 617218 318476 624934
rect 313558 617125 313742 617159
rect 314016 617125 314200 617159
rect 314474 617125 314658 617159
rect 314932 617125 315116 617159
rect 315390 617125 315574 617159
rect 315848 617125 316032 617159
rect 316306 617125 316490 617159
rect 316764 617125 316948 617159
rect 317222 617125 317406 617159
rect 317680 617125 317864 617159
rect 318138 617125 318322 617159
rect 312804 616608 313204 616708
rect 319362 617218 319396 624934
rect 319820 617218 319854 624934
rect 320278 617218 320312 624934
rect 320736 617218 320770 624934
rect 321194 617218 321228 624934
rect 321652 617218 321686 624934
rect 322110 617218 322144 624934
rect 322568 617218 322602 624934
rect 323026 617218 323060 624934
rect 323484 617218 323518 624934
rect 323942 617218 323976 624934
rect 319516 617125 319700 617159
rect 319974 617125 320158 617159
rect 320432 617125 320616 617159
rect 320890 617125 321074 617159
rect 321348 617125 321532 617159
rect 321806 617125 321990 617159
rect 322264 617125 322448 617159
rect 322722 617125 322906 617159
rect 323180 617125 323364 617159
rect 323638 617125 323822 617159
rect 318714 616608 319114 616708
rect 324862 617218 324896 624934
rect 325320 617218 325354 624934
rect 325778 617218 325812 624934
rect 326236 617218 326270 624934
rect 326694 617218 326728 624934
rect 327152 617218 327186 624934
rect 327610 617218 327644 624934
rect 328068 617218 328102 624934
rect 328526 617218 328560 624934
rect 328984 617218 329018 624934
rect 329442 617218 329476 624934
rect 329900 617218 329934 624934
rect 325016 617125 325200 617159
rect 325474 617125 325658 617159
rect 325932 617125 326116 617159
rect 326390 617125 326574 617159
rect 326848 617125 327032 617159
rect 327306 617125 327490 617159
rect 327764 617125 327948 617159
rect 328222 617125 328406 617159
rect 328680 617125 328864 617159
rect 329138 617125 329322 617159
rect 329596 617125 329780 617159
rect 324214 616608 324614 616708
rect 335032 624772 335038 624794
rect 335038 624772 335066 624794
rect 335032 624760 335066 624772
rect 335132 624760 335166 624794
rect 335232 624760 335266 624794
rect 335332 624772 335364 624794
rect 335364 624772 335366 624794
rect 335432 624772 335454 624794
rect 335454 624772 335466 624794
rect 335532 624772 335544 624794
rect 335544 624772 335566 624794
rect 335332 624760 335366 624772
rect 335432 624760 335466 624772
rect 335532 624760 335566 624772
rect 335032 624682 335038 624694
rect 335038 624682 335066 624694
rect 335032 624660 335066 624682
rect 335132 624660 335166 624694
rect 335232 624660 335266 624694
rect 335332 624682 335364 624694
rect 335364 624682 335366 624694
rect 335432 624682 335454 624694
rect 335454 624682 335466 624694
rect 335532 624682 335544 624694
rect 335544 624682 335566 624694
rect 335332 624660 335366 624682
rect 335432 624660 335466 624682
rect 335532 624660 335566 624682
rect 335032 624592 335038 624594
rect 335038 624592 335066 624594
rect 335032 624560 335066 624592
rect 335132 624560 335166 624594
rect 335232 624560 335266 624594
rect 335332 624592 335364 624594
rect 335364 624592 335366 624594
rect 335432 624592 335454 624594
rect 335454 624592 335466 624594
rect 335532 624592 335544 624594
rect 335544 624592 335566 624594
rect 335332 624560 335366 624592
rect 335432 624560 335466 624592
rect 335532 624560 335566 624592
rect 335032 624460 335066 624494
rect 335132 624460 335166 624494
rect 335232 624460 335266 624494
rect 335332 624460 335366 624494
rect 335432 624460 335466 624494
rect 335532 624460 335566 624494
rect 335032 624360 335066 624394
rect 335132 624360 335166 624394
rect 335232 624360 335266 624394
rect 335332 624360 335366 624394
rect 335432 624360 335466 624394
rect 335532 624360 335566 624394
rect 335032 624266 335066 624294
rect 335032 624260 335038 624266
rect 335038 624260 335066 624266
rect 335132 624260 335166 624294
rect 335232 624260 335266 624294
rect 335332 624266 335366 624294
rect 335432 624266 335466 624294
rect 335532 624266 335566 624294
rect 335332 624260 335364 624266
rect 335364 624260 335366 624266
rect 335432 624260 335454 624266
rect 335454 624260 335466 624266
rect 335532 624260 335544 624266
rect 335544 624260 335566 624266
rect 336320 624772 336326 624794
rect 336326 624772 336354 624794
rect 336320 624760 336354 624772
rect 336420 624760 336454 624794
rect 336520 624760 336554 624794
rect 336620 624772 336652 624794
rect 336652 624772 336654 624794
rect 336720 624772 336742 624794
rect 336742 624772 336754 624794
rect 336820 624772 336832 624794
rect 336832 624772 336854 624794
rect 336620 624760 336654 624772
rect 336720 624760 336754 624772
rect 336820 624760 336854 624772
rect 336320 624682 336326 624694
rect 336326 624682 336354 624694
rect 336320 624660 336354 624682
rect 336420 624660 336454 624694
rect 336520 624660 336554 624694
rect 336620 624682 336652 624694
rect 336652 624682 336654 624694
rect 336720 624682 336742 624694
rect 336742 624682 336754 624694
rect 336820 624682 336832 624694
rect 336832 624682 336854 624694
rect 336620 624660 336654 624682
rect 336720 624660 336754 624682
rect 336820 624660 336854 624682
rect 336320 624592 336326 624594
rect 336326 624592 336354 624594
rect 336320 624560 336354 624592
rect 336420 624560 336454 624594
rect 336520 624560 336554 624594
rect 336620 624592 336652 624594
rect 336652 624592 336654 624594
rect 336720 624592 336742 624594
rect 336742 624592 336754 624594
rect 336820 624592 336832 624594
rect 336832 624592 336854 624594
rect 336620 624560 336654 624592
rect 336720 624560 336754 624592
rect 336820 624560 336854 624592
rect 336320 624460 336354 624494
rect 336420 624460 336454 624494
rect 336520 624460 336554 624494
rect 336620 624460 336654 624494
rect 336720 624460 336754 624494
rect 336820 624460 336854 624494
rect 336320 624360 336354 624394
rect 336420 624360 336454 624394
rect 336520 624360 336554 624394
rect 336620 624360 336654 624394
rect 336720 624360 336754 624394
rect 336820 624360 336854 624394
rect 336320 624266 336354 624294
rect 336320 624260 336326 624266
rect 336326 624260 336354 624266
rect 336420 624260 336454 624294
rect 336520 624260 336554 624294
rect 336620 624266 336654 624294
rect 336720 624266 336754 624294
rect 336820 624266 336854 624294
rect 336620 624260 336652 624266
rect 336652 624260 336654 624266
rect 336720 624260 336742 624266
rect 336742 624260 336754 624266
rect 336820 624260 336832 624266
rect 336832 624260 336854 624266
rect 337608 624772 337614 624794
rect 337614 624772 337642 624794
rect 337608 624760 337642 624772
rect 337708 624760 337742 624794
rect 337808 624760 337842 624794
rect 337908 624772 337940 624794
rect 337940 624772 337942 624794
rect 338008 624772 338030 624794
rect 338030 624772 338042 624794
rect 338108 624772 338120 624794
rect 338120 624772 338142 624794
rect 337908 624760 337942 624772
rect 338008 624760 338042 624772
rect 338108 624760 338142 624772
rect 337608 624682 337614 624694
rect 337614 624682 337642 624694
rect 337608 624660 337642 624682
rect 337708 624660 337742 624694
rect 337808 624660 337842 624694
rect 337908 624682 337940 624694
rect 337940 624682 337942 624694
rect 338008 624682 338030 624694
rect 338030 624682 338042 624694
rect 338108 624682 338120 624694
rect 338120 624682 338142 624694
rect 337908 624660 337942 624682
rect 338008 624660 338042 624682
rect 338108 624660 338142 624682
rect 337608 624592 337614 624594
rect 337614 624592 337642 624594
rect 337608 624560 337642 624592
rect 337708 624560 337742 624594
rect 337808 624560 337842 624594
rect 337908 624592 337940 624594
rect 337940 624592 337942 624594
rect 338008 624592 338030 624594
rect 338030 624592 338042 624594
rect 338108 624592 338120 624594
rect 338120 624592 338142 624594
rect 337908 624560 337942 624592
rect 338008 624560 338042 624592
rect 338108 624560 338142 624592
rect 337608 624460 337642 624494
rect 337708 624460 337742 624494
rect 337808 624460 337842 624494
rect 337908 624460 337942 624494
rect 338008 624460 338042 624494
rect 338108 624460 338142 624494
rect 337608 624360 337642 624394
rect 337708 624360 337742 624394
rect 337808 624360 337842 624394
rect 337908 624360 337942 624394
rect 338008 624360 338042 624394
rect 338108 624360 338142 624394
rect 337608 624266 337642 624294
rect 337608 624260 337614 624266
rect 337614 624260 337642 624266
rect 337708 624260 337742 624294
rect 337808 624260 337842 624294
rect 337908 624266 337942 624294
rect 338008 624266 338042 624294
rect 338108 624266 338142 624294
rect 337908 624260 337940 624266
rect 337940 624260 337942 624266
rect 338008 624260 338030 624266
rect 338030 624260 338042 624266
rect 338108 624260 338120 624266
rect 338120 624260 338142 624266
rect 338896 624772 338902 624794
rect 338902 624772 338930 624794
rect 338896 624760 338930 624772
rect 338996 624760 339030 624794
rect 339096 624760 339130 624794
rect 339196 624772 339228 624794
rect 339228 624772 339230 624794
rect 339296 624772 339318 624794
rect 339318 624772 339330 624794
rect 339396 624772 339408 624794
rect 339408 624772 339430 624794
rect 339196 624760 339230 624772
rect 339296 624760 339330 624772
rect 339396 624760 339430 624772
rect 338896 624682 338902 624694
rect 338902 624682 338930 624694
rect 338896 624660 338930 624682
rect 338996 624660 339030 624694
rect 339096 624660 339130 624694
rect 339196 624682 339228 624694
rect 339228 624682 339230 624694
rect 339296 624682 339318 624694
rect 339318 624682 339330 624694
rect 339396 624682 339408 624694
rect 339408 624682 339430 624694
rect 339196 624660 339230 624682
rect 339296 624660 339330 624682
rect 339396 624660 339430 624682
rect 338896 624592 338902 624594
rect 338902 624592 338930 624594
rect 338896 624560 338930 624592
rect 338996 624560 339030 624594
rect 339096 624560 339130 624594
rect 339196 624592 339228 624594
rect 339228 624592 339230 624594
rect 339296 624592 339318 624594
rect 339318 624592 339330 624594
rect 339396 624592 339408 624594
rect 339408 624592 339430 624594
rect 339196 624560 339230 624592
rect 339296 624560 339330 624592
rect 339396 624560 339430 624592
rect 338896 624460 338930 624494
rect 338996 624460 339030 624494
rect 339096 624460 339130 624494
rect 339196 624460 339230 624494
rect 339296 624460 339330 624494
rect 339396 624460 339430 624494
rect 338896 624360 338930 624394
rect 338996 624360 339030 624394
rect 339096 624360 339130 624394
rect 339196 624360 339230 624394
rect 339296 624360 339330 624394
rect 339396 624360 339430 624394
rect 338896 624266 338930 624294
rect 338896 624260 338902 624266
rect 338902 624260 338930 624266
rect 338996 624260 339030 624294
rect 339096 624260 339130 624294
rect 339196 624266 339230 624294
rect 339296 624266 339330 624294
rect 339396 624266 339430 624294
rect 339196 624260 339228 624266
rect 339228 624260 339230 624266
rect 339296 624260 339318 624266
rect 339318 624260 339330 624266
rect 339396 624260 339408 624266
rect 339408 624260 339430 624266
rect 340184 624772 340190 624794
rect 340190 624772 340218 624794
rect 340184 624760 340218 624772
rect 340284 624760 340318 624794
rect 340384 624760 340418 624794
rect 340484 624772 340516 624794
rect 340516 624772 340518 624794
rect 340584 624772 340606 624794
rect 340606 624772 340618 624794
rect 340684 624772 340696 624794
rect 340696 624772 340718 624794
rect 340484 624760 340518 624772
rect 340584 624760 340618 624772
rect 340684 624760 340718 624772
rect 340184 624682 340190 624694
rect 340190 624682 340218 624694
rect 340184 624660 340218 624682
rect 340284 624660 340318 624694
rect 340384 624660 340418 624694
rect 340484 624682 340516 624694
rect 340516 624682 340518 624694
rect 340584 624682 340606 624694
rect 340606 624682 340618 624694
rect 340684 624682 340696 624694
rect 340696 624682 340718 624694
rect 340484 624660 340518 624682
rect 340584 624660 340618 624682
rect 340684 624660 340718 624682
rect 340184 624592 340190 624594
rect 340190 624592 340218 624594
rect 340184 624560 340218 624592
rect 340284 624560 340318 624594
rect 340384 624560 340418 624594
rect 340484 624592 340516 624594
rect 340516 624592 340518 624594
rect 340584 624592 340606 624594
rect 340606 624592 340618 624594
rect 340684 624592 340696 624594
rect 340696 624592 340718 624594
rect 340484 624560 340518 624592
rect 340584 624560 340618 624592
rect 340684 624560 340718 624592
rect 340184 624460 340218 624494
rect 340284 624460 340318 624494
rect 340384 624460 340418 624494
rect 340484 624460 340518 624494
rect 340584 624460 340618 624494
rect 340684 624460 340718 624494
rect 340184 624360 340218 624394
rect 340284 624360 340318 624394
rect 340384 624360 340418 624394
rect 340484 624360 340518 624394
rect 340584 624360 340618 624394
rect 340684 624360 340718 624394
rect 340184 624266 340218 624294
rect 340184 624260 340190 624266
rect 340190 624260 340218 624266
rect 340284 624260 340318 624294
rect 340384 624260 340418 624294
rect 340484 624266 340518 624294
rect 340584 624266 340618 624294
rect 340684 624266 340718 624294
rect 340484 624260 340516 624266
rect 340516 624260 340518 624266
rect 340584 624260 340606 624266
rect 340606 624260 340618 624266
rect 340684 624260 340696 624266
rect 340696 624260 340718 624266
rect 335032 623484 335038 623506
rect 335038 623484 335066 623506
rect 335032 623472 335066 623484
rect 335132 623472 335166 623506
rect 335232 623472 335266 623506
rect 335332 623484 335364 623506
rect 335364 623484 335366 623506
rect 335432 623484 335454 623506
rect 335454 623484 335466 623506
rect 335532 623484 335544 623506
rect 335544 623484 335566 623506
rect 335332 623472 335366 623484
rect 335432 623472 335466 623484
rect 335532 623472 335566 623484
rect 335032 623394 335038 623406
rect 335038 623394 335066 623406
rect 335032 623372 335066 623394
rect 335132 623372 335166 623406
rect 335232 623372 335266 623406
rect 335332 623394 335364 623406
rect 335364 623394 335366 623406
rect 335432 623394 335454 623406
rect 335454 623394 335466 623406
rect 335532 623394 335544 623406
rect 335544 623394 335566 623406
rect 335332 623372 335366 623394
rect 335432 623372 335466 623394
rect 335532 623372 335566 623394
rect 335032 623304 335038 623306
rect 335038 623304 335066 623306
rect 335032 623272 335066 623304
rect 335132 623272 335166 623306
rect 335232 623272 335266 623306
rect 335332 623304 335364 623306
rect 335364 623304 335366 623306
rect 335432 623304 335454 623306
rect 335454 623304 335466 623306
rect 335532 623304 335544 623306
rect 335544 623304 335566 623306
rect 335332 623272 335366 623304
rect 335432 623272 335466 623304
rect 335532 623272 335566 623304
rect 335032 623172 335066 623206
rect 335132 623172 335166 623206
rect 335232 623172 335266 623206
rect 335332 623172 335366 623206
rect 335432 623172 335466 623206
rect 335532 623172 335566 623206
rect 335032 623072 335066 623106
rect 335132 623072 335166 623106
rect 335232 623072 335266 623106
rect 335332 623072 335366 623106
rect 335432 623072 335466 623106
rect 335532 623072 335566 623106
rect 335032 622978 335066 623006
rect 335032 622972 335038 622978
rect 335038 622972 335066 622978
rect 335132 622972 335166 623006
rect 335232 622972 335266 623006
rect 335332 622978 335366 623006
rect 335432 622978 335466 623006
rect 335532 622978 335566 623006
rect 335332 622972 335364 622978
rect 335364 622972 335366 622978
rect 335432 622972 335454 622978
rect 335454 622972 335466 622978
rect 335532 622972 335544 622978
rect 335544 622972 335566 622978
rect 336320 623484 336326 623506
rect 336326 623484 336354 623506
rect 336320 623472 336354 623484
rect 336420 623472 336454 623506
rect 336520 623472 336554 623506
rect 336620 623484 336652 623506
rect 336652 623484 336654 623506
rect 336720 623484 336742 623506
rect 336742 623484 336754 623506
rect 336820 623484 336832 623506
rect 336832 623484 336854 623506
rect 336620 623472 336654 623484
rect 336720 623472 336754 623484
rect 336820 623472 336854 623484
rect 336320 623394 336326 623406
rect 336326 623394 336354 623406
rect 336320 623372 336354 623394
rect 336420 623372 336454 623406
rect 336520 623372 336554 623406
rect 336620 623394 336652 623406
rect 336652 623394 336654 623406
rect 336720 623394 336742 623406
rect 336742 623394 336754 623406
rect 336820 623394 336832 623406
rect 336832 623394 336854 623406
rect 336620 623372 336654 623394
rect 336720 623372 336754 623394
rect 336820 623372 336854 623394
rect 336320 623304 336326 623306
rect 336326 623304 336354 623306
rect 336320 623272 336354 623304
rect 336420 623272 336454 623306
rect 336520 623272 336554 623306
rect 336620 623304 336652 623306
rect 336652 623304 336654 623306
rect 336720 623304 336742 623306
rect 336742 623304 336754 623306
rect 336820 623304 336832 623306
rect 336832 623304 336854 623306
rect 336620 623272 336654 623304
rect 336720 623272 336754 623304
rect 336820 623272 336854 623304
rect 336320 623172 336354 623206
rect 336420 623172 336454 623206
rect 336520 623172 336554 623206
rect 336620 623172 336654 623206
rect 336720 623172 336754 623206
rect 336820 623172 336854 623206
rect 336320 623072 336354 623106
rect 336420 623072 336454 623106
rect 336520 623072 336554 623106
rect 336620 623072 336654 623106
rect 336720 623072 336754 623106
rect 336820 623072 336854 623106
rect 336320 622978 336354 623006
rect 336320 622972 336326 622978
rect 336326 622972 336354 622978
rect 336420 622972 336454 623006
rect 336520 622972 336554 623006
rect 336620 622978 336654 623006
rect 336720 622978 336754 623006
rect 336820 622978 336854 623006
rect 336620 622972 336652 622978
rect 336652 622972 336654 622978
rect 336720 622972 336742 622978
rect 336742 622972 336754 622978
rect 336820 622972 336832 622978
rect 336832 622972 336854 622978
rect 337608 623484 337614 623506
rect 337614 623484 337642 623506
rect 337608 623472 337642 623484
rect 337708 623472 337742 623506
rect 337808 623472 337842 623506
rect 337908 623484 337940 623506
rect 337940 623484 337942 623506
rect 338008 623484 338030 623506
rect 338030 623484 338042 623506
rect 338108 623484 338120 623506
rect 338120 623484 338142 623506
rect 337908 623472 337942 623484
rect 338008 623472 338042 623484
rect 338108 623472 338142 623484
rect 337608 623394 337614 623406
rect 337614 623394 337642 623406
rect 337608 623372 337642 623394
rect 337708 623372 337742 623406
rect 337808 623372 337842 623406
rect 337908 623394 337940 623406
rect 337940 623394 337942 623406
rect 338008 623394 338030 623406
rect 338030 623394 338042 623406
rect 338108 623394 338120 623406
rect 338120 623394 338142 623406
rect 337908 623372 337942 623394
rect 338008 623372 338042 623394
rect 338108 623372 338142 623394
rect 337608 623304 337614 623306
rect 337614 623304 337642 623306
rect 337608 623272 337642 623304
rect 337708 623272 337742 623306
rect 337808 623272 337842 623306
rect 337908 623304 337940 623306
rect 337940 623304 337942 623306
rect 338008 623304 338030 623306
rect 338030 623304 338042 623306
rect 338108 623304 338120 623306
rect 338120 623304 338142 623306
rect 337908 623272 337942 623304
rect 338008 623272 338042 623304
rect 338108 623272 338142 623304
rect 337608 623172 337642 623206
rect 337708 623172 337742 623206
rect 337808 623172 337842 623206
rect 337908 623172 337942 623206
rect 338008 623172 338042 623206
rect 338108 623172 338142 623206
rect 337608 623072 337642 623106
rect 337708 623072 337742 623106
rect 337808 623072 337842 623106
rect 337908 623072 337942 623106
rect 338008 623072 338042 623106
rect 338108 623072 338142 623106
rect 337608 622978 337642 623006
rect 337608 622972 337614 622978
rect 337614 622972 337642 622978
rect 337708 622972 337742 623006
rect 337808 622972 337842 623006
rect 337908 622978 337942 623006
rect 338008 622978 338042 623006
rect 338108 622978 338142 623006
rect 337908 622972 337940 622978
rect 337940 622972 337942 622978
rect 338008 622972 338030 622978
rect 338030 622972 338042 622978
rect 338108 622972 338120 622978
rect 338120 622972 338142 622978
rect 338896 623484 338902 623506
rect 338902 623484 338930 623506
rect 338896 623472 338930 623484
rect 338996 623472 339030 623506
rect 339096 623472 339130 623506
rect 339196 623484 339228 623506
rect 339228 623484 339230 623506
rect 339296 623484 339318 623506
rect 339318 623484 339330 623506
rect 339396 623484 339408 623506
rect 339408 623484 339430 623506
rect 339196 623472 339230 623484
rect 339296 623472 339330 623484
rect 339396 623472 339430 623484
rect 338896 623394 338902 623406
rect 338902 623394 338930 623406
rect 338896 623372 338930 623394
rect 338996 623372 339030 623406
rect 339096 623372 339130 623406
rect 339196 623394 339228 623406
rect 339228 623394 339230 623406
rect 339296 623394 339318 623406
rect 339318 623394 339330 623406
rect 339396 623394 339408 623406
rect 339408 623394 339430 623406
rect 339196 623372 339230 623394
rect 339296 623372 339330 623394
rect 339396 623372 339430 623394
rect 338896 623304 338902 623306
rect 338902 623304 338930 623306
rect 338896 623272 338930 623304
rect 338996 623272 339030 623306
rect 339096 623272 339130 623306
rect 339196 623304 339228 623306
rect 339228 623304 339230 623306
rect 339296 623304 339318 623306
rect 339318 623304 339330 623306
rect 339396 623304 339408 623306
rect 339408 623304 339430 623306
rect 339196 623272 339230 623304
rect 339296 623272 339330 623304
rect 339396 623272 339430 623304
rect 338896 623172 338930 623206
rect 338996 623172 339030 623206
rect 339096 623172 339130 623206
rect 339196 623172 339230 623206
rect 339296 623172 339330 623206
rect 339396 623172 339430 623206
rect 338896 623072 338930 623106
rect 338996 623072 339030 623106
rect 339096 623072 339130 623106
rect 339196 623072 339230 623106
rect 339296 623072 339330 623106
rect 339396 623072 339430 623106
rect 338896 622978 338930 623006
rect 338896 622972 338902 622978
rect 338902 622972 338930 622978
rect 338996 622972 339030 623006
rect 339096 622972 339130 623006
rect 339196 622978 339230 623006
rect 339296 622978 339330 623006
rect 339396 622978 339430 623006
rect 339196 622972 339228 622978
rect 339228 622972 339230 622978
rect 339296 622972 339318 622978
rect 339318 622972 339330 622978
rect 339396 622972 339408 622978
rect 339408 622972 339430 622978
rect 340184 623484 340190 623506
rect 340190 623484 340218 623506
rect 340184 623472 340218 623484
rect 340284 623472 340318 623506
rect 340384 623472 340418 623506
rect 340484 623484 340516 623506
rect 340516 623484 340518 623506
rect 340584 623484 340606 623506
rect 340606 623484 340618 623506
rect 340684 623484 340696 623506
rect 340696 623484 340718 623506
rect 340484 623472 340518 623484
rect 340584 623472 340618 623484
rect 340684 623472 340718 623484
rect 340184 623394 340190 623406
rect 340190 623394 340218 623406
rect 340184 623372 340218 623394
rect 340284 623372 340318 623406
rect 340384 623372 340418 623406
rect 340484 623394 340516 623406
rect 340516 623394 340518 623406
rect 340584 623394 340606 623406
rect 340606 623394 340618 623406
rect 340684 623394 340696 623406
rect 340696 623394 340718 623406
rect 340484 623372 340518 623394
rect 340584 623372 340618 623394
rect 340684 623372 340718 623394
rect 340184 623304 340190 623306
rect 340190 623304 340218 623306
rect 340184 623272 340218 623304
rect 340284 623272 340318 623306
rect 340384 623272 340418 623306
rect 340484 623304 340516 623306
rect 340516 623304 340518 623306
rect 340584 623304 340606 623306
rect 340606 623304 340618 623306
rect 340684 623304 340696 623306
rect 340696 623304 340718 623306
rect 340484 623272 340518 623304
rect 340584 623272 340618 623304
rect 340684 623272 340718 623304
rect 340184 623172 340218 623206
rect 340284 623172 340318 623206
rect 340384 623172 340418 623206
rect 340484 623172 340518 623206
rect 340584 623172 340618 623206
rect 340684 623172 340718 623206
rect 340184 623072 340218 623106
rect 340284 623072 340318 623106
rect 340384 623072 340418 623106
rect 340484 623072 340518 623106
rect 340584 623072 340618 623106
rect 340684 623072 340718 623106
rect 340184 622978 340218 623006
rect 340184 622972 340190 622978
rect 340190 622972 340218 622978
rect 340284 622972 340318 623006
rect 340384 622972 340418 623006
rect 340484 622978 340518 623006
rect 340584 622978 340618 623006
rect 340684 622978 340718 623006
rect 340484 622972 340516 622978
rect 340516 622972 340518 622978
rect 340584 622972 340606 622978
rect 340606 622972 340618 622978
rect 340684 622972 340696 622978
rect 340696 622972 340718 622978
rect 335032 622196 335038 622218
rect 335038 622196 335066 622218
rect 335032 622184 335066 622196
rect 335132 622184 335166 622218
rect 335232 622184 335266 622218
rect 335332 622196 335364 622218
rect 335364 622196 335366 622218
rect 335432 622196 335454 622218
rect 335454 622196 335466 622218
rect 335532 622196 335544 622218
rect 335544 622196 335566 622218
rect 335332 622184 335366 622196
rect 335432 622184 335466 622196
rect 335532 622184 335566 622196
rect 335032 622106 335038 622118
rect 335038 622106 335066 622118
rect 335032 622084 335066 622106
rect 335132 622084 335166 622118
rect 335232 622084 335266 622118
rect 335332 622106 335364 622118
rect 335364 622106 335366 622118
rect 335432 622106 335454 622118
rect 335454 622106 335466 622118
rect 335532 622106 335544 622118
rect 335544 622106 335566 622118
rect 335332 622084 335366 622106
rect 335432 622084 335466 622106
rect 335532 622084 335566 622106
rect 335032 622016 335038 622018
rect 335038 622016 335066 622018
rect 335032 621984 335066 622016
rect 335132 621984 335166 622018
rect 335232 621984 335266 622018
rect 335332 622016 335364 622018
rect 335364 622016 335366 622018
rect 335432 622016 335454 622018
rect 335454 622016 335466 622018
rect 335532 622016 335544 622018
rect 335544 622016 335566 622018
rect 335332 621984 335366 622016
rect 335432 621984 335466 622016
rect 335532 621984 335566 622016
rect 335032 621884 335066 621918
rect 335132 621884 335166 621918
rect 335232 621884 335266 621918
rect 335332 621884 335366 621918
rect 335432 621884 335466 621918
rect 335532 621884 335566 621918
rect 335032 621784 335066 621818
rect 335132 621784 335166 621818
rect 335232 621784 335266 621818
rect 335332 621784 335366 621818
rect 335432 621784 335466 621818
rect 335532 621784 335566 621818
rect 335032 621690 335066 621718
rect 335032 621684 335038 621690
rect 335038 621684 335066 621690
rect 335132 621684 335166 621718
rect 335232 621684 335266 621718
rect 335332 621690 335366 621718
rect 335432 621690 335466 621718
rect 335532 621690 335566 621718
rect 335332 621684 335364 621690
rect 335364 621684 335366 621690
rect 335432 621684 335454 621690
rect 335454 621684 335466 621690
rect 335532 621684 335544 621690
rect 335544 621684 335566 621690
rect 336320 622196 336326 622218
rect 336326 622196 336354 622218
rect 336320 622184 336354 622196
rect 336420 622184 336454 622218
rect 336520 622184 336554 622218
rect 336620 622196 336652 622218
rect 336652 622196 336654 622218
rect 336720 622196 336742 622218
rect 336742 622196 336754 622218
rect 336820 622196 336832 622218
rect 336832 622196 336854 622218
rect 336620 622184 336654 622196
rect 336720 622184 336754 622196
rect 336820 622184 336854 622196
rect 336320 622106 336326 622118
rect 336326 622106 336354 622118
rect 336320 622084 336354 622106
rect 336420 622084 336454 622118
rect 336520 622084 336554 622118
rect 336620 622106 336652 622118
rect 336652 622106 336654 622118
rect 336720 622106 336742 622118
rect 336742 622106 336754 622118
rect 336820 622106 336832 622118
rect 336832 622106 336854 622118
rect 336620 622084 336654 622106
rect 336720 622084 336754 622106
rect 336820 622084 336854 622106
rect 336320 622016 336326 622018
rect 336326 622016 336354 622018
rect 336320 621984 336354 622016
rect 336420 621984 336454 622018
rect 336520 621984 336554 622018
rect 336620 622016 336652 622018
rect 336652 622016 336654 622018
rect 336720 622016 336742 622018
rect 336742 622016 336754 622018
rect 336820 622016 336832 622018
rect 336832 622016 336854 622018
rect 336620 621984 336654 622016
rect 336720 621984 336754 622016
rect 336820 621984 336854 622016
rect 336320 621884 336354 621918
rect 336420 621884 336454 621918
rect 336520 621884 336554 621918
rect 336620 621884 336654 621918
rect 336720 621884 336754 621918
rect 336820 621884 336854 621918
rect 336320 621784 336354 621818
rect 336420 621784 336454 621818
rect 336520 621784 336554 621818
rect 336620 621784 336654 621818
rect 336720 621784 336754 621818
rect 336820 621784 336854 621818
rect 336320 621690 336354 621718
rect 336320 621684 336326 621690
rect 336326 621684 336354 621690
rect 336420 621684 336454 621718
rect 336520 621684 336554 621718
rect 336620 621690 336654 621718
rect 336720 621690 336754 621718
rect 336820 621690 336854 621718
rect 336620 621684 336652 621690
rect 336652 621684 336654 621690
rect 336720 621684 336742 621690
rect 336742 621684 336754 621690
rect 336820 621684 336832 621690
rect 336832 621684 336854 621690
rect 337608 622196 337614 622218
rect 337614 622196 337642 622218
rect 337608 622184 337642 622196
rect 337708 622184 337742 622218
rect 337808 622184 337842 622218
rect 337908 622196 337940 622218
rect 337940 622196 337942 622218
rect 338008 622196 338030 622218
rect 338030 622196 338042 622218
rect 338108 622196 338120 622218
rect 338120 622196 338142 622218
rect 337908 622184 337942 622196
rect 338008 622184 338042 622196
rect 338108 622184 338142 622196
rect 337608 622106 337614 622118
rect 337614 622106 337642 622118
rect 337608 622084 337642 622106
rect 337708 622084 337742 622118
rect 337808 622084 337842 622118
rect 337908 622106 337940 622118
rect 337940 622106 337942 622118
rect 338008 622106 338030 622118
rect 338030 622106 338042 622118
rect 338108 622106 338120 622118
rect 338120 622106 338142 622118
rect 337908 622084 337942 622106
rect 338008 622084 338042 622106
rect 338108 622084 338142 622106
rect 337608 622016 337614 622018
rect 337614 622016 337642 622018
rect 337608 621984 337642 622016
rect 337708 621984 337742 622018
rect 337808 621984 337842 622018
rect 337908 622016 337940 622018
rect 337940 622016 337942 622018
rect 338008 622016 338030 622018
rect 338030 622016 338042 622018
rect 338108 622016 338120 622018
rect 338120 622016 338142 622018
rect 337908 621984 337942 622016
rect 338008 621984 338042 622016
rect 338108 621984 338142 622016
rect 337608 621884 337642 621918
rect 337708 621884 337742 621918
rect 337808 621884 337842 621918
rect 337908 621884 337942 621918
rect 338008 621884 338042 621918
rect 338108 621884 338142 621918
rect 337608 621784 337642 621818
rect 337708 621784 337742 621818
rect 337808 621784 337842 621818
rect 337908 621784 337942 621818
rect 338008 621784 338042 621818
rect 338108 621784 338142 621818
rect 337608 621690 337642 621718
rect 337608 621684 337614 621690
rect 337614 621684 337642 621690
rect 337708 621684 337742 621718
rect 337808 621684 337842 621718
rect 337908 621690 337942 621718
rect 338008 621690 338042 621718
rect 338108 621690 338142 621718
rect 337908 621684 337940 621690
rect 337940 621684 337942 621690
rect 338008 621684 338030 621690
rect 338030 621684 338042 621690
rect 338108 621684 338120 621690
rect 338120 621684 338142 621690
rect 338896 622196 338902 622218
rect 338902 622196 338930 622218
rect 338896 622184 338930 622196
rect 338996 622184 339030 622218
rect 339096 622184 339130 622218
rect 339196 622196 339228 622218
rect 339228 622196 339230 622218
rect 339296 622196 339318 622218
rect 339318 622196 339330 622218
rect 339396 622196 339408 622218
rect 339408 622196 339430 622218
rect 339196 622184 339230 622196
rect 339296 622184 339330 622196
rect 339396 622184 339430 622196
rect 338896 622106 338902 622118
rect 338902 622106 338930 622118
rect 338896 622084 338930 622106
rect 338996 622084 339030 622118
rect 339096 622084 339130 622118
rect 339196 622106 339228 622118
rect 339228 622106 339230 622118
rect 339296 622106 339318 622118
rect 339318 622106 339330 622118
rect 339396 622106 339408 622118
rect 339408 622106 339430 622118
rect 339196 622084 339230 622106
rect 339296 622084 339330 622106
rect 339396 622084 339430 622106
rect 338896 622016 338902 622018
rect 338902 622016 338930 622018
rect 338896 621984 338930 622016
rect 338996 621984 339030 622018
rect 339096 621984 339130 622018
rect 339196 622016 339228 622018
rect 339228 622016 339230 622018
rect 339296 622016 339318 622018
rect 339318 622016 339330 622018
rect 339396 622016 339408 622018
rect 339408 622016 339430 622018
rect 339196 621984 339230 622016
rect 339296 621984 339330 622016
rect 339396 621984 339430 622016
rect 338896 621884 338930 621918
rect 338996 621884 339030 621918
rect 339096 621884 339130 621918
rect 339196 621884 339230 621918
rect 339296 621884 339330 621918
rect 339396 621884 339430 621918
rect 338896 621784 338930 621818
rect 338996 621784 339030 621818
rect 339096 621784 339130 621818
rect 339196 621784 339230 621818
rect 339296 621784 339330 621818
rect 339396 621784 339430 621818
rect 338896 621690 338930 621718
rect 338896 621684 338902 621690
rect 338902 621684 338930 621690
rect 338996 621684 339030 621718
rect 339096 621684 339130 621718
rect 339196 621690 339230 621718
rect 339296 621690 339330 621718
rect 339396 621690 339430 621718
rect 339196 621684 339228 621690
rect 339228 621684 339230 621690
rect 339296 621684 339318 621690
rect 339318 621684 339330 621690
rect 339396 621684 339408 621690
rect 339408 621684 339430 621690
rect 340184 622196 340190 622218
rect 340190 622196 340218 622218
rect 340184 622184 340218 622196
rect 340284 622184 340318 622218
rect 340384 622184 340418 622218
rect 340484 622196 340516 622218
rect 340516 622196 340518 622218
rect 340584 622196 340606 622218
rect 340606 622196 340618 622218
rect 340684 622196 340696 622218
rect 340696 622196 340718 622218
rect 340484 622184 340518 622196
rect 340584 622184 340618 622196
rect 340684 622184 340718 622196
rect 340184 622106 340190 622118
rect 340190 622106 340218 622118
rect 340184 622084 340218 622106
rect 340284 622084 340318 622118
rect 340384 622084 340418 622118
rect 340484 622106 340516 622118
rect 340516 622106 340518 622118
rect 340584 622106 340606 622118
rect 340606 622106 340618 622118
rect 340684 622106 340696 622118
rect 340696 622106 340718 622118
rect 340484 622084 340518 622106
rect 340584 622084 340618 622106
rect 340684 622084 340718 622106
rect 340184 622016 340190 622018
rect 340190 622016 340218 622018
rect 340184 621984 340218 622016
rect 340284 621984 340318 622018
rect 340384 621984 340418 622018
rect 340484 622016 340516 622018
rect 340516 622016 340518 622018
rect 340584 622016 340606 622018
rect 340606 622016 340618 622018
rect 340684 622016 340696 622018
rect 340696 622016 340718 622018
rect 340484 621984 340518 622016
rect 340584 621984 340618 622016
rect 340684 621984 340718 622016
rect 340184 621884 340218 621918
rect 340284 621884 340318 621918
rect 340384 621884 340418 621918
rect 340484 621884 340518 621918
rect 340584 621884 340618 621918
rect 340684 621884 340718 621918
rect 340184 621784 340218 621818
rect 340284 621784 340318 621818
rect 340384 621784 340418 621818
rect 340484 621784 340518 621818
rect 340584 621784 340618 621818
rect 340684 621784 340718 621818
rect 340184 621690 340218 621718
rect 340184 621684 340190 621690
rect 340190 621684 340218 621690
rect 340284 621684 340318 621718
rect 340384 621684 340418 621718
rect 340484 621690 340518 621718
rect 340584 621690 340618 621718
rect 340684 621690 340718 621718
rect 340484 621684 340516 621690
rect 340516 621684 340518 621690
rect 340584 621684 340606 621690
rect 340606 621684 340618 621690
rect 340684 621684 340696 621690
rect 340696 621684 340718 621690
rect 335032 620908 335038 620930
rect 335038 620908 335066 620930
rect 335032 620896 335066 620908
rect 335132 620896 335166 620930
rect 335232 620896 335266 620930
rect 335332 620908 335364 620930
rect 335364 620908 335366 620930
rect 335432 620908 335454 620930
rect 335454 620908 335466 620930
rect 335532 620908 335544 620930
rect 335544 620908 335566 620930
rect 335332 620896 335366 620908
rect 335432 620896 335466 620908
rect 335532 620896 335566 620908
rect 335032 620818 335038 620830
rect 335038 620818 335066 620830
rect 335032 620796 335066 620818
rect 335132 620796 335166 620830
rect 335232 620796 335266 620830
rect 335332 620818 335364 620830
rect 335364 620818 335366 620830
rect 335432 620818 335454 620830
rect 335454 620818 335466 620830
rect 335532 620818 335544 620830
rect 335544 620818 335566 620830
rect 335332 620796 335366 620818
rect 335432 620796 335466 620818
rect 335532 620796 335566 620818
rect 335032 620728 335038 620730
rect 335038 620728 335066 620730
rect 335032 620696 335066 620728
rect 335132 620696 335166 620730
rect 335232 620696 335266 620730
rect 335332 620728 335364 620730
rect 335364 620728 335366 620730
rect 335432 620728 335454 620730
rect 335454 620728 335466 620730
rect 335532 620728 335544 620730
rect 335544 620728 335566 620730
rect 335332 620696 335366 620728
rect 335432 620696 335466 620728
rect 335532 620696 335566 620728
rect 335032 620596 335066 620630
rect 335132 620596 335166 620630
rect 335232 620596 335266 620630
rect 335332 620596 335366 620630
rect 335432 620596 335466 620630
rect 335532 620596 335566 620630
rect 335032 620496 335066 620530
rect 335132 620496 335166 620530
rect 335232 620496 335266 620530
rect 335332 620496 335366 620530
rect 335432 620496 335466 620530
rect 335532 620496 335566 620530
rect 335032 620402 335066 620430
rect 335032 620396 335038 620402
rect 335038 620396 335066 620402
rect 335132 620396 335166 620430
rect 335232 620396 335266 620430
rect 335332 620402 335366 620430
rect 335432 620402 335466 620430
rect 335532 620402 335566 620430
rect 335332 620396 335364 620402
rect 335364 620396 335366 620402
rect 335432 620396 335454 620402
rect 335454 620396 335466 620402
rect 335532 620396 335544 620402
rect 335544 620396 335566 620402
rect 336320 620908 336326 620930
rect 336326 620908 336354 620930
rect 336320 620896 336354 620908
rect 336420 620896 336454 620930
rect 336520 620896 336554 620930
rect 336620 620908 336652 620930
rect 336652 620908 336654 620930
rect 336720 620908 336742 620930
rect 336742 620908 336754 620930
rect 336820 620908 336832 620930
rect 336832 620908 336854 620930
rect 336620 620896 336654 620908
rect 336720 620896 336754 620908
rect 336820 620896 336854 620908
rect 336320 620818 336326 620830
rect 336326 620818 336354 620830
rect 336320 620796 336354 620818
rect 336420 620796 336454 620830
rect 336520 620796 336554 620830
rect 336620 620818 336652 620830
rect 336652 620818 336654 620830
rect 336720 620818 336742 620830
rect 336742 620818 336754 620830
rect 336820 620818 336832 620830
rect 336832 620818 336854 620830
rect 336620 620796 336654 620818
rect 336720 620796 336754 620818
rect 336820 620796 336854 620818
rect 336320 620728 336326 620730
rect 336326 620728 336354 620730
rect 336320 620696 336354 620728
rect 336420 620696 336454 620730
rect 336520 620696 336554 620730
rect 336620 620728 336652 620730
rect 336652 620728 336654 620730
rect 336720 620728 336742 620730
rect 336742 620728 336754 620730
rect 336820 620728 336832 620730
rect 336832 620728 336854 620730
rect 336620 620696 336654 620728
rect 336720 620696 336754 620728
rect 336820 620696 336854 620728
rect 336320 620596 336354 620630
rect 336420 620596 336454 620630
rect 336520 620596 336554 620630
rect 336620 620596 336654 620630
rect 336720 620596 336754 620630
rect 336820 620596 336854 620630
rect 336320 620496 336354 620530
rect 336420 620496 336454 620530
rect 336520 620496 336554 620530
rect 336620 620496 336654 620530
rect 336720 620496 336754 620530
rect 336820 620496 336854 620530
rect 336320 620402 336354 620430
rect 336320 620396 336326 620402
rect 336326 620396 336354 620402
rect 336420 620396 336454 620430
rect 336520 620396 336554 620430
rect 336620 620402 336654 620430
rect 336720 620402 336754 620430
rect 336820 620402 336854 620430
rect 336620 620396 336652 620402
rect 336652 620396 336654 620402
rect 336720 620396 336742 620402
rect 336742 620396 336754 620402
rect 336820 620396 336832 620402
rect 336832 620396 336854 620402
rect 337608 620908 337614 620930
rect 337614 620908 337642 620930
rect 337608 620896 337642 620908
rect 337708 620896 337742 620930
rect 337808 620896 337842 620930
rect 337908 620908 337940 620930
rect 337940 620908 337942 620930
rect 338008 620908 338030 620930
rect 338030 620908 338042 620930
rect 338108 620908 338120 620930
rect 338120 620908 338142 620930
rect 337908 620896 337942 620908
rect 338008 620896 338042 620908
rect 338108 620896 338142 620908
rect 337608 620818 337614 620830
rect 337614 620818 337642 620830
rect 337608 620796 337642 620818
rect 337708 620796 337742 620830
rect 337808 620796 337842 620830
rect 337908 620818 337940 620830
rect 337940 620818 337942 620830
rect 338008 620818 338030 620830
rect 338030 620818 338042 620830
rect 338108 620818 338120 620830
rect 338120 620818 338142 620830
rect 337908 620796 337942 620818
rect 338008 620796 338042 620818
rect 338108 620796 338142 620818
rect 337608 620728 337614 620730
rect 337614 620728 337642 620730
rect 337608 620696 337642 620728
rect 337708 620696 337742 620730
rect 337808 620696 337842 620730
rect 337908 620728 337940 620730
rect 337940 620728 337942 620730
rect 338008 620728 338030 620730
rect 338030 620728 338042 620730
rect 338108 620728 338120 620730
rect 338120 620728 338142 620730
rect 337908 620696 337942 620728
rect 338008 620696 338042 620728
rect 338108 620696 338142 620728
rect 337608 620596 337642 620630
rect 337708 620596 337742 620630
rect 337808 620596 337842 620630
rect 337908 620596 337942 620630
rect 338008 620596 338042 620630
rect 338108 620596 338142 620630
rect 337608 620496 337642 620530
rect 337708 620496 337742 620530
rect 337808 620496 337842 620530
rect 337908 620496 337942 620530
rect 338008 620496 338042 620530
rect 338108 620496 338142 620530
rect 337608 620402 337642 620430
rect 337608 620396 337614 620402
rect 337614 620396 337642 620402
rect 337708 620396 337742 620430
rect 337808 620396 337842 620430
rect 337908 620402 337942 620430
rect 338008 620402 338042 620430
rect 338108 620402 338142 620430
rect 337908 620396 337940 620402
rect 337940 620396 337942 620402
rect 338008 620396 338030 620402
rect 338030 620396 338042 620402
rect 338108 620396 338120 620402
rect 338120 620396 338142 620402
rect 338896 620908 338902 620930
rect 338902 620908 338930 620930
rect 338896 620896 338930 620908
rect 338996 620896 339030 620930
rect 339096 620896 339130 620930
rect 339196 620908 339228 620930
rect 339228 620908 339230 620930
rect 339296 620908 339318 620930
rect 339318 620908 339330 620930
rect 339396 620908 339408 620930
rect 339408 620908 339430 620930
rect 339196 620896 339230 620908
rect 339296 620896 339330 620908
rect 339396 620896 339430 620908
rect 338896 620818 338902 620830
rect 338902 620818 338930 620830
rect 338896 620796 338930 620818
rect 338996 620796 339030 620830
rect 339096 620796 339130 620830
rect 339196 620818 339228 620830
rect 339228 620818 339230 620830
rect 339296 620818 339318 620830
rect 339318 620818 339330 620830
rect 339396 620818 339408 620830
rect 339408 620818 339430 620830
rect 339196 620796 339230 620818
rect 339296 620796 339330 620818
rect 339396 620796 339430 620818
rect 338896 620728 338902 620730
rect 338902 620728 338930 620730
rect 338896 620696 338930 620728
rect 338996 620696 339030 620730
rect 339096 620696 339130 620730
rect 339196 620728 339228 620730
rect 339228 620728 339230 620730
rect 339296 620728 339318 620730
rect 339318 620728 339330 620730
rect 339396 620728 339408 620730
rect 339408 620728 339430 620730
rect 339196 620696 339230 620728
rect 339296 620696 339330 620728
rect 339396 620696 339430 620728
rect 338896 620596 338930 620630
rect 338996 620596 339030 620630
rect 339096 620596 339130 620630
rect 339196 620596 339230 620630
rect 339296 620596 339330 620630
rect 339396 620596 339430 620630
rect 338896 620496 338930 620530
rect 338996 620496 339030 620530
rect 339096 620496 339130 620530
rect 339196 620496 339230 620530
rect 339296 620496 339330 620530
rect 339396 620496 339430 620530
rect 338896 620402 338930 620430
rect 338896 620396 338902 620402
rect 338902 620396 338930 620402
rect 338996 620396 339030 620430
rect 339096 620396 339130 620430
rect 339196 620402 339230 620430
rect 339296 620402 339330 620430
rect 339396 620402 339430 620430
rect 339196 620396 339228 620402
rect 339228 620396 339230 620402
rect 339296 620396 339318 620402
rect 339318 620396 339330 620402
rect 339396 620396 339408 620402
rect 339408 620396 339430 620402
rect 340184 620908 340190 620930
rect 340190 620908 340218 620930
rect 340184 620896 340218 620908
rect 340284 620896 340318 620930
rect 340384 620896 340418 620930
rect 340484 620908 340516 620930
rect 340516 620908 340518 620930
rect 340584 620908 340606 620930
rect 340606 620908 340618 620930
rect 340684 620908 340696 620930
rect 340696 620908 340718 620930
rect 340484 620896 340518 620908
rect 340584 620896 340618 620908
rect 340684 620896 340718 620908
rect 340184 620818 340190 620830
rect 340190 620818 340218 620830
rect 340184 620796 340218 620818
rect 340284 620796 340318 620830
rect 340384 620796 340418 620830
rect 340484 620818 340516 620830
rect 340516 620818 340518 620830
rect 340584 620818 340606 620830
rect 340606 620818 340618 620830
rect 340684 620818 340696 620830
rect 340696 620818 340718 620830
rect 340484 620796 340518 620818
rect 340584 620796 340618 620818
rect 340684 620796 340718 620818
rect 340184 620728 340190 620730
rect 340190 620728 340218 620730
rect 340184 620696 340218 620728
rect 340284 620696 340318 620730
rect 340384 620696 340418 620730
rect 340484 620728 340516 620730
rect 340516 620728 340518 620730
rect 340584 620728 340606 620730
rect 340606 620728 340618 620730
rect 340684 620728 340696 620730
rect 340696 620728 340718 620730
rect 340484 620696 340518 620728
rect 340584 620696 340618 620728
rect 340684 620696 340718 620728
rect 340184 620596 340218 620630
rect 340284 620596 340318 620630
rect 340384 620596 340418 620630
rect 340484 620596 340518 620630
rect 340584 620596 340618 620630
rect 340684 620596 340718 620630
rect 340184 620496 340218 620530
rect 340284 620496 340318 620530
rect 340384 620496 340418 620530
rect 340484 620496 340518 620530
rect 340584 620496 340618 620530
rect 340684 620496 340718 620530
rect 340184 620402 340218 620430
rect 340184 620396 340190 620402
rect 340190 620396 340218 620402
rect 340284 620396 340318 620430
rect 340384 620396 340418 620430
rect 340484 620402 340518 620430
rect 340584 620402 340618 620430
rect 340684 620402 340718 620430
rect 340484 620396 340516 620402
rect 340516 620396 340518 620402
rect 340584 620396 340606 620402
rect 340606 620396 340618 620402
rect 340684 620396 340696 620402
rect 340696 620396 340718 620402
rect 335032 619620 335038 619642
rect 335038 619620 335066 619642
rect 335032 619608 335066 619620
rect 335132 619608 335166 619642
rect 335232 619608 335266 619642
rect 335332 619620 335364 619642
rect 335364 619620 335366 619642
rect 335432 619620 335454 619642
rect 335454 619620 335466 619642
rect 335532 619620 335544 619642
rect 335544 619620 335566 619642
rect 335332 619608 335366 619620
rect 335432 619608 335466 619620
rect 335532 619608 335566 619620
rect 335032 619530 335038 619542
rect 335038 619530 335066 619542
rect 335032 619508 335066 619530
rect 335132 619508 335166 619542
rect 335232 619508 335266 619542
rect 335332 619530 335364 619542
rect 335364 619530 335366 619542
rect 335432 619530 335454 619542
rect 335454 619530 335466 619542
rect 335532 619530 335544 619542
rect 335544 619530 335566 619542
rect 335332 619508 335366 619530
rect 335432 619508 335466 619530
rect 335532 619508 335566 619530
rect 335032 619440 335038 619442
rect 335038 619440 335066 619442
rect 335032 619408 335066 619440
rect 335132 619408 335166 619442
rect 335232 619408 335266 619442
rect 335332 619440 335364 619442
rect 335364 619440 335366 619442
rect 335432 619440 335454 619442
rect 335454 619440 335466 619442
rect 335532 619440 335544 619442
rect 335544 619440 335566 619442
rect 335332 619408 335366 619440
rect 335432 619408 335466 619440
rect 335532 619408 335566 619440
rect 335032 619308 335066 619342
rect 335132 619308 335166 619342
rect 335232 619308 335266 619342
rect 335332 619308 335366 619342
rect 335432 619308 335466 619342
rect 335532 619308 335566 619342
rect 335032 619208 335066 619242
rect 335132 619208 335166 619242
rect 335232 619208 335266 619242
rect 335332 619208 335366 619242
rect 335432 619208 335466 619242
rect 335532 619208 335566 619242
rect 335032 619114 335066 619142
rect 335032 619108 335038 619114
rect 335038 619108 335066 619114
rect 335132 619108 335166 619142
rect 335232 619108 335266 619142
rect 335332 619114 335366 619142
rect 335432 619114 335466 619142
rect 335532 619114 335566 619142
rect 335332 619108 335364 619114
rect 335364 619108 335366 619114
rect 335432 619108 335454 619114
rect 335454 619108 335466 619114
rect 335532 619108 335544 619114
rect 335544 619108 335566 619114
rect 336320 619620 336326 619642
rect 336326 619620 336354 619642
rect 336320 619608 336354 619620
rect 336420 619608 336454 619642
rect 336520 619608 336554 619642
rect 336620 619620 336652 619642
rect 336652 619620 336654 619642
rect 336720 619620 336742 619642
rect 336742 619620 336754 619642
rect 336820 619620 336832 619642
rect 336832 619620 336854 619642
rect 336620 619608 336654 619620
rect 336720 619608 336754 619620
rect 336820 619608 336854 619620
rect 336320 619530 336326 619542
rect 336326 619530 336354 619542
rect 336320 619508 336354 619530
rect 336420 619508 336454 619542
rect 336520 619508 336554 619542
rect 336620 619530 336652 619542
rect 336652 619530 336654 619542
rect 336720 619530 336742 619542
rect 336742 619530 336754 619542
rect 336820 619530 336832 619542
rect 336832 619530 336854 619542
rect 336620 619508 336654 619530
rect 336720 619508 336754 619530
rect 336820 619508 336854 619530
rect 336320 619440 336326 619442
rect 336326 619440 336354 619442
rect 336320 619408 336354 619440
rect 336420 619408 336454 619442
rect 336520 619408 336554 619442
rect 336620 619440 336652 619442
rect 336652 619440 336654 619442
rect 336720 619440 336742 619442
rect 336742 619440 336754 619442
rect 336820 619440 336832 619442
rect 336832 619440 336854 619442
rect 336620 619408 336654 619440
rect 336720 619408 336754 619440
rect 336820 619408 336854 619440
rect 336320 619308 336354 619342
rect 336420 619308 336454 619342
rect 336520 619308 336554 619342
rect 336620 619308 336654 619342
rect 336720 619308 336754 619342
rect 336820 619308 336854 619342
rect 336320 619208 336354 619242
rect 336420 619208 336454 619242
rect 336520 619208 336554 619242
rect 336620 619208 336654 619242
rect 336720 619208 336754 619242
rect 336820 619208 336854 619242
rect 336320 619114 336354 619142
rect 336320 619108 336326 619114
rect 336326 619108 336354 619114
rect 336420 619108 336454 619142
rect 336520 619108 336554 619142
rect 336620 619114 336654 619142
rect 336720 619114 336754 619142
rect 336820 619114 336854 619142
rect 336620 619108 336652 619114
rect 336652 619108 336654 619114
rect 336720 619108 336742 619114
rect 336742 619108 336754 619114
rect 336820 619108 336832 619114
rect 336832 619108 336854 619114
rect 337608 619620 337614 619642
rect 337614 619620 337642 619642
rect 337608 619608 337642 619620
rect 337708 619608 337742 619642
rect 337808 619608 337842 619642
rect 337908 619620 337940 619642
rect 337940 619620 337942 619642
rect 338008 619620 338030 619642
rect 338030 619620 338042 619642
rect 338108 619620 338120 619642
rect 338120 619620 338142 619642
rect 337908 619608 337942 619620
rect 338008 619608 338042 619620
rect 338108 619608 338142 619620
rect 337608 619530 337614 619542
rect 337614 619530 337642 619542
rect 337608 619508 337642 619530
rect 337708 619508 337742 619542
rect 337808 619508 337842 619542
rect 337908 619530 337940 619542
rect 337940 619530 337942 619542
rect 338008 619530 338030 619542
rect 338030 619530 338042 619542
rect 338108 619530 338120 619542
rect 338120 619530 338142 619542
rect 337908 619508 337942 619530
rect 338008 619508 338042 619530
rect 338108 619508 338142 619530
rect 337608 619440 337614 619442
rect 337614 619440 337642 619442
rect 337608 619408 337642 619440
rect 337708 619408 337742 619442
rect 337808 619408 337842 619442
rect 337908 619440 337940 619442
rect 337940 619440 337942 619442
rect 338008 619440 338030 619442
rect 338030 619440 338042 619442
rect 338108 619440 338120 619442
rect 338120 619440 338142 619442
rect 337908 619408 337942 619440
rect 338008 619408 338042 619440
rect 338108 619408 338142 619440
rect 337608 619308 337642 619342
rect 337708 619308 337742 619342
rect 337808 619308 337842 619342
rect 337908 619308 337942 619342
rect 338008 619308 338042 619342
rect 338108 619308 338142 619342
rect 337608 619208 337642 619242
rect 337708 619208 337742 619242
rect 337808 619208 337842 619242
rect 337908 619208 337942 619242
rect 338008 619208 338042 619242
rect 338108 619208 338142 619242
rect 337608 619114 337642 619142
rect 337608 619108 337614 619114
rect 337614 619108 337642 619114
rect 337708 619108 337742 619142
rect 337808 619108 337842 619142
rect 337908 619114 337942 619142
rect 338008 619114 338042 619142
rect 338108 619114 338142 619142
rect 337908 619108 337940 619114
rect 337940 619108 337942 619114
rect 338008 619108 338030 619114
rect 338030 619108 338042 619114
rect 338108 619108 338120 619114
rect 338120 619108 338142 619114
rect 338896 619620 338902 619642
rect 338902 619620 338930 619642
rect 338896 619608 338930 619620
rect 338996 619608 339030 619642
rect 339096 619608 339130 619642
rect 339196 619620 339228 619642
rect 339228 619620 339230 619642
rect 339296 619620 339318 619642
rect 339318 619620 339330 619642
rect 339396 619620 339408 619642
rect 339408 619620 339430 619642
rect 339196 619608 339230 619620
rect 339296 619608 339330 619620
rect 339396 619608 339430 619620
rect 338896 619530 338902 619542
rect 338902 619530 338930 619542
rect 338896 619508 338930 619530
rect 338996 619508 339030 619542
rect 339096 619508 339130 619542
rect 339196 619530 339228 619542
rect 339228 619530 339230 619542
rect 339296 619530 339318 619542
rect 339318 619530 339330 619542
rect 339396 619530 339408 619542
rect 339408 619530 339430 619542
rect 339196 619508 339230 619530
rect 339296 619508 339330 619530
rect 339396 619508 339430 619530
rect 338896 619440 338902 619442
rect 338902 619440 338930 619442
rect 338896 619408 338930 619440
rect 338996 619408 339030 619442
rect 339096 619408 339130 619442
rect 339196 619440 339228 619442
rect 339228 619440 339230 619442
rect 339296 619440 339318 619442
rect 339318 619440 339330 619442
rect 339396 619440 339408 619442
rect 339408 619440 339430 619442
rect 339196 619408 339230 619440
rect 339296 619408 339330 619440
rect 339396 619408 339430 619440
rect 338896 619308 338930 619342
rect 338996 619308 339030 619342
rect 339096 619308 339130 619342
rect 339196 619308 339230 619342
rect 339296 619308 339330 619342
rect 339396 619308 339430 619342
rect 338896 619208 338930 619242
rect 338996 619208 339030 619242
rect 339096 619208 339130 619242
rect 339196 619208 339230 619242
rect 339296 619208 339330 619242
rect 339396 619208 339430 619242
rect 338896 619114 338930 619142
rect 338896 619108 338902 619114
rect 338902 619108 338930 619114
rect 338996 619108 339030 619142
rect 339096 619108 339130 619142
rect 339196 619114 339230 619142
rect 339296 619114 339330 619142
rect 339396 619114 339430 619142
rect 339196 619108 339228 619114
rect 339228 619108 339230 619114
rect 339296 619108 339318 619114
rect 339318 619108 339330 619114
rect 339396 619108 339408 619114
rect 339408 619108 339430 619114
rect 340184 619620 340190 619642
rect 340190 619620 340218 619642
rect 340184 619608 340218 619620
rect 340284 619608 340318 619642
rect 340384 619608 340418 619642
rect 340484 619620 340516 619642
rect 340516 619620 340518 619642
rect 340584 619620 340606 619642
rect 340606 619620 340618 619642
rect 340684 619620 340696 619642
rect 340696 619620 340718 619642
rect 340484 619608 340518 619620
rect 340584 619608 340618 619620
rect 340684 619608 340718 619620
rect 340184 619530 340190 619542
rect 340190 619530 340218 619542
rect 340184 619508 340218 619530
rect 340284 619508 340318 619542
rect 340384 619508 340418 619542
rect 340484 619530 340516 619542
rect 340516 619530 340518 619542
rect 340584 619530 340606 619542
rect 340606 619530 340618 619542
rect 340684 619530 340696 619542
rect 340696 619530 340718 619542
rect 340484 619508 340518 619530
rect 340584 619508 340618 619530
rect 340684 619508 340718 619530
rect 340184 619440 340190 619442
rect 340190 619440 340218 619442
rect 340184 619408 340218 619440
rect 340284 619408 340318 619442
rect 340384 619408 340418 619442
rect 340484 619440 340516 619442
rect 340516 619440 340518 619442
rect 340584 619440 340606 619442
rect 340606 619440 340618 619442
rect 340684 619440 340696 619442
rect 340696 619440 340718 619442
rect 340484 619408 340518 619440
rect 340584 619408 340618 619440
rect 340684 619408 340718 619440
rect 340184 619308 340218 619342
rect 340284 619308 340318 619342
rect 340384 619308 340418 619342
rect 340484 619308 340518 619342
rect 340584 619308 340618 619342
rect 340684 619308 340718 619342
rect 340184 619208 340218 619242
rect 340284 619208 340318 619242
rect 340384 619208 340418 619242
rect 340484 619208 340518 619242
rect 340584 619208 340618 619242
rect 340684 619208 340718 619242
rect 340184 619114 340218 619142
rect 340184 619108 340190 619114
rect 340190 619108 340218 619114
rect 340284 619108 340318 619142
rect 340384 619108 340418 619142
rect 340484 619114 340518 619142
rect 340584 619114 340618 619142
rect 340684 619114 340718 619142
rect 340484 619108 340516 619114
rect 340516 619108 340518 619114
rect 340584 619108 340606 619114
rect 340606 619108 340618 619114
rect 340684 619108 340696 619114
rect 340696 619108 340718 619114
rect 335032 618332 335038 618354
rect 335038 618332 335066 618354
rect 335032 618320 335066 618332
rect 335132 618320 335166 618354
rect 335232 618320 335266 618354
rect 335332 618332 335364 618354
rect 335364 618332 335366 618354
rect 335432 618332 335454 618354
rect 335454 618332 335466 618354
rect 335532 618332 335544 618354
rect 335544 618332 335566 618354
rect 335332 618320 335366 618332
rect 335432 618320 335466 618332
rect 335532 618320 335566 618332
rect 335032 618242 335038 618254
rect 335038 618242 335066 618254
rect 335032 618220 335066 618242
rect 335132 618220 335166 618254
rect 335232 618220 335266 618254
rect 335332 618242 335364 618254
rect 335364 618242 335366 618254
rect 335432 618242 335454 618254
rect 335454 618242 335466 618254
rect 335532 618242 335544 618254
rect 335544 618242 335566 618254
rect 335332 618220 335366 618242
rect 335432 618220 335466 618242
rect 335532 618220 335566 618242
rect 335032 618152 335038 618154
rect 335038 618152 335066 618154
rect 335032 618120 335066 618152
rect 335132 618120 335166 618154
rect 335232 618120 335266 618154
rect 335332 618152 335364 618154
rect 335364 618152 335366 618154
rect 335432 618152 335454 618154
rect 335454 618152 335466 618154
rect 335532 618152 335544 618154
rect 335544 618152 335566 618154
rect 335332 618120 335366 618152
rect 335432 618120 335466 618152
rect 335532 618120 335566 618152
rect 335032 618020 335066 618054
rect 335132 618020 335166 618054
rect 335232 618020 335266 618054
rect 335332 618020 335366 618054
rect 335432 618020 335466 618054
rect 335532 618020 335566 618054
rect 335032 617920 335066 617954
rect 335132 617920 335166 617954
rect 335232 617920 335266 617954
rect 335332 617920 335366 617954
rect 335432 617920 335466 617954
rect 335532 617920 335566 617954
rect 335032 617826 335066 617854
rect 335032 617820 335038 617826
rect 335038 617820 335066 617826
rect 335132 617820 335166 617854
rect 335232 617820 335266 617854
rect 335332 617826 335366 617854
rect 335432 617826 335466 617854
rect 335532 617826 335566 617854
rect 335332 617820 335364 617826
rect 335364 617820 335366 617826
rect 335432 617820 335454 617826
rect 335454 617820 335466 617826
rect 335532 617820 335544 617826
rect 335544 617820 335566 617826
rect 336320 618332 336326 618354
rect 336326 618332 336354 618354
rect 336320 618320 336354 618332
rect 336420 618320 336454 618354
rect 336520 618320 336554 618354
rect 336620 618332 336652 618354
rect 336652 618332 336654 618354
rect 336720 618332 336742 618354
rect 336742 618332 336754 618354
rect 336820 618332 336832 618354
rect 336832 618332 336854 618354
rect 336620 618320 336654 618332
rect 336720 618320 336754 618332
rect 336820 618320 336854 618332
rect 336320 618242 336326 618254
rect 336326 618242 336354 618254
rect 336320 618220 336354 618242
rect 336420 618220 336454 618254
rect 336520 618220 336554 618254
rect 336620 618242 336652 618254
rect 336652 618242 336654 618254
rect 336720 618242 336742 618254
rect 336742 618242 336754 618254
rect 336820 618242 336832 618254
rect 336832 618242 336854 618254
rect 336620 618220 336654 618242
rect 336720 618220 336754 618242
rect 336820 618220 336854 618242
rect 336320 618152 336326 618154
rect 336326 618152 336354 618154
rect 336320 618120 336354 618152
rect 336420 618120 336454 618154
rect 336520 618120 336554 618154
rect 336620 618152 336652 618154
rect 336652 618152 336654 618154
rect 336720 618152 336742 618154
rect 336742 618152 336754 618154
rect 336820 618152 336832 618154
rect 336832 618152 336854 618154
rect 336620 618120 336654 618152
rect 336720 618120 336754 618152
rect 336820 618120 336854 618152
rect 336320 618020 336354 618054
rect 336420 618020 336454 618054
rect 336520 618020 336554 618054
rect 336620 618020 336654 618054
rect 336720 618020 336754 618054
rect 336820 618020 336854 618054
rect 336320 617920 336354 617954
rect 336420 617920 336454 617954
rect 336520 617920 336554 617954
rect 336620 617920 336654 617954
rect 336720 617920 336754 617954
rect 336820 617920 336854 617954
rect 336320 617826 336354 617854
rect 336320 617820 336326 617826
rect 336326 617820 336354 617826
rect 336420 617820 336454 617854
rect 336520 617820 336554 617854
rect 336620 617826 336654 617854
rect 336720 617826 336754 617854
rect 336820 617826 336854 617854
rect 336620 617820 336652 617826
rect 336652 617820 336654 617826
rect 336720 617820 336742 617826
rect 336742 617820 336754 617826
rect 336820 617820 336832 617826
rect 336832 617820 336854 617826
rect 337608 618332 337614 618354
rect 337614 618332 337642 618354
rect 337608 618320 337642 618332
rect 337708 618320 337742 618354
rect 337808 618320 337842 618354
rect 337908 618332 337940 618354
rect 337940 618332 337942 618354
rect 338008 618332 338030 618354
rect 338030 618332 338042 618354
rect 338108 618332 338120 618354
rect 338120 618332 338142 618354
rect 337908 618320 337942 618332
rect 338008 618320 338042 618332
rect 338108 618320 338142 618332
rect 337608 618242 337614 618254
rect 337614 618242 337642 618254
rect 337608 618220 337642 618242
rect 337708 618220 337742 618254
rect 337808 618220 337842 618254
rect 337908 618242 337940 618254
rect 337940 618242 337942 618254
rect 338008 618242 338030 618254
rect 338030 618242 338042 618254
rect 338108 618242 338120 618254
rect 338120 618242 338142 618254
rect 337908 618220 337942 618242
rect 338008 618220 338042 618242
rect 338108 618220 338142 618242
rect 337608 618152 337614 618154
rect 337614 618152 337642 618154
rect 337608 618120 337642 618152
rect 337708 618120 337742 618154
rect 337808 618120 337842 618154
rect 337908 618152 337940 618154
rect 337940 618152 337942 618154
rect 338008 618152 338030 618154
rect 338030 618152 338042 618154
rect 338108 618152 338120 618154
rect 338120 618152 338142 618154
rect 337908 618120 337942 618152
rect 338008 618120 338042 618152
rect 338108 618120 338142 618152
rect 337608 618020 337642 618054
rect 337708 618020 337742 618054
rect 337808 618020 337842 618054
rect 337908 618020 337942 618054
rect 338008 618020 338042 618054
rect 338108 618020 338142 618054
rect 337608 617920 337642 617954
rect 337708 617920 337742 617954
rect 337808 617920 337842 617954
rect 337908 617920 337942 617954
rect 338008 617920 338042 617954
rect 338108 617920 338142 617954
rect 337608 617826 337642 617854
rect 337608 617820 337614 617826
rect 337614 617820 337642 617826
rect 337708 617820 337742 617854
rect 337808 617820 337842 617854
rect 337908 617826 337942 617854
rect 338008 617826 338042 617854
rect 338108 617826 338142 617854
rect 337908 617820 337940 617826
rect 337940 617820 337942 617826
rect 338008 617820 338030 617826
rect 338030 617820 338042 617826
rect 338108 617820 338120 617826
rect 338120 617820 338142 617826
rect 338896 618332 338902 618354
rect 338902 618332 338930 618354
rect 338896 618320 338930 618332
rect 338996 618320 339030 618354
rect 339096 618320 339130 618354
rect 339196 618332 339228 618354
rect 339228 618332 339230 618354
rect 339296 618332 339318 618354
rect 339318 618332 339330 618354
rect 339396 618332 339408 618354
rect 339408 618332 339430 618354
rect 339196 618320 339230 618332
rect 339296 618320 339330 618332
rect 339396 618320 339430 618332
rect 338896 618242 338902 618254
rect 338902 618242 338930 618254
rect 338896 618220 338930 618242
rect 338996 618220 339030 618254
rect 339096 618220 339130 618254
rect 339196 618242 339228 618254
rect 339228 618242 339230 618254
rect 339296 618242 339318 618254
rect 339318 618242 339330 618254
rect 339396 618242 339408 618254
rect 339408 618242 339430 618254
rect 339196 618220 339230 618242
rect 339296 618220 339330 618242
rect 339396 618220 339430 618242
rect 338896 618152 338902 618154
rect 338902 618152 338930 618154
rect 338896 618120 338930 618152
rect 338996 618120 339030 618154
rect 339096 618120 339130 618154
rect 339196 618152 339228 618154
rect 339228 618152 339230 618154
rect 339296 618152 339318 618154
rect 339318 618152 339330 618154
rect 339396 618152 339408 618154
rect 339408 618152 339430 618154
rect 339196 618120 339230 618152
rect 339296 618120 339330 618152
rect 339396 618120 339430 618152
rect 338896 618020 338930 618054
rect 338996 618020 339030 618054
rect 339096 618020 339130 618054
rect 339196 618020 339230 618054
rect 339296 618020 339330 618054
rect 339396 618020 339430 618054
rect 338896 617920 338930 617954
rect 338996 617920 339030 617954
rect 339096 617920 339130 617954
rect 339196 617920 339230 617954
rect 339296 617920 339330 617954
rect 339396 617920 339430 617954
rect 338896 617826 338930 617854
rect 338896 617820 338902 617826
rect 338902 617820 338930 617826
rect 338996 617820 339030 617854
rect 339096 617820 339130 617854
rect 339196 617826 339230 617854
rect 339296 617826 339330 617854
rect 339396 617826 339430 617854
rect 339196 617820 339228 617826
rect 339228 617820 339230 617826
rect 339296 617820 339318 617826
rect 339318 617820 339330 617826
rect 339396 617820 339408 617826
rect 339408 617820 339430 617826
rect 340184 618332 340190 618354
rect 340190 618332 340218 618354
rect 340184 618320 340218 618332
rect 340284 618320 340318 618354
rect 340384 618320 340418 618354
rect 340484 618332 340516 618354
rect 340516 618332 340518 618354
rect 340584 618332 340606 618354
rect 340606 618332 340618 618354
rect 340684 618332 340696 618354
rect 340696 618332 340718 618354
rect 340484 618320 340518 618332
rect 340584 618320 340618 618332
rect 340684 618320 340718 618332
rect 340184 618242 340190 618254
rect 340190 618242 340218 618254
rect 340184 618220 340218 618242
rect 340284 618220 340318 618254
rect 340384 618220 340418 618254
rect 340484 618242 340516 618254
rect 340516 618242 340518 618254
rect 340584 618242 340606 618254
rect 340606 618242 340618 618254
rect 340684 618242 340696 618254
rect 340696 618242 340718 618254
rect 340484 618220 340518 618242
rect 340584 618220 340618 618242
rect 340684 618220 340718 618242
rect 340184 618152 340190 618154
rect 340190 618152 340218 618154
rect 340184 618120 340218 618152
rect 340284 618120 340318 618154
rect 340384 618120 340418 618154
rect 340484 618152 340516 618154
rect 340516 618152 340518 618154
rect 340584 618152 340606 618154
rect 340606 618152 340618 618154
rect 340684 618152 340696 618154
rect 340696 618152 340718 618154
rect 340484 618120 340518 618152
rect 340584 618120 340618 618152
rect 340684 618120 340718 618152
rect 340184 618020 340218 618054
rect 340284 618020 340318 618054
rect 340384 618020 340418 618054
rect 340484 618020 340518 618054
rect 340584 618020 340618 618054
rect 340684 618020 340718 618054
rect 340184 617920 340218 617954
rect 340284 617920 340318 617954
rect 340384 617920 340418 617954
rect 340484 617920 340518 617954
rect 340584 617920 340618 617954
rect 340684 617920 340718 617954
rect 340184 617826 340218 617854
rect 340184 617820 340190 617826
rect 340190 617820 340218 617826
rect 340284 617820 340318 617854
rect 340384 617820 340418 617854
rect 340484 617826 340518 617854
rect 340584 617826 340618 617854
rect 340684 617826 340718 617854
rect 340484 617820 340516 617826
rect 340516 617820 340518 617826
rect 340584 617820 340606 617826
rect 340606 617820 340618 617826
rect 340684 617820 340696 617826
rect 340696 617820 340718 617826
rect 330170 616606 330570 616706
rect 298876 615448 298976 615474
rect 299100 615448 299200 615474
rect 299324 615448 299424 615474
rect 299548 615448 299648 615474
rect 299772 615448 299872 615474
rect 299996 615448 300096 615474
rect 300220 615448 300320 615474
rect 300444 615448 300544 615474
rect 300668 615448 300768 615474
rect 300892 615448 300992 615474
rect 301116 615448 301216 615474
rect 301340 615448 301440 615474
rect 301564 615448 301664 615474
rect 301788 615448 301888 615474
rect 302012 615448 302112 615474
rect 302236 615448 302336 615474
rect 302460 615448 302560 615474
rect 302684 615448 302784 615474
rect 302908 615448 303008 615474
rect 303132 615448 303232 615474
rect 303356 615448 303456 615474
rect 303580 615448 303680 615474
rect 303804 615448 303904 615474
rect 304028 615448 304128 615474
rect 304252 615448 304352 615474
rect 304476 615448 304576 615474
rect 304700 615448 304800 615474
rect 304924 615448 305024 615474
rect 305148 615448 305248 615474
rect 305372 615448 305472 615474
rect 309346 615448 309446 615474
rect 309570 615448 309670 615474
rect 309794 615448 309894 615474
rect 310018 615448 310118 615474
rect 310242 615448 310342 615474
rect 310466 615448 310566 615474
rect 310690 615448 310790 615474
rect 310914 615448 311014 615474
rect 311138 615448 311238 615474
rect 311362 615448 311462 615474
rect 311586 615448 311686 615474
rect 311810 615448 311910 615474
rect 312034 615448 312134 615474
rect 312258 615448 312358 615474
rect 312482 615448 312582 615474
rect 312706 615448 312806 615474
rect 312930 615448 313030 615474
rect 313154 615448 313254 615474
rect 313378 615448 313478 615474
rect 313602 615448 313702 615474
rect 313826 615448 313926 615474
rect 314050 615448 314150 615474
rect 314274 615448 314374 615474
rect 314498 615448 314598 615474
rect 314722 615448 314822 615474
rect 314946 615448 315046 615474
rect 315170 615448 315270 615474
rect 315394 615448 315494 615474
rect 315618 615448 315718 615474
rect 315842 615448 315942 615474
rect 335616 615448 335716 615494
rect 335840 615448 335940 615494
rect 336064 615448 336164 615494
rect 336288 615448 336388 615494
rect 336512 615448 336612 615494
rect 336736 615448 336836 615494
rect 336960 615448 337060 615494
rect 337184 615448 337284 615494
rect 337408 615448 337508 615494
rect 337632 615448 337732 615494
rect 337856 615448 337956 615494
rect 338080 615448 338180 615494
rect 338304 615448 338404 615494
rect 338528 615448 338628 615494
rect 338752 615448 338852 615494
rect 338976 615448 339076 615494
rect 339200 615448 339300 615494
rect 339424 615448 339524 615494
rect 339648 615448 339748 615494
rect 339872 615448 339972 615494
rect 340096 615448 340196 615494
rect 340320 615448 340420 615494
rect 340544 615448 340644 615494
rect 340768 615448 340868 615494
rect 340992 615448 341092 615494
rect 298876 615374 298976 615448
rect 299100 615374 299200 615448
rect 299324 615374 299424 615448
rect 299548 615374 299648 615448
rect 299772 615374 299872 615448
rect 299996 615374 300096 615448
rect 300220 615374 300320 615448
rect 300444 615374 300544 615448
rect 300668 615374 300768 615448
rect 300892 615374 300992 615448
rect 301116 615374 301216 615448
rect 301340 615374 301440 615448
rect 301564 615374 301664 615448
rect 301788 615374 301888 615448
rect 302012 615374 302112 615448
rect 302236 615374 302336 615448
rect 302460 615374 302560 615448
rect 302684 615374 302784 615448
rect 302908 615374 303008 615448
rect 303132 615374 303232 615448
rect 303356 615374 303456 615448
rect 303580 615374 303680 615448
rect 303804 615374 303904 615448
rect 304028 615374 304128 615448
rect 304252 615374 304352 615448
rect 304476 615374 304576 615448
rect 304700 615374 304800 615448
rect 304924 615374 305024 615448
rect 305148 615374 305248 615448
rect 305372 615374 305472 615448
rect 309346 615374 309446 615448
rect 309570 615374 309670 615448
rect 309794 615374 309894 615448
rect 310018 615374 310118 615448
rect 310242 615374 310342 615448
rect 310466 615374 310566 615448
rect 310690 615374 310790 615448
rect 310914 615374 311014 615448
rect 311138 615374 311238 615448
rect 311362 615374 311462 615448
rect 311586 615374 311686 615448
rect 311810 615374 311910 615448
rect 312034 615374 312134 615448
rect 312258 615374 312358 615448
rect 312482 615374 312582 615448
rect 312706 615374 312806 615448
rect 312930 615374 313030 615448
rect 313154 615374 313254 615448
rect 313378 615374 313478 615448
rect 313602 615374 313702 615448
rect 313826 615374 313926 615448
rect 314050 615374 314150 615448
rect 314274 615374 314374 615448
rect 314498 615374 314598 615448
rect 314722 615374 314822 615448
rect 314946 615374 315046 615448
rect 315170 615374 315270 615448
rect 315394 615374 315494 615448
rect 315618 615374 315718 615448
rect 315842 615374 315942 615448
rect 335616 615394 335716 615448
rect 335840 615394 335940 615448
rect 336064 615394 336164 615448
rect 336288 615394 336388 615448
rect 336512 615394 336612 615448
rect 336736 615394 336836 615448
rect 336960 615394 337060 615448
rect 337184 615394 337284 615448
rect 337408 615394 337508 615448
rect 337632 615394 337732 615448
rect 337856 615394 337956 615448
rect 338080 615394 338180 615448
rect 338304 615394 338404 615448
rect 338528 615394 338628 615448
rect 338752 615394 338852 615448
rect 338976 615394 339076 615448
rect 339200 615394 339300 615448
rect 339424 615394 339524 615448
rect 339648 615394 339748 615448
rect 339872 615394 339972 615448
rect 340096 615394 340196 615448
rect 340320 615394 340420 615448
rect 340544 615394 340644 615448
rect 340768 615394 340868 615448
rect 340992 615394 341088 615448
rect 341088 615394 341092 615448
rect 341216 615394 341316 615494
rect 341440 615394 341540 615494
rect 341664 615394 341764 615494
rect 341888 615394 341988 615494
rect 342130 637896 342230 637996
rect 342354 637896 342454 637996
rect 342578 637896 342678 637996
rect 342802 637896 342902 637996
rect 343026 637896 343112 637996
rect 343112 637896 343126 637996
rect 342130 637672 342230 637772
rect 342354 637672 342454 637772
rect 342578 637672 342678 637772
rect 342802 637672 342902 637772
rect 343026 637672 343112 637772
rect 343112 637672 343126 637772
rect 342130 637448 342230 637548
rect 342354 637448 342454 637548
rect 342578 637448 342678 637548
rect 342802 637448 342902 637548
rect 343026 637448 343112 637548
rect 343112 637448 343126 637548
rect 342130 637224 342230 637324
rect 342354 637224 342454 637324
rect 342578 637224 342678 637324
rect 342802 637224 342902 637324
rect 343026 637224 343112 637324
rect 343112 637224 343126 637324
rect 342130 637000 342230 637100
rect 342354 637000 342454 637100
rect 342578 637000 342678 637100
rect 342802 637000 342902 637100
rect 343026 637000 343112 637100
rect 343112 637000 343126 637100
rect 342130 636776 342230 636876
rect 342354 636776 342454 636876
rect 342578 636776 342678 636876
rect 342802 636776 342902 636876
rect 343026 636776 343112 636876
rect 343112 636776 343126 636876
rect 342130 636552 342230 636652
rect 342354 636552 342454 636652
rect 342578 636552 342678 636652
rect 342802 636552 342902 636652
rect 343026 636552 343112 636652
rect 343112 636552 343126 636652
rect 342130 636328 342230 636428
rect 342354 636328 342454 636428
rect 342578 636328 342678 636428
rect 342802 636328 342902 636428
rect 343026 636328 343112 636428
rect 343112 636328 343126 636428
rect 342130 636104 342230 636204
rect 342354 636104 342454 636204
rect 342578 636104 342678 636204
rect 342802 636104 342902 636204
rect 343026 636104 343112 636204
rect 343112 636104 343126 636204
rect 342130 635880 342230 635980
rect 342354 635880 342454 635980
rect 342578 635880 342678 635980
rect 342802 635880 342902 635980
rect 343026 635880 343112 635980
rect 343112 635880 343126 635980
rect 342130 635656 342230 635756
rect 342354 635656 342454 635756
rect 342578 635656 342678 635756
rect 342802 635656 342902 635756
rect 343026 635656 343112 635756
rect 343112 635656 343126 635756
rect 342130 635432 342230 635532
rect 342354 635432 342454 635532
rect 342578 635432 342678 635532
rect 342802 635432 342902 635532
rect 343026 635432 343112 635532
rect 343112 635432 343126 635532
rect 342130 635208 342230 635308
rect 342354 635208 342454 635308
rect 342578 635208 342678 635308
rect 342802 635208 342902 635308
rect 343026 635208 343112 635308
rect 343112 635208 343126 635308
rect 342130 634984 342230 635084
rect 342354 634984 342454 635084
rect 342578 634984 342678 635084
rect 342802 634984 342902 635084
rect 343026 634984 343112 635084
rect 343112 634984 343126 635084
rect 342130 634760 342230 634860
rect 342354 634760 342454 634860
rect 342578 634760 342678 634860
rect 342802 634760 342902 634860
rect 343026 634760 343112 634860
rect 343112 634760 343126 634860
rect 342130 634536 342230 634636
rect 342354 634536 342454 634636
rect 342578 634536 342678 634636
rect 342802 634536 342902 634636
rect 343026 634536 343112 634636
rect 343112 634536 343126 634636
rect 342130 634312 342230 634412
rect 342354 634312 342454 634412
rect 342578 634312 342678 634412
rect 342802 634312 342902 634412
rect 343026 634312 343112 634412
rect 343112 634312 343126 634412
rect 342130 634088 342230 634188
rect 342354 634088 342454 634188
rect 342578 634088 342678 634188
rect 342802 634088 342902 634188
rect 343026 634088 343112 634188
rect 343112 634088 343126 634188
rect 342130 633864 342230 633964
rect 342354 633864 342454 633964
rect 342578 633864 342678 633964
rect 342802 633864 342902 633964
rect 343026 633864 343112 633964
rect 343112 633864 343126 633964
rect 342130 633640 342230 633740
rect 342354 633640 342454 633740
rect 342578 633640 342678 633740
rect 342802 633640 342902 633740
rect 343026 633640 343112 633740
rect 343112 633640 343126 633740
rect 342130 633416 342230 633516
rect 342354 633416 342454 633516
rect 342578 633416 342678 633516
rect 342802 633416 342902 633516
rect 343026 633416 343112 633516
rect 343112 633416 343126 633516
rect 342130 633192 342230 633292
rect 342354 633192 342454 633292
rect 342578 633192 342678 633292
rect 342802 633192 342902 633292
rect 343026 633192 343112 633292
rect 343112 633192 343126 633292
rect 342130 632968 342230 633068
rect 342354 632968 342454 633068
rect 342578 632968 342678 633068
rect 342802 632968 342902 633068
rect 343026 632968 343112 633068
rect 343112 632968 343126 633068
rect 342130 632744 342230 632844
rect 342354 632744 342454 632844
rect 342578 632744 342678 632844
rect 342802 632744 342902 632844
rect 343026 632744 343112 632844
rect 343112 632744 343126 632844
rect 342130 632520 342230 632620
rect 342354 632520 342454 632620
rect 342578 632520 342678 632620
rect 342802 632520 342902 632620
rect 343026 632520 343112 632620
rect 343112 632520 343126 632620
rect 342130 632296 342230 632396
rect 342354 632296 342454 632396
rect 342578 632296 342678 632396
rect 342802 632296 342902 632396
rect 343026 632296 343112 632396
rect 343112 632296 343126 632396
rect 342130 632072 342230 632172
rect 342354 632072 342454 632172
rect 342578 632072 342678 632172
rect 342802 632072 342902 632172
rect 343026 632072 343112 632172
rect 343112 632072 343126 632172
rect 342130 631848 342230 631948
rect 342354 631848 342454 631948
rect 342578 631848 342678 631948
rect 342802 631848 342902 631948
rect 343026 631848 343112 631948
rect 343112 631848 343126 631948
rect 342130 631624 342230 631724
rect 342354 631624 342454 631724
rect 342578 631624 342678 631724
rect 342802 631624 342902 631724
rect 343026 631624 343112 631724
rect 343112 631624 343126 631724
rect 342130 631400 342230 631500
rect 342354 631400 342454 631500
rect 342578 631400 342678 631500
rect 342802 631400 342902 631500
rect 343026 631400 343112 631500
rect 343112 631400 343126 631500
rect 342130 624496 342230 624596
rect 342354 624496 342454 624596
rect 342578 624496 342678 624596
rect 342802 624496 342902 624596
rect 343026 624496 343112 624596
rect 343112 624496 343126 624596
rect 342130 624272 342230 624372
rect 342354 624272 342454 624372
rect 342578 624272 342678 624372
rect 342802 624272 342902 624372
rect 343026 624272 343112 624372
rect 343112 624272 343126 624372
rect 342130 624048 342230 624148
rect 342354 624048 342454 624148
rect 342578 624048 342678 624148
rect 342802 624048 342902 624148
rect 343026 624048 343112 624148
rect 343112 624048 343126 624148
rect 342130 623824 342230 623924
rect 342354 623824 342454 623924
rect 342578 623824 342678 623924
rect 342802 623824 342902 623924
rect 343026 623824 343112 623924
rect 343112 623824 343126 623924
rect 342130 623600 342230 623700
rect 342354 623600 342454 623700
rect 342578 623600 342678 623700
rect 342802 623600 342902 623700
rect 343026 623600 343112 623700
rect 343112 623600 343126 623700
rect 342130 623376 342230 623476
rect 342354 623376 342454 623476
rect 342578 623376 342678 623476
rect 342802 623376 342902 623476
rect 343026 623376 343112 623476
rect 343112 623376 343126 623476
rect 342130 623152 342230 623252
rect 342354 623152 342454 623252
rect 342578 623152 342678 623252
rect 342802 623152 342902 623252
rect 343026 623152 343112 623252
rect 343112 623152 343126 623252
rect 342130 622928 342230 623028
rect 342354 622928 342454 623028
rect 342578 622928 342678 623028
rect 342802 622928 342902 623028
rect 343026 622928 343112 623028
rect 343112 622928 343126 623028
rect 342130 622704 342230 622804
rect 342354 622704 342454 622804
rect 342578 622704 342678 622804
rect 342802 622704 342902 622804
rect 343026 622704 343112 622804
rect 343112 622704 343126 622804
rect 342130 622480 342230 622580
rect 342354 622480 342454 622580
rect 342578 622480 342678 622580
rect 342802 622480 342902 622580
rect 343026 622480 343112 622580
rect 343112 622480 343126 622580
rect 342130 622256 342230 622356
rect 342354 622256 342454 622356
rect 342578 622256 342678 622356
rect 342802 622256 342902 622356
rect 343026 622256 343112 622356
rect 343112 622256 343126 622356
rect 342130 622032 342230 622132
rect 342354 622032 342454 622132
rect 342578 622032 342678 622132
rect 342802 622032 342902 622132
rect 343026 622032 343112 622132
rect 343112 622032 343126 622132
rect 342130 621808 342230 621908
rect 342354 621808 342454 621908
rect 342578 621808 342678 621908
rect 342802 621808 342902 621908
rect 343026 621808 343112 621908
rect 343112 621808 343126 621908
rect 342130 621584 342230 621684
rect 342354 621584 342454 621684
rect 342578 621584 342678 621684
rect 342802 621584 342902 621684
rect 343026 621584 343112 621684
rect 343112 621584 343126 621684
rect 342130 621360 342230 621460
rect 342354 621360 342454 621460
rect 342578 621360 342678 621460
rect 342802 621360 342902 621460
rect 343026 621360 343112 621460
rect 343112 621360 343126 621460
rect 342130 621136 342230 621236
rect 342354 621136 342454 621236
rect 342578 621136 342678 621236
rect 342802 621136 342902 621236
rect 343026 621136 343112 621236
rect 343112 621136 343126 621236
rect 342130 620912 342230 621012
rect 342354 620912 342454 621012
rect 342578 620912 342678 621012
rect 342802 620912 342902 621012
rect 343026 620912 343112 621012
rect 343112 620912 343126 621012
rect 342130 620688 342230 620788
rect 342354 620688 342454 620788
rect 342578 620688 342678 620788
rect 342802 620688 342902 620788
rect 343026 620688 343112 620788
rect 343112 620688 343126 620788
rect 342130 620464 342230 620564
rect 342354 620464 342454 620564
rect 342578 620464 342678 620564
rect 342802 620464 342902 620564
rect 343026 620464 343112 620564
rect 343112 620464 343126 620564
rect 342130 620240 342230 620340
rect 342354 620240 342454 620340
rect 342578 620240 342678 620340
rect 342802 620240 342902 620340
rect 343026 620240 343112 620340
rect 343112 620240 343126 620340
rect 342130 620016 342230 620116
rect 342354 620016 342454 620116
rect 342578 620016 342678 620116
rect 342802 620016 342902 620116
rect 343026 620016 343112 620116
rect 343112 620016 343126 620116
rect 342130 619792 342230 619892
rect 342354 619792 342454 619892
rect 342578 619792 342678 619892
rect 342802 619792 342902 619892
rect 343026 619792 343112 619892
rect 343112 619792 343126 619892
rect 342130 619568 342230 619668
rect 342354 619568 342454 619668
rect 342578 619568 342678 619668
rect 342802 619568 342902 619668
rect 343026 619568 343112 619668
rect 343112 619568 343126 619668
rect 342130 619344 342230 619444
rect 342354 619344 342454 619444
rect 342578 619344 342678 619444
rect 342802 619344 342902 619444
rect 343026 619344 343112 619444
rect 343112 619344 343126 619444
rect 342130 619120 342230 619220
rect 342354 619120 342454 619220
rect 342578 619120 342678 619220
rect 342802 619120 342902 619220
rect 343026 619120 343112 619220
rect 343112 619120 343126 619220
rect 342130 618896 342230 618996
rect 342354 618896 342454 618996
rect 342578 618896 342678 618996
rect 342802 618896 342902 618996
rect 343026 618896 343112 618996
rect 343112 618896 343126 618996
rect 342130 618672 342230 618772
rect 342354 618672 342454 618772
rect 342578 618672 342678 618772
rect 342802 618672 342902 618772
rect 343026 618672 343112 618772
rect 343112 618672 343126 618772
rect 342130 618448 342230 618548
rect 342354 618448 342454 618548
rect 342578 618448 342678 618548
rect 342802 618448 342902 618548
rect 343026 618448 343112 618548
rect 343112 618448 343126 618548
rect 342130 618224 342230 618324
rect 342354 618224 342454 618324
rect 342578 618224 342678 618324
rect 342802 618224 342902 618324
rect 343026 618224 343112 618324
rect 343112 618224 343126 618324
rect 342130 618000 342230 618100
rect 342354 618000 342454 618100
rect 342578 618000 342678 618100
rect 342802 618000 342902 618100
rect 343026 618000 343112 618100
rect 343112 618000 343126 618100
rect 342112 615394 342212 615494
rect 298876 615150 298976 615250
rect 299100 615150 299200 615250
rect 299324 615150 299424 615250
rect 299548 615150 299648 615250
rect 299772 615150 299872 615250
rect 299996 615150 300096 615250
rect 300220 615150 300320 615250
rect 300444 615150 300544 615250
rect 300668 615150 300768 615250
rect 300892 615150 300992 615250
rect 301116 615150 301216 615250
rect 301340 615150 301440 615250
rect 301564 615150 301664 615250
rect 301788 615150 301888 615250
rect 302012 615150 302112 615250
rect 302236 615150 302336 615250
rect 302460 615150 302560 615250
rect 302684 615150 302784 615250
rect 302908 615150 303008 615250
rect 303132 615150 303232 615250
rect 303356 615150 303456 615250
rect 303580 615150 303680 615250
rect 303804 615150 303904 615250
rect 304028 615150 304128 615250
rect 304252 615150 304352 615250
rect 304476 615150 304576 615250
rect 304700 615150 304800 615250
rect 304924 615150 305024 615250
rect 305148 615150 305248 615250
rect 305372 615150 305472 615250
rect 309346 615150 309446 615250
rect 309570 615150 309670 615250
rect 309794 615150 309894 615250
rect 310018 615150 310118 615250
rect 310242 615150 310342 615250
rect 310466 615150 310566 615250
rect 310690 615150 310790 615250
rect 310914 615150 311014 615250
rect 311138 615150 311238 615250
rect 311362 615150 311462 615250
rect 311586 615150 311686 615250
rect 311810 615150 311910 615250
rect 312034 615150 312134 615250
rect 312258 615150 312358 615250
rect 312482 615150 312582 615250
rect 312706 615150 312806 615250
rect 312930 615150 313030 615250
rect 313154 615150 313254 615250
rect 313378 615150 313478 615250
rect 313602 615150 313702 615250
rect 313826 615150 313926 615250
rect 314050 615150 314150 615250
rect 314274 615150 314374 615250
rect 314498 615150 314598 615250
rect 314722 615150 314822 615250
rect 314946 615150 315046 615250
rect 315170 615150 315270 615250
rect 315394 615150 315494 615250
rect 315618 615150 315718 615250
rect 315842 615150 315942 615250
rect 335616 615170 335716 615270
rect 335840 615170 335940 615270
rect 336064 615170 336164 615270
rect 336288 615170 336388 615270
rect 336512 615170 336612 615270
rect 336736 615170 336836 615270
rect 336960 615170 337060 615270
rect 337184 615170 337284 615270
rect 337408 615170 337508 615270
rect 337632 615170 337732 615270
rect 337856 615170 337956 615270
rect 338080 615170 338180 615270
rect 338304 615170 338404 615270
rect 338528 615170 338628 615270
rect 338752 615170 338852 615270
rect 338976 615170 339076 615270
rect 339200 615170 339300 615270
rect 339424 615170 339524 615270
rect 339648 615170 339748 615270
rect 339872 615170 339972 615270
rect 340096 615170 340196 615270
rect 340320 615170 340420 615270
rect 340544 615170 340644 615270
rect 340768 615170 340868 615270
rect 340992 615170 341088 615270
rect 341088 615170 341092 615270
rect 341216 615170 341316 615270
rect 341440 615170 341540 615270
rect 341664 615170 341764 615270
rect 341888 615170 341988 615270
rect 342112 615170 342212 615270
rect 298876 614926 298976 615026
rect 299100 614926 299200 615026
rect 299324 614926 299424 615026
rect 299548 614926 299648 615026
rect 299772 614926 299872 615026
rect 299996 614926 300096 615026
rect 300220 614926 300320 615026
rect 300444 614926 300544 615026
rect 300668 614926 300768 615026
rect 300892 614926 300992 615026
rect 301116 614926 301216 615026
rect 301340 614926 301440 615026
rect 301564 614926 301664 615026
rect 301788 614926 301888 615026
rect 302012 614926 302112 615026
rect 302236 614926 302336 615026
rect 302460 614926 302560 615026
rect 302684 614926 302784 615026
rect 302908 614926 303008 615026
rect 303132 614926 303232 615026
rect 303356 614926 303456 615026
rect 303580 614926 303680 615026
rect 303804 614926 303904 615026
rect 304028 614926 304128 615026
rect 304252 614926 304352 615026
rect 304476 614926 304576 615026
rect 304700 614926 304800 615026
rect 304924 614926 305024 615026
rect 305148 614926 305248 615026
rect 305372 614926 305472 615026
rect 309346 614926 309446 615026
rect 309570 614926 309670 615026
rect 309794 614926 309894 615026
rect 310018 614926 310118 615026
rect 310242 614926 310342 615026
rect 310466 614926 310566 615026
rect 310690 614926 310790 615026
rect 310914 614926 311014 615026
rect 311138 614926 311238 615026
rect 311362 614926 311462 615026
rect 311586 614926 311686 615026
rect 311810 614926 311910 615026
rect 312034 614926 312134 615026
rect 312258 614926 312358 615026
rect 312482 614926 312582 615026
rect 312706 614926 312806 615026
rect 312930 614926 313030 615026
rect 313154 614926 313254 615026
rect 313378 614926 313478 615026
rect 313602 614926 313702 615026
rect 313826 614926 313926 615026
rect 314050 614926 314150 615026
rect 314274 614926 314374 615026
rect 314498 614926 314598 615026
rect 314722 614926 314822 615026
rect 314946 614926 315046 615026
rect 315170 614926 315270 615026
rect 315394 614926 315494 615026
rect 315618 614926 315718 615026
rect 315842 614926 315942 615026
rect 335616 614946 335716 615046
rect 335840 614946 335940 615046
rect 336064 614946 336164 615046
rect 336288 614946 336388 615046
rect 336512 614946 336612 615046
rect 336736 614946 336836 615046
rect 336960 614946 337060 615046
rect 337184 614946 337284 615046
rect 337408 614946 337508 615046
rect 337632 614946 337732 615046
rect 337856 614946 337956 615046
rect 338080 614946 338180 615046
rect 338304 614946 338404 615046
rect 338528 614946 338628 615046
rect 338752 614946 338852 615046
rect 338976 614946 339076 615046
rect 339200 614946 339300 615046
rect 339424 614946 339524 615046
rect 339648 614946 339748 615046
rect 339872 614946 339972 615046
rect 340096 614946 340196 615046
rect 340320 614946 340420 615046
rect 340544 614946 340644 615046
rect 340768 614946 340868 615046
rect 340992 614946 341088 615046
rect 341088 614946 341092 615046
rect 341216 614946 341316 615046
rect 341440 614946 341540 615046
rect 341664 614946 341764 615046
rect 341888 614946 341988 615046
rect 342112 614946 342212 615046
rect 298876 614702 298976 614802
rect 299100 614702 299200 614802
rect 299324 614702 299424 614802
rect 299548 614702 299648 614802
rect 299772 614702 299872 614802
rect 299996 614702 300096 614802
rect 300220 614702 300320 614802
rect 300444 614702 300544 614802
rect 300668 614702 300768 614802
rect 300892 614702 300992 614802
rect 301116 614702 301216 614802
rect 301340 614702 301440 614802
rect 301564 614702 301664 614802
rect 301788 614702 301888 614802
rect 302012 614702 302112 614802
rect 302236 614702 302336 614802
rect 302460 614702 302560 614802
rect 302684 614702 302784 614802
rect 302908 614702 303008 614802
rect 303132 614702 303232 614802
rect 303356 614702 303456 614802
rect 303580 614702 303680 614802
rect 303804 614702 303904 614802
rect 304028 614702 304128 614802
rect 304252 614702 304352 614802
rect 304476 614702 304576 614802
rect 304700 614702 304800 614802
rect 304924 614702 305024 614802
rect 305148 614702 305248 614802
rect 305372 614702 305472 614802
rect 309346 614702 309446 614802
rect 309570 614702 309670 614802
rect 309794 614702 309894 614802
rect 310018 614702 310118 614802
rect 310242 614702 310342 614802
rect 310466 614702 310566 614802
rect 310690 614702 310790 614802
rect 310914 614702 311014 614802
rect 311138 614702 311238 614802
rect 311362 614702 311462 614802
rect 311586 614702 311686 614802
rect 311810 614702 311910 614802
rect 312034 614702 312134 614802
rect 312258 614702 312358 614802
rect 312482 614702 312582 614802
rect 312706 614702 312806 614802
rect 312930 614702 313030 614802
rect 313154 614702 313254 614802
rect 313378 614702 313478 614802
rect 313602 614702 313702 614802
rect 313826 614702 313926 614802
rect 314050 614702 314150 614802
rect 314274 614702 314374 614802
rect 314498 614702 314598 614802
rect 314722 614702 314822 614802
rect 314946 614702 315046 614802
rect 315170 614702 315270 614802
rect 315394 614702 315494 614802
rect 315618 614702 315718 614802
rect 315842 614702 315942 614802
rect 335616 614722 335716 614822
rect 335840 614722 335940 614822
rect 336064 614722 336164 614822
rect 336288 614722 336388 614822
rect 336512 614722 336612 614822
rect 336736 614722 336836 614822
rect 336960 614722 337060 614822
rect 337184 614722 337284 614822
rect 337408 614722 337508 614822
rect 337632 614722 337732 614822
rect 337856 614722 337956 614822
rect 338080 614722 338180 614822
rect 338304 614722 338404 614822
rect 338528 614722 338628 614822
rect 338752 614722 338852 614822
rect 338976 614722 339076 614822
rect 339200 614722 339300 614822
rect 339424 614722 339524 614822
rect 339648 614722 339748 614822
rect 339872 614722 339972 614822
rect 340096 614722 340196 614822
rect 340320 614722 340420 614822
rect 340544 614722 340644 614822
rect 340768 614722 340868 614822
rect 340992 614722 341088 614822
rect 341088 614722 341092 614822
rect 341216 614722 341316 614822
rect 341440 614722 341540 614822
rect 341664 614722 341764 614822
rect 341888 614722 341988 614822
rect 342112 614722 342212 614822
rect 298876 614478 298976 614578
rect 299100 614478 299200 614578
rect 299324 614478 299424 614578
rect 299548 614478 299648 614578
rect 299772 614478 299872 614578
rect 299996 614478 300096 614578
rect 300220 614478 300320 614578
rect 300444 614478 300544 614578
rect 300668 614478 300768 614578
rect 300892 614478 300992 614578
rect 301116 614478 301216 614578
rect 301340 614478 301440 614578
rect 301564 614478 301664 614578
rect 301788 614478 301888 614578
rect 302012 614478 302112 614578
rect 302236 614478 302336 614578
rect 302460 614478 302560 614578
rect 302684 614478 302784 614578
rect 302908 614478 303008 614578
rect 303132 614478 303232 614578
rect 303356 614478 303456 614578
rect 303580 614478 303680 614578
rect 303804 614478 303904 614578
rect 304028 614478 304128 614578
rect 304252 614478 304352 614578
rect 304476 614478 304576 614578
rect 304700 614478 304800 614578
rect 304924 614478 305024 614578
rect 305148 614478 305248 614578
rect 305372 614478 305472 614578
rect 309346 614478 309446 614578
rect 309570 614478 309670 614578
rect 309794 614478 309894 614578
rect 310018 614478 310118 614578
rect 310242 614478 310342 614578
rect 310466 614478 310566 614578
rect 310690 614478 310790 614578
rect 310914 614478 311014 614578
rect 311138 614478 311238 614578
rect 311362 614478 311462 614578
rect 311586 614478 311686 614578
rect 311810 614478 311910 614578
rect 312034 614478 312134 614578
rect 312258 614478 312358 614578
rect 312482 614478 312582 614578
rect 312706 614478 312806 614578
rect 312930 614478 313030 614578
rect 313154 614478 313254 614578
rect 313378 614478 313478 614578
rect 313602 614478 313702 614578
rect 313826 614478 313926 614578
rect 314050 614478 314150 614578
rect 314274 614478 314374 614578
rect 314498 614478 314598 614578
rect 314722 614478 314822 614578
rect 314946 614478 315046 614578
rect 315170 614478 315270 614578
rect 315394 614478 315494 614578
rect 315618 614478 315718 614578
rect 315842 614478 315942 614578
rect 335616 614498 335716 614598
rect 335840 614498 335940 614598
rect 336064 614498 336164 614598
rect 336288 614498 336388 614598
rect 336512 614498 336612 614598
rect 336736 614498 336836 614598
rect 336960 614498 337060 614598
rect 337184 614498 337284 614598
rect 337408 614498 337508 614598
rect 337632 614498 337732 614598
rect 337856 614498 337956 614598
rect 338080 614498 338180 614598
rect 338304 614498 338404 614598
rect 338528 614498 338628 614598
rect 338752 614498 338852 614598
rect 338976 614498 339076 614598
rect 339200 614498 339300 614598
rect 339424 614498 339524 614598
rect 339648 614498 339748 614598
rect 339872 614498 339972 614598
rect 340096 614498 340196 614598
rect 340320 614498 340420 614598
rect 340544 614498 340644 614598
rect 340768 614498 340868 614598
rect 340992 614498 341088 614598
rect 341088 614498 341092 614598
rect 341216 614498 341316 614598
rect 341440 614498 341540 614598
rect 341664 614498 341764 614598
rect 341888 614498 341988 614598
rect 342112 614498 342212 614598
<< metal1 >>
rect 298836 642694 305496 642724
rect 298836 642594 298876 642694
rect 298976 642594 299100 642694
rect 299200 642594 299324 642694
rect 299424 642594 299548 642694
rect 299648 642594 299772 642694
rect 299872 642594 299996 642694
rect 300096 642594 300220 642694
rect 300320 642594 300444 642694
rect 300544 642594 300668 642694
rect 300768 642594 300892 642694
rect 300992 642594 301116 642694
rect 301216 642594 301340 642694
rect 301440 642594 301564 642694
rect 301664 642594 301788 642694
rect 301888 642594 302012 642694
rect 302112 642594 302236 642694
rect 302336 642594 302460 642694
rect 302560 642594 302684 642694
rect 302784 642594 302908 642694
rect 303008 642594 303132 642694
rect 303232 642594 303356 642694
rect 303456 642594 303580 642694
rect 303680 642594 303804 642694
rect 303904 642594 304028 642694
rect 304128 642594 304252 642694
rect 304352 642594 304476 642694
rect 304576 642594 304700 642694
rect 304800 642594 304924 642694
rect 305024 642594 305148 642694
rect 305248 642594 305372 642694
rect 305472 642594 305496 642694
rect 298836 642470 305496 642594
rect 298836 642370 298876 642470
rect 298976 642370 299100 642470
rect 299200 642370 299324 642470
rect 299424 642370 299548 642470
rect 299648 642370 299772 642470
rect 299872 642370 299996 642470
rect 300096 642370 300220 642470
rect 300320 642370 300444 642470
rect 300544 642370 300668 642470
rect 300768 642370 300892 642470
rect 300992 642370 301116 642470
rect 301216 642370 301340 642470
rect 301440 642370 301564 642470
rect 301664 642370 301788 642470
rect 301888 642370 302012 642470
rect 302112 642370 302236 642470
rect 302336 642370 302460 642470
rect 302560 642370 302684 642470
rect 302784 642370 302908 642470
rect 303008 642370 303132 642470
rect 303232 642370 303356 642470
rect 303456 642370 303580 642470
rect 303680 642370 303804 642470
rect 303904 642370 304028 642470
rect 304128 642370 304252 642470
rect 304352 642370 304476 642470
rect 304576 642370 304700 642470
rect 304800 642370 304924 642470
rect 305024 642370 305148 642470
rect 305248 642370 305372 642470
rect 305472 642370 305496 642470
rect 298836 642246 305496 642370
rect 298836 642146 298876 642246
rect 298976 642146 299100 642246
rect 299200 642146 299324 642246
rect 299424 642146 299548 642246
rect 299648 642146 299772 642246
rect 299872 642146 299996 642246
rect 300096 642146 300220 642246
rect 300320 642146 300444 642246
rect 300544 642146 300668 642246
rect 300768 642146 300892 642246
rect 300992 642146 301116 642246
rect 301216 642146 301340 642246
rect 301440 642146 301564 642246
rect 301664 642146 301788 642246
rect 301888 642146 302012 642246
rect 302112 642146 302236 642246
rect 302336 642146 302460 642246
rect 302560 642146 302684 642246
rect 302784 642146 302908 642246
rect 303008 642146 303132 642246
rect 303232 642146 303356 642246
rect 303456 642146 303580 642246
rect 303680 642146 303804 642246
rect 303904 642146 304028 642246
rect 304128 642146 304252 642246
rect 304352 642146 304476 642246
rect 304576 642146 304700 642246
rect 304800 642146 304924 642246
rect 305024 642146 305148 642246
rect 305248 642146 305372 642246
rect 305472 642146 305496 642246
rect 298836 642022 305496 642146
rect 298836 641922 298876 642022
rect 298976 641922 299100 642022
rect 299200 641922 299324 642022
rect 299424 641922 299548 642022
rect 299648 641922 299772 642022
rect 299872 641922 299996 642022
rect 300096 641922 300220 642022
rect 300320 641922 300444 642022
rect 300544 641922 300668 642022
rect 300768 641922 300892 642022
rect 300992 641922 301116 642022
rect 301216 641922 301340 642022
rect 301440 641922 301564 642022
rect 301664 641922 301788 642022
rect 301888 641922 302012 642022
rect 302112 641922 302236 642022
rect 302336 641922 302460 642022
rect 302560 641922 302684 642022
rect 302784 641922 302908 642022
rect 303008 641922 303132 642022
rect 303232 641922 303356 642022
rect 303456 641922 303580 642022
rect 303680 641922 303804 642022
rect 303904 641922 304028 642022
rect 304128 641922 304252 642022
rect 304352 641922 304476 642022
rect 304576 641922 304700 642022
rect 304800 641922 304924 642022
rect 305024 641922 305148 642022
rect 305248 641922 305372 642022
rect 305472 641922 305496 642022
rect 298836 641798 305496 641922
rect 298836 641698 298876 641798
rect 298976 641698 299100 641798
rect 299200 641698 299324 641798
rect 299424 641698 299548 641798
rect 299648 641698 299772 641798
rect 299872 641698 299996 641798
rect 300096 641698 300220 641798
rect 300320 641698 300444 641798
rect 300544 641698 300668 641798
rect 300768 641698 300892 641798
rect 300992 641698 301116 641798
rect 301216 641698 301340 641798
rect 301440 641698 301564 641798
rect 301664 641698 301788 641798
rect 301888 641698 302012 641798
rect 302112 641698 302236 641798
rect 302336 641698 302460 641798
rect 302560 641698 302684 641798
rect 302784 641698 302908 641798
rect 303008 641698 303132 641798
rect 303232 641698 303356 641798
rect 303456 641698 303580 641798
rect 303680 641698 303804 641798
rect 303904 641698 304028 641798
rect 304128 641698 304252 641798
rect 304352 641698 304476 641798
rect 304576 641698 304700 641798
rect 304800 641698 304924 641798
rect 305024 641698 305148 641798
rect 305248 641698 305372 641798
rect 305472 641698 305496 641798
rect 298836 641664 305496 641698
rect 309306 642694 315966 642724
rect 309306 642594 309346 642694
rect 309446 642594 309570 642694
rect 309670 642594 309794 642694
rect 309894 642594 310018 642694
rect 310118 642594 310242 642694
rect 310342 642594 310466 642694
rect 310566 642594 310690 642694
rect 310790 642594 310914 642694
rect 311014 642594 311138 642694
rect 311238 642594 311362 642694
rect 311462 642594 311586 642694
rect 311686 642594 311810 642694
rect 311910 642594 312034 642694
rect 312134 642594 312258 642694
rect 312358 642594 312482 642694
rect 312582 642594 312706 642694
rect 312806 642594 312930 642694
rect 313030 642594 313154 642694
rect 313254 642594 313378 642694
rect 313478 642594 313602 642694
rect 313702 642594 313826 642694
rect 313926 642594 314050 642694
rect 314150 642594 314274 642694
rect 314374 642594 314498 642694
rect 314598 642594 314722 642694
rect 314822 642594 314946 642694
rect 315046 642594 315170 642694
rect 315270 642594 315394 642694
rect 315494 642594 315618 642694
rect 315718 642594 315842 642694
rect 315942 642594 315966 642694
rect 309306 642470 315966 642594
rect 309306 642370 309346 642470
rect 309446 642370 309570 642470
rect 309670 642370 309794 642470
rect 309894 642370 310018 642470
rect 310118 642370 310242 642470
rect 310342 642370 310466 642470
rect 310566 642370 310690 642470
rect 310790 642370 310914 642470
rect 311014 642370 311138 642470
rect 311238 642370 311362 642470
rect 311462 642370 311586 642470
rect 311686 642370 311810 642470
rect 311910 642370 312034 642470
rect 312134 642370 312258 642470
rect 312358 642370 312482 642470
rect 312582 642370 312706 642470
rect 312806 642370 312930 642470
rect 313030 642370 313154 642470
rect 313254 642370 313378 642470
rect 313478 642370 313602 642470
rect 313702 642370 313826 642470
rect 313926 642370 314050 642470
rect 314150 642370 314274 642470
rect 314374 642370 314498 642470
rect 314598 642370 314722 642470
rect 314822 642370 314946 642470
rect 315046 642370 315170 642470
rect 315270 642370 315394 642470
rect 315494 642370 315618 642470
rect 315718 642370 315842 642470
rect 315942 642370 315966 642470
rect 309306 642246 315966 642370
rect 309306 642146 309346 642246
rect 309446 642146 309570 642246
rect 309670 642146 309794 642246
rect 309894 642146 310018 642246
rect 310118 642146 310242 642246
rect 310342 642146 310466 642246
rect 310566 642146 310690 642246
rect 310790 642146 310914 642246
rect 311014 642146 311138 642246
rect 311238 642146 311362 642246
rect 311462 642146 311586 642246
rect 311686 642146 311810 642246
rect 311910 642146 312034 642246
rect 312134 642146 312258 642246
rect 312358 642146 312482 642246
rect 312582 642146 312706 642246
rect 312806 642146 312930 642246
rect 313030 642146 313154 642246
rect 313254 642146 313378 642246
rect 313478 642146 313602 642246
rect 313702 642146 313826 642246
rect 313926 642146 314050 642246
rect 314150 642146 314274 642246
rect 314374 642146 314498 642246
rect 314598 642146 314722 642246
rect 314822 642146 314946 642246
rect 315046 642146 315170 642246
rect 315270 642146 315394 642246
rect 315494 642146 315618 642246
rect 315718 642146 315842 642246
rect 315942 642146 315966 642246
rect 309306 642022 315966 642146
rect 309306 641922 309346 642022
rect 309446 641922 309570 642022
rect 309670 641922 309794 642022
rect 309894 641922 310018 642022
rect 310118 641922 310242 642022
rect 310342 641922 310466 642022
rect 310566 641922 310690 642022
rect 310790 641922 310914 642022
rect 311014 641922 311138 642022
rect 311238 641922 311362 642022
rect 311462 641922 311586 642022
rect 311686 641922 311810 642022
rect 311910 641922 312034 642022
rect 312134 641922 312258 642022
rect 312358 641922 312482 642022
rect 312582 641922 312706 642022
rect 312806 641922 312930 642022
rect 313030 641922 313154 642022
rect 313254 641922 313378 642022
rect 313478 641922 313602 642022
rect 313702 641922 313826 642022
rect 313926 641922 314050 642022
rect 314150 641922 314274 642022
rect 314374 641922 314498 642022
rect 314598 641922 314722 642022
rect 314822 641922 314946 642022
rect 315046 641922 315170 642022
rect 315270 641922 315394 642022
rect 315494 641922 315618 642022
rect 315718 641922 315842 642022
rect 315942 641922 315966 642022
rect 309306 641798 315966 641922
rect 309306 641698 309346 641798
rect 309446 641698 309570 641798
rect 309670 641698 309794 641798
rect 309894 641698 310018 641798
rect 310118 641698 310242 641798
rect 310342 641698 310466 641798
rect 310566 641698 310690 641798
rect 310790 641698 310914 641798
rect 311014 641698 311138 641798
rect 311238 641698 311362 641798
rect 311462 641698 311586 641798
rect 311686 641698 311810 641798
rect 311910 641698 312034 641798
rect 312134 641698 312258 641798
rect 312358 641698 312482 641798
rect 312582 641698 312706 641798
rect 312806 641698 312930 641798
rect 313030 641698 313154 641798
rect 313254 641698 313378 641798
rect 313478 641698 313602 641798
rect 313702 641698 313826 641798
rect 313926 641698 314050 641798
rect 314150 641698 314274 641798
rect 314374 641698 314498 641798
rect 314598 641698 314722 641798
rect 314822 641698 314946 641798
rect 315046 641698 315170 641798
rect 315270 641698 315394 641798
rect 315494 641698 315618 641798
rect 315718 641698 315842 641798
rect 315942 641698 315966 641798
rect 309306 641664 315966 641698
rect 335576 642714 342236 642744
rect 335576 642614 335616 642714
rect 335716 642614 335840 642714
rect 335940 642614 336064 642714
rect 336164 642614 336288 642714
rect 336388 642614 336512 642714
rect 336612 642614 336736 642714
rect 336836 642614 336960 642714
rect 337060 642614 337184 642714
rect 337284 642614 337408 642714
rect 337508 642614 337632 642714
rect 337732 642614 337856 642714
rect 337956 642614 338080 642714
rect 338180 642614 338304 642714
rect 338404 642614 338528 642714
rect 338628 642614 338752 642714
rect 338852 642614 338976 642714
rect 339076 642614 339200 642714
rect 339300 642614 339424 642714
rect 339524 642614 339648 642714
rect 339748 642614 339872 642714
rect 339972 642614 340096 642714
rect 340196 642614 340320 642714
rect 340420 642614 340544 642714
rect 340644 642614 340768 642714
rect 340868 642614 340992 642714
rect 341092 642614 341216 642714
rect 341316 642614 341440 642714
rect 341540 642614 341664 642714
rect 341764 642614 341888 642714
rect 341988 642614 342112 642714
rect 342212 642614 342236 642714
rect 335576 642490 342236 642614
rect 335576 642390 335616 642490
rect 335716 642390 335840 642490
rect 335940 642390 336064 642490
rect 336164 642390 336288 642490
rect 336388 642390 336512 642490
rect 336612 642390 336736 642490
rect 336836 642390 336960 642490
rect 337060 642390 337184 642490
rect 337284 642390 337408 642490
rect 337508 642390 337632 642490
rect 337732 642390 337856 642490
rect 337956 642390 338080 642490
rect 338180 642390 338304 642490
rect 338404 642390 338528 642490
rect 338628 642390 338752 642490
rect 338852 642390 338976 642490
rect 339076 642390 339200 642490
rect 339300 642390 339424 642490
rect 339524 642390 339648 642490
rect 339748 642390 339872 642490
rect 339972 642390 340096 642490
rect 340196 642390 340320 642490
rect 340420 642390 340544 642490
rect 340644 642390 340768 642490
rect 340868 642390 340992 642490
rect 341092 642390 341216 642490
rect 341316 642390 341440 642490
rect 341540 642390 341664 642490
rect 341764 642390 341888 642490
rect 341988 642390 342112 642490
rect 342212 642390 342236 642490
rect 335576 642266 342236 642390
rect 335576 642166 335616 642266
rect 335716 642166 335840 642266
rect 335940 642166 336064 642266
rect 336164 642166 336288 642266
rect 336388 642166 336512 642266
rect 336612 642166 336736 642266
rect 336836 642166 336960 642266
rect 337060 642166 337184 642266
rect 337284 642166 337408 642266
rect 337508 642166 337632 642266
rect 337732 642166 337856 642266
rect 337956 642166 338080 642266
rect 338180 642166 338304 642266
rect 338404 642166 338528 642266
rect 338628 642166 338752 642266
rect 338852 642166 338976 642266
rect 339076 642166 339200 642266
rect 339300 642166 339424 642266
rect 339524 642166 339648 642266
rect 339748 642166 339872 642266
rect 339972 642166 340096 642266
rect 340196 642166 340320 642266
rect 340420 642166 340544 642266
rect 340644 642166 340768 642266
rect 340868 642166 340992 642266
rect 341092 642166 341216 642266
rect 341316 642166 341440 642266
rect 341540 642166 341664 642266
rect 341764 642166 341888 642266
rect 341988 642166 342112 642266
rect 342212 642166 342236 642266
rect 335576 642042 342236 642166
rect 335576 641942 335616 642042
rect 335716 641942 335840 642042
rect 335940 641942 336064 642042
rect 336164 641942 336288 642042
rect 336388 641942 336512 642042
rect 336612 641942 336736 642042
rect 336836 641942 336960 642042
rect 337060 641942 337184 642042
rect 337284 641942 337408 642042
rect 337508 641942 337632 642042
rect 337732 641942 337856 642042
rect 337956 641942 338080 642042
rect 338180 641942 338304 642042
rect 338404 641942 338528 642042
rect 338628 641942 338752 642042
rect 338852 641942 338976 642042
rect 339076 641942 339200 642042
rect 339300 641942 339424 642042
rect 339524 641942 339648 642042
rect 339748 641942 339872 642042
rect 339972 641942 340096 642042
rect 340196 641942 340320 642042
rect 340420 641942 340544 642042
rect 340644 641942 340768 642042
rect 340868 641942 340992 642042
rect 341092 641942 341216 642042
rect 341316 641942 341440 642042
rect 341540 641942 341664 642042
rect 341764 641942 341888 642042
rect 341988 641942 342112 642042
rect 342212 641942 342236 642042
rect 335576 641818 342236 641942
rect 335576 641718 335616 641818
rect 335716 641718 335840 641818
rect 335940 641718 336064 641818
rect 336164 641718 336288 641818
rect 336388 641718 336512 641818
rect 336612 641718 336736 641818
rect 336836 641718 336960 641818
rect 337060 641718 337184 641818
rect 337284 641718 337408 641818
rect 337508 641718 337632 641818
rect 337732 641718 337856 641818
rect 337956 641718 338080 641818
rect 338180 641718 338304 641818
rect 338404 641718 338528 641818
rect 338628 641718 338752 641818
rect 338852 641718 338976 641818
rect 339076 641718 339200 641818
rect 339300 641718 339424 641818
rect 339524 641718 339648 641818
rect 339748 641718 339872 641818
rect 339972 641718 340096 641818
rect 340196 641718 340320 641818
rect 340420 641718 340544 641818
rect 340644 641718 340768 641818
rect 340868 641718 340992 641818
rect 341092 641718 341216 641818
rect 341316 641718 341440 641818
rect 341540 641718 341664 641818
rect 341764 641718 341888 641818
rect 341988 641718 342112 641818
rect 342212 641718 342236 641818
rect 335576 641684 342236 641718
rect 300652 640572 311908 640578
rect 300652 639746 300658 640572
rect 311902 639746 311908 640572
rect 300652 639740 311908 639746
rect 323918 639032 326112 639038
rect 323918 638474 323924 639032
rect 324482 638474 325548 639032
rect 326106 638474 326112 639032
rect 323918 638468 326112 638474
rect 329464 639032 332662 639038
rect 329464 638474 329638 639032
rect 330196 638474 332092 639032
rect 332650 638474 332662 639032
rect 329464 638468 332662 638474
rect 317362 638232 323658 638238
rect 297820 637996 298880 638020
rect 297820 637896 297850 637996
rect 297950 637896 298074 637996
rect 298174 637896 298298 637996
rect 298398 637896 298522 637996
rect 298622 637896 298746 637996
rect 298846 637896 298880 637996
rect 297820 637772 298880 637896
rect 297820 637672 297850 637772
rect 297950 637672 298074 637772
rect 298174 637672 298298 637772
rect 298398 637672 298522 637772
rect 298622 637672 298746 637772
rect 298846 637672 298880 637772
rect 297820 637548 298880 637672
rect 317362 637674 317368 638232
rect 317926 637674 323094 638232
rect 323652 637674 323658 638232
rect 317362 637668 323658 637674
rect 326238 638232 329384 638238
rect 326238 637674 326366 638232
rect 326924 637674 328820 638232
rect 329378 637674 329384 638232
rect 326238 637668 329384 637674
rect 331154 638232 334292 638238
rect 331154 637674 331274 638232
rect 331832 637674 333728 638232
rect 334286 637674 334292 638232
rect 331154 637668 334292 637674
rect 342100 637996 343160 638020
rect 342100 637896 342130 637996
rect 342230 637896 342354 637996
rect 342454 637896 342578 637996
rect 342678 637896 342802 637996
rect 342902 637896 343026 637996
rect 343126 637896 343160 637996
rect 342100 637772 343160 637896
rect 342100 637672 342130 637772
rect 342230 637672 342354 637772
rect 342454 637672 342578 637772
rect 342678 637672 342802 637772
rect 342902 637672 343026 637772
rect 343126 637672 343160 637772
rect 297820 637448 297850 637548
rect 297950 637448 298074 637548
rect 298174 637448 298298 637548
rect 298398 637448 298522 637548
rect 298622 637448 298746 637548
rect 298846 637448 298880 637548
rect 342100 637548 343160 637672
rect 317362 637494 317932 637500
rect 297820 637324 298880 637448
rect 297820 637224 297850 637324
rect 297950 637224 298074 637324
rect 298174 637224 298298 637324
rect 298398 637224 298522 637324
rect 298622 637224 298746 637324
rect 298846 637224 298880 637324
rect 297820 637100 298880 637224
rect 297820 637000 297850 637100
rect 297950 637000 298074 637100
rect 298174 637000 298298 637100
rect 298398 637000 298522 637100
rect 298622 637000 298746 637100
rect 298846 637000 298880 637100
rect 316548 637482 317110 637488
rect 316548 637085 316560 637482
rect 317098 637085 317110 637482
rect 316548 637079 317110 637085
rect 317362 637074 317368 637494
rect 317926 637074 317932 637494
rect 317362 637068 317932 637074
rect 318180 637494 318750 637500
rect 318180 637074 318186 637494
rect 318744 637074 318750 637494
rect 319002 637482 319564 637488
rect 319002 637085 319014 637482
rect 319552 637085 319564 637482
rect 342100 637448 342130 637548
rect 342230 637448 342354 637548
rect 342454 637448 342578 637548
rect 342678 637448 342802 637548
rect 342902 637448 343026 637548
rect 343126 637448 343160 637548
rect 322270 637432 322840 637438
rect 319002 637079 319564 637085
rect 321456 637420 322018 637426
rect 318180 637068 318750 637074
rect 321456 637023 321468 637420
rect 322006 637023 322018 637420
rect 321456 637017 322018 637023
rect 322270 637012 322276 637432
rect 322834 637012 322840 637432
rect 322270 637006 322840 637012
rect 323088 637432 323658 637438
rect 323088 637012 323094 637432
rect 323652 637012 323658 637432
rect 323088 637006 323658 637012
rect 323906 637432 324476 637438
rect 323906 637012 323912 637432
rect 324470 637012 324476 637432
rect 323906 637006 324476 637012
rect 324724 637432 325294 637438
rect 324724 637012 324730 637432
rect 325288 637012 325294 637432
rect 324724 637006 325294 637012
rect 325542 637432 326112 637438
rect 325542 637012 325548 637432
rect 326106 637012 326112 637432
rect 325542 637006 326112 637012
rect 326360 637432 326930 637438
rect 326360 637012 326366 637432
rect 326924 637012 326930 637432
rect 326360 637006 326930 637012
rect 327178 637432 327748 637438
rect 327178 637012 327184 637432
rect 327742 637012 327748 637432
rect 327178 637006 327748 637012
rect 327996 637432 328566 637438
rect 327996 637012 328002 637432
rect 328560 637012 328566 637432
rect 327996 637006 328566 637012
rect 328814 637432 329384 637438
rect 328814 637012 328820 637432
rect 329378 637012 329384 637432
rect 328814 637006 329384 637012
rect 329632 637432 330202 637438
rect 329632 637012 329638 637432
rect 330196 637012 330202 637432
rect 329632 637006 330202 637012
rect 330450 637432 331020 637438
rect 330450 637012 330456 637432
rect 331014 637012 331020 637432
rect 330450 637006 331020 637012
rect 331268 637432 331838 637438
rect 331268 637012 331274 637432
rect 331832 637012 331838 637432
rect 331268 637006 331838 637012
rect 332086 637432 332656 637438
rect 332086 637012 332092 637432
rect 332650 637012 332656 637432
rect 332086 637006 332656 637012
rect 332904 637432 333474 637438
rect 332904 637012 332910 637432
rect 333468 637012 333474 637432
rect 332904 637006 333474 637012
rect 333722 637432 334292 637438
rect 333722 637012 333728 637432
rect 334286 637012 334292 637432
rect 334544 637420 335106 637426
rect 334544 637023 334556 637420
rect 335094 637023 335106 637420
rect 334544 637017 335106 637023
rect 342100 637324 343160 637448
rect 342100 637224 342130 637324
rect 342230 637224 342354 637324
rect 342454 637224 342578 637324
rect 342678 637224 342802 637324
rect 342902 637224 343026 637324
rect 343126 637224 343160 637324
rect 342100 637100 343160 637224
rect 333722 637006 334292 637012
rect 297820 636876 298880 637000
rect 297820 636776 297850 636876
rect 297950 636776 298074 636876
rect 298174 636776 298298 636876
rect 298398 636776 298522 636876
rect 298622 636776 298746 636876
rect 298846 636776 298880 636876
rect 342100 637000 342130 637100
rect 342230 637000 342354 637100
rect 342454 637000 342578 637100
rect 342678 637000 342802 637100
rect 342902 637000 343026 637100
rect 343126 637000 343160 637100
rect 342100 636876 343160 637000
rect 342100 636776 342130 636876
rect 342230 636776 342354 636876
rect 342454 636776 342578 636876
rect 342678 636776 342802 636876
rect 342902 636776 343026 636876
rect 343126 636776 343160 636876
rect 297820 636652 298880 636776
rect 297820 636552 297850 636652
rect 297950 636552 298074 636652
rect 298174 636552 298298 636652
rect 298398 636552 298522 636652
rect 298622 636552 298746 636652
rect 298846 636552 298880 636652
rect 297820 636428 298880 636552
rect 297820 636328 297850 636428
rect 297950 636328 298074 636428
rect 298174 636328 298298 636428
rect 298398 636328 298522 636428
rect 298622 636328 298746 636428
rect 298846 636328 298880 636428
rect 297820 636204 298880 636328
rect 318178 636770 322840 636776
rect 318178 636278 318186 636770
rect 318744 636278 322276 636770
rect 318178 636212 322276 636278
rect 322834 636212 322840 636770
rect 318178 636206 322840 636212
rect 324724 636770 327748 636776
rect 324724 636212 324730 636770
rect 325288 636212 327184 636770
rect 327742 636212 327748 636770
rect 324724 636206 327748 636212
rect 330450 636770 333474 636776
rect 330450 636212 330456 636770
rect 331014 636212 332910 636770
rect 333468 636212 333474 636770
rect 330450 636206 333474 636212
rect 342100 636652 343160 636776
rect 342100 636552 342130 636652
rect 342230 636552 342354 636652
rect 342454 636552 342578 636652
rect 342678 636552 342802 636652
rect 342902 636552 343026 636652
rect 343126 636552 343160 636652
rect 342100 636428 343160 636552
rect 342100 636328 342130 636428
rect 342230 636328 342354 636428
rect 342454 636328 342578 636428
rect 342678 636328 342802 636428
rect 342902 636328 343026 636428
rect 343126 636328 343160 636428
rect 297820 636104 297850 636204
rect 297950 636104 298074 636204
rect 298174 636104 298298 636204
rect 298398 636104 298522 636204
rect 298622 636104 298746 636204
rect 298846 636104 298880 636204
rect 297820 635980 298880 636104
rect 342100 636204 343160 636328
rect 342100 636104 342130 636204
rect 342230 636104 342354 636204
rect 342454 636104 342578 636204
rect 342678 636104 342802 636204
rect 342902 636104 343026 636204
rect 343126 636104 343160 636204
rect 297820 635880 297850 635980
rect 297950 635880 298074 635980
rect 298174 635880 298298 635980
rect 298398 635880 298522 635980
rect 298622 635880 298746 635980
rect 298846 635880 298880 635980
rect 297820 635756 298880 635880
rect 297820 635656 297850 635756
rect 297950 635656 298074 635756
rect 298174 635656 298298 635756
rect 298398 635656 298522 635756
rect 298622 635656 298746 635756
rect 298846 635656 298880 635756
rect 313276 636096 313838 636102
rect 313276 635699 313288 636096
rect 313826 635699 313838 636096
rect 313276 635693 313838 635699
rect 314094 636096 314656 636102
rect 314094 635699 314106 636096
rect 314644 635699 314656 636096
rect 314094 635693 314656 635699
rect 314912 636096 315474 636102
rect 314912 635699 314924 636096
rect 315462 635699 315474 636096
rect 314912 635693 315474 635699
rect 342100 635980 343160 636104
rect 342100 635880 342130 635980
rect 342230 635880 342354 635980
rect 342454 635880 342578 635980
rect 342678 635880 342802 635980
rect 342902 635880 343026 635980
rect 343126 635880 343160 635980
rect 342100 635756 343160 635880
rect 297820 635532 298880 635656
rect 297820 635432 297850 635532
rect 297950 635432 298074 635532
rect 298174 635432 298298 635532
rect 298398 635432 298522 635532
rect 298622 635432 298746 635532
rect 298846 635432 298880 635532
rect 297820 635308 298880 635432
rect 297820 635208 297850 635308
rect 297950 635208 298074 635308
rect 298174 635208 298298 635308
rect 298398 635208 298522 635308
rect 298622 635208 298746 635308
rect 298846 635208 298880 635308
rect 297820 635084 298880 635208
rect 297820 634984 297850 635084
rect 297950 634984 298074 635084
rect 298174 634984 298298 635084
rect 298398 634984 298522 635084
rect 298622 634984 298746 635084
rect 298846 634984 298880 635084
rect 297820 634860 298880 634984
rect 297820 634760 297850 634860
rect 297950 634760 298074 634860
rect 298174 634760 298298 634860
rect 298398 634760 298522 634860
rect 298622 634760 298746 634860
rect 298846 634760 298880 634860
rect 297820 634636 298880 634760
rect 297820 634536 297850 634636
rect 297950 634536 298074 634636
rect 298174 634536 298298 634636
rect 298398 634536 298522 634636
rect 298622 634536 298746 634636
rect 298846 634536 298880 634636
rect 297820 634412 298880 634536
rect 297820 634312 297850 634412
rect 297950 634312 298074 634412
rect 298174 634312 298298 634412
rect 298398 634312 298522 634412
rect 298622 634312 298746 634412
rect 298846 634312 298880 634412
rect 297820 634188 298880 634312
rect 297820 634088 297850 634188
rect 297950 634088 298074 634188
rect 298174 634088 298298 634188
rect 298398 634088 298522 634188
rect 298622 634088 298746 634188
rect 298846 634088 298880 634188
rect 297820 633964 298880 634088
rect 297820 633864 297850 633964
rect 297950 633864 298074 633964
rect 298174 633864 298298 633964
rect 298398 633864 298522 633964
rect 298622 633864 298746 633964
rect 298846 633864 298880 633964
rect 297820 633740 298880 633864
rect 297820 633640 297850 633740
rect 297950 633640 298074 633740
rect 298174 633640 298298 633740
rect 298398 633640 298522 633740
rect 298622 633640 298746 633740
rect 298846 633640 298880 633740
rect 297820 633516 298880 633640
rect 297820 633416 297850 633516
rect 297950 633416 298074 633516
rect 298174 633416 298298 633516
rect 298398 633416 298522 633516
rect 298622 633416 298746 633516
rect 298846 633416 298880 633516
rect 297820 633292 298880 633416
rect 297820 633192 297850 633292
rect 297950 633192 298074 633292
rect 298174 633192 298298 633292
rect 298398 633192 298522 633292
rect 298622 633192 298746 633292
rect 298846 633192 298880 633292
rect 297820 633068 298880 633192
rect 297820 632968 297850 633068
rect 297950 632968 298074 633068
rect 298174 632968 298298 633068
rect 298398 632968 298522 633068
rect 298622 632968 298746 633068
rect 298846 632968 298880 633068
rect 297820 632844 298880 632968
rect 297820 632744 297850 632844
rect 297950 632744 298074 632844
rect 298174 632744 298298 632844
rect 298398 632744 298522 632844
rect 298622 632744 298746 632844
rect 298846 632744 298880 632844
rect 342100 635656 342130 635756
rect 342230 635656 342354 635756
rect 342454 635656 342578 635756
rect 342678 635656 342802 635756
rect 342902 635656 343026 635756
rect 343126 635656 343160 635756
rect 342100 635532 343160 635656
rect 342100 635432 342130 635532
rect 342230 635432 342354 635532
rect 342454 635432 342578 635532
rect 342678 635432 342802 635532
rect 342902 635432 343026 635532
rect 343126 635432 343160 635532
rect 342100 635308 343160 635432
rect 342100 635208 342130 635308
rect 342230 635208 342354 635308
rect 342454 635208 342578 635308
rect 342678 635208 342802 635308
rect 342902 635208 343026 635308
rect 343126 635208 343160 635308
rect 342100 635084 343160 635208
rect 342100 634984 342130 635084
rect 342230 634984 342354 635084
rect 342454 634984 342578 635084
rect 342678 634984 342802 635084
rect 342902 634984 343026 635084
rect 343126 634984 343160 635084
rect 342100 634860 343160 634984
rect 342100 634760 342130 634860
rect 342230 634760 342354 634860
rect 342454 634760 342578 634860
rect 342678 634760 342802 634860
rect 342902 634760 343026 634860
rect 343126 634760 343160 634860
rect 342100 634636 343160 634760
rect 342100 634536 342130 634636
rect 342230 634536 342354 634636
rect 342454 634536 342578 634636
rect 342678 634536 342802 634636
rect 342902 634536 343026 634636
rect 343126 634536 343160 634636
rect 342100 634412 343160 634536
rect 342100 634312 342130 634412
rect 342230 634312 342354 634412
rect 342454 634312 342578 634412
rect 342678 634312 342802 634412
rect 342902 634312 343026 634412
rect 343126 634312 343160 634412
rect 342100 634188 343160 634312
rect 342100 634088 342130 634188
rect 342230 634088 342354 634188
rect 342454 634088 342578 634188
rect 342678 634088 342802 634188
rect 342902 634088 343026 634188
rect 343126 634088 343160 634188
rect 342100 633964 343160 634088
rect 342100 633864 342130 633964
rect 342230 633864 342354 633964
rect 342454 633864 342578 633964
rect 342678 633864 342802 633964
rect 342902 633864 343026 633964
rect 343126 633864 343160 633964
rect 342100 633740 343160 633864
rect 342100 633640 342130 633740
rect 342230 633640 342354 633740
rect 342454 633640 342578 633740
rect 342678 633640 342802 633740
rect 342902 633640 343026 633740
rect 343126 633640 343160 633740
rect 342100 633516 343160 633640
rect 342100 633416 342130 633516
rect 342230 633416 342354 633516
rect 342454 633416 342578 633516
rect 342678 633416 342802 633516
rect 342902 633416 343026 633516
rect 343126 633416 343160 633516
rect 342100 633292 343160 633416
rect 342100 633192 342130 633292
rect 342230 633192 342354 633292
rect 342454 633192 342578 633292
rect 342678 633192 342802 633292
rect 342902 633192 343026 633292
rect 343126 633192 343160 633292
rect 342100 633068 343160 633192
rect 342100 632968 342130 633068
rect 342230 632968 342354 633068
rect 342454 632968 342578 633068
rect 342678 632968 342802 633068
rect 342902 632968 343026 633068
rect 343126 632968 343160 633068
rect 342100 632844 343160 632968
rect 297820 632620 298880 632744
rect 297820 632520 297850 632620
rect 297950 632520 298074 632620
rect 298174 632520 298298 632620
rect 298398 632520 298522 632620
rect 298622 632520 298746 632620
rect 298846 632520 298880 632620
rect 297820 632396 298880 632520
rect 297820 632296 297850 632396
rect 297950 632296 298074 632396
rect 298174 632296 298298 632396
rect 298398 632296 298522 632396
rect 298622 632296 298746 632396
rect 298846 632296 298880 632396
rect 315722 632751 321218 632768
rect 315722 632740 316560 632751
rect 297820 632172 298880 632296
rect 297820 632072 297850 632172
rect 297950 632072 298074 632172
rect 298174 632072 298298 632172
rect 298398 632072 298522 632172
rect 298622 632072 298746 632172
rect 298846 632072 298880 632172
rect 297820 631948 298880 632072
rect 297820 631848 297850 631948
rect 297950 631848 298074 631948
rect 298174 631848 298298 631948
rect 298398 631848 298522 631948
rect 298622 631848 298746 631948
rect 298846 631848 298880 631948
rect 313276 632341 313838 632347
rect 313276 631944 313288 632341
rect 313826 631944 313838 632341
rect 313276 631938 313838 631944
rect 314090 632341 314660 632358
rect 314090 631944 314106 632341
rect 314644 631944 314660 632341
rect 297820 631724 298880 631848
rect 297820 631624 297850 631724
rect 297950 631624 298074 631724
rect 298174 631624 298298 631724
rect 298398 631624 298522 631724
rect 298622 631624 298746 631724
rect 298846 631624 298880 631724
rect 297820 631500 298880 631624
rect 297820 631400 297850 631500
rect 297950 631400 298074 631500
rect 298174 631400 298298 631500
rect 298398 631400 298522 631500
rect 298622 631400 298746 631500
rect 298846 631400 298880 631500
rect 297820 631360 298880 631400
rect 314090 631502 314660 631944
rect 314912 632341 315474 632347
rect 314912 631944 314924 632341
rect 315462 631944 315474 632341
rect 314912 631938 315474 631944
rect 315722 631674 315744 632740
rect 316238 632354 316560 632740
rect 317098 632354 317378 632751
rect 317916 632354 318196 632751
rect 318734 632354 319014 632751
rect 319552 632738 321218 632751
rect 319552 632354 320696 632738
rect 316238 631686 320696 632354
rect 321208 631686 321218 632738
rect 342100 632744 342130 632844
rect 342230 632744 342354 632844
rect 342454 632744 342578 632844
rect 342678 632744 342802 632844
rect 342902 632744 343026 632844
rect 343126 632744 343160 632844
rect 342100 632620 343160 632744
rect 342100 632520 342130 632620
rect 342230 632520 342354 632620
rect 342454 632520 342578 632620
rect 342678 632520 342802 632620
rect 342902 632520 343026 632620
rect 343126 632520 343160 632620
rect 342100 632396 343160 632520
rect 323088 632296 326930 632302
rect 323088 631738 323094 632296
rect 323652 631738 326366 632296
rect 326924 631738 326930 632296
rect 323088 631732 326930 631738
rect 328820 632296 331838 632302
rect 329378 631738 331274 632296
rect 331832 631738 331838 632296
rect 328820 631732 331838 631738
rect 342100 632296 342130 632396
rect 342230 632296 342354 632396
rect 342454 632296 342578 632396
rect 342678 632296 342802 632396
rect 342902 632296 343026 632396
rect 343126 632296 343160 632396
rect 342100 632172 343160 632296
rect 342100 632072 342130 632172
rect 342230 632072 342354 632172
rect 342454 632072 342578 632172
rect 342678 632072 342802 632172
rect 342902 632072 343026 632172
rect 343126 632072 343160 632172
rect 342100 631948 343160 632072
rect 342100 631848 342130 631948
rect 342230 631848 342354 631948
rect 342454 631848 342578 631948
rect 342678 631848 342802 631948
rect 342902 631848 343026 631948
rect 343126 631848 343160 631948
rect 316238 631674 321218 631686
rect 315722 631632 321218 631674
rect 342100 631724 343160 631848
rect 342100 631624 342130 631724
rect 342230 631624 342354 631724
rect 342454 631624 342578 631724
rect 342678 631624 342802 631724
rect 342902 631624 343026 631724
rect 343126 631624 343160 631724
rect 314090 631496 324476 631502
rect 314090 630938 323912 631496
rect 324470 630938 324476 631496
rect 314090 630932 324476 630938
rect 325542 631496 330202 631502
rect 325542 630938 325548 631496
rect 326106 630938 329638 631496
rect 330196 630938 330202 631496
rect 342100 631500 343160 631624
rect 342100 631400 342130 631500
rect 342230 631400 342354 631500
rect 342454 631400 342578 631500
rect 342678 631400 342802 631500
rect 342902 631400 343026 631500
rect 343126 631400 343160 631500
rect 342100 631360 343160 631400
rect 325542 630932 330202 630938
rect 322270 630696 322840 630702
rect 321456 630685 322018 630691
rect 321456 630288 321468 630685
rect 322006 630288 322018 630685
rect 321456 630282 322018 630288
rect 322270 630276 322276 630696
rect 322834 630276 322840 630696
rect 322270 630270 322840 630276
rect 323088 630696 323658 630702
rect 323088 630276 323094 630696
rect 323652 630276 323658 630696
rect 323088 630270 323658 630276
rect 323906 630696 324476 630702
rect 323906 630276 323912 630696
rect 324470 630276 324476 630696
rect 323906 630270 324476 630276
rect 324724 630696 325294 630702
rect 324724 630276 324730 630696
rect 325288 630276 325294 630696
rect 324724 630270 325294 630276
rect 325542 630696 326112 630702
rect 325542 630276 325548 630696
rect 326106 630276 326112 630696
rect 325542 630270 326112 630276
rect 326360 630696 326930 630702
rect 326360 630276 326366 630696
rect 326924 630276 326930 630696
rect 326360 630270 326930 630276
rect 327178 630696 327748 630702
rect 327178 630276 327184 630696
rect 327742 630276 327748 630696
rect 327178 630270 327748 630276
rect 327918 630696 328622 630702
rect 327918 630664 328002 630696
rect 327918 630146 327924 630664
rect 328560 630664 328622 630696
rect 328616 630146 328622 630664
rect 328814 630696 329384 630702
rect 328814 630276 328820 630696
rect 329378 630276 329384 630696
rect 328814 630270 329384 630276
rect 329632 630696 330202 630702
rect 329632 630276 329638 630696
rect 330196 630276 330202 630696
rect 329632 630270 330202 630276
rect 330450 630696 331020 630702
rect 330450 630276 330456 630696
rect 331014 630276 331020 630696
rect 330450 630270 331020 630276
rect 331268 630696 331838 630702
rect 331268 630276 331274 630696
rect 331832 630276 331838 630696
rect 331268 630270 331838 630276
rect 332008 630696 332712 630702
rect 322270 630034 325294 630040
rect 322270 629476 322276 630034
rect 322834 629476 324730 630034
rect 325288 629476 325294 630034
rect 322270 629470 325294 629476
rect 327178 630034 331020 630040
rect 327178 629476 327184 630034
rect 327742 629476 330456 630034
rect 331014 629476 331020 630034
rect 327178 629470 331020 629476
rect 332008 630004 332014 630696
rect 332706 630004 332712 630696
rect 332008 629006 332712 630004
rect 319314 628868 332712 629006
rect 319314 628668 319400 628868
rect 319600 628668 319834 628868
rect 320034 628668 320268 628868
rect 320468 628668 320702 628868
rect 320902 628668 321136 628868
rect 321336 628668 321570 628868
rect 321770 628668 322004 628868
rect 322204 628668 322438 628868
rect 322638 628668 322872 628868
rect 323072 628668 323306 628868
rect 323506 628668 323740 628868
rect 323940 628668 324140 628868
rect 324340 628668 324540 628868
rect 324740 628668 324940 628868
rect 325140 628668 325340 628868
rect 325540 628668 325740 628868
rect 325940 628668 326140 628868
rect 326340 628668 326540 628868
rect 326740 628668 326940 628868
rect 327140 628668 327340 628868
rect 327540 628668 328940 628868
rect 329140 628668 329340 628868
rect 329540 628668 329740 628868
rect 329940 628668 330140 628868
rect 330340 628668 330540 628868
rect 330740 628668 330940 628868
rect 331140 628668 331340 628868
rect 331540 628668 331740 628868
rect 331940 628668 332140 628868
rect 332340 628668 332712 628868
rect 319314 628434 332712 628668
rect 319314 628234 319400 628434
rect 319600 628234 319834 628434
rect 320034 628234 320268 628434
rect 320468 628234 320702 628434
rect 320902 628234 321136 628434
rect 321336 628234 321570 628434
rect 321770 628234 322004 628434
rect 322204 628234 322438 628434
rect 322638 628234 322872 628434
rect 323072 628234 323306 628434
rect 323506 628234 323740 628434
rect 323940 628314 332712 628434
rect 332826 630696 333530 630702
rect 332826 630004 332832 630696
rect 333524 630004 333530 630696
rect 323940 628234 324014 628314
rect 319314 628000 324014 628234
rect 319314 627800 319400 628000
rect 319600 627800 319834 628000
rect 320034 627800 320268 628000
rect 320468 627800 320702 628000
rect 320902 627800 321136 628000
rect 321336 627800 321570 628000
rect 321770 627800 322004 628000
rect 322204 627800 322438 628000
rect 322638 627800 322872 628000
rect 323072 627800 323306 628000
rect 323506 627800 323740 628000
rect 323940 627800 324014 628000
rect 313814 627366 315814 627408
rect 313814 626916 313820 627366
rect 315808 626916 315814 627366
rect 312296 626610 312428 626616
rect 312296 626196 312302 626610
rect 312422 626196 312428 626610
rect 311840 625904 311972 626190
rect 311840 625612 311846 625904
rect 311966 625612 311972 625904
rect 304304 624894 310792 624906
rect 297820 624596 298878 624606
rect 297820 624496 297850 624596
rect 297950 624496 298074 624596
rect 298174 624496 298298 624596
rect 298398 624496 298522 624596
rect 298622 624496 298746 624596
rect 298846 624496 298878 624596
rect 297820 624372 298878 624496
rect 297820 624272 297850 624372
rect 297950 624272 298074 624372
rect 298174 624272 298298 624372
rect 298398 624272 298522 624372
rect 298622 624272 298746 624372
rect 298846 624272 298878 624372
rect 304304 624550 304316 624894
rect 310780 624550 310792 624894
rect 304304 624358 310792 624550
rect 304304 624338 305040 624358
rect 305028 624324 305040 624338
rect 310416 624338 310792 624358
rect 310416 624324 310428 624338
rect 305028 624318 310428 624324
rect 297820 624148 298878 624272
rect 297820 624048 297850 624148
rect 297950 624048 298074 624148
rect 298174 624048 298298 624148
rect 298398 624048 298522 624148
rect 298622 624048 298746 624148
rect 298846 624048 298878 624148
rect 297820 623924 298878 624048
rect 302950 624204 304996 624216
rect 302950 624184 304956 624204
rect 302950 624114 302972 624184
rect 303032 624114 303044 624184
rect 303104 624114 303116 624184
rect 303176 624114 303188 624184
rect 303248 624114 303260 624184
rect 303320 624114 303332 624184
rect 303392 624114 303404 624184
rect 303464 624114 303476 624184
rect 303536 624114 304956 624184
rect 302950 624090 304956 624114
rect 302950 624020 302972 624090
rect 303032 624020 303044 624090
rect 303104 624020 303116 624090
rect 303176 624020 303188 624090
rect 303248 624020 303260 624090
rect 303320 624020 303332 624090
rect 303392 624020 303404 624090
rect 303464 624020 303476 624090
rect 303536 624020 304956 624090
rect 304990 624020 304996 624204
rect 302950 624008 304996 624020
rect 297820 623824 297850 623924
rect 297950 623824 298074 623924
rect 298174 623824 298298 623924
rect 298398 623824 298522 623924
rect 298622 623824 298746 623924
rect 298846 623824 298878 623924
rect 305028 623900 310428 623906
rect 297820 623700 298878 623824
rect 297820 623600 297850 623700
rect 297950 623600 298074 623700
rect 298174 623600 298298 623700
rect 298398 623600 298522 623700
rect 298622 623600 298746 623700
rect 298846 623600 298878 623700
rect 297820 623476 298878 623600
rect 297820 623376 297850 623476
rect 297950 623376 298074 623476
rect 298174 623376 298298 623476
rect 298398 623376 298522 623476
rect 298622 623376 298746 623476
rect 298846 623376 298878 623476
rect 297820 623252 298878 623376
rect 297820 623152 297850 623252
rect 297950 623152 298074 623252
rect 298174 623152 298298 623252
rect 298398 623152 298522 623252
rect 298622 623152 298746 623252
rect 298846 623152 298878 623252
rect 297820 623028 298878 623152
rect 297820 622928 297850 623028
rect 297950 622928 298074 623028
rect 298174 622928 298298 623028
rect 298398 622928 298522 623028
rect 298622 622928 298746 623028
rect 298846 622928 298878 623028
rect 297820 622804 298878 622928
rect 297820 622704 297850 622804
rect 297950 622704 298074 622804
rect 298174 622704 298298 622804
rect 298398 622704 298522 622804
rect 298622 622704 298746 622804
rect 298846 622704 298878 622804
rect 297820 622580 298878 622704
rect 297820 622480 297850 622580
rect 297950 622480 298074 622580
rect 298174 622480 298298 622580
rect 298398 622480 298522 622580
rect 298622 622480 298746 622580
rect 298846 622480 298878 622580
rect 297820 622356 298878 622480
rect 297820 622256 297850 622356
rect 297950 622256 298074 622356
rect 298174 622256 298298 622356
rect 298398 622256 298522 622356
rect 298622 622256 298746 622356
rect 298846 622256 298878 622356
rect 297820 622132 298878 622256
rect 297820 622032 297850 622132
rect 297950 622032 298074 622132
rect 298174 622032 298298 622132
rect 298398 622032 298522 622132
rect 298622 622032 298746 622132
rect 298846 622032 298878 622132
rect 297820 621908 298878 622032
rect 297820 621808 297850 621908
rect 297950 621808 298074 621908
rect 298174 621808 298298 621908
rect 298398 621808 298522 621908
rect 298622 621808 298746 621908
rect 298846 621808 298878 621908
rect 297820 621684 298878 621808
rect 297820 621584 297850 621684
rect 297950 621584 298074 621684
rect 298174 621584 298298 621684
rect 298398 621584 298522 621684
rect 298622 621584 298746 621684
rect 298846 621584 298878 621684
rect 297820 621460 298878 621584
rect 297820 621360 297850 621460
rect 297950 621360 298074 621460
rect 298174 621360 298298 621460
rect 298398 621360 298522 621460
rect 298622 621360 298746 621460
rect 298846 621360 298878 621460
rect 297820 621236 298878 621360
rect 304310 623866 305040 623900
rect 310416 623866 310786 623900
rect 304310 623544 310786 623866
rect 297820 621136 297850 621236
rect 297950 621136 298074 621236
rect 298174 621136 298298 621236
rect 298398 621136 298522 621236
rect 298622 621136 298746 621236
rect 298846 621136 298878 621236
rect 301286 621226 301362 621238
rect 301286 621174 301298 621226
rect 301350 621174 301362 621226
rect 301286 621162 301362 621174
rect 302202 621226 302278 621238
rect 302202 621174 302214 621226
rect 302266 621174 302278 621226
rect 302202 621162 302278 621174
rect 297820 621012 298878 621136
rect 300534 621110 300742 621116
rect 300980 621110 301212 621122
rect 300534 621076 300546 621110
rect 300730 621076 300742 621110
rect 300534 621070 300742 621076
rect 300844 621076 301004 621110
rect 301188 621076 301212 621110
rect 300844 621038 300888 621076
rect 300980 621058 301212 621076
rect 297820 620912 297850 621012
rect 297950 620912 298074 621012
rect 298174 620912 298298 621012
rect 298398 620912 298522 621012
rect 298622 620912 298746 621012
rect 298846 620912 298878 621012
rect 297820 620788 298878 620912
rect 297820 620688 297850 620788
rect 297950 620688 298074 620788
rect 298174 620688 298298 620788
rect 298398 620688 298522 620788
rect 298622 620688 298746 620788
rect 298846 620688 298878 620788
rect 297820 620564 298878 620688
rect 300386 621026 300432 621038
rect 300386 620650 300392 621026
rect 300426 620650 300432 621026
rect 300386 620638 300432 620650
rect 300844 621026 300890 621038
rect 300844 620650 300850 621026
rect 300884 620650 300890 621026
rect 297820 620464 297850 620564
rect 297950 620464 298074 620564
rect 298174 620464 298298 620564
rect 298398 620464 298522 620564
rect 298622 620464 298746 620564
rect 298846 620464 298878 620564
rect 300844 620508 300890 620650
rect 301302 621026 301348 621162
rect 301450 621110 301658 621116
rect 301450 621076 301462 621110
rect 301646 621076 301658 621110
rect 301450 621070 301658 621076
rect 301908 621110 302116 621116
rect 301908 621076 301920 621110
rect 302104 621076 302116 621110
rect 301908 621070 302116 621076
rect 301302 620650 301308 621026
rect 301342 620650 301348 621026
rect 301302 620638 301348 620650
rect 301760 621026 301806 621038
rect 301760 620650 301766 621026
rect 301800 620650 301806 621026
rect 297820 620340 298878 620464
rect 300834 620502 300898 620508
rect 300834 620450 300840 620502
rect 300892 620450 300898 620502
rect 300834 620444 300898 620450
rect 297820 620240 297850 620340
rect 297950 620240 298074 620340
rect 298174 620240 298298 620340
rect 298398 620240 298522 620340
rect 298622 620240 298746 620340
rect 298846 620240 298878 620340
rect 301760 620302 301806 620650
rect 302218 621026 302264 621162
rect 302344 621110 302576 621122
rect 302824 621110 303032 621116
rect 302344 621076 302378 621110
rect 302562 621076 302722 621110
rect 302344 621058 302576 621076
rect 302218 620650 302224 621026
rect 302258 620650 302264 621026
rect 302218 620638 302264 620650
rect 302676 621026 302722 621076
rect 302824 621076 302836 621110
rect 303020 621076 303032 621110
rect 302824 621070 303032 621076
rect 302676 620650 302682 621026
rect 302716 620650 302722 621026
rect 302676 620514 302722 620650
rect 303134 621026 303180 621038
rect 303134 620650 303140 621026
rect 303174 620650 303180 621026
rect 303134 620638 303180 620650
rect 302668 620508 302732 620514
rect 302668 620456 302674 620508
rect 302726 620456 302732 620508
rect 302668 620450 302732 620456
rect 303274 620508 303480 620514
rect 303274 620450 303280 620508
rect 303474 620450 303480 620508
rect 297820 620116 298878 620240
rect 301752 620296 301816 620302
rect 301752 620244 301758 620296
rect 301810 620244 301816 620296
rect 301752 620238 301816 620244
rect 297820 620016 297850 620116
rect 297950 620016 298074 620116
rect 298174 620016 298298 620116
rect 298398 620016 298522 620116
rect 298622 620016 298746 620116
rect 298846 620016 298878 620116
rect 297820 619892 298878 620016
rect 297820 619792 297850 619892
rect 297950 619792 298074 619892
rect 298174 619792 298298 619892
rect 298398 619792 298522 619892
rect 298622 619792 298746 619892
rect 298846 619792 298878 619892
rect 297820 619668 298878 619792
rect 297820 619568 297850 619668
rect 297950 619568 298074 619668
rect 298174 619568 298298 619668
rect 298398 619568 298522 619668
rect 298622 619568 298746 619668
rect 298846 619568 298878 619668
rect 297820 619444 298878 619568
rect 297820 619344 297850 619444
rect 297950 619344 298074 619444
rect 298174 619344 298298 619444
rect 298398 619344 298522 619444
rect 298622 619344 298746 619444
rect 298846 619344 298878 619444
rect 297820 619220 298878 619344
rect 297820 619120 297850 619220
rect 297950 619120 298074 619220
rect 298174 619120 298298 619220
rect 298398 619120 298522 619220
rect 298622 619120 298746 619220
rect 298846 619120 298878 619220
rect 297820 618996 298878 619120
rect 297820 618896 297850 618996
rect 297950 618896 298074 618996
rect 298174 618896 298298 618996
rect 298398 618896 298522 618996
rect 298622 618896 298746 618996
rect 298846 618896 298878 618996
rect 297820 618772 298878 618896
rect 297820 618672 297850 618772
rect 297950 618672 298074 618772
rect 298174 618672 298298 618772
rect 298398 618672 298522 618772
rect 298622 618672 298746 618772
rect 298846 618672 298878 618772
rect 297820 618548 298878 618672
rect 297820 618448 297850 618548
rect 297950 618448 298074 618548
rect 298174 618448 298298 618548
rect 298398 618448 298522 618548
rect 298622 618448 298746 618548
rect 298846 618448 298878 618548
rect 297820 618324 298878 618448
rect 297820 618224 297850 618324
rect 297950 618224 298074 618324
rect 298174 618224 298298 618324
rect 298398 618224 298522 618324
rect 298622 618224 298746 618324
rect 298846 618224 298878 618324
rect 297820 618100 298878 618224
rect 297820 618000 297850 618100
rect 297950 618000 298074 618100
rect 298174 618000 298298 618100
rect 298398 618000 298522 618100
rect 298622 618000 298746 618100
rect 298846 618000 298878 618100
rect 297820 617980 298878 618000
rect 302938 619648 303070 619660
rect 302938 617306 302954 619648
rect 303054 617306 303070 619648
rect 302938 617058 303070 617306
rect 302938 616954 302964 617058
rect 303016 616954 303070 617058
rect 302938 616944 303070 616954
rect 303274 616864 303480 620450
rect 304310 620136 304518 623544
rect 306620 622492 306804 622512
rect 306620 622438 306640 622492
rect 306784 622438 306804 622492
rect 306048 622352 306232 622372
rect 306048 622298 306068 622352
rect 306212 622298 306232 622352
rect 306048 622238 306232 622298
rect 306620 622238 306804 622438
rect 307764 622492 307948 622512
rect 307764 622438 307784 622492
rect 307928 622438 307948 622492
rect 307192 622352 307376 622372
rect 307192 622298 307212 622352
rect 307356 622298 307376 622352
rect 307192 622238 307376 622298
rect 307764 622238 307948 622438
rect 308908 622492 309092 622512
rect 308908 622438 308928 622492
rect 309072 622438 309092 622492
rect 308336 622352 308520 622372
rect 308336 622298 308356 622352
rect 308500 622298 308520 622352
rect 308336 622238 308520 622298
rect 308908 622238 309092 622438
rect 304764 622232 305820 622238
rect 304764 622198 305476 622232
rect 305660 622198 305820 622232
rect 304764 622192 305820 622198
rect 306036 622232 306244 622238
rect 306036 622198 306048 622232
rect 306232 622198 306244 622232
rect 306036 622192 306244 622198
rect 306608 622232 306816 622238
rect 306608 622198 306620 622232
rect 306804 622198 306816 622232
rect 306608 622192 306816 622198
rect 307180 622232 307388 622238
rect 307180 622198 307192 622232
rect 307376 622198 307388 622232
rect 307180 622192 307388 622198
rect 307752 622232 307960 622238
rect 307752 622198 307764 622232
rect 307948 622198 307960 622232
rect 307752 622192 307960 622198
rect 308324 622232 308532 622238
rect 308324 622198 308336 622232
rect 308520 622198 308532 622232
rect 308324 622192 308532 622198
rect 308896 622232 309104 622238
rect 308896 622198 308908 622232
rect 309092 622198 309104 622232
rect 308896 622192 309104 622198
rect 309320 622232 310376 622238
rect 309320 622198 309480 622232
rect 309664 622198 310376 622232
rect 309320 622192 310376 622198
rect 304764 622164 304878 622192
rect 304754 622148 304886 622164
rect 304754 620550 304770 622148
rect 304870 620550 304886 622148
rect 304754 620532 304886 620550
rect 305316 622148 305362 622192
rect 305316 620372 305322 622148
rect 305356 620372 305362 622148
rect 305316 620360 305362 620372
rect 305774 622148 305820 622192
rect 305774 620372 305780 622148
rect 305814 620372 305820 622148
rect 305774 620360 305820 620372
rect 305888 622148 305934 622160
rect 305888 620372 305894 622148
rect 305928 620372 305934 622148
rect 305888 620360 305934 620372
rect 306346 622148 306392 622160
rect 306346 620372 306352 622148
rect 306386 620372 306392 622148
rect 306346 620360 306392 620372
rect 306460 622148 306506 622160
rect 306460 620372 306466 622148
rect 306500 620372 306506 622148
rect 306460 620360 306506 620372
rect 306918 622148 306964 622160
rect 306918 620372 306924 622148
rect 306958 620372 306964 622148
rect 306918 620360 306964 620372
rect 307032 622148 307078 622160
rect 307032 620372 307038 622148
rect 307072 620372 307078 622148
rect 307032 620360 307078 620372
rect 307490 622148 307536 622160
rect 307490 620372 307496 622148
rect 307530 620372 307536 622148
rect 307490 620360 307536 620372
rect 307604 622148 307650 622160
rect 307604 620372 307610 622148
rect 307644 620372 307650 622148
rect 307604 620360 307650 620372
rect 308062 622148 308108 622160
rect 308062 620372 308068 622148
rect 308102 620372 308108 622148
rect 308062 620360 308108 620372
rect 308176 622148 308222 622160
rect 308176 620372 308182 622148
rect 308216 620372 308222 622148
rect 308176 620360 308222 620372
rect 308634 622148 308680 622160
rect 308634 620372 308640 622148
rect 308674 620372 308680 622148
rect 308634 620360 308680 620372
rect 308748 622148 308794 622160
rect 308748 620372 308754 622148
rect 308788 620372 308794 622148
rect 308748 620360 308794 620372
rect 309206 622148 309252 622160
rect 309206 620372 309212 622148
rect 309246 620372 309252 622148
rect 309206 620360 309252 620372
rect 309320 622148 309366 622192
rect 309320 620372 309326 622148
rect 309360 620372 309366 622148
rect 309320 620360 309366 620372
rect 309778 622148 309824 622192
rect 310262 622164 310376 622192
rect 309778 620372 309784 622148
rect 309818 620372 309824 622148
rect 310254 622148 310386 622164
rect 310254 620550 310270 622148
rect 310370 620550 310386 622148
rect 310254 620532 310386 620550
rect 309778 620360 309824 620372
rect 304310 619882 304436 620136
rect 304488 619882 304518 620136
rect 303590 619829 304094 619836
rect 303590 619795 303750 619829
rect 303934 619795 304094 619829
rect 303590 619788 304094 619795
rect 304310 619829 304518 619882
rect 304310 619795 304322 619829
rect 304506 619795 304518 619829
rect 304310 619788 304518 619795
rect 304870 620136 305078 620142
rect 304870 619882 304996 620136
rect 305048 619882 305078 620136
rect 304870 619835 305078 619882
rect 305430 620136 305638 620142
rect 305430 619882 305556 620136
rect 305608 619882 305638 620136
rect 305430 619835 305638 619882
rect 304870 619829 305090 619835
rect 304870 619795 304894 619829
rect 305078 619795 305090 619829
rect 304870 619789 305090 619795
rect 305430 619829 305662 619835
rect 305430 619795 305466 619829
rect 305650 619795 305662 619829
rect 305430 619789 305662 619795
rect 305892 619830 305926 620360
rect 306352 620296 306386 620360
rect 306326 620286 306398 620296
rect 306326 620182 306336 620286
rect 306388 620182 306398 620286
rect 306326 620172 306398 620182
rect 306464 620142 306498 620360
rect 306924 620296 306958 620360
rect 306898 620286 306970 620296
rect 306898 620182 306908 620286
rect 306960 620182 306970 620286
rect 306898 620172 306970 620182
rect 306450 620136 306514 620142
rect 306450 619882 306456 620136
rect 306508 619882 306514 620136
rect 306450 619876 306514 619882
rect 306028 619846 306248 619848
rect 306028 619835 306034 619846
rect 306026 619830 306034 619835
rect 305892 619790 306034 619830
rect 306242 619826 306248 619846
rect 304870 619788 305078 619789
rect 305430 619788 305638 619789
rect 303590 619736 303636 619788
rect 303590 617180 303596 619736
rect 303630 617180 303636 619736
rect 303590 617068 303636 617180
rect 304048 619736 304094 619788
rect 305892 619748 305926 619790
rect 306026 619789 306034 619790
rect 306028 619788 306034 619789
rect 306242 619790 306338 619826
rect 306242 619788 306248 619790
rect 306028 619778 306248 619788
rect 306464 619748 306498 619876
rect 306600 619842 306820 619848
rect 306600 619835 306606 619842
rect 306598 619789 306606 619835
rect 306600 619784 306606 619789
rect 306814 619784 306820 619842
rect 306600 619778 306820 619784
rect 307036 619830 307070 620360
rect 307496 620296 307530 620360
rect 307470 620286 307542 620296
rect 307470 620182 307480 620286
rect 307532 620182 307542 620286
rect 307470 620172 307542 620182
rect 307608 620142 307642 620360
rect 308068 620296 308102 620360
rect 308042 620286 308114 620296
rect 308042 620182 308052 620286
rect 308104 620182 308114 620286
rect 308042 620172 308114 620182
rect 307594 620136 307658 620142
rect 307594 619882 307600 620136
rect 307652 619882 307658 620136
rect 307594 619876 307658 619882
rect 307172 619846 307392 619852
rect 307172 619835 307178 619846
rect 307170 619830 307178 619835
rect 307036 619794 307178 619830
rect 307386 619830 307392 619846
rect 307036 619748 307070 619794
rect 307170 619789 307178 619794
rect 307172 619788 307178 619789
rect 307386 619794 307482 619830
rect 307386 619788 307392 619794
rect 307172 619782 307392 619788
rect 307608 619748 307642 619876
rect 307744 619846 307964 619852
rect 307744 619835 307750 619846
rect 307742 619789 307750 619835
rect 307744 619788 307750 619789
rect 307958 619788 307964 619846
rect 307744 619782 307964 619788
rect 308180 619830 308214 620360
rect 308640 620296 308674 620360
rect 308614 620286 308686 620296
rect 308614 620182 308624 620286
rect 308676 620182 308686 620286
rect 308614 620172 308686 620182
rect 308752 620142 308786 620360
rect 309212 620296 309246 620360
rect 309186 620286 309258 620296
rect 309186 620182 309196 620286
rect 309248 620182 309258 620286
rect 309186 620172 309258 620182
rect 308738 620136 308802 620142
rect 308738 619882 308744 620136
rect 308796 619882 308802 620136
rect 308738 619876 308802 619882
rect 309458 620136 309666 620142
rect 309458 619882 309544 620136
rect 309596 619882 309666 620136
rect 308316 619846 308536 619852
rect 308316 619835 308322 619846
rect 308314 619830 308322 619835
rect 308180 619794 308322 619830
rect 308530 619830 308536 619846
rect 308180 619748 308214 619794
rect 308314 619789 308322 619794
rect 308316 619788 308322 619789
rect 308530 619794 308626 619830
rect 308530 619788 308536 619794
rect 308316 619782 308536 619788
rect 308752 619748 308786 619876
rect 308888 619846 309108 619852
rect 308888 619835 308894 619846
rect 308886 619789 308894 619835
rect 308888 619788 308894 619789
rect 309102 619788 309108 619846
rect 309458 619829 309666 619882
rect 309458 619795 309470 619829
rect 309654 619795 309666 619829
rect 309458 619788 309666 619795
rect 310018 620136 310226 620142
rect 310018 619882 310104 620136
rect 310156 619882 310226 620136
rect 310018 619835 310226 619882
rect 310578 620136 310786 623544
rect 311840 622372 311972 625612
rect 312296 622512 312428 626196
rect 313814 626502 315814 626916
rect 313814 626214 313820 626502
rect 315808 626214 315814 626502
rect 313814 625008 315814 626214
rect 316514 625902 318514 625914
rect 316514 625614 316520 625902
rect 318508 625614 318514 625902
rect 316514 625008 318514 625614
rect 313854 624946 313894 625008
rect 314774 624946 314814 625008
rect 315694 624946 315734 625008
rect 312296 622432 312302 622512
rect 312422 622432 312428 622512
rect 312296 622426 312428 622432
rect 313398 624934 313444 624946
rect 311840 622292 311846 622372
rect 311956 622292 311972 622372
rect 311840 622286 311972 622292
rect 310578 619882 310664 620136
rect 310716 619882 310786 620136
rect 310578 619835 310786 619882
rect 312708 620136 313188 620142
rect 312708 619882 312714 620136
rect 313182 619882 313188 620136
rect 310018 619829 310238 619835
rect 310018 619795 310042 619829
rect 310226 619795 310238 619829
rect 310018 619789 310238 619795
rect 310578 619829 310810 619835
rect 310578 619795 310614 619829
rect 310798 619795 310810 619829
rect 310578 619789 310810 619795
rect 311026 619829 311530 619836
rect 311026 619795 311186 619829
rect 311370 619795 311530 619829
rect 310018 619788 310226 619789
rect 310578 619788 310786 619789
rect 311026 619788 311530 619795
rect 308888 619782 309108 619788
rect 304048 617180 304054 619736
rect 304088 617180 304094 619736
rect 304048 617068 304094 617180
rect 304162 619736 304208 619748
rect 304162 617180 304168 619736
rect 304202 617180 304208 619736
rect 304162 617168 304208 617180
rect 304620 619736 304666 619748
rect 304620 617180 304626 619736
rect 304660 617180 304666 619736
rect 304620 617168 304666 617180
rect 304734 619736 304780 619748
rect 304734 617180 304740 619736
rect 304774 617180 304780 619736
rect 304734 617168 304780 617180
rect 305192 619736 305238 619748
rect 305192 617180 305198 619736
rect 305232 619732 305238 619736
rect 305306 619736 305352 619748
rect 305232 617180 305240 619732
rect 305192 617168 305240 617180
rect 305306 617180 305312 619736
rect 305346 617180 305352 619736
rect 305306 617168 305352 617180
rect 305764 619736 305810 619748
rect 305764 617180 305770 619736
rect 305804 619732 305810 619736
rect 305878 619736 305926 619748
rect 305804 617180 305820 619732
rect 305764 617168 305820 617180
rect 305878 617180 305884 619736
rect 305918 619732 305926 619736
rect 306336 619736 306382 619748
rect 305918 617180 305924 619732
rect 305878 617168 305924 617180
rect 306336 617180 306342 619736
rect 306376 619732 306382 619736
rect 306450 619736 306498 619748
rect 306908 619736 306954 619748
rect 306376 617180 306384 619732
rect 306336 617168 306384 617180
rect 306450 617180 306456 619736
rect 306490 617180 306496 619736
rect 306450 617168 306496 617180
rect 306908 617180 306914 619736
rect 306948 619732 306954 619736
rect 307022 619736 307070 619748
rect 307480 619736 307526 619748
rect 306948 617180 306956 619732
rect 306908 617168 306956 617180
rect 307022 617180 307028 619736
rect 307062 617180 307068 619736
rect 307022 617168 307068 617180
rect 307480 617180 307486 619736
rect 307520 617180 307526 619736
rect 307480 617168 307526 617180
rect 307594 619736 307642 619748
rect 308052 619736 308098 619748
rect 307594 617180 307600 619736
rect 307634 617180 307640 619736
rect 307594 617168 307640 617180
rect 308052 617180 308058 619736
rect 308092 617180 308098 619736
rect 308052 617168 308098 617180
rect 308166 619736 308214 619748
rect 308624 619736 308670 619748
rect 308166 617180 308172 619736
rect 308206 617180 308212 619736
rect 308166 617168 308212 617180
rect 308624 617180 308630 619736
rect 308664 617180 308670 619736
rect 308624 617168 308670 617180
rect 308738 619736 308786 619748
rect 309196 619736 309242 619748
rect 308738 617180 308744 619736
rect 308778 617180 308784 619736
rect 308738 617168 308784 617180
rect 309196 617180 309202 619736
rect 309236 617180 309242 619736
rect 309196 617168 309242 617180
rect 309310 619736 309356 619748
rect 309310 617180 309316 619736
rect 309350 617180 309356 619736
rect 309310 617168 309356 617180
rect 309768 619736 309814 619748
rect 309768 617180 309774 619736
rect 309808 617180 309814 619736
rect 309768 617168 309814 617180
rect 309882 619736 309928 619748
rect 309882 617180 309888 619736
rect 309922 617180 309928 619736
rect 309882 617168 309928 617180
rect 310340 619736 310386 619748
rect 310340 617180 310346 619736
rect 310380 617180 310386 619736
rect 310340 617168 310386 617180
rect 310454 619736 310500 619748
rect 310454 617180 310460 619736
rect 310494 617180 310500 619736
rect 310454 617168 310500 617180
rect 310912 619736 310958 619748
rect 310912 617180 310918 619736
rect 310952 617180 310958 619736
rect 310912 617168 310958 617180
rect 311026 619736 311072 619788
rect 311026 617180 311032 619736
rect 311066 617180 311072 619736
rect 303576 617058 303648 617068
rect 303576 616954 303586 617058
rect 303638 616954 303648 617058
rect 303576 616944 303648 616954
rect 304034 617058 304106 617068
rect 304034 616954 304044 617058
rect 304096 616954 304106 617058
rect 304034 616944 304106 616954
rect 304164 616868 304206 617168
rect 304626 617068 304660 617168
rect 304610 617058 304682 617068
rect 304610 616954 304620 617058
rect 304672 616954 304682 617058
rect 304610 616944 304682 616954
rect 304736 616868 304778 617168
rect 305198 617068 305240 617168
rect 305182 617058 305254 617068
rect 305182 616954 305192 617058
rect 305244 616954 305254 617058
rect 305182 616944 305254 616954
rect 305308 616868 305350 617168
rect 305770 617068 305820 617168
rect 306342 617068 306384 617168
rect 306914 617068 306956 617168
rect 307486 617068 307520 617168
rect 308058 617068 308092 617168
rect 308630 617068 308664 617168
rect 309202 617068 309236 617168
rect 305754 617058 305826 617068
rect 305754 616954 305764 617058
rect 305816 616954 305826 617058
rect 305754 616944 305826 616954
rect 306326 617058 306398 617068
rect 306326 616954 306336 617058
rect 306388 616954 306398 617058
rect 306326 616944 306398 616954
rect 306898 617058 306970 617068
rect 306898 616954 306908 617058
rect 306960 616954 306970 617058
rect 306898 616944 306970 616954
rect 307470 617058 307542 617068
rect 307470 616954 307480 617058
rect 307532 616954 307542 617058
rect 307470 616944 307542 616954
rect 308042 617058 308114 617068
rect 308042 616954 308052 617058
rect 308104 616954 308114 617058
rect 308042 616944 308114 616954
rect 308614 617058 308686 617068
rect 308614 616954 308624 617058
rect 308676 616954 308686 617058
rect 308614 616944 308686 616954
rect 309186 617058 309254 617068
rect 309186 616954 309196 617058
rect 309248 616954 309254 617058
rect 309186 616944 309254 616954
rect 309312 616868 309354 617168
rect 309774 617068 309808 617168
rect 309758 617058 309826 617068
rect 309758 616954 309768 617058
rect 309820 616954 309826 617058
rect 309758 616944 309826 616954
rect 309884 616868 309926 617168
rect 310346 617068 310380 617168
rect 310330 617058 310398 617068
rect 310330 616954 310340 617058
rect 310392 616954 310398 617058
rect 310330 616944 310398 616954
rect 310456 616868 310498 617168
rect 310918 617068 310952 617168
rect 311026 617068 311072 617180
rect 311484 619736 311530 619788
rect 311484 617180 311490 619736
rect 311524 617180 311530 619736
rect 311484 617068 311530 617180
rect 312066 619648 312198 619660
rect 312066 617306 312082 619648
rect 312182 617306 312198 619648
rect 310902 617058 310970 617068
rect 310902 616954 310912 617058
rect 310964 616954 310970 617058
rect 310902 616944 310970 616954
rect 311012 617058 311084 617068
rect 311012 616954 311022 617058
rect 311074 616954 311084 617058
rect 311012 616944 311084 616954
rect 311470 617058 311542 617068
rect 311470 616954 311480 617058
rect 311532 616954 311542 617058
rect 311470 616944 311542 616954
rect 312066 617058 312198 617306
rect 312066 616954 312092 617058
rect 312144 616954 312198 617058
rect 312066 616944 312198 616954
rect 312708 617042 313188 619882
rect 312708 616894 312714 617042
rect 313182 616894 313188 617042
rect 312708 616888 313188 616894
rect 313398 617218 313404 624934
rect 313438 617218 313444 624934
rect 313854 624934 313902 624946
rect 313854 624908 313862 624934
rect 313398 617166 313444 617218
rect 313856 617218 313862 624908
rect 313896 617218 313902 624934
rect 313856 617202 313902 617218
rect 314314 624934 314360 624946
rect 314314 617218 314320 624934
rect 314354 617218 314360 624934
rect 314314 617206 314360 617218
rect 314772 624934 314818 624946
rect 314772 617218 314778 624934
rect 314812 617218 314818 624934
rect 314772 617206 314818 617218
rect 315230 624934 315276 624946
rect 315230 617218 315236 624934
rect 315270 617218 315276 624934
rect 315230 617206 315276 617218
rect 315688 624934 315734 624946
rect 315688 617218 315694 624934
rect 315728 617218 315734 624934
rect 315688 617206 315734 617218
rect 316146 624934 316192 624946
rect 316146 617218 316152 624934
rect 316186 617228 316192 624934
rect 316594 624934 316654 625008
rect 316594 624928 316610 624934
rect 316186 617218 316194 617228
rect 316146 617206 316194 617218
rect 316604 617218 316610 624928
rect 316644 624928 316654 624934
rect 317062 624934 317108 624946
rect 316644 617218 316650 624928
rect 317062 617228 317068 624934
rect 316604 617206 316650 617218
rect 317054 617218 317068 617228
rect 317102 617218 317108 624934
rect 317514 624934 317574 625008
rect 317514 624908 317526 624934
rect 317054 617206 317108 617218
rect 317520 617218 317526 624908
rect 317560 624908 317574 624934
rect 317978 624934 318024 624946
rect 317560 617218 317566 624908
rect 317978 617228 317984 624934
rect 317520 617206 317566 617218
rect 317974 617218 317984 617228
rect 318018 617218 318024 624934
rect 318434 624934 318494 625008
rect 319314 625006 324014 627800
rect 331482 628146 332430 628152
rect 331482 627628 331490 628146
rect 332424 627628 332430 628146
rect 327514 627366 329514 627408
rect 327514 626916 327520 627366
rect 329508 626916 329514 627366
rect 327514 626502 329514 626916
rect 327514 626214 327520 626502
rect 329508 626214 329514 626502
rect 324814 625902 326814 625914
rect 324814 625614 324820 625902
rect 326808 625614 326814 625902
rect 324814 625008 326814 625614
rect 327514 625008 329514 626214
rect 318434 624908 318442 624934
rect 317974 617206 318024 617218
rect 318436 617218 318442 624908
rect 318476 624908 318494 624934
rect 319354 624946 319394 625006
rect 320274 624946 320314 625006
rect 321194 624946 321234 625006
rect 322114 624946 322154 625006
rect 319354 624934 319402 624946
rect 319354 624928 319362 624934
rect 318476 617218 318482 624908
rect 318436 617206 318482 617218
rect 319356 617218 319362 624928
rect 319396 617218 319402 624934
rect 319356 617206 319402 617218
rect 319814 624934 319860 624946
rect 319814 617218 319820 624934
rect 319854 617218 319860 624934
rect 319814 617206 319860 617218
rect 320272 624934 320318 624946
rect 320272 617218 320278 624934
rect 320312 617218 320318 624934
rect 320272 617206 320318 617218
rect 320730 624934 320776 624946
rect 320730 617218 320736 624934
rect 320770 617218 320776 624934
rect 320730 617206 320776 617218
rect 321188 624934 321234 624946
rect 321188 617218 321194 624934
rect 321228 617218 321234 624934
rect 321188 617206 321234 617218
rect 321646 624934 321692 624946
rect 321646 617218 321652 624934
rect 321686 617228 321692 624934
rect 322104 624934 322154 624946
rect 321686 617218 321694 617228
rect 321646 617206 321694 617218
rect 322104 617218 322110 624934
rect 322144 624908 322154 624934
rect 322562 624934 322608 624946
rect 322144 617218 322150 624908
rect 322562 617228 322568 624934
rect 322104 617206 322150 617218
rect 322554 617218 322568 617228
rect 322602 617218 322608 624934
rect 323014 624934 323074 625006
rect 323014 624908 323026 624934
rect 322554 617206 322608 617218
rect 323020 617218 323026 624908
rect 323060 624908 323074 624934
rect 323478 624934 323524 624946
rect 323060 617218 323066 624908
rect 323478 617228 323484 624934
rect 323020 617206 323066 617218
rect 323474 617218 323484 617228
rect 323518 617218 323524 624934
rect 323934 624934 323994 625006
rect 323934 624908 323942 624934
rect 323474 617206 323524 617218
rect 323936 617218 323942 624908
rect 323976 624908 323994 624934
rect 324854 624946 324894 625008
rect 325774 624946 325814 625008
rect 326694 624946 326734 625008
rect 324854 624934 324902 624946
rect 324854 624908 324862 624934
rect 323976 617218 323982 624908
rect 323936 617206 323982 617218
rect 324856 617218 324862 624908
rect 324896 617218 324902 624934
rect 324856 617206 324902 617218
rect 325314 624934 325360 624946
rect 325314 617218 325320 624934
rect 325354 617218 325360 624934
rect 325314 617206 325360 617218
rect 325772 624934 325818 624946
rect 325772 617218 325778 624934
rect 325812 617218 325818 624934
rect 325772 617206 325818 617218
rect 326230 624934 326276 624946
rect 326230 617218 326236 624934
rect 326270 617218 326276 624934
rect 326230 617206 326276 617218
rect 326688 624934 326734 624946
rect 326688 617218 326694 624934
rect 326728 617218 326734 624934
rect 326688 617206 326734 617218
rect 327146 624934 327192 624946
rect 327146 617218 327152 624934
rect 327186 617228 327192 624934
rect 327594 624934 327654 625008
rect 327594 624908 327610 624934
rect 327186 617218 327194 617228
rect 327146 617206 327194 617218
rect 327604 617218 327610 624908
rect 327644 624908 327654 624934
rect 328062 624934 328108 624946
rect 327644 617218 327650 624908
rect 328062 617228 328068 624934
rect 327604 617206 327650 617218
rect 328054 617218 328068 617228
rect 328102 617218 328108 624934
rect 328514 624934 328574 625008
rect 329434 624946 329474 625008
rect 328514 624928 328526 624934
rect 328054 617206 328108 617218
rect 328520 617218 328526 624928
rect 328560 624928 328574 624934
rect 328978 624934 329024 624946
rect 328560 617218 328566 624928
rect 328978 617228 328984 624934
rect 328520 617206 328566 617218
rect 328974 617218 328984 617228
rect 329018 617218 329024 624934
rect 329434 624934 329482 624946
rect 329434 624928 329442 624934
rect 328974 617206 329024 617218
rect 329436 617218 329442 624928
rect 329476 617218 329482 624934
rect 313398 617165 313546 617166
rect 313738 617165 313856 617166
rect 314014 617165 314194 617168
rect 313398 617159 313856 617165
rect 313398 617125 313558 617159
rect 313742 617125 313856 617159
rect 303274 616750 303280 616864
rect 303474 616750 303480 616864
rect 303274 616744 303480 616750
rect 304150 616858 304222 616868
rect 304150 616754 304160 616858
rect 304212 616754 304222 616858
rect 304150 616744 304222 616754
rect 304722 616858 304794 616868
rect 304722 616754 304732 616858
rect 304784 616754 304794 616858
rect 304722 616744 304794 616754
rect 305294 616858 305366 616868
rect 305294 616754 305304 616858
rect 305356 616754 305366 616858
rect 309298 616858 309370 616868
rect 305294 616744 305366 616754
rect 306524 616802 308978 616818
rect 306524 616702 306536 616802
rect 308878 616702 308978 616802
rect 309298 616754 309308 616858
rect 309360 616754 309370 616858
rect 309298 616744 309370 616754
rect 309870 616858 309942 616868
rect 309870 616754 309880 616858
rect 309932 616754 309942 616858
rect 309870 616744 309942 616754
rect 310442 616858 310514 616868
rect 310442 616754 310452 616858
rect 310504 616754 310514 616858
rect 313398 616808 313856 617125
rect 314004 617159 314212 617165
rect 314004 617125 314016 617159
rect 314200 617125 314212 617159
rect 314004 617119 314212 617125
rect 314014 617028 314194 617119
rect 314014 616908 314034 617028
rect 314174 616908 314194 617028
rect 314014 616888 314194 616908
rect 314314 616848 314354 617206
rect 314474 617165 314654 617168
rect 314934 617165 315114 617168
rect 314462 617159 314670 617165
rect 314462 617125 314474 617159
rect 314658 617125 314670 617159
rect 314462 617119 314670 617125
rect 314920 617159 315128 617165
rect 314920 617125 314932 617159
rect 315116 617125 315128 617159
rect 314920 617119 315128 617125
rect 314474 617028 314654 617119
rect 314474 616908 314494 617028
rect 314634 616908 314654 617028
rect 314474 616888 314654 616908
rect 314934 617028 315114 617119
rect 314934 616908 314954 617028
rect 315094 616908 315114 617028
rect 314934 616888 315114 616908
rect 315234 616848 315274 617206
rect 315394 617165 315574 617168
rect 315854 617165 316034 617168
rect 315378 617159 315586 617165
rect 315378 617125 315390 617159
rect 315574 617125 315586 617159
rect 315378 617119 315586 617125
rect 315836 617159 316044 617165
rect 315836 617125 315848 617159
rect 316032 617125 316044 617159
rect 315836 617119 316044 617125
rect 315394 617028 315574 617119
rect 315394 616908 315414 617028
rect 315554 616908 315574 617028
rect 315394 616888 315574 616908
rect 315854 617028 316034 617119
rect 315854 616908 315874 617028
rect 316014 616908 316034 617028
rect 315854 616888 316034 616908
rect 316154 616848 316194 617206
rect 316314 617165 316494 617168
rect 316774 617165 316954 617168
rect 316294 617159 316502 617165
rect 316294 617125 316306 617159
rect 316490 617125 316502 617159
rect 316294 617119 316502 617125
rect 316752 617159 316960 617165
rect 316752 617125 316764 617159
rect 316948 617125 316960 617159
rect 316752 617119 316960 617125
rect 316314 617028 316494 617119
rect 316314 616908 316334 617028
rect 316474 616908 316494 617028
rect 316314 616888 316494 616908
rect 316774 617028 316954 617119
rect 316774 616908 316794 617028
rect 316934 616908 316954 617028
rect 316774 616888 316954 616908
rect 317054 616848 317094 617206
rect 317234 617165 317414 617168
rect 317694 617165 317874 617168
rect 317210 617159 317418 617165
rect 317210 617125 317222 617159
rect 317406 617125 317418 617159
rect 317210 617119 317418 617125
rect 317668 617159 317876 617165
rect 317668 617125 317680 617159
rect 317864 617125 317876 617159
rect 317668 617119 317876 617125
rect 317234 617028 317414 617119
rect 317234 616908 317254 617028
rect 317394 616908 317414 617028
rect 317234 616888 317414 616908
rect 317694 617028 317874 617119
rect 317694 616908 317714 617028
rect 317854 616908 317874 617028
rect 317694 616888 317874 616908
rect 317974 616848 318014 617206
rect 318154 617165 318334 617168
rect 319514 617165 319694 617168
rect 318126 617159 318334 617165
rect 318126 617125 318138 617159
rect 318322 617125 318334 617159
rect 318126 617119 318334 617125
rect 319504 617159 319712 617165
rect 319504 617125 319516 617159
rect 319700 617125 319712 617159
rect 319504 617119 319712 617125
rect 318154 617028 318334 617119
rect 318154 616908 318174 617028
rect 318314 616908 318334 617028
rect 318154 616888 318334 616908
rect 319514 617028 319694 617119
rect 319514 616908 319534 617028
rect 319674 616908 319694 617028
rect 319514 616888 319694 616908
rect 319814 616848 319854 617206
rect 319974 617165 320154 617168
rect 320434 617165 320614 617168
rect 319962 617159 320170 617165
rect 319962 617125 319974 617159
rect 320158 617125 320170 617159
rect 319962 617119 320170 617125
rect 320420 617159 320628 617165
rect 320420 617125 320432 617159
rect 320616 617125 320628 617159
rect 320420 617119 320628 617125
rect 319974 617028 320154 617119
rect 319974 616908 319994 617028
rect 320134 616908 320154 617028
rect 319974 616888 320154 616908
rect 320434 617028 320614 617119
rect 320434 616908 320454 617028
rect 320594 616908 320614 617028
rect 320434 616888 320614 616908
rect 320734 616848 320774 617206
rect 320894 617165 321074 617168
rect 321354 617165 321534 617168
rect 320878 617159 321086 617165
rect 320878 617125 320890 617159
rect 321074 617125 321086 617159
rect 320878 617119 321086 617125
rect 321336 617159 321544 617165
rect 321336 617125 321348 617159
rect 321532 617125 321544 617159
rect 321336 617119 321544 617125
rect 320894 617028 321074 617119
rect 320894 616908 320914 617028
rect 321054 616908 321074 617028
rect 320894 616888 321074 616908
rect 321354 617028 321534 617119
rect 321354 616908 321374 617028
rect 321514 616908 321534 617028
rect 321354 616888 321534 616908
rect 321654 616848 321694 617206
rect 321814 617165 321994 617168
rect 322274 617165 322454 617168
rect 321794 617159 322002 617165
rect 321794 617125 321806 617159
rect 321990 617125 322002 617159
rect 321794 617119 322002 617125
rect 322252 617159 322460 617165
rect 322252 617125 322264 617159
rect 322448 617125 322460 617159
rect 322252 617119 322460 617125
rect 321814 617028 321994 617119
rect 321814 616908 321834 617028
rect 321974 616908 321994 617028
rect 321814 616888 321994 616908
rect 322274 617028 322454 617119
rect 322274 616908 322294 617028
rect 322434 616908 322454 617028
rect 322274 616888 322454 616908
rect 322554 616848 322594 617206
rect 322734 617165 322914 617168
rect 323194 617165 323374 617168
rect 322710 617159 322918 617165
rect 322710 617125 322722 617159
rect 322906 617125 322918 617159
rect 322710 617119 322918 617125
rect 323168 617159 323376 617165
rect 323168 617125 323180 617159
rect 323364 617125 323376 617159
rect 323168 617119 323376 617125
rect 322734 617028 322914 617119
rect 322734 616908 322754 617028
rect 322894 616908 322914 617028
rect 322734 616888 322914 616908
rect 323194 617028 323374 617119
rect 323194 616908 323214 617028
rect 323354 616908 323374 617028
rect 323194 616888 323374 616908
rect 323474 616848 323514 617206
rect 323654 617165 323834 617168
rect 325014 617165 325194 617168
rect 323626 617159 323834 617165
rect 323626 617125 323638 617159
rect 323822 617125 323834 617159
rect 323626 617119 323834 617125
rect 325004 617159 325212 617165
rect 325004 617125 325016 617159
rect 325200 617125 325212 617159
rect 325004 617119 325212 617125
rect 323654 617028 323834 617119
rect 323654 616908 323674 617028
rect 323814 616908 323834 617028
rect 323654 616888 323834 616908
rect 325014 617028 325194 617119
rect 325014 616908 325034 617028
rect 325174 616908 325194 617028
rect 325014 616888 325194 616908
rect 325314 616848 325354 617206
rect 325474 617165 325654 617168
rect 325934 617165 326114 617168
rect 325462 617159 325670 617165
rect 325462 617125 325474 617159
rect 325658 617125 325670 617159
rect 325462 617119 325670 617125
rect 325920 617159 326128 617165
rect 325920 617125 325932 617159
rect 326116 617125 326128 617159
rect 325920 617119 326128 617125
rect 325474 617028 325654 617119
rect 325474 616908 325494 617028
rect 325634 616908 325654 617028
rect 325474 616888 325654 616908
rect 325934 617028 326114 617119
rect 325934 616908 325954 617028
rect 326094 616908 326114 617028
rect 325934 616888 326114 616908
rect 326234 616848 326274 617206
rect 326394 617165 326574 617168
rect 326854 617165 327034 617168
rect 326378 617159 326586 617165
rect 326378 617125 326390 617159
rect 326574 617125 326586 617159
rect 326378 617119 326586 617125
rect 326836 617159 327044 617165
rect 326836 617125 326848 617159
rect 327032 617125 327044 617159
rect 326836 617119 327044 617125
rect 326394 617028 326574 617119
rect 326394 616908 326414 617028
rect 326554 616908 326574 617028
rect 326394 616888 326574 616908
rect 326854 617028 327034 617119
rect 326854 616908 326874 617028
rect 327014 616908 327034 617028
rect 326854 616888 327034 616908
rect 327154 616848 327194 617206
rect 327314 617165 327494 617168
rect 327774 617165 327954 617168
rect 327294 617159 327502 617165
rect 327294 617125 327306 617159
rect 327490 617125 327502 617159
rect 327294 617119 327502 617125
rect 327752 617159 327960 617165
rect 327752 617125 327764 617159
rect 327948 617125 327960 617159
rect 327752 617119 327960 617125
rect 327314 617028 327494 617119
rect 327314 616908 327334 617028
rect 327474 616908 327494 617028
rect 327314 616888 327494 616908
rect 327774 617028 327954 617119
rect 327774 616908 327794 617028
rect 327934 616908 327954 617028
rect 327774 616888 327954 616908
rect 328054 616848 328094 617206
rect 328234 617165 328414 617168
rect 328694 617165 328874 617168
rect 328210 617159 328418 617165
rect 328210 617125 328222 617159
rect 328406 617125 328418 617159
rect 328210 617119 328418 617125
rect 328668 617159 328876 617165
rect 328668 617125 328680 617159
rect 328864 617125 328876 617159
rect 328668 617119 328876 617125
rect 328234 617028 328414 617119
rect 328234 616908 328254 617028
rect 328394 616908 328414 617028
rect 328234 616888 328414 616908
rect 328694 617028 328874 617119
rect 328694 616908 328714 617028
rect 328854 616908 328874 617028
rect 328694 616888 328874 616908
rect 328974 616848 329014 617206
rect 329436 617202 329482 617218
rect 329894 624934 329940 624946
rect 329894 617218 329900 624934
rect 329934 617218 329940 624934
rect 331482 618668 332430 627628
rect 332826 627366 333530 630004
rect 332826 626916 332832 627366
rect 333524 626916 333530 627366
rect 332826 623578 333530 626916
rect 333644 630696 334348 630702
rect 333644 630004 333650 630696
rect 334342 630004 334348 630696
rect 334544 630685 335106 630691
rect 334544 630288 334556 630685
rect 335094 630288 335106 630685
rect 334544 630282 335106 630288
rect 333644 625902 334348 630004
rect 333644 625614 333652 625902
rect 334342 625614 334348 625902
rect 333644 625608 334348 625614
rect 334944 627370 340788 627424
rect 334944 627336 335032 627370
rect 335066 627336 335132 627370
rect 335166 627336 335232 627370
rect 335266 627336 335332 627370
rect 335366 627336 335432 627370
rect 335466 627336 335532 627370
rect 335566 627336 336320 627370
rect 336354 627336 336420 627370
rect 336454 627336 336520 627370
rect 336554 627336 336620 627370
rect 336654 627336 336720 627370
rect 336754 627336 336820 627370
rect 336854 627336 337608 627370
rect 337642 627336 337708 627370
rect 337742 627336 337808 627370
rect 337842 627336 337908 627370
rect 337942 627336 338008 627370
rect 338042 627336 338108 627370
rect 338142 627336 338896 627370
rect 338930 627336 338996 627370
rect 339030 627336 339096 627370
rect 339130 627336 339196 627370
rect 339230 627336 339296 627370
rect 339330 627336 339396 627370
rect 339430 627336 340184 627370
rect 340218 627336 340284 627370
rect 340318 627336 340384 627370
rect 340418 627336 340484 627370
rect 340518 627336 340584 627370
rect 340618 627336 340684 627370
rect 340718 627336 340788 627370
rect 334944 627270 340788 627336
rect 334944 627236 335032 627270
rect 335066 627236 335132 627270
rect 335166 627236 335232 627270
rect 335266 627236 335332 627270
rect 335366 627236 335432 627270
rect 335466 627236 335532 627270
rect 335566 627236 336320 627270
rect 336354 627236 336420 627270
rect 336454 627236 336520 627270
rect 336554 627236 336620 627270
rect 336654 627236 336720 627270
rect 336754 627236 336820 627270
rect 336854 627236 337608 627270
rect 337642 627236 337708 627270
rect 337742 627236 337808 627270
rect 337842 627236 337908 627270
rect 337942 627236 338008 627270
rect 338042 627236 338108 627270
rect 338142 627236 338896 627270
rect 338930 627236 338996 627270
rect 339030 627236 339096 627270
rect 339130 627236 339196 627270
rect 339230 627236 339296 627270
rect 339330 627236 339396 627270
rect 339430 627236 340184 627270
rect 340218 627236 340284 627270
rect 340318 627236 340384 627270
rect 340418 627236 340484 627270
rect 340518 627236 340584 627270
rect 340618 627236 340684 627270
rect 340718 627236 340788 627270
rect 334944 627170 340788 627236
rect 334944 627136 335032 627170
rect 335066 627136 335132 627170
rect 335166 627136 335232 627170
rect 335266 627136 335332 627170
rect 335366 627136 335432 627170
rect 335466 627136 335532 627170
rect 335566 627136 336320 627170
rect 336354 627136 336420 627170
rect 336454 627136 336520 627170
rect 336554 627136 336620 627170
rect 336654 627136 336720 627170
rect 336754 627136 336820 627170
rect 336854 627136 337608 627170
rect 337642 627136 337708 627170
rect 337742 627136 337808 627170
rect 337842 627136 337908 627170
rect 337942 627136 338008 627170
rect 338042 627136 338108 627170
rect 338142 627136 338896 627170
rect 338930 627136 338996 627170
rect 339030 627136 339096 627170
rect 339130 627136 339196 627170
rect 339230 627136 339296 627170
rect 339330 627136 339396 627170
rect 339430 627136 340184 627170
rect 340218 627136 340284 627170
rect 340318 627136 340384 627170
rect 340418 627136 340484 627170
rect 340518 627136 340584 627170
rect 340618 627136 340684 627170
rect 340718 627136 340788 627170
rect 334944 627070 340788 627136
rect 334944 627036 335032 627070
rect 335066 627036 335132 627070
rect 335166 627036 335232 627070
rect 335266 627036 335332 627070
rect 335366 627036 335432 627070
rect 335466 627036 335532 627070
rect 335566 627036 336320 627070
rect 336354 627036 336420 627070
rect 336454 627036 336520 627070
rect 336554 627036 336620 627070
rect 336654 627036 336720 627070
rect 336754 627036 336820 627070
rect 336854 627036 337608 627070
rect 337642 627036 337708 627070
rect 337742 627036 337808 627070
rect 337842 627036 337908 627070
rect 337942 627036 338008 627070
rect 338042 627036 338108 627070
rect 338142 627036 338896 627070
rect 338930 627036 338996 627070
rect 339030 627036 339096 627070
rect 339130 627036 339196 627070
rect 339230 627036 339296 627070
rect 339330 627036 339396 627070
rect 339430 627036 340184 627070
rect 340218 627036 340284 627070
rect 340318 627036 340384 627070
rect 340418 627036 340484 627070
rect 340518 627036 340584 627070
rect 340618 627036 340684 627070
rect 340718 627036 340788 627070
rect 334944 626970 340788 627036
rect 334944 626936 335032 626970
rect 335066 626936 335132 626970
rect 335166 626936 335232 626970
rect 335266 626936 335332 626970
rect 335366 626936 335432 626970
rect 335466 626936 335532 626970
rect 335566 626936 336320 626970
rect 336354 626936 336420 626970
rect 336454 626936 336520 626970
rect 336554 626936 336620 626970
rect 336654 626936 336720 626970
rect 336754 626936 336820 626970
rect 336854 626936 337608 626970
rect 337642 626936 337708 626970
rect 337742 626936 337808 626970
rect 337842 626936 337908 626970
rect 337942 626936 338008 626970
rect 338042 626936 338108 626970
rect 338142 626936 338896 626970
rect 338930 626936 338996 626970
rect 339030 626936 339096 626970
rect 339130 626936 339196 626970
rect 339230 626936 339296 626970
rect 339330 626936 339396 626970
rect 339430 626936 340184 626970
rect 340218 626936 340284 626970
rect 340318 626936 340384 626970
rect 340418 626936 340484 626970
rect 340518 626936 340584 626970
rect 340618 626936 340684 626970
rect 340718 626936 340788 626970
rect 334944 626870 340788 626936
rect 334944 626836 335032 626870
rect 335066 626836 335132 626870
rect 335166 626836 335232 626870
rect 335266 626836 335332 626870
rect 335366 626836 335432 626870
rect 335466 626836 335532 626870
rect 335566 626836 336320 626870
rect 336354 626836 336420 626870
rect 336454 626836 336520 626870
rect 336554 626836 336620 626870
rect 336654 626836 336720 626870
rect 336754 626836 336820 626870
rect 336854 626836 337608 626870
rect 337642 626836 337708 626870
rect 337742 626836 337808 626870
rect 337842 626836 337908 626870
rect 337942 626836 338008 626870
rect 338042 626836 338108 626870
rect 338142 626836 338896 626870
rect 338930 626836 338996 626870
rect 339030 626836 339096 626870
rect 339130 626836 339196 626870
rect 339230 626836 339296 626870
rect 339330 626836 339396 626870
rect 339430 626836 340184 626870
rect 340218 626836 340284 626870
rect 340318 626836 340384 626870
rect 340418 626836 340484 626870
rect 340518 626836 340584 626870
rect 340618 626836 340684 626870
rect 340718 626836 340788 626870
rect 334944 626082 340788 626836
rect 334944 626048 335032 626082
rect 335066 626048 335132 626082
rect 335166 626048 335232 626082
rect 335266 626048 335332 626082
rect 335366 626048 335432 626082
rect 335466 626048 335532 626082
rect 335566 626048 336320 626082
rect 336354 626048 336420 626082
rect 336454 626048 336520 626082
rect 336554 626048 336620 626082
rect 336654 626048 336720 626082
rect 336754 626048 336820 626082
rect 336854 626048 337608 626082
rect 337642 626048 337708 626082
rect 337742 626048 337808 626082
rect 337842 626048 337908 626082
rect 337942 626048 338008 626082
rect 338042 626048 338108 626082
rect 338142 626048 338896 626082
rect 338930 626048 338996 626082
rect 339030 626048 339096 626082
rect 339130 626048 339196 626082
rect 339230 626048 339296 626082
rect 339330 626048 339396 626082
rect 339430 626048 340184 626082
rect 340218 626048 340284 626082
rect 340318 626048 340384 626082
rect 340418 626048 340484 626082
rect 340518 626048 340584 626082
rect 340618 626048 340684 626082
rect 340718 626048 340788 626082
rect 334944 625982 340788 626048
rect 334944 625948 335032 625982
rect 335066 625948 335132 625982
rect 335166 625948 335232 625982
rect 335266 625948 335332 625982
rect 335366 625948 335432 625982
rect 335466 625948 335532 625982
rect 335566 625948 336320 625982
rect 336354 625948 336420 625982
rect 336454 625948 336520 625982
rect 336554 625948 336620 625982
rect 336654 625948 336720 625982
rect 336754 625948 336820 625982
rect 336854 625948 337608 625982
rect 337642 625948 337708 625982
rect 337742 625948 337808 625982
rect 337842 625948 337908 625982
rect 337942 625948 338008 625982
rect 338042 625948 338108 625982
rect 338142 625948 338896 625982
rect 338930 625948 338996 625982
rect 339030 625948 339096 625982
rect 339130 625948 339196 625982
rect 339230 625948 339296 625982
rect 339330 625948 339396 625982
rect 339430 625948 340184 625982
rect 340218 625948 340284 625982
rect 340318 625948 340384 625982
rect 340418 625948 340484 625982
rect 340518 625948 340584 625982
rect 340618 625948 340684 625982
rect 340718 625948 340788 625982
rect 334944 625882 340788 625948
rect 334944 625848 335032 625882
rect 335066 625848 335132 625882
rect 335166 625848 335232 625882
rect 335266 625848 335332 625882
rect 335366 625848 335432 625882
rect 335466 625848 335532 625882
rect 335566 625848 336320 625882
rect 336354 625848 336420 625882
rect 336454 625848 336520 625882
rect 336554 625848 336620 625882
rect 336654 625848 336720 625882
rect 336754 625848 336820 625882
rect 336854 625848 337608 625882
rect 337642 625848 337708 625882
rect 337742 625848 337808 625882
rect 337842 625848 337908 625882
rect 337942 625848 338008 625882
rect 338042 625848 338108 625882
rect 338142 625848 338896 625882
rect 338930 625848 338996 625882
rect 339030 625848 339096 625882
rect 339130 625848 339196 625882
rect 339230 625848 339296 625882
rect 339330 625848 339396 625882
rect 339430 625848 340184 625882
rect 340218 625848 340284 625882
rect 340318 625848 340384 625882
rect 340418 625848 340484 625882
rect 340518 625848 340584 625882
rect 340618 625848 340684 625882
rect 340718 625848 340788 625882
rect 334944 625782 340788 625848
rect 334944 625748 335032 625782
rect 335066 625748 335132 625782
rect 335166 625748 335232 625782
rect 335266 625748 335332 625782
rect 335366 625748 335432 625782
rect 335466 625748 335532 625782
rect 335566 625748 336320 625782
rect 336354 625748 336420 625782
rect 336454 625748 336520 625782
rect 336554 625748 336620 625782
rect 336654 625748 336720 625782
rect 336754 625748 336820 625782
rect 336854 625748 337608 625782
rect 337642 625748 337708 625782
rect 337742 625748 337808 625782
rect 337842 625748 337908 625782
rect 337942 625748 338008 625782
rect 338042 625748 338108 625782
rect 338142 625748 338896 625782
rect 338930 625748 338996 625782
rect 339030 625748 339096 625782
rect 339130 625748 339196 625782
rect 339230 625748 339296 625782
rect 339330 625748 339396 625782
rect 339430 625748 340184 625782
rect 340218 625748 340284 625782
rect 340318 625748 340384 625782
rect 340418 625748 340484 625782
rect 340518 625748 340584 625782
rect 340618 625748 340684 625782
rect 340718 625748 340788 625782
rect 334944 625682 340788 625748
rect 334944 625648 335032 625682
rect 335066 625648 335132 625682
rect 335166 625648 335232 625682
rect 335266 625648 335332 625682
rect 335366 625648 335432 625682
rect 335466 625648 335532 625682
rect 335566 625648 336320 625682
rect 336354 625648 336420 625682
rect 336454 625648 336520 625682
rect 336554 625648 336620 625682
rect 336654 625648 336720 625682
rect 336754 625648 336820 625682
rect 336854 625648 337608 625682
rect 337642 625648 337708 625682
rect 337742 625648 337808 625682
rect 337842 625648 337908 625682
rect 337942 625648 338008 625682
rect 338042 625648 338108 625682
rect 338142 625648 338896 625682
rect 338930 625648 338996 625682
rect 339030 625648 339096 625682
rect 339130 625648 339196 625682
rect 339230 625648 339296 625682
rect 339330 625648 339396 625682
rect 339430 625648 340184 625682
rect 340218 625648 340284 625682
rect 340318 625648 340384 625682
rect 340418 625648 340484 625682
rect 340518 625648 340584 625682
rect 340618 625648 340684 625682
rect 340718 625648 340788 625682
rect 332826 622886 332832 623578
rect 333524 622886 333530 623578
rect 332826 622878 333530 622886
rect 334944 625582 340788 625648
rect 334944 625548 335032 625582
rect 335066 625548 335132 625582
rect 335166 625548 335232 625582
rect 335266 625548 335332 625582
rect 335366 625548 335432 625582
rect 335466 625548 335532 625582
rect 335566 625548 336320 625582
rect 336354 625548 336420 625582
rect 336454 625548 336520 625582
rect 336554 625548 336620 625582
rect 336654 625548 336720 625582
rect 336754 625548 336820 625582
rect 336854 625548 337608 625582
rect 337642 625548 337708 625582
rect 337742 625548 337808 625582
rect 337842 625548 337908 625582
rect 337942 625548 338008 625582
rect 338042 625548 338108 625582
rect 338142 625548 338896 625582
rect 338930 625548 338996 625582
rect 339030 625548 339096 625582
rect 339130 625548 339196 625582
rect 339230 625548 339296 625582
rect 339330 625548 339396 625582
rect 339430 625548 340184 625582
rect 340218 625548 340284 625582
rect 340318 625548 340384 625582
rect 340418 625548 340484 625582
rect 340518 625548 340584 625582
rect 340618 625548 340684 625582
rect 340718 625548 340788 625582
rect 334944 624794 340788 625548
rect 334944 624760 335032 624794
rect 335066 624760 335132 624794
rect 335166 624760 335232 624794
rect 335266 624760 335332 624794
rect 335366 624760 335432 624794
rect 335466 624760 335532 624794
rect 335566 624760 336320 624794
rect 336354 624760 336420 624794
rect 336454 624760 336520 624794
rect 336554 624760 336620 624794
rect 336654 624760 336720 624794
rect 336754 624760 336820 624794
rect 336854 624760 337608 624794
rect 337642 624760 337708 624794
rect 337742 624760 337808 624794
rect 337842 624760 337908 624794
rect 337942 624760 338008 624794
rect 338042 624760 338108 624794
rect 338142 624760 338896 624794
rect 338930 624760 338996 624794
rect 339030 624760 339096 624794
rect 339130 624760 339196 624794
rect 339230 624760 339296 624794
rect 339330 624760 339396 624794
rect 339430 624760 340184 624794
rect 340218 624760 340284 624794
rect 340318 624760 340384 624794
rect 340418 624760 340484 624794
rect 340518 624760 340584 624794
rect 340618 624760 340684 624794
rect 340718 624760 340788 624794
rect 334944 624694 340788 624760
rect 334944 624660 335032 624694
rect 335066 624660 335132 624694
rect 335166 624660 335232 624694
rect 335266 624660 335332 624694
rect 335366 624660 335432 624694
rect 335466 624660 335532 624694
rect 335566 624660 336320 624694
rect 336354 624660 336420 624694
rect 336454 624660 336520 624694
rect 336554 624660 336620 624694
rect 336654 624660 336720 624694
rect 336754 624660 336820 624694
rect 336854 624660 337608 624694
rect 337642 624660 337708 624694
rect 337742 624660 337808 624694
rect 337842 624660 337908 624694
rect 337942 624660 338008 624694
rect 338042 624660 338108 624694
rect 338142 624660 338896 624694
rect 338930 624660 338996 624694
rect 339030 624660 339096 624694
rect 339130 624660 339196 624694
rect 339230 624660 339296 624694
rect 339330 624660 339396 624694
rect 339430 624660 340184 624694
rect 340218 624660 340284 624694
rect 340318 624660 340384 624694
rect 340418 624660 340484 624694
rect 340518 624660 340584 624694
rect 340618 624660 340684 624694
rect 340718 624660 340788 624694
rect 334944 624594 340788 624660
rect 334944 624560 335032 624594
rect 335066 624560 335132 624594
rect 335166 624560 335232 624594
rect 335266 624560 335332 624594
rect 335366 624560 335432 624594
rect 335466 624560 335532 624594
rect 335566 624560 336320 624594
rect 336354 624560 336420 624594
rect 336454 624560 336520 624594
rect 336554 624560 336620 624594
rect 336654 624560 336720 624594
rect 336754 624560 336820 624594
rect 336854 624560 337608 624594
rect 337642 624560 337708 624594
rect 337742 624560 337808 624594
rect 337842 624560 337908 624594
rect 337942 624560 338008 624594
rect 338042 624560 338108 624594
rect 338142 624560 338896 624594
rect 338930 624560 338996 624594
rect 339030 624560 339096 624594
rect 339130 624560 339196 624594
rect 339230 624560 339296 624594
rect 339330 624560 339396 624594
rect 339430 624560 340184 624594
rect 340218 624560 340284 624594
rect 340318 624560 340384 624594
rect 340418 624560 340484 624594
rect 340518 624560 340584 624594
rect 340618 624560 340684 624594
rect 340718 624560 340788 624594
rect 334944 624494 340788 624560
rect 334944 624460 335032 624494
rect 335066 624460 335132 624494
rect 335166 624460 335232 624494
rect 335266 624460 335332 624494
rect 335366 624460 335432 624494
rect 335466 624460 335532 624494
rect 335566 624460 336320 624494
rect 336354 624460 336420 624494
rect 336454 624460 336520 624494
rect 336554 624460 336620 624494
rect 336654 624460 336720 624494
rect 336754 624460 336820 624494
rect 336854 624460 337608 624494
rect 337642 624460 337708 624494
rect 337742 624460 337808 624494
rect 337842 624460 337908 624494
rect 337942 624460 338008 624494
rect 338042 624460 338108 624494
rect 338142 624460 338896 624494
rect 338930 624460 338996 624494
rect 339030 624460 339096 624494
rect 339130 624460 339196 624494
rect 339230 624460 339296 624494
rect 339330 624460 339396 624494
rect 339430 624460 340184 624494
rect 340218 624460 340284 624494
rect 340318 624460 340384 624494
rect 340418 624460 340484 624494
rect 340518 624460 340584 624494
rect 340618 624460 340684 624494
rect 340718 624460 340788 624494
rect 334944 624394 340788 624460
rect 334944 624360 335032 624394
rect 335066 624360 335132 624394
rect 335166 624360 335232 624394
rect 335266 624360 335332 624394
rect 335366 624360 335432 624394
rect 335466 624360 335532 624394
rect 335566 624360 336320 624394
rect 336354 624360 336420 624394
rect 336454 624360 336520 624394
rect 336554 624360 336620 624394
rect 336654 624360 336720 624394
rect 336754 624360 336820 624394
rect 336854 624360 337608 624394
rect 337642 624360 337708 624394
rect 337742 624360 337808 624394
rect 337842 624360 337908 624394
rect 337942 624360 338008 624394
rect 338042 624360 338108 624394
rect 338142 624360 338896 624394
rect 338930 624360 338996 624394
rect 339030 624360 339096 624394
rect 339130 624360 339196 624394
rect 339230 624360 339296 624394
rect 339330 624360 339396 624394
rect 339430 624360 340184 624394
rect 340218 624360 340284 624394
rect 340318 624360 340384 624394
rect 340418 624360 340484 624394
rect 340518 624360 340584 624394
rect 340618 624360 340684 624394
rect 340718 624360 340788 624394
rect 334944 624294 340788 624360
rect 334944 624260 335032 624294
rect 335066 624260 335132 624294
rect 335166 624260 335232 624294
rect 335266 624260 335332 624294
rect 335366 624260 335432 624294
rect 335466 624260 335532 624294
rect 335566 624260 336320 624294
rect 336354 624260 336420 624294
rect 336454 624260 336520 624294
rect 336554 624260 336620 624294
rect 336654 624260 336720 624294
rect 336754 624260 336820 624294
rect 336854 624260 337608 624294
rect 337642 624260 337708 624294
rect 337742 624260 337808 624294
rect 337842 624260 337908 624294
rect 337942 624260 338008 624294
rect 338042 624260 338108 624294
rect 338142 624260 338896 624294
rect 338930 624260 338996 624294
rect 339030 624260 339096 624294
rect 339130 624260 339196 624294
rect 339230 624260 339296 624294
rect 339330 624260 339396 624294
rect 339430 624260 340184 624294
rect 340218 624260 340284 624294
rect 340318 624260 340384 624294
rect 340418 624260 340484 624294
rect 340518 624260 340584 624294
rect 340618 624260 340684 624294
rect 340718 624260 340788 624294
rect 334944 623642 340788 624260
rect 334944 623506 337458 623642
rect 334944 623472 335032 623506
rect 335066 623472 335132 623506
rect 335166 623472 335232 623506
rect 335266 623472 335332 623506
rect 335366 623472 335432 623506
rect 335466 623472 335532 623506
rect 335566 623472 336320 623506
rect 336354 623472 336420 623506
rect 336454 623472 336520 623506
rect 336554 623472 336620 623506
rect 336654 623472 336720 623506
rect 336754 623472 336820 623506
rect 336854 623472 337458 623506
rect 334944 623406 337458 623472
rect 334944 623372 335032 623406
rect 335066 623372 335132 623406
rect 335166 623372 335232 623406
rect 335266 623372 335332 623406
rect 335366 623372 335432 623406
rect 335466 623372 335532 623406
rect 335566 623372 336320 623406
rect 336354 623372 336420 623406
rect 336454 623372 336520 623406
rect 336554 623372 336620 623406
rect 336654 623372 336720 623406
rect 336754 623372 336820 623406
rect 336854 623372 337458 623406
rect 334944 623306 337458 623372
rect 334944 623272 335032 623306
rect 335066 623272 335132 623306
rect 335166 623272 335232 623306
rect 335266 623272 335332 623306
rect 335366 623272 335432 623306
rect 335466 623272 335532 623306
rect 335566 623272 336320 623306
rect 336354 623272 336420 623306
rect 336454 623272 336520 623306
rect 336554 623272 336620 623306
rect 336654 623272 336720 623306
rect 336754 623272 336820 623306
rect 336854 623272 337458 623306
rect 334944 623206 337458 623272
rect 334944 623172 335032 623206
rect 335066 623172 335132 623206
rect 335166 623172 335232 623206
rect 335266 623172 335332 623206
rect 335366 623172 335432 623206
rect 335466 623172 335532 623206
rect 335566 623172 336320 623206
rect 336354 623172 336420 623206
rect 336454 623172 336520 623206
rect 336554 623172 336620 623206
rect 336654 623172 336720 623206
rect 336754 623172 336820 623206
rect 336854 623172 337458 623206
rect 334944 623106 337458 623172
rect 334944 623072 335032 623106
rect 335066 623072 335132 623106
rect 335166 623072 335232 623106
rect 335266 623072 335332 623106
rect 335366 623072 335432 623106
rect 335466 623072 335532 623106
rect 335566 623072 336320 623106
rect 336354 623072 336420 623106
rect 336454 623072 336520 623106
rect 336554 623072 336620 623106
rect 336654 623072 336720 623106
rect 336754 623072 336820 623106
rect 336854 623072 337458 623106
rect 334944 623006 337458 623072
rect 334944 622972 335032 623006
rect 335066 622972 335132 623006
rect 335166 622972 335232 623006
rect 335266 622972 335332 623006
rect 335366 622972 335432 623006
rect 335466 622972 335532 623006
rect 335566 622972 336320 623006
rect 336354 622972 336420 623006
rect 336454 622972 336520 623006
rect 336554 622972 336620 623006
rect 336654 622972 336720 623006
rect 336754 622972 336820 623006
rect 336854 622972 337458 623006
rect 331482 617732 331488 618668
rect 332424 617732 332430 618668
rect 331482 617726 332430 617732
rect 334944 622824 337458 622972
rect 337516 623578 338220 623584
rect 337516 622886 337522 623578
rect 338214 622886 338220 623578
rect 337516 622880 338220 622886
rect 338278 623506 340788 623642
rect 338278 623472 338896 623506
rect 338930 623472 338996 623506
rect 339030 623472 339096 623506
rect 339130 623472 339196 623506
rect 339230 623472 339296 623506
rect 339330 623472 339396 623506
rect 339430 623472 340184 623506
rect 340218 623472 340284 623506
rect 340318 623472 340384 623506
rect 340418 623472 340484 623506
rect 340518 623472 340584 623506
rect 340618 623472 340684 623506
rect 340718 623472 340788 623506
rect 338278 623406 340788 623472
rect 338278 623372 338896 623406
rect 338930 623372 338996 623406
rect 339030 623372 339096 623406
rect 339130 623372 339196 623406
rect 339230 623372 339296 623406
rect 339330 623372 339396 623406
rect 339430 623372 340184 623406
rect 340218 623372 340284 623406
rect 340318 623372 340384 623406
rect 340418 623372 340484 623406
rect 340518 623372 340584 623406
rect 340618 623372 340684 623406
rect 340718 623372 340788 623406
rect 338278 623306 340788 623372
rect 338278 623272 338896 623306
rect 338930 623272 338996 623306
rect 339030 623272 339096 623306
rect 339130 623272 339196 623306
rect 339230 623272 339296 623306
rect 339330 623272 339396 623306
rect 339430 623272 340184 623306
rect 340218 623272 340284 623306
rect 340318 623272 340384 623306
rect 340418 623272 340484 623306
rect 340518 623272 340584 623306
rect 340618 623272 340684 623306
rect 340718 623272 340788 623306
rect 338278 623206 340788 623272
rect 338278 623172 338896 623206
rect 338930 623172 338996 623206
rect 339030 623172 339096 623206
rect 339130 623172 339196 623206
rect 339230 623172 339296 623206
rect 339330 623172 339396 623206
rect 339430 623172 340184 623206
rect 340218 623172 340284 623206
rect 340318 623172 340384 623206
rect 340418 623172 340484 623206
rect 340518 623172 340584 623206
rect 340618 623172 340684 623206
rect 340718 623172 340788 623206
rect 338278 623106 340788 623172
rect 338278 623072 338896 623106
rect 338930 623072 338996 623106
rect 339030 623072 339096 623106
rect 339130 623072 339196 623106
rect 339230 623072 339296 623106
rect 339330 623072 339396 623106
rect 339430 623072 340184 623106
rect 340218 623072 340284 623106
rect 340318 623072 340384 623106
rect 340418 623072 340484 623106
rect 340518 623072 340584 623106
rect 340618 623072 340684 623106
rect 340718 623072 340788 623106
rect 338278 623006 340788 623072
rect 338278 622972 338896 623006
rect 338930 622972 338996 623006
rect 339030 622972 339096 623006
rect 339130 622972 339196 623006
rect 339230 622972 339296 623006
rect 339330 622972 339396 623006
rect 339430 622972 340184 623006
rect 340218 622972 340284 623006
rect 340318 622972 340384 623006
rect 340418 622972 340484 623006
rect 340518 622972 340584 623006
rect 340618 622972 340684 623006
rect 340718 622972 340788 623006
rect 338278 622824 340788 622972
rect 334944 622218 340788 622824
rect 334944 622184 335032 622218
rect 335066 622184 335132 622218
rect 335166 622184 335232 622218
rect 335266 622184 335332 622218
rect 335366 622184 335432 622218
rect 335466 622184 335532 622218
rect 335566 622184 336320 622218
rect 336354 622184 336420 622218
rect 336454 622184 336520 622218
rect 336554 622184 336620 622218
rect 336654 622184 336720 622218
rect 336754 622184 336820 622218
rect 336854 622184 337608 622218
rect 337642 622184 337708 622218
rect 337742 622184 337808 622218
rect 337842 622184 337908 622218
rect 337942 622184 338008 622218
rect 338042 622184 338108 622218
rect 338142 622184 338896 622218
rect 338930 622184 338996 622218
rect 339030 622184 339096 622218
rect 339130 622184 339196 622218
rect 339230 622184 339296 622218
rect 339330 622184 339396 622218
rect 339430 622184 340184 622218
rect 340218 622184 340284 622218
rect 340318 622184 340384 622218
rect 340418 622184 340484 622218
rect 340518 622184 340584 622218
rect 340618 622184 340684 622218
rect 340718 622184 340788 622218
rect 334944 622118 340788 622184
rect 334944 622084 335032 622118
rect 335066 622084 335132 622118
rect 335166 622084 335232 622118
rect 335266 622084 335332 622118
rect 335366 622084 335432 622118
rect 335466 622084 335532 622118
rect 335566 622084 336320 622118
rect 336354 622084 336420 622118
rect 336454 622084 336520 622118
rect 336554 622084 336620 622118
rect 336654 622084 336720 622118
rect 336754 622084 336820 622118
rect 336854 622084 337608 622118
rect 337642 622084 337708 622118
rect 337742 622084 337808 622118
rect 337842 622084 337908 622118
rect 337942 622084 338008 622118
rect 338042 622084 338108 622118
rect 338142 622084 338896 622118
rect 338930 622084 338996 622118
rect 339030 622084 339096 622118
rect 339130 622084 339196 622118
rect 339230 622084 339296 622118
rect 339330 622084 339396 622118
rect 339430 622084 340184 622118
rect 340218 622084 340284 622118
rect 340318 622084 340384 622118
rect 340418 622084 340484 622118
rect 340518 622084 340584 622118
rect 340618 622084 340684 622118
rect 340718 622084 340788 622118
rect 334944 622018 340788 622084
rect 334944 621984 335032 622018
rect 335066 621984 335132 622018
rect 335166 621984 335232 622018
rect 335266 621984 335332 622018
rect 335366 621984 335432 622018
rect 335466 621984 335532 622018
rect 335566 621984 336320 622018
rect 336354 621984 336420 622018
rect 336454 621984 336520 622018
rect 336554 621984 336620 622018
rect 336654 621984 336720 622018
rect 336754 621984 336820 622018
rect 336854 621984 337608 622018
rect 337642 621984 337708 622018
rect 337742 621984 337808 622018
rect 337842 621984 337908 622018
rect 337942 621984 338008 622018
rect 338042 621984 338108 622018
rect 338142 621984 338896 622018
rect 338930 621984 338996 622018
rect 339030 621984 339096 622018
rect 339130 621984 339196 622018
rect 339230 621984 339296 622018
rect 339330 621984 339396 622018
rect 339430 621984 340184 622018
rect 340218 621984 340284 622018
rect 340318 621984 340384 622018
rect 340418 621984 340484 622018
rect 340518 621984 340584 622018
rect 340618 621984 340684 622018
rect 340718 621984 340788 622018
rect 334944 621918 340788 621984
rect 334944 621884 335032 621918
rect 335066 621884 335132 621918
rect 335166 621884 335232 621918
rect 335266 621884 335332 621918
rect 335366 621884 335432 621918
rect 335466 621884 335532 621918
rect 335566 621884 336320 621918
rect 336354 621884 336420 621918
rect 336454 621884 336520 621918
rect 336554 621884 336620 621918
rect 336654 621884 336720 621918
rect 336754 621884 336820 621918
rect 336854 621884 337608 621918
rect 337642 621884 337708 621918
rect 337742 621884 337808 621918
rect 337842 621884 337908 621918
rect 337942 621884 338008 621918
rect 338042 621884 338108 621918
rect 338142 621884 338896 621918
rect 338930 621884 338996 621918
rect 339030 621884 339096 621918
rect 339130 621884 339196 621918
rect 339230 621884 339296 621918
rect 339330 621884 339396 621918
rect 339430 621884 340184 621918
rect 340218 621884 340284 621918
rect 340318 621884 340384 621918
rect 340418 621884 340484 621918
rect 340518 621884 340584 621918
rect 340618 621884 340684 621918
rect 340718 621884 340788 621918
rect 334944 621818 340788 621884
rect 334944 621784 335032 621818
rect 335066 621784 335132 621818
rect 335166 621784 335232 621818
rect 335266 621784 335332 621818
rect 335366 621784 335432 621818
rect 335466 621784 335532 621818
rect 335566 621784 336320 621818
rect 336354 621784 336420 621818
rect 336454 621784 336520 621818
rect 336554 621784 336620 621818
rect 336654 621784 336720 621818
rect 336754 621784 336820 621818
rect 336854 621784 337608 621818
rect 337642 621784 337708 621818
rect 337742 621784 337808 621818
rect 337842 621784 337908 621818
rect 337942 621784 338008 621818
rect 338042 621784 338108 621818
rect 338142 621784 338896 621818
rect 338930 621784 338996 621818
rect 339030 621784 339096 621818
rect 339130 621784 339196 621818
rect 339230 621784 339296 621818
rect 339330 621784 339396 621818
rect 339430 621784 340184 621818
rect 340218 621784 340284 621818
rect 340318 621784 340384 621818
rect 340418 621784 340484 621818
rect 340518 621784 340584 621818
rect 340618 621784 340684 621818
rect 340718 621784 340788 621818
rect 334944 621718 340788 621784
rect 334944 621684 335032 621718
rect 335066 621684 335132 621718
rect 335166 621684 335232 621718
rect 335266 621684 335332 621718
rect 335366 621684 335432 621718
rect 335466 621684 335532 621718
rect 335566 621684 336320 621718
rect 336354 621684 336420 621718
rect 336454 621684 336520 621718
rect 336554 621684 336620 621718
rect 336654 621684 336720 621718
rect 336754 621684 336820 621718
rect 336854 621684 337608 621718
rect 337642 621684 337708 621718
rect 337742 621684 337808 621718
rect 337842 621684 337908 621718
rect 337942 621684 338008 621718
rect 338042 621684 338108 621718
rect 338142 621684 338896 621718
rect 338930 621684 338996 621718
rect 339030 621684 339096 621718
rect 339130 621684 339196 621718
rect 339230 621684 339296 621718
rect 339330 621684 339396 621718
rect 339430 621684 340184 621718
rect 340218 621684 340284 621718
rect 340318 621684 340384 621718
rect 340418 621684 340484 621718
rect 340518 621684 340584 621718
rect 340618 621684 340684 621718
rect 340718 621684 340788 621718
rect 334944 620930 340788 621684
rect 334944 620896 335032 620930
rect 335066 620896 335132 620930
rect 335166 620896 335232 620930
rect 335266 620896 335332 620930
rect 335366 620896 335432 620930
rect 335466 620896 335532 620930
rect 335566 620896 336320 620930
rect 336354 620896 336420 620930
rect 336454 620896 336520 620930
rect 336554 620896 336620 620930
rect 336654 620896 336720 620930
rect 336754 620896 336820 620930
rect 336854 620896 337608 620930
rect 337642 620896 337708 620930
rect 337742 620896 337808 620930
rect 337842 620896 337908 620930
rect 337942 620896 338008 620930
rect 338042 620896 338108 620930
rect 338142 620896 338896 620930
rect 338930 620896 338996 620930
rect 339030 620896 339096 620930
rect 339130 620896 339196 620930
rect 339230 620896 339296 620930
rect 339330 620896 339396 620930
rect 339430 620896 340184 620930
rect 340218 620896 340284 620930
rect 340318 620896 340384 620930
rect 340418 620896 340484 620930
rect 340518 620896 340584 620930
rect 340618 620896 340684 620930
rect 340718 620896 340788 620930
rect 334944 620830 340788 620896
rect 334944 620796 335032 620830
rect 335066 620796 335132 620830
rect 335166 620796 335232 620830
rect 335266 620796 335332 620830
rect 335366 620796 335432 620830
rect 335466 620796 335532 620830
rect 335566 620796 336320 620830
rect 336354 620796 336420 620830
rect 336454 620796 336520 620830
rect 336554 620796 336620 620830
rect 336654 620796 336720 620830
rect 336754 620796 336820 620830
rect 336854 620796 337608 620830
rect 337642 620796 337708 620830
rect 337742 620796 337808 620830
rect 337842 620796 337908 620830
rect 337942 620796 338008 620830
rect 338042 620796 338108 620830
rect 338142 620796 338896 620830
rect 338930 620796 338996 620830
rect 339030 620796 339096 620830
rect 339130 620796 339196 620830
rect 339230 620796 339296 620830
rect 339330 620796 339396 620830
rect 339430 620796 340184 620830
rect 340218 620796 340284 620830
rect 340318 620796 340384 620830
rect 340418 620796 340484 620830
rect 340518 620796 340584 620830
rect 340618 620796 340684 620830
rect 340718 620796 340788 620830
rect 334944 620730 340788 620796
rect 334944 620696 335032 620730
rect 335066 620696 335132 620730
rect 335166 620696 335232 620730
rect 335266 620696 335332 620730
rect 335366 620696 335432 620730
rect 335466 620696 335532 620730
rect 335566 620696 336320 620730
rect 336354 620696 336420 620730
rect 336454 620696 336520 620730
rect 336554 620696 336620 620730
rect 336654 620696 336720 620730
rect 336754 620696 336820 620730
rect 336854 620696 337608 620730
rect 337642 620696 337708 620730
rect 337742 620696 337808 620730
rect 337842 620696 337908 620730
rect 337942 620696 338008 620730
rect 338042 620696 338108 620730
rect 338142 620696 338896 620730
rect 338930 620696 338996 620730
rect 339030 620696 339096 620730
rect 339130 620696 339196 620730
rect 339230 620696 339296 620730
rect 339330 620696 339396 620730
rect 339430 620696 340184 620730
rect 340218 620696 340284 620730
rect 340318 620696 340384 620730
rect 340418 620696 340484 620730
rect 340518 620696 340584 620730
rect 340618 620696 340684 620730
rect 340718 620696 340788 620730
rect 334944 620630 340788 620696
rect 334944 620596 335032 620630
rect 335066 620596 335132 620630
rect 335166 620596 335232 620630
rect 335266 620596 335332 620630
rect 335366 620596 335432 620630
rect 335466 620596 335532 620630
rect 335566 620596 336320 620630
rect 336354 620596 336420 620630
rect 336454 620596 336520 620630
rect 336554 620596 336620 620630
rect 336654 620596 336720 620630
rect 336754 620596 336820 620630
rect 336854 620596 337608 620630
rect 337642 620596 337708 620630
rect 337742 620596 337808 620630
rect 337842 620596 337908 620630
rect 337942 620596 338008 620630
rect 338042 620596 338108 620630
rect 338142 620596 338896 620630
rect 338930 620596 338996 620630
rect 339030 620596 339096 620630
rect 339130 620596 339196 620630
rect 339230 620596 339296 620630
rect 339330 620596 339396 620630
rect 339430 620596 340184 620630
rect 340218 620596 340284 620630
rect 340318 620596 340384 620630
rect 340418 620596 340484 620630
rect 340518 620596 340584 620630
rect 340618 620596 340684 620630
rect 340718 620596 340788 620630
rect 334944 620530 340788 620596
rect 334944 620496 335032 620530
rect 335066 620496 335132 620530
rect 335166 620496 335232 620530
rect 335266 620496 335332 620530
rect 335366 620496 335432 620530
rect 335466 620496 335532 620530
rect 335566 620496 336320 620530
rect 336354 620496 336420 620530
rect 336454 620496 336520 620530
rect 336554 620496 336620 620530
rect 336654 620496 336720 620530
rect 336754 620496 336820 620530
rect 336854 620496 337608 620530
rect 337642 620496 337708 620530
rect 337742 620496 337808 620530
rect 337842 620496 337908 620530
rect 337942 620496 338008 620530
rect 338042 620496 338108 620530
rect 338142 620496 338896 620530
rect 338930 620496 338996 620530
rect 339030 620496 339096 620530
rect 339130 620496 339196 620530
rect 339230 620496 339296 620530
rect 339330 620496 339396 620530
rect 339430 620496 340184 620530
rect 340218 620496 340284 620530
rect 340318 620496 340384 620530
rect 340418 620496 340484 620530
rect 340518 620496 340584 620530
rect 340618 620496 340684 620530
rect 340718 620496 340788 620530
rect 334944 620430 340788 620496
rect 334944 620396 335032 620430
rect 335066 620396 335132 620430
rect 335166 620396 335232 620430
rect 335266 620396 335332 620430
rect 335366 620396 335432 620430
rect 335466 620396 335532 620430
rect 335566 620396 336320 620430
rect 336354 620396 336420 620430
rect 336454 620396 336520 620430
rect 336554 620396 336620 620430
rect 336654 620396 336720 620430
rect 336754 620396 336820 620430
rect 336854 620396 337608 620430
rect 337642 620396 337708 620430
rect 337742 620396 337808 620430
rect 337842 620396 337908 620430
rect 337942 620396 338008 620430
rect 338042 620396 338108 620430
rect 338142 620396 338896 620430
rect 338930 620396 338996 620430
rect 339030 620396 339096 620430
rect 339130 620396 339196 620430
rect 339230 620396 339296 620430
rect 339330 620396 339396 620430
rect 339430 620396 340184 620430
rect 340218 620396 340284 620430
rect 340318 620396 340384 620430
rect 340418 620396 340484 620430
rect 340518 620396 340584 620430
rect 340618 620396 340684 620430
rect 340718 620396 340788 620430
rect 334944 619642 340788 620396
rect 334944 619608 335032 619642
rect 335066 619608 335132 619642
rect 335166 619608 335232 619642
rect 335266 619608 335332 619642
rect 335366 619608 335432 619642
rect 335466 619608 335532 619642
rect 335566 619608 336320 619642
rect 336354 619608 336420 619642
rect 336454 619608 336520 619642
rect 336554 619608 336620 619642
rect 336654 619608 336720 619642
rect 336754 619608 336820 619642
rect 336854 619608 337608 619642
rect 337642 619608 337708 619642
rect 337742 619608 337808 619642
rect 337842 619608 337908 619642
rect 337942 619608 338008 619642
rect 338042 619608 338108 619642
rect 338142 619608 338896 619642
rect 338930 619608 338996 619642
rect 339030 619608 339096 619642
rect 339130 619608 339196 619642
rect 339230 619608 339296 619642
rect 339330 619608 339396 619642
rect 339430 619608 340184 619642
rect 340218 619608 340284 619642
rect 340318 619608 340384 619642
rect 340418 619608 340484 619642
rect 340518 619608 340584 619642
rect 340618 619608 340684 619642
rect 340718 619608 340788 619642
rect 334944 619542 340788 619608
rect 334944 619508 335032 619542
rect 335066 619508 335132 619542
rect 335166 619508 335232 619542
rect 335266 619508 335332 619542
rect 335366 619508 335432 619542
rect 335466 619508 335532 619542
rect 335566 619508 336320 619542
rect 336354 619508 336420 619542
rect 336454 619508 336520 619542
rect 336554 619508 336620 619542
rect 336654 619508 336720 619542
rect 336754 619508 336820 619542
rect 336854 619508 337608 619542
rect 337642 619508 337708 619542
rect 337742 619508 337808 619542
rect 337842 619508 337908 619542
rect 337942 619508 338008 619542
rect 338042 619508 338108 619542
rect 338142 619508 338896 619542
rect 338930 619508 338996 619542
rect 339030 619508 339096 619542
rect 339130 619508 339196 619542
rect 339230 619508 339296 619542
rect 339330 619508 339396 619542
rect 339430 619508 340184 619542
rect 340218 619508 340284 619542
rect 340318 619508 340384 619542
rect 340418 619508 340484 619542
rect 340518 619508 340584 619542
rect 340618 619508 340684 619542
rect 340718 619508 340788 619542
rect 334944 619442 340788 619508
rect 334944 619408 335032 619442
rect 335066 619408 335132 619442
rect 335166 619408 335232 619442
rect 335266 619408 335332 619442
rect 335366 619408 335432 619442
rect 335466 619408 335532 619442
rect 335566 619408 336320 619442
rect 336354 619408 336420 619442
rect 336454 619408 336520 619442
rect 336554 619408 336620 619442
rect 336654 619408 336720 619442
rect 336754 619408 336820 619442
rect 336854 619408 337608 619442
rect 337642 619408 337708 619442
rect 337742 619408 337808 619442
rect 337842 619408 337908 619442
rect 337942 619408 338008 619442
rect 338042 619408 338108 619442
rect 338142 619408 338896 619442
rect 338930 619408 338996 619442
rect 339030 619408 339096 619442
rect 339130 619408 339196 619442
rect 339230 619408 339296 619442
rect 339330 619408 339396 619442
rect 339430 619408 340184 619442
rect 340218 619408 340284 619442
rect 340318 619408 340384 619442
rect 340418 619408 340484 619442
rect 340518 619408 340584 619442
rect 340618 619408 340684 619442
rect 340718 619408 340788 619442
rect 334944 619342 340788 619408
rect 334944 619308 335032 619342
rect 335066 619308 335132 619342
rect 335166 619308 335232 619342
rect 335266 619308 335332 619342
rect 335366 619308 335432 619342
rect 335466 619308 335532 619342
rect 335566 619308 336320 619342
rect 336354 619308 336420 619342
rect 336454 619308 336520 619342
rect 336554 619308 336620 619342
rect 336654 619308 336720 619342
rect 336754 619308 336820 619342
rect 336854 619308 337608 619342
rect 337642 619308 337708 619342
rect 337742 619308 337808 619342
rect 337842 619308 337908 619342
rect 337942 619308 338008 619342
rect 338042 619308 338108 619342
rect 338142 619308 338896 619342
rect 338930 619308 338996 619342
rect 339030 619308 339096 619342
rect 339130 619308 339196 619342
rect 339230 619308 339296 619342
rect 339330 619308 339396 619342
rect 339430 619308 340184 619342
rect 340218 619308 340284 619342
rect 340318 619308 340384 619342
rect 340418 619308 340484 619342
rect 340518 619308 340584 619342
rect 340618 619308 340684 619342
rect 340718 619308 340788 619342
rect 334944 619242 340788 619308
rect 334944 619208 335032 619242
rect 335066 619208 335132 619242
rect 335166 619208 335232 619242
rect 335266 619208 335332 619242
rect 335366 619208 335432 619242
rect 335466 619208 335532 619242
rect 335566 619208 336320 619242
rect 336354 619208 336420 619242
rect 336454 619208 336520 619242
rect 336554 619208 336620 619242
rect 336654 619208 336720 619242
rect 336754 619208 336820 619242
rect 336854 619208 337608 619242
rect 337642 619208 337708 619242
rect 337742 619208 337808 619242
rect 337842 619208 337908 619242
rect 337942 619208 338008 619242
rect 338042 619208 338108 619242
rect 338142 619208 338896 619242
rect 338930 619208 338996 619242
rect 339030 619208 339096 619242
rect 339130 619208 339196 619242
rect 339230 619208 339296 619242
rect 339330 619208 339396 619242
rect 339430 619208 340184 619242
rect 340218 619208 340284 619242
rect 340318 619208 340384 619242
rect 340418 619208 340484 619242
rect 340518 619208 340584 619242
rect 340618 619208 340684 619242
rect 340718 619208 340788 619242
rect 334944 619142 340788 619208
rect 334944 619108 335032 619142
rect 335066 619108 335132 619142
rect 335166 619108 335232 619142
rect 335266 619108 335332 619142
rect 335366 619108 335432 619142
rect 335466 619108 335532 619142
rect 335566 619108 336320 619142
rect 336354 619108 336420 619142
rect 336454 619108 336520 619142
rect 336554 619108 336620 619142
rect 336654 619108 336720 619142
rect 336754 619108 336820 619142
rect 336854 619108 337608 619142
rect 337642 619108 337708 619142
rect 337742 619108 337808 619142
rect 337842 619108 337908 619142
rect 337942 619108 338008 619142
rect 338042 619108 338108 619142
rect 338142 619108 338896 619142
rect 338930 619108 338996 619142
rect 339030 619108 339096 619142
rect 339130 619108 339196 619142
rect 339230 619108 339296 619142
rect 339330 619108 339396 619142
rect 339430 619108 340184 619142
rect 340218 619108 340284 619142
rect 340318 619108 340384 619142
rect 340418 619108 340484 619142
rect 340518 619108 340584 619142
rect 340618 619108 340684 619142
rect 340718 619108 340788 619142
rect 334944 618422 340788 619108
rect 334944 618414 336240 618422
rect 334944 617738 334946 618414
rect 335628 617746 336240 618414
rect 336922 618354 340788 618422
rect 336922 618320 337608 618354
rect 337642 618320 337708 618354
rect 337742 618320 337808 618354
rect 337842 618320 337908 618354
rect 337942 618320 338008 618354
rect 338042 618320 338108 618354
rect 338142 618320 338896 618354
rect 338930 618320 338996 618354
rect 339030 618320 339096 618354
rect 339130 618320 339196 618354
rect 339230 618320 339296 618354
rect 339330 618320 339396 618354
rect 339430 618320 340184 618354
rect 340218 618320 340284 618354
rect 340318 618320 340384 618354
rect 340418 618320 340484 618354
rect 340518 618320 340584 618354
rect 340618 618320 340684 618354
rect 340718 618320 340788 618354
rect 336922 618254 340788 618320
rect 336922 618220 337608 618254
rect 337642 618220 337708 618254
rect 337742 618220 337808 618254
rect 337842 618220 337908 618254
rect 337942 618220 338008 618254
rect 338042 618220 338108 618254
rect 338142 618220 338896 618254
rect 338930 618220 338996 618254
rect 339030 618220 339096 618254
rect 339130 618220 339196 618254
rect 339230 618220 339296 618254
rect 339330 618220 339396 618254
rect 339430 618220 340184 618254
rect 340218 618220 340284 618254
rect 340318 618220 340384 618254
rect 340418 618220 340484 618254
rect 340518 618220 340584 618254
rect 340618 618220 340684 618254
rect 340718 618220 340788 618254
rect 336922 618154 340788 618220
rect 336922 618120 337608 618154
rect 337642 618120 337708 618154
rect 337742 618120 337808 618154
rect 337842 618120 337908 618154
rect 337942 618120 338008 618154
rect 338042 618120 338108 618154
rect 338142 618120 338896 618154
rect 338930 618120 338996 618154
rect 339030 618120 339096 618154
rect 339130 618120 339196 618154
rect 339230 618120 339296 618154
rect 339330 618120 339396 618154
rect 339430 618120 340184 618154
rect 340218 618120 340284 618154
rect 340318 618120 340384 618154
rect 340418 618120 340484 618154
rect 340518 618120 340584 618154
rect 340618 618120 340684 618154
rect 340718 618120 340788 618154
rect 336922 618054 340788 618120
rect 336922 618020 337608 618054
rect 337642 618020 337708 618054
rect 337742 618020 337808 618054
rect 337842 618020 337908 618054
rect 337942 618020 338008 618054
rect 338042 618020 338108 618054
rect 338142 618020 338896 618054
rect 338930 618020 338996 618054
rect 339030 618020 339096 618054
rect 339130 618020 339196 618054
rect 339230 618020 339296 618054
rect 339330 618020 339396 618054
rect 339430 618020 340184 618054
rect 340218 618020 340284 618054
rect 340318 618020 340384 618054
rect 340418 618020 340484 618054
rect 340518 618020 340584 618054
rect 340618 618020 340684 618054
rect 340718 618020 340788 618054
rect 336922 617954 340788 618020
rect 342100 624596 343158 624606
rect 342100 624496 342130 624596
rect 342230 624496 342354 624596
rect 342454 624496 342578 624596
rect 342678 624496 342802 624596
rect 342902 624496 343026 624596
rect 343126 624496 343158 624596
rect 342100 624372 343158 624496
rect 342100 624272 342130 624372
rect 342230 624272 342354 624372
rect 342454 624272 342578 624372
rect 342678 624272 342802 624372
rect 342902 624272 343026 624372
rect 343126 624272 343158 624372
rect 342100 624148 343158 624272
rect 342100 624048 342130 624148
rect 342230 624048 342354 624148
rect 342454 624048 342578 624148
rect 342678 624048 342802 624148
rect 342902 624048 343026 624148
rect 343126 624048 343158 624148
rect 342100 623924 343158 624048
rect 342100 623824 342130 623924
rect 342230 623824 342354 623924
rect 342454 623824 342578 623924
rect 342678 623824 342802 623924
rect 342902 623824 343026 623924
rect 343126 623824 343158 623924
rect 342100 623700 343158 623824
rect 342100 623600 342130 623700
rect 342230 623600 342354 623700
rect 342454 623600 342578 623700
rect 342678 623600 342802 623700
rect 342902 623600 343026 623700
rect 343126 623600 343158 623700
rect 342100 623476 343158 623600
rect 342100 623376 342130 623476
rect 342230 623376 342354 623476
rect 342454 623376 342578 623476
rect 342678 623376 342802 623476
rect 342902 623376 343026 623476
rect 343126 623376 343158 623476
rect 342100 623252 343158 623376
rect 342100 623152 342130 623252
rect 342230 623152 342354 623252
rect 342454 623152 342578 623252
rect 342678 623152 342802 623252
rect 342902 623152 343026 623252
rect 343126 623152 343158 623252
rect 342100 623028 343158 623152
rect 342100 622928 342130 623028
rect 342230 622928 342354 623028
rect 342454 622928 342578 623028
rect 342678 622928 342802 623028
rect 342902 622928 343026 623028
rect 343126 622928 343158 623028
rect 342100 622804 343158 622928
rect 342100 622704 342130 622804
rect 342230 622704 342354 622804
rect 342454 622704 342578 622804
rect 342678 622704 342802 622804
rect 342902 622704 343026 622804
rect 343126 622704 343158 622804
rect 342100 622580 343158 622704
rect 342100 622480 342130 622580
rect 342230 622480 342354 622580
rect 342454 622480 342578 622580
rect 342678 622480 342802 622580
rect 342902 622480 343026 622580
rect 343126 622480 343158 622580
rect 342100 622356 343158 622480
rect 342100 622256 342130 622356
rect 342230 622256 342354 622356
rect 342454 622256 342578 622356
rect 342678 622256 342802 622356
rect 342902 622256 343026 622356
rect 343126 622256 343158 622356
rect 342100 622132 343158 622256
rect 342100 622032 342130 622132
rect 342230 622032 342354 622132
rect 342454 622032 342578 622132
rect 342678 622032 342802 622132
rect 342902 622032 343026 622132
rect 343126 622032 343158 622132
rect 342100 621908 343158 622032
rect 342100 621808 342130 621908
rect 342230 621808 342354 621908
rect 342454 621808 342578 621908
rect 342678 621808 342802 621908
rect 342902 621808 343026 621908
rect 343126 621808 343158 621908
rect 342100 621684 343158 621808
rect 342100 621584 342130 621684
rect 342230 621584 342354 621684
rect 342454 621584 342578 621684
rect 342678 621584 342802 621684
rect 342902 621584 343026 621684
rect 343126 621584 343158 621684
rect 342100 621460 343158 621584
rect 342100 621360 342130 621460
rect 342230 621360 342354 621460
rect 342454 621360 342578 621460
rect 342678 621360 342802 621460
rect 342902 621360 343026 621460
rect 343126 621360 343158 621460
rect 342100 621236 343158 621360
rect 342100 621136 342130 621236
rect 342230 621136 342354 621236
rect 342454 621136 342578 621236
rect 342678 621136 342802 621236
rect 342902 621136 343026 621236
rect 343126 621136 343158 621236
rect 342100 621012 343158 621136
rect 342100 620912 342130 621012
rect 342230 620912 342354 621012
rect 342454 620912 342578 621012
rect 342678 620912 342802 621012
rect 342902 620912 343026 621012
rect 343126 620912 343158 621012
rect 342100 620788 343158 620912
rect 342100 620688 342130 620788
rect 342230 620688 342354 620788
rect 342454 620688 342578 620788
rect 342678 620688 342802 620788
rect 342902 620688 343026 620788
rect 343126 620688 343158 620788
rect 342100 620564 343158 620688
rect 342100 620464 342130 620564
rect 342230 620464 342354 620564
rect 342454 620464 342578 620564
rect 342678 620464 342802 620564
rect 342902 620464 343026 620564
rect 343126 620464 343158 620564
rect 342100 620340 343158 620464
rect 342100 620240 342130 620340
rect 342230 620240 342354 620340
rect 342454 620240 342578 620340
rect 342678 620240 342802 620340
rect 342902 620240 343026 620340
rect 343126 620240 343158 620340
rect 342100 620116 343158 620240
rect 342100 620016 342130 620116
rect 342230 620016 342354 620116
rect 342454 620016 342578 620116
rect 342678 620016 342802 620116
rect 342902 620016 343026 620116
rect 343126 620016 343158 620116
rect 342100 619892 343158 620016
rect 342100 619792 342130 619892
rect 342230 619792 342354 619892
rect 342454 619792 342578 619892
rect 342678 619792 342802 619892
rect 342902 619792 343026 619892
rect 343126 619792 343158 619892
rect 342100 619668 343158 619792
rect 342100 619568 342130 619668
rect 342230 619568 342354 619668
rect 342454 619568 342578 619668
rect 342678 619568 342802 619668
rect 342902 619568 343026 619668
rect 343126 619568 343158 619668
rect 342100 619444 343158 619568
rect 342100 619344 342130 619444
rect 342230 619344 342354 619444
rect 342454 619344 342578 619444
rect 342678 619344 342802 619444
rect 342902 619344 343026 619444
rect 343126 619344 343158 619444
rect 342100 619220 343158 619344
rect 342100 619120 342130 619220
rect 342230 619120 342354 619220
rect 342454 619120 342578 619220
rect 342678 619120 342802 619220
rect 342902 619120 343026 619220
rect 343126 619120 343158 619220
rect 342100 618996 343158 619120
rect 342100 618896 342130 618996
rect 342230 618896 342354 618996
rect 342454 618896 342578 618996
rect 342678 618896 342802 618996
rect 342902 618896 343026 618996
rect 343126 618896 343158 618996
rect 342100 618772 343158 618896
rect 342100 618672 342130 618772
rect 342230 618672 342354 618772
rect 342454 618672 342578 618772
rect 342678 618672 342802 618772
rect 342902 618672 343026 618772
rect 343126 618672 343158 618772
rect 342100 618548 343158 618672
rect 342100 618448 342130 618548
rect 342230 618448 342354 618548
rect 342454 618448 342578 618548
rect 342678 618448 342802 618548
rect 342902 618448 343026 618548
rect 343126 618448 343158 618548
rect 342100 618324 343158 618448
rect 342100 618224 342130 618324
rect 342230 618224 342354 618324
rect 342454 618224 342578 618324
rect 342678 618224 342802 618324
rect 342902 618224 343026 618324
rect 343126 618224 343158 618324
rect 342100 618100 343158 618224
rect 342100 618000 342130 618100
rect 342230 618000 342354 618100
rect 342454 618000 342578 618100
rect 342678 618000 342802 618100
rect 342902 618000 343026 618100
rect 343126 618000 343158 618100
rect 342100 617980 343158 618000
rect 336922 617920 337608 617954
rect 337642 617920 337708 617954
rect 337742 617920 337808 617954
rect 337842 617920 337908 617954
rect 337942 617920 338008 617954
rect 338042 617920 338108 617954
rect 338142 617920 338896 617954
rect 338930 617920 338996 617954
rect 339030 617920 339096 617954
rect 339130 617920 339196 617954
rect 339230 617920 339296 617954
rect 339330 617920 339396 617954
rect 339430 617920 340184 617954
rect 340218 617920 340284 617954
rect 340318 617920 340384 617954
rect 340418 617920 340484 617954
rect 340518 617920 340584 617954
rect 340618 617920 340684 617954
rect 340718 617920 340788 617954
rect 336922 617854 340788 617920
rect 336922 617820 337608 617854
rect 337642 617820 337708 617854
rect 337742 617820 337808 617854
rect 337842 617820 337908 617854
rect 337942 617820 338008 617854
rect 338042 617820 338108 617854
rect 338142 617820 338896 617854
rect 338930 617820 338996 617854
rect 339030 617820 339096 617854
rect 339130 617820 339196 617854
rect 339230 617820 339296 617854
rect 339330 617820 339396 617854
rect 339430 617820 340184 617854
rect 340218 617820 340284 617854
rect 340318 617820 340384 617854
rect 340418 617820 340484 617854
rect 340518 617820 340584 617854
rect 340618 617820 340684 617854
rect 340718 617820 340788 617854
rect 336922 617746 340788 617820
rect 335628 617738 340788 617746
rect 334944 617724 340788 617738
rect 329154 617165 329334 617168
rect 329894 617166 329940 617218
rect 329126 617159 329334 617165
rect 329126 617125 329138 617159
rect 329322 617125 329334 617159
rect 329126 617119 329334 617125
rect 329154 617028 329334 617119
rect 329154 616908 329174 617028
rect 329314 616908 329334 617028
rect 329154 616888 329334 616908
rect 329482 617159 329940 617166
rect 329482 617125 329596 617159
rect 329780 617125 329940 617159
rect 310442 616744 310514 616754
rect 306524 616686 308978 616702
rect 312704 616708 313856 616808
rect 314274 616828 314394 616848
rect 314274 616748 314294 616828
rect 314374 616748 314394 616828
rect 314274 616728 314394 616748
rect 315194 616828 315314 616848
rect 315194 616748 315214 616828
rect 315294 616748 315314 616828
rect 315194 616728 315314 616748
rect 316114 616828 316234 616848
rect 316114 616748 316134 616828
rect 316214 616748 316234 616828
rect 316114 616728 316234 616748
rect 317034 616828 317154 616848
rect 317034 616748 317054 616828
rect 317134 616748 317154 616828
rect 317034 616728 317154 616748
rect 317954 616828 318074 616848
rect 317954 616748 317974 616828
rect 318054 616748 318074 616828
rect 319774 616828 319894 616848
rect 317954 616728 318074 616748
rect 312704 616608 312804 616708
rect 313204 616608 313856 616708
rect 312704 616508 313856 616608
rect 318614 616708 319214 616808
rect 319774 616748 319794 616828
rect 319874 616748 319894 616828
rect 319774 616728 319894 616748
rect 320694 616828 320814 616848
rect 320694 616748 320714 616828
rect 320794 616748 320814 616828
rect 320694 616728 320814 616748
rect 321614 616828 321734 616848
rect 321614 616748 321634 616828
rect 321714 616748 321734 616828
rect 321614 616728 321734 616748
rect 322534 616828 322654 616848
rect 322534 616748 322554 616828
rect 322634 616748 322654 616828
rect 322534 616728 322654 616748
rect 323454 616828 323574 616848
rect 323454 616748 323474 616828
rect 323554 616748 323574 616828
rect 325274 616828 325394 616848
rect 323454 616728 323574 616748
rect 318614 616608 318714 616708
rect 319114 616608 319214 616708
rect 318614 616508 319214 616608
rect 324114 616708 324714 616808
rect 325274 616748 325294 616828
rect 325374 616748 325394 616828
rect 325274 616728 325394 616748
rect 326194 616828 326314 616848
rect 326194 616748 326214 616828
rect 326294 616748 326314 616828
rect 326194 616728 326314 616748
rect 327114 616828 327234 616848
rect 327114 616748 327134 616828
rect 327214 616748 327234 616828
rect 327114 616728 327234 616748
rect 328034 616828 328154 616848
rect 328034 616748 328054 616828
rect 328134 616748 328154 616828
rect 328034 616728 328154 616748
rect 328954 616828 329074 616848
rect 328954 616748 328974 616828
rect 329054 616748 329074 616828
rect 328954 616728 329074 616748
rect 329482 616806 329940 617125
rect 324114 616608 324214 616708
rect 324614 616608 324714 616708
rect 324114 616508 324714 616608
rect 329482 616706 330670 616806
rect 329482 616606 330170 616706
rect 330570 616606 330670 616706
rect 329482 616506 330670 616606
rect 298836 615474 305496 615504
rect 298836 615374 298876 615474
rect 298976 615374 299100 615474
rect 299200 615374 299324 615474
rect 299424 615374 299548 615474
rect 299648 615374 299772 615474
rect 299872 615374 299996 615474
rect 300096 615374 300220 615474
rect 300320 615374 300444 615474
rect 300544 615374 300668 615474
rect 300768 615374 300892 615474
rect 300992 615374 301116 615474
rect 301216 615374 301340 615474
rect 301440 615374 301564 615474
rect 301664 615374 301788 615474
rect 301888 615374 302012 615474
rect 302112 615374 302236 615474
rect 302336 615374 302460 615474
rect 302560 615374 302684 615474
rect 302784 615374 302908 615474
rect 303008 615374 303132 615474
rect 303232 615374 303356 615474
rect 303456 615374 303580 615474
rect 303680 615374 303804 615474
rect 303904 615374 304028 615474
rect 304128 615374 304252 615474
rect 304352 615374 304476 615474
rect 304576 615374 304700 615474
rect 304800 615374 304924 615474
rect 305024 615374 305148 615474
rect 305248 615374 305372 615474
rect 305472 615374 305496 615474
rect 298836 615250 305496 615374
rect 298836 615150 298876 615250
rect 298976 615150 299100 615250
rect 299200 615150 299324 615250
rect 299424 615150 299548 615250
rect 299648 615150 299772 615250
rect 299872 615150 299996 615250
rect 300096 615150 300220 615250
rect 300320 615150 300444 615250
rect 300544 615150 300668 615250
rect 300768 615150 300892 615250
rect 300992 615150 301116 615250
rect 301216 615150 301340 615250
rect 301440 615150 301564 615250
rect 301664 615150 301788 615250
rect 301888 615150 302012 615250
rect 302112 615150 302236 615250
rect 302336 615150 302460 615250
rect 302560 615150 302684 615250
rect 302784 615150 302908 615250
rect 303008 615150 303132 615250
rect 303232 615150 303356 615250
rect 303456 615150 303580 615250
rect 303680 615150 303804 615250
rect 303904 615150 304028 615250
rect 304128 615150 304252 615250
rect 304352 615150 304476 615250
rect 304576 615150 304700 615250
rect 304800 615150 304924 615250
rect 305024 615150 305148 615250
rect 305248 615150 305372 615250
rect 305472 615150 305496 615250
rect 298836 615026 305496 615150
rect 298836 614926 298876 615026
rect 298976 614926 299100 615026
rect 299200 614926 299324 615026
rect 299424 614926 299548 615026
rect 299648 614926 299772 615026
rect 299872 614926 299996 615026
rect 300096 614926 300220 615026
rect 300320 614926 300444 615026
rect 300544 614926 300668 615026
rect 300768 614926 300892 615026
rect 300992 614926 301116 615026
rect 301216 614926 301340 615026
rect 301440 614926 301564 615026
rect 301664 614926 301788 615026
rect 301888 614926 302012 615026
rect 302112 614926 302236 615026
rect 302336 614926 302460 615026
rect 302560 614926 302684 615026
rect 302784 614926 302908 615026
rect 303008 614926 303132 615026
rect 303232 614926 303356 615026
rect 303456 614926 303580 615026
rect 303680 614926 303804 615026
rect 303904 614926 304028 615026
rect 304128 614926 304252 615026
rect 304352 614926 304476 615026
rect 304576 614926 304700 615026
rect 304800 614926 304924 615026
rect 305024 614926 305148 615026
rect 305248 614926 305372 615026
rect 305472 614926 305496 615026
rect 298836 614802 305496 614926
rect 298836 614702 298876 614802
rect 298976 614702 299100 614802
rect 299200 614702 299324 614802
rect 299424 614702 299548 614802
rect 299648 614702 299772 614802
rect 299872 614702 299996 614802
rect 300096 614702 300220 614802
rect 300320 614702 300444 614802
rect 300544 614702 300668 614802
rect 300768 614702 300892 614802
rect 300992 614702 301116 614802
rect 301216 614702 301340 614802
rect 301440 614702 301564 614802
rect 301664 614702 301788 614802
rect 301888 614702 302012 614802
rect 302112 614702 302236 614802
rect 302336 614702 302460 614802
rect 302560 614702 302684 614802
rect 302784 614702 302908 614802
rect 303008 614702 303132 614802
rect 303232 614702 303356 614802
rect 303456 614702 303580 614802
rect 303680 614702 303804 614802
rect 303904 614702 304028 614802
rect 304128 614702 304252 614802
rect 304352 614702 304476 614802
rect 304576 614702 304700 614802
rect 304800 614702 304924 614802
rect 305024 614702 305148 614802
rect 305248 614702 305372 614802
rect 305472 614702 305496 614802
rect 298836 614578 305496 614702
rect 298836 614478 298876 614578
rect 298976 614478 299100 614578
rect 299200 614478 299324 614578
rect 299424 614478 299548 614578
rect 299648 614478 299772 614578
rect 299872 614478 299996 614578
rect 300096 614478 300220 614578
rect 300320 614478 300444 614578
rect 300544 614478 300668 614578
rect 300768 614478 300892 614578
rect 300992 614478 301116 614578
rect 301216 614478 301340 614578
rect 301440 614478 301564 614578
rect 301664 614478 301788 614578
rect 301888 614478 302012 614578
rect 302112 614478 302236 614578
rect 302336 614478 302460 614578
rect 302560 614478 302684 614578
rect 302784 614478 302908 614578
rect 303008 614478 303132 614578
rect 303232 614478 303356 614578
rect 303456 614478 303580 614578
rect 303680 614478 303804 614578
rect 303904 614478 304028 614578
rect 304128 614478 304252 614578
rect 304352 614478 304476 614578
rect 304576 614478 304700 614578
rect 304800 614478 304924 614578
rect 305024 614478 305148 614578
rect 305248 614478 305372 614578
rect 305472 614478 305496 614578
rect 298836 614444 305496 614478
rect 309306 615474 315966 615504
rect 309306 615374 309346 615474
rect 309446 615374 309570 615474
rect 309670 615374 309794 615474
rect 309894 615374 310018 615474
rect 310118 615374 310242 615474
rect 310342 615374 310466 615474
rect 310566 615374 310690 615474
rect 310790 615374 310914 615474
rect 311014 615374 311138 615474
rect 311238 615374 311362 615474
rect 311462 615374 311586 615474
rect 311686 615374 311810 615474
rect 311910 615374 312034 615474
rect 312134 615374 312258 615474
rect 312358 615374 312482 615474
rect 312582 615374 312706 615474
rect 312806 615374 312930 615474
rect 313030 615374 313154 615474
rect 313254 615374 313378 615474
rect 313478 615374 313602 615474
rect 313702 615374 313826 615474
rect 313926 615374 314050 615474
rect 314150 615374 314274 615474
rect 314374 615374 314498 615474
rect 314598 615374 314722 615474
rect 314822 615374 314946 615474
rect 315046 615374 315170 615474
rect 315270 615374 315394 615474
rect 315494 615374 315618 615474
rect 315718 615374 315842 615474
rect 315942 615374 315966 615474
rect 309306 615250 315966 615374
rect 309306 615150 309346 615250
rect 309446 615150 309570 615250
rect 309670 615150 309794 615250
rect 309894 615150 310018 615250
rect 310118 615150 310242 615250
rect 310342 615150 310466 615250
rect 310566 615150 310690 615250
rect 310790 615150 310914 615250
rect 311014 615150 311138 615250
rect 311238 615150 311362 615250
rect 311462 615150 311586 615250
rect 311686 615150 311810 615250
rect 311910 615150 312034 615250
rect 312134 615150 312258 615250
rect 312358 615150 312482 615250
rect 312582 615150 312706 615250
rect 312806 615150 312930 615250
rect 313030 615150 313154 615250
rect 313254 615150 313378 615250
rect 313478 615150 313602 615250
rect 313702 615150 313826 615250
rect 313926 615150 314050 615250
rect 314150 615150 314274 615250
rect 314374 615150 314498 615250
rect 314598 615150 314722 615250
rect 314822 615150 314946 615250
rect 315046 615150 315170 615250
rect 315270 615150 315394 615250
rect 315494 615150 315618 615250
rect 315718 615150 315842 615250
rect 315942 615150 315966 615250
rect 309306 615026 315966 615150
rect 309306 614926 309346 615026
rect 309446 614926 309570 615026
rect 309670 614926 309794 615026
rect 309894 614926 310018 615026
rect 310118 614926 310242 615026
rect 310342 614926 310466 615026
rect 310566 614926 310690 615026
rect 310790 614926 310914 615026
rect 311014 614926 311138 615026
rect 311238 614926 311362 615026
rect 311462 614926 311586 615026
rect 311686 614926 311810 615026
rect 311910 614926 312034 615026
rect 312134 614926 312258 615026
rect 312358 614926 312482 615026
rect 312582 614926 312706 615026
rect 312806 614926 312930 615026
rect 313030 614926 313154 615026
rect 313254 614926 313378 615026
rect 313478 614926 313602 615026
rect 313702 614926 313826 615026
rect 313926 614926 314050 615026
rect 314150 614926 314274 615026
rect 314374 614926 314498 615026
rect 314598 614926 314722 615026
rect 314822 614926 314946 615026
rect 315046 614926 315170 615026
rect 315270 614926 315394 615026
rect 315494 614926 315618 615026
rect 315718 614926 315842 615026
rect 315942 614926 315966 615026
rect 309306 614802 315966 614926
rect 309306 614702 309346 614802
rect 309446 614702 309570 614802
rect 309670 614702 309794 614802
rect 309894 614702 310018 614802
rect 310118 614702 310242 614802
rect 310342 614702 310466 614802
rect 310566 614702 310690 614802
rect 310790 614702 310914 614802
rect 311014 614702 311138 614802
rect 311238 614702 311362 614802
rect 311462 614702 311586 614802
rect 311686 614702 311810 614802
rect 311910 614702 312034 614802
rect 312134 614702 312258 614802
rect 312358 614702 312482 614802
rect 312582 614702 312706 614802
rect 312806 614702 312930 614802
rect 313030 614702 313154 614802
rect 313254 614702 313378 614802
rect 313478 614702 313602 614802
rect 313702 614702 313826 614802
rect 313926 614702 314050 614802
rect 314150 614702 314274 614802
rect 314374 614702 314498 614802
rect 314598 614702 314722 614802
rect 314822 614702 314946 614802
rect 315046 614702 315170 614802
rect 315270 614702 315394 614802
rect 315494 614702 315618 614802
rect 315718 614702 315842 614802
rect 315942 614702 315966 614802
rect 309306 614578 315966 614702
rect 309306 614478 309346 614578
rect 309446 614478 309570 614578
rect 309670 614478 309794 614578
rect 309894 614478 310018 614578
rect 310118 614478 310242 614578
rect 310342 614478 310466 614578
rect 310566 614478 310690 614578
rect 310790 614478 310914 614578
rect 311014 614478 311138 614578
rect 311238 614478 311362 614578
rect 311462 614478 311586 614578
rect 311686 614478 311810 614578
rect 311910 614478 312034 614578
rect 312134 614478 312258 614578
rect 312358 614478 312482 614578
rect 312582 614478 312706 614578
rect 312806 614478 312930 614578
rect 313030 614478 313154 614578
rect 313254 614478 313378 614578
rect 313478 614478 313602 614578
rect 313702 614478 313826 614578
rect 313926 614478 314050 614578
rect 314150 614478 314274 614578
rect 314374 614478 314498 614578
rect 314598 614478 314722 614578
rect 314822 614478 314946 614578
rect 315046 614478 315170 614578
rect 315270 614478 315394 614578
rect 315494 614478 315618 614578
rect 315718 614478 315842 614578
rect 315942 614478 315966 614578
rect 309306 614444 315966 614478
rect 335576 615494 342236 615524
rect 335576 615394 335616 615494
rect 335716 615394 335840 615494
rect 335940 615394 336064 615494
rect 336164 615394 336288 615494
rect 336388 615394 336512 615494
rect 336612 615394 336736 615494
rect 336836 615394 336960 615494
rect 337060 615394 337184 615494
rect 337284 615394 337408 615494
rect 337508 615394 337632 615494
rect 337732 615394 337856 615494
rect 337956 615394 338080 615494
rect 338180 615394 338304 615494
rect 338404 615394 338528 615494
rect 338628 615394 338752 615494
rect 338852 615394 338976 615494
rect 339076 615394 339200 615494
rect 339300 615394 339424 615494
rect 339524 615394 339648 615494
rect 339748 615394 339872 615494
rect 339972 615394 340096 615494
rect 340196 615394 340320 615494
rect 340420 615394 340544 615494
rect 340644 615394 340768 615494
rect 340868 615394 340992 615494
rect 341092 615394 341216 615494
rect 341316 615394 341440 615494
rect 341540 615394 341664 615494
rect 341764 615394 341888 615494
rect 341988 615394 342112 615494
rect 342212 615394 342236 615494
rect 335576 615270 342236 615394
rect 335576 615170 335616 615270
rect 335716 615170 335840 615270
rect 335940 615170 336064 615270
rect 336164 615170 336288 615270
rect 336388 615170 336512 615270
rect 336612 615170 336736 615270
rect 336836 615170 336960 615270
rect 337060 615170 337184 615270
rect 337284 615170 337408 615270
rect 337508 615170 337632 615270
rect 337732 615170 337856 615270
rect 337956 615170 338080 615270
rect 338180 615170 338304 615270
rect 338404 615170 338528 615270
rect 338628 615170 338752 615270
rect 338852 615170 338976 615270
rect 339076 615170 339200 615270
rect 339300 615170 339424 615270
rect 339524 615170 339648 615270
rect 339748 615170 339872 615270
rect 339972 615170 340096 615270
rect 340196 615170 340320 615270
rect 340420 615170 340544 615270
rect 340644 615170 340768 615270
rect 340868 615170 340992 615270
rect 341092 615170 341216 615270
rect 341316 615170 341440 615270
rect 341540 615170 341664 615270
rect 341764 615170 341888 615270
rect 341988 615170 342112 615270
rect 342212 615170 342236 615270
rect 335576 615046 342236 615170
rect 335576 614946 335616 615046
rect 335716 614946 335840 615046
rect 335940 614946 336064 615046
rect 336164 614946 336288 615046
rect 336388 614946 336512 615046
rect 336612 614946 336736 615046
rect 336836 614946 336960 615046
rect 337060 614946 337184 615046
rect 337284 614946 337408 615046
rect 337508 614946 337632 615046
rect 337732 614946 337856 615046
rect 337956 614946 338080 615046
rect 338180 614946 338304 615046
rect 338404 614946 338528 615046
rect 338628 614946 338752 615046
rect 338852 614946 338976 615046
rect 339076 614946 339200 615046
rect 339300 614946 339424 615046
rect 339524 614946 339648 615046
rect 339748 614946 339872 615046
rect 339972 614946 340096 615046
rect 340196 614946 340320 615046
rect 340420 614946 340544 615046
rect 340644 614946 340768 615046
rect 340868 614946 340992 615046
rect 341092 614946 341216 615046
rect 341316 614946 341440 615046
rect 341540 614946 341664 615046
rect 341764 614946 341888 615046
rect 341988 614946 342112 615046
rect 342212 614946 342236 615046
rect 335576 614822 342236 614946
rect 335576 614722 335616 614822
rect 335716 614722 335840 614822
rect 335940 614722 336064 614822
rect 336164 614722 336288 614822
rect 336388 614722 336512 614822
rect 336612 614722 336736 614822
rect 336836 614722 336960 614822
rect 337060 614722 337184 614822
rect 337284 614722 337408 614822
rect 337508 614722 337632 614822
rect 337732 614722 337856 614822
rect 337956 614722 338080 614822
rect 338180 614722 338304 614822
rect 338404 614722 338528 614822
rect 338628 614722 338752 614822
rect 338852 614722 338976 614822
rect 339076 614722 339200 614822
rect 339300 614722 339424 614822
rect 339524 614722 339648 614822
rect 339748 614722 339872 614822
rect 339972 614722 340096 614822
rect 340196 614722 340320 614822
rect 340420 614722 340544 614822
rect 340644 614722 340768 614822
rect 340868 614722 340992 614822
rect 341092 614722 341216 614822
rect 341316 614722 341440 614822
rect 341540 614722 341664 614822
rect 341764 614722 341888 614822
rect 341988 614722 342112 614822
rect 342212 614722 342236 614822
rect 335576 614598 342236 614722
rect 335576 614498 335616 614598
rect 335716 614498 335840 614598
rect 335940 614498 336064 614598
rect 336164 614498 336288 614598
rect 336388 614498 336512 614598
rect 336612 614498 336736 614598
rect 336836 614498 336960 614598
rect 337060 614498 337184 614598
rect 337284 614498 337408 614598
rect 337508 614498 337632 614598
rect 337732 614498 337856 614598
rect 337956 614498 338080 614598
rect 338180 614498 338304 614598
rect 338404 614498 338528 614598
rect 338628 614498 338752 614598
rect 338852 614498 338976 614598
rect 339076 614498 339200 614598
rect 339300 614498 339424 614598
rect 339524 614498 339648 614598
rect 339748 614498 339872 614598
rect 339972 614498 340096 614598
rect 340196 614498 340320 614598
rect 340420 614498 340544 614598
rect 340644 614498 340768 614598
rect 340868 614498 340992 614598
rect 341092 614498 341216 614598
rect 341316 614498 341440 614598
rect 341540 614498 341664 614598
rect 341764 614498 341888 614598
rect 341988 614498 342112 614598
rect 342212 614498 342236 614598
rect 335576 614464 342236 614498
<< via1 >>
rect 298876 642594 298976 642694
rect 299100 642594 299200 642694
rect 299324 642594 299424 642694
rect 299548 642594 299648 642694
rect 299772 642594 299872 642694
rect 299996 642594 300096 642694
rect 300220 642594 300320 642694
rect 300444 642594 300544 642694
rect 300668 642594 300768 642694
rect 300892 642594 300992 642694
rect 301116 642594 301216 642694
rect 301340 642594 301440 642694
rect 301564 642594 301664 642694
rect 301788 642594 301888 642694
rect 302012 642594 302112 642694
rect 302236 642594 302336 642694
rect 302460 642594 302560 642694
rect 302684 642594 302784 642694
rect 302908 642594 303008 642694
rect 303132 642594 303232 642694
rect 303356 642594 303456 642694
rect 303580 642594 303680 642694
rect 303804 642594 303904 642694
rect 304028 642594 304128 642694
rect 304252 642594 304352 642694
rect 304476 642594 304576 642694
rect 304700 642594 304800 642694
rect 304924 642594 305024 642694
rect 305148 642594 305248 642694
rect 305372 642594 305472 642694
rect 298876 642370 298976 642470
rect 299100 642370 299200 642470
rect 299324 642370 299424 642470
rect 299548 642370 299648 642470
rect 299772 642370 299872 642470
rect 299996 642370 300096 642470
rect 300220 642370 300320 642470
rect 300444 642370 300544 642470
rect 300668 642370 300768 642470
rect 300892 642370 300992 642470
rect 301116 642370 301216 642470
rect 301340 642370 301440 642470
rect 301564 642370 301664 642470
rect 301788 642370 301888 642470
rect 302012 642370 302112 642470
rect 302236 642370 302336 642470
rect 302460 642370 302560 642470
rect 302684 642370 302784 642470
rect 302908 642370 303008 642470
rect 303132 642370 303232 642470
rect 303356 642370 303456 642470
rect 303580 642370 303680 642470
rect 303804 642370 303904 642470
rect 304028 642370 304128 642470
rect 304252 642370 304352 642470
rect 304476 642370 304576 642470
rect 304700 642370 304800 642470
rect 304924 642370 305024 642470
rect 305148 642370 305248 642470
rect 305372 642370 305472 642470
rect 298876 642146 298976 642246
rect 299100 642146 299200 642246
rect 299324 642146 299424 642246
rect 299548 642146 299648 642246
rect 299772 642146 299872 642246
rect 299996 642146 300096 642246
rect 300220 642146 300320 642246
rect 300444 642146 300544 642246
rect 300668 642146 300768 642246
rect 300892 642146 300992 642246
rect 301116 642146 301216 642246
rect 301340 642146 301440 642246
rect 301564 642146 301664 642246
rect 301788 642146 301888 642246
rect 302012 642146 302112 642246
rect 302236 642146 302336 642246
rect 302460 642146 302560 642246
rect 302684 642146 302784 642246
rect 302908 642146 303008 642246
rect 303132 642146 303232 642246
rect 303356 642146 303456 642246
rect 303580 642146 303680 642246
rect 303804 642146 303904 642246
rect 304028 642146 304128 642246
rect 304252 642146 304352 642246
rect 304476 642146 304576 642246
rect 304700 642146 304800 642246
rect 304924 642146 305024 642246
rect 305148 642146 305248 642246
rect 305372 642146 305472 642246
rect 298876 641922 298976 642022
rect 299100 641922 299200 642022
rect 299324 641922 299424 642022
rect 299548 641922 299648 642022
rect 299772 641922 299872 642022
rect 299996 641922 300096 642022
rect 300220 641922 300320 642022
rect 300444 641922 300544 642022
rect 300668 641922 300768 642022
rect 300892 641922 300992 642022
rect 301116 641922 301216 642022
rect 301340 641922 301440 642022
rect 301564 641922 301664 642022
rect 301788 641922 301888 642022
rect 302012 641922 302112 642022
rect 302236 641922 302336 642022
rect 302460 641922 302560 642022
rect 302684 641922 302784 642022
rect 302908 641922 303008 642022
rect 303132 641922 303232 642022
rect 303356 641922 303456 642022
rect 303580 641922 303680 642022
rect 303804 641922 303904 642022
rect 304028 641922 304128 642022
rect 304252 641922 304352 642022
rect 304476 641922 304576 642022
rect 304700 641922 304800 642022
rect 304924 641922 305024 642022
rect 305148 641922 305248 642022
rect 305372 641922 305472 642022
rect 298876 641698 298976 641798
rect 299100 641698 299200 641798
rect 299324 641698 299424 641798
rect 299548 641698 299648 641798
rect 299772 641698 299872 641798
rect 299996 641698 300096 641798
rect 300220 641698 300320 641798
rect 300444 641698 300544 641798
rect 300668 641698 300768 641798
rect 300892 641698 300992 641798
rect 301116 641698 301216 641798
rect 301340 641698 301440 641798
rect 301564 641698 301664 641798
rect 301788 641698 301888 641798
rect 302012 641698 302112 641798
rect 302236 641698 302336 641798
rect 302460 641698 302560 641798
rect 302684 641698 302784 641798
rect 302908 641698 303008 641798
rect 303132 641698 303232 641798
rect 303356 641698 303456 641798
rect 303580 641698 303680 641798
rect 303804 641698 303904 641798
rect 304028 641698 304128 641798
rect 304252 641698 304352 641798
rect 304476 641698 304576 641798
rect 304700 641698 304800 641798
rect 304924 641698 305024 641798
rect 305148 641698 305248 641798
rect 305372 641698 305472 641798
rect 309346 642594 309446 642694
rect 309570 642594 309670 642694
rect 309794 642594 309894 642694
rect 310018 642594 310118 642694
rect 310242 642594 310342 642694
rect 310466 642594 310566 642694
rect 310690 642594 310790 642694
rect 310914 642594 311014 642694
rect 311138 642594 311238 642694
rect 311362 642594 311462 642694
rect 311586 642594 311686 642694
rect 311810 642594 311910 642694
rect 312034 642594 312134 642694
rect 312258 642594 312358 642694
rect 312482 642594 312582 642694
rect 312706 642594 312806 642694
rect 312930 642594 313030 642694
rect 313154 642594 313254 642694
rect 313378 642594 313478 642694
rect 313602 642594 313702 642694
rect 313826 642594 313926 642694
rect 314050 642594 314150 642694
rect 314274 642594 314374 642694
rect 314498 642594 314598 642694
rect 314722 642594 314822 642694
rect 314946 642594 315046 642694
rect 315170 642594 315270 642694
rect 315394 642594 315494 642694
rect 315618 642594 315718 642694
rect 315842 642594 315942 642694
rect 309346 642370 309446 642470
rect 309570 642370 309670 642470
rect 309794 642370 309894 642470
rect 310018 642370 310118 642470
rect 310242 642370 310342 642470
rect 310466 642370 310566 642470
rect 310690 642370 310790 642470
rect 310914 642370 311014 642470
rect 311138 642370 311238 642470
rect 311362 642370 311462 642470
rect 311586 642370 311686 642470
rect 311810 642370 311910 642470
rect 312034 642370 312134 642470
rect 312258 642370 312358 642470
rect 312482 642370 312582 642470
rect 312706 642370 312806 642470
rect 312930 642370 313030 642470
rect 313154 642370 313254 642470
rect 313378 642370 313478 642470
rect 313602 642370 313702 642470
rect 313826 642370 313926 642470
rect 314050 642370 314150 642470
rect 314274 642370 314374 642470
rect 314498 642370 314598 642470
rect 314722 642370 314822 642470
rect 314946 642370 315046 642470
rect 315170 642370 315270 642470
rect 315394 642370 315494 642470
rect 315618 642370 315718 642470
rect 315842 642370 315942 642470
rect 309346 642146 309446 642246
rect 309570 642146 309670 642246
rect 309794 642146 309894 642246
rect 310018 642146 310118 642246
rect 310242 642146 310342 642246
rect 310466 642146 310566 642246
rect 310690 642146 310790 642246
rect 310914 642146 311014 642246
rect 311138 642146 311238 642246
rect 311362 642146 311462 642246
rect 311586 642146 311686 642246
rect 311810 642146 311910 642246
rect 312034 642146 312134 642246
rect 312258 642146 312358 642246
rect 312482 642146 312582 642246
rect 312706 642146 312806 642246
rect 312930 642146 313030 642246
rect 313154 642146 313254 642246
rect 313378 642146 313478 642246
rect 313602 642146 313702 642246
rect 313826 642146 313926 642246
rect 314050 642146 314150 642246
rect 314274 642146 314374 642246
rect 314498 642146 314598 642246
rect 314722 642146 314822 642246
rect 314946 642146 315046 642246
rect 315170 642146 315270 642246
rect 315394 642146 315494 642246
rect 315618 642146 315718 642246
rect 315842 642146 315942 642246
rect 309346 641922 309446 642022
rect 309570 641922 309670 642022
rect 309794 641922 309894 642022
rect 310018 641922 310118 642022
rect 310242 641922 310342 642022
rect 310466 641922 310566 642022
rect 310690 641922 310790 642022
rect 310914 641922 311014 642022
rect 311138 641922 311238 642022
rect 311362 641922 311462 642022
rect 311586 641922 311686 642022
rect 311810 641922 311910 642022
rect 312034 641922 312134 642022
rect 312258 641922 312358 642022
rect 312482 641922 312582 642022
rect 312706 641922 312806 642022
rect 312930 641922 313030 642022
rect 313154 641922 313254 642022
rect 313378 641922 313478 642022
rect 313602 641922 313702 642022
rect 313826 641922 313926 642022
rect 314050 641922 314150 642022
rect 314274 641922 314374 642022
rect 314498 641922 314598 642022
rect 314722 641922 314822 642022
rect 314946 641922 315046 642022
rect 315170 641922 315270 642022
rect 315394 641922 315494 642022
rect 315618 641922 315718 642022
rect 315842 641922 315942 642022
rect 309346 641698 309446 641798
rect 309570 641698 309670 641798
rect 309794 641698 309894 641798
rect 310018 641698 310118 641798
rect 310242 641698 310342 641798
rect 310466 641698 310566 641798
rect 310690 641698 310790 641798
rect 310914 641698 311014 641798
rect 311138 641698 311238 641798
rect 311362 641698 311462 641798
rect 311586 641698 311686 641798
rect 311810 641698 311910 641798
rect 312034 641698 312134 641798
rect 312258 641698 312358 641798
rect 312482 641698 312582 641798
rect 312706 641698 312806 641798
rect 312930 641698 313030 641798
rect 313154 641698 313254 641798
rect 313378 641698 313478 641798
rect 313602 641698 313702 641798
rect 313826 641698 313926 641798
rect 314050 641698 314150 641798
rect 314274 641698 314374 641798
rect 314498 641698 314598 641798
rect 314722 641698 314822 641798
rect 314946 641698 315046 641798
rect 315170 641698 315270 641798
rect 315394 641698 315494 641798
rect 315618 641698 315718 641798
rect 315842 641698 315942 641798
rect 335616 642614 335716 642714
rect 335840 642614 335940 642714
rect 336064 642614 336164 642714
rect 336288 642614 336388 642714
rect 336512 642614 336612 642714
rect 336736 642614 336836 642714
rect 336960 642614 337060 642714
rect 337184 642614 337284 642714
rect 337408 642614 337508 642714
rect 337632 642614 337732 642714
rect 337856 642614 337956 642714
rect 338080 642614 338180 642714
rect 338304 642614 338404 642714
rect 338528 642614 338628 642714
rect 338752 642614 338852 642714
rect 338976 642614 339076 642714
rect 339200 642614 339300 642714
rect 339424 642614 339524 642714
rect 339648 642614 339748 642714
rect 339872 642614 339972 642714
rect 340096 642614 340196 642714
rect 340320 642614 340420 642714
rect 340544 642614 340644 642714
rect 340768 642614 340868 642714
rect 340992 642614 341092 642714
rect 341216 642614 341316 642714
rect 341440 642614 341540 642714
rect 341664 642614 341764 642714
rect 341888 642614 341988 642714
rect 342112 642614 342212 642714
rect 335616 642390 335716 642490
rect 335840 642390 335940 642490
rect 336064 642390 336164 642490
rect 336288 642390 336388 642490
rect 336512 642390 336612 642490
rect 336736 642390 336836 642490
rect 336960 642390 337060 642490
rect 337184 642390 337284 642490
rect 337408 642390 337508 642490
rect 337632 642390 337732 642490
rect 337856 642390 337956 642490
rect 338080 642390 338180 642490
rect 338304 642390 338404 642490
rect 338528 642390 338628 642490
rect 338752 642390 338852 642490
rect 338976 642390 339076 642490
rect 339200 642390 339300 642490
rect 339424 642390 339524 642490
rect 339648 642390 339748 642490
rect 339872 642390 339972 642490
rect 340096 642390 340196 642490
rect 340320 642390 340420 642490
rect 340544 642390 340644 642490
rect 340768 642390 340868 642490
rect 340992 642390 341092 642490
rect 341216 642390 341316 642490
rect 341440 642390 341540 642490
rect 341664 642390 341764 642490
rect 341888 642390 341988 642490
rect 342112 642390 342212 642490
rect 335616 642166 335716 642266
rect 335840 642166 335940 642266
rect 336064 642166 336164 642266
rect 336288 642166 336388 642266
rect 336512 642166 336612 642266
rect 336736 642166 336836 642266
rect 336960 642166 337060 642266
rect 337184 642166 337284 642266
rect 337408 642166 337508 642266
rect 337632 642166 337732 642266
rect 337856 642166 337956 642266
rect 338080 642166 338180 642266
rect 338304 642166 338404 642266
rect 338528 642166 338628 642266
rect 338752 642166 338852 642266
rect 338976 642166 339076 642266
rect 339200 642166 339300 642266
rect 339424 642166 339524 642266
rect 339648 642166 339748 642266
rect 339872 642166 339972 642266
rect 340096 642166 340196 642266
rect 340320 642166 340420 642266
rect 340544 642166 340644 642266
rect 340768 642166 340868 642266
rect 340992 642166 341092 642266
rect 341216 642166 341316 642266
rect 341440 642166 341540 642266
rect 341664 642166 341764 642266
rect 341888 642166 341988 642266
rect 342112 642166 342212 642266
rect 335616 641942 335716 642042
rect 335840 641942 335940 642042
rect 336064 641942 336164 642042
rect 336288 641942 336388 642042
rect 336512 641942 336612 642042
rect 336736 641942 336836 642042
rect 336960 641942 337060 642042
rect 337184 641942 337284 642042
rect 337408 641942 337508 642042
rect 337632 641942 337732 642042
rect 337856 641942 337956 642042
rect 338080 641942 338180 642042
rect 338304 641942 338404 642042
rect 338528 641942 338628 642042
rect 338752 641942 338852 642042
rect 338976 641942 339076 642042
rect 339200 641942 339300 642042
rect 339424 641942 339524 642042
rect 339648 641942 339748 642042
rect 339872 641942 339972 642042
rect 340096 641942 340196 642042
rect 340320 641942 340420 642042
rect 340544 641942 340644 642042
rect 340768 641942 340868 642042
rect 340992 641942 341092 642042
rect 341216 641942 341316 642042
rect 341440 641942 341540 642042
rect 341664 641942 341764 642042
rect 341888 641942 341988 642042
rect 342112 641942 342212 642042
rect 335616 641718 335716 641818
rect 335840 641718 335940 641818
rect 336064 641718 336164 641818
rect 336288 641718 336388 641818
rect 336512 641718 336612 641818
rect 336736 641718 336836 641818
rect 336960 641718 337060 641818
rect 337184 641718 337284 641818
rect 337408 641718 337508 641818
rect 337632 641718 337732 641818
rect 337856 641718 337956 641818
rect 338080 641718 338180 641818
rect 338304 641718 338404 641818
rect 338528 641718 338628 641818
rect 338752 641718 338852 641818
rect 338976 641718 339076 641818
rect 339200 641718 339300 641818
rect 339424 641718 339524 641818
rect 339648 641718 339748 641818
rect 339872 641718 339972 641818
rect 340096 641718 340196 641818
rect 340320 641718 340420 641818
rect 340544 641718 340644 641818
rect 340768 641718 340868 641818
rect 340992 641718 341092 641818
rect 341216 641718 341316 641818
rect 341440 641718 341540 641818
rect 341664 641718 341764 641818
rect 341888 641718 341988 641818
rect 342112 641718 342212 641818
rect 300658 640558 311902 640572
rect 300658 639760 300672 640558
rect 300672 639760 311888 640558
rect 311888 639760 311902 640558
rect 300658 639746 311902 639760
rect 323924 638474 324482 639032
rect 325548 638474 326106 639032
rect 329638 638474 330196 639032
rect 332092 638474 332650 639032
rect 297850 637896 297950 637996
rect 298074 637896 298174 637996
rect 298298 637896 298398 637996
rect 298522 637896 298622 637996
rect 298746 637896 298846 637996
rect 297850 637672 297950 637772
rect 298074 637672 298174 637772
rect 298298 637672 298398 637772
rect 298522 637672 298622 637772
rect 298746 637672 298846 637772
rect 317368 637674 317926 638232
rect 323094 637674 323652 638232
rect 326366 637674 326924 638232
rect 328820 637674 329378 638232
rect 331274 637674 331832 638232
rect 333728 637674 334286 638232
rect 342130 637896 342230 637996
rect 342354 637896 342454 637996
rect 342578 637896 342678 637996
rect 342802 637896 342902 637996
rect 343026 637896 343126 637996
rect 342130 637672 342230 637772
rect 342354 637672 342454 637772
rect 342578 637672 342678 637772
rect 342802 637672 342902 637772
rect 343026 637672 343126 637772
rect 297850 637448 297950 637548
rect 298074 637448 298174 637548
rect 298298 637448 298398 637548
rect 298522 637448 298622 637548
rect 298746 637448 298846 637548
rect 297850 637224 297950 637324
rect 298074 637224 298174 637324
rect 298298 637224 298398 637324
rect 298522 637224 298622 637324
rect 298746 637224 298846 637324
rect 297850 637000 297950 637100
rect 298074 637000 298174 637100
rect 298298 637000 298398 637100
rect 298522 637000 298622 637100
rect 298746 637000 298846 637100
rect 317368 637482 317926 637494
rect 317368 637085 317378 637482
rect 317378 637085 317916 637482
rect 317916 637085 317926 637482
rect 317368 637074 317926 637085
rect 318186 637482 318744 637494
rect 318186 637085 318196 637482
rect 318196 637085 318734 637482
rect 318734 637085 318744 637482
rect 318186 637074 318744 637085
rect 342130 637448 342230 637548
rect 342354 637448 342454 637548
rect 342578 637448 342678 637548
rect 342802 637448 342902 637548
rect 343026 637448 343126 637548
rect 322276 637420 322834 637432
rect 322276 637023 322286 637420
rect 322286 637023 322824 637420
rect 322824 637023 322834 637420
rect 322276 637012 322834 637023
rect 323094 637420 323652 637432
rect 323094 637023 323104 637420
rect 323104 637023 323642 637420
rect 323642 637023 323652 637420
rect 323094 637012 323652 637023
rect 323912 637420 324470 637432
rect 323912 637023 323922 637420
rect 323922 637023 324460 637420
rect 324460 637023 324470 637420
rect 323912 637012 324470 637023
rect 324730 637420 325288 637432
rect 324730 637023 324740 637420
rect 324740 637023 325278 637420
rect 325278 637023 325288 637420
rect 324730 637012 325288 637023
rect 325548 637420 326106 637432
rect 325548 637023 325558 637420
rect 325558 637023 326096 637420
rect 326096 637023 326106 637420
rect 325548 637012 326106 637023
rect 326366 637420 326924 637432
rect 326366 637023 326376 637420
rect 326376 637023 326914 637420
rect 326914 637023 326924 637420
rect 326366 637012 326924 637023
rect 327184 637420 327742 637432
rect 327184 637023 327194 637420
rect 327194 637023 327732 637420
rect 327732 637023 327742 637420
rect 327184 637012 327742 637023
rect 328002 637420 328560 637432
rect 328002 637023 328012 637420
rect 328012 637023 328550 637420
rect 328550 637023 328560 637420
rect 328002 637012 328560 637023
rect 328820 637420 329378 637432
rect 328820 637023 328830 637420
rect 328830 637023 329368 637420
rect 329368 637023 329378 637420
rect 328820 637012 329378 637023
rect 329638 637420 330196 637432
rect 329638 637023 329648 637420
rect 329648 637023 330186 637420
rect 330186 637023 330196 637420
rect 329638 637012 330196 637023
rect 330456 637420 331014 637432
rect 330456 637023 330466 637420
rect 330466 637023 331004 637420
rect 331004 637023 331014 637420
rect 330456 637012 331014 637023
rect 331274 637420 331832 637432
rect 331274 637023 331284 637420
rect 331284 637023 331822 637420
rect 331822 637023 331832 637420
rect 331274 637012 331832 637023
rect 332092 637420 332650 637432
rect 332092 637023 332102 637420
rect 332102 637023 332640 637420
rect 332640 637023 332650 637420
rect 332092 637012 332650 637023
rect 332910 637420 333468 637432
rect 332910 637023 332920 637420
rect 332920 637023 333458 637420
rect 333458 637023 333468 637420
rect 332910 637012 333468 637023
rect 333728 637420 334286 637432
rect 333728 637023 333738 637420
rect 333738 637023 334276 637420
rect 334276 637023 334286 637420
rect 333728 637012 334286 637023
rect 342130 637224 342230 637324
rect 342354 637224 342454 637324
rect 342578 637224 342678 637324
rect 342802 637224 342902 637324
rect 343026 637224 343126 637324
rect 297850 636776 297950 636876
rect 298074 636776 298174 636876
rect 298298 636776 298398 636876
rect 298522 636776 298622 636876
rect 298746 636776 298846 636876
rect 342130 637000 342230 637100
rect 342354 637000 342454 637100
rect 342578 637000 342678 637100
rect 342802 637000 342902 637100
rect 343026 637000 343126 637100
rect 342130 636776 342230 636876
rect 342354 636776 342454 636876
rect 342578 636776 342678 636876
rect 342802 636776 342902 636876
rect 343026 636776 343126 636876
rect 297850 636552 297950 636652
rect 298074 636552 298174 636652
rect 298298 636552 298398 636652
rect 298522 636552 298622 636652
rect 298746 636552 298846 636652
rect 297850 636328 297950 636428
rect 298074 636328 298174 636428
rect 298298 636328 298398 636428
rect 298522 636328 298622 636428
rect 298746 636328 298846 636428
rect 318186 636278 318744 636770
rect 322276 636212 322834 636770
rect 324730 636212 325288 636770
rect 327184 636212 327742 636770
rect 330456 636212 331014 636770
rect 332910 636212 333468 636770
rect 342130 636552 342230 636652
rect 342354 636552 342454 636652
rect 342578 636552 342678 636652
rect 342802 636552 342902 636652
rect 343026 636552 343126 636652
rect 342130 636328 342230 636428
rect 342354 636328 342454 636428
rect 342578 636328 342678 636428
rect 342802 636328 342902 636428
rect 343026 636328 343126 636428
rect 297850 636104 297950 636204
rect 298074 636104 298174 636204
rect 298298 636104 298398 636204
rect 298522 636104 298622 636204
rect 298746 636104 298846 636204
rect 342130 636104 342230 636204
rect 342354 636104 342454 636204
rect 342578 636104 342678 636204
rect 342802 636104 342902 636204
rect 343026 636104 343126 636204
rect 297850 635880 297950 635980
rect 298074 635880 298174 635980
rect 298298 635880 298398 635980
rect 298522 635880 298622 635980
rect 298746 635880 298846 635980
rect 297850 635656 297950 635756
rect 298074 635656 298174 635756
rect 298298 635656 298398 635756
rect 298522 635656 298622 635756
rect 298746 635656 298846 635756
rect 342130 635880 342230 635980
rect 342354 635880 342454 635980
rect 342578 635880 342678 635980
rect 342802 635880 342902 635980
rect 343026 635880 343126 635980
rect 297850 635432 297950 635532
rect 298074 635432 298174 635532
rect 298298 635432 298398 635532
rect 298522 635432 298622 635532
rect 298746 635432 298846 635532
rect 297850 635208 297950 635308
rect 298074 635208 298174 635308
rect 298298 635208 298398 635308
rect 298522 635208 298622 635308
rect 298746 635208 298846 635308
rect 297850 634984 297950 635084
rect 298074 634984 298174 635084
rect 298298 634984 298398 635084
rect 298522 634984 298622 635084
rect 298746 634984 298846 635084
rect 297850 634760 297950 634860
rect 298074 634760 298174 634860
rect 298298 634760 298398 634860
rect 298522 634760 298622 634860
rect 298746 634760 298846 634860
rect 297850 634536 297950 634636
rect 298074 634536 298174 634636
rect 298298 634536 298398 634636
rect 298522 634536 298622 634636
rect 298746 634536 298846 634636
rect 297850 634312 297950 634412
rect 298074 634312 298174 634412
rect 298298 634312 298398 634412
rect 298522 634312 298622 634412
rect 298746 634312 298846 634412
rect 297850 634088 297950 634188
rect 298074 634088 298174 634188
rect 298298 634088 298398 634188
rect 298522 634088 298622 634188
rect 298746 634088 298846 634188
rect 297850 633864 297950 633964
rect 298074 633864 298174 633964
rect 298298 633864 298398 633964
rect 298522 633864 298622 633964
rect 298746 633864 298846 633964
rect 297850 633640 297950 633740
rect 298074 633640 298174 633740
rect 298298 633640 298398 633740
rect 298522 633640 298622 633740
rect 298746 633640 298846 633740
rect 297850 633416 297950 633516
rect 298074 633416 298174 633516
rect 298298 633416 298398 633516
rect 298522 633416 298622 633516
rect 298746 633416 298846 633516
rect 297850 633192 297950 633292
rect 298074 633192 298174 633292
rect 298298 633192 298398 633292
rect 298522 633192 298622 633292
rect 298746 633192 298846 633292
rect 297850 632968 297950 633068
rect 298074 632968 298174 633068
rect 298298 632968 298398 633068
rect 298522 632968 298622 633068
rect 298746 632968 298846 633068
rect 297850 632744 297950 632844
rect 298074 632744 298174 632844
rect 298298 632744 298398 632844
rect 298522 632744 298622 632844
rect 298746 632744 298846 632844
rect 342130 635656 342230 635756
rect 342354 635656 342454 635756
rect 342578 635656 342678 635756
rect 342802 635656 342902 635756
rect 343026 635656 343126 635756
rect 342130 635432 342230 635532
rect 342354 635432 342454 635532
rect 342578 635432 342678 635532
rect 342802 635432 342902 635532
rect 343026 635432 343126 635532
rect 342130 635208 342230 635308
rect 342354 635208 342454 635308
rect 342578 635208 342678 635308
rect 342802 635208 342902 635308
rect 343026 635208 343126 635308
rect 342130 634984 342230 635084
rect 342354 634984 342454 635084
rect 342578 634984 342678 635084
rect 342802 634984 342902 635084
rect 343026 634984 343126 635084
rect 342130 634760 342230 634860
rect 342354 634760 342454 634860
rect 342578 634760 342678 634860
rect 342802 634760 342902 634860
rect 343026 634760 343126 634860
rect 342130 634536 342230 634636
rect 342354 634536 342454 634636
rect 342578 634536 342678 634636
rect 342802 634536 342902 634636
rect 343026 634536 343126 634636
rect 342130 634312 342230 634412
rect 342354 634312 342454 634412
rect 342578 634312 342678 634412
rect 342802 634312 342902 634412
rect 343026 634312 343126 634412
rect 342130 634088 342230 634188
rect 342354 634088 342454 634188
rect 342578 634088 342678 634188
rect 342802 634088 342902 634188
rect 343026 634088 343126 634188
rect 342130 633864 342230 633964
rect 342354 633864 342454 633964
rect 342578 633864 342678 633964
rect 342802 633864 342902 633964
rect 343026 633864 343126 633964
rect 342130 633640 342230 633740
rect 342354 633640 342454 633740
rect 342578 633640 342678 633740
rect 342802 633640 342902 633740
rect 343026 633640 343126 633740
rect 342130 633416 342230 633516
rect 342354 633416 342454 633516
rect 342578 633416 342678 633516
rect 342802 633416 342902 633516
rect 343026 633416 343126 633516
rect 342130 633192 342230 633292
rect 342354 633192 342454 633292
rect 342578 633192 342678 633292
rect 342802 633192 342902 633292
rect 343026 633192 343126 633292
rect 342130 632968 342230 633068
rect 342354 632968 342454 633068
rect 342578 632968 342678 633068
rect 342802 632968 342902 633068
rect 343026 632968 343126 633068
rect 297850 632520 297950 632620
rect 298074 632520 298174 632620
rect 298298 632520 298398 632620
rect 298522 632520 298622 632620
rect 298746 632520 298846 632620
rect 297850 632296 297950 632396
rect 298074 632296 298174 632396
rect 298298 632296 298398 632396
rect 298522 632296 298622 632396
rect 298746 632296 298846 632396
rect 297850 632072 297950 632172
rect 298074 632072 298174 632172
rect 298298 632072 298398 632172
rect 298522 632072 298622 632172
rect 298746 632072 298846 632172
rect 297850 631848 297950 631948
rect 298074 631848 298174 631948
rect 298298 631848 298398 631948
rect 298522 631848 298622 631948
rect 298746 631848 298846 631948
rect 297850 631624 297950 631724
rect 298074 631624 298174 631724
rect 298298 631624 298398 631724
rect 298522 631624 298622 631724
rect 298746 631624 298846 631724
rect 297850 631400 297950 631500
rect 298074 631400 298174 631500
rect 298298 631400 298398 631500
rect 298522 631400 298622 631500
rect 298746 631400 298846 631500
rect 342130 632744 342230 632844
rect 342354 632744 342454 632844
rect 342578 632744 342678 632844
rect 342802 632744 342902 632844
rect 343026 632744 343126 632844
rect 342130 632520 342230 632620
rect 342354 632520 342454 632620
rect 342578 632520 342678 632620
rect 342802 632520 342902 632620
rect 343026 632520 343126 632620
rect 323094 631738 323652 632296
rect 326366 631738 326924 632296
rect 328820 631738 329378 632296
rect 331274 631738 331832 632296
rect 342130 632296 342230 632396
rect 342354 632296 342454 632396
rect 342578 632296 342678 632396
rect 342802 632296 342902 632396
rect 343026 632296 343126 632396
rect 342130 632072 342230 632172
rect 342354 632072 342454 632172
rect 342578 632072 342678 632172
rect 342802 632072 342902 632172
rect 343026 632072 343126 632172
rect 342130 631848 342230 631948
rect 342354 631848 342454 631948
rect 342578 631848 342678 631948
rect 342802 631848 342902 631948
rect 343026 631848 343126 631948
rect 342130 631624 342230 631724
rect 342354 631624 342454 631724
rect 342578 631624 342678 631724
rect 342802 631624 342902 631724
rect 343026 631624 343126 631724
rect 323912 630938 324470 631496
rect 325548 630938 326106 631496
rect 329638 630938 330196 631496
rect 342130 631400 342230 631500
rect 342354 631400 342454 631500
rect 342578 631400 342678 631500
rect 342802 631400 342902 631500
rect 343026 631400 343126 631500
rect 322276 630685 322834 630696
rect 322276 630287 322286 630685
rect 322286 630287 322824 630685
rect 322824 630287 322834 630685
rect 322276 630276 322834 630287
rect 323094 630685 323652 630696
rect 323094 630288 323104 630685
rect 323104 630288 323642 630685
rect 323642 630288 323652 630685
rect 323094 630276 323652 630288
rect 323912 630685 324470 630696
rect 323912 630288 323922 630685
rect 323922 630288 324460 630685
rect 324460 630288 324470 630685
rect 323912 630276 324470 630288
rect 324730 630685 325288 630696
rect 324730 630287 324740 630685
rect 324740 630287 325278 630685
rect 325278 630287 325288 630685
rect 324730 630276 325288 630287
rect 325548 630685 326106 630696
rect 325548 630288 325558 630685
rect 325558 630288 326096 630685
rect 326096 630288 326106 630685
rect 325548 630276 326106 630288
rect 326366 630685 326924 630696
rect 326366 630288 326376 630685
rect 326376 630288 326914 630685
rect 326914 630288 326924 630685
rect 326366 630276 326924 630288
rect 327184 630685 327742 630696
rect 327184 630287 327194 630685
rect 327194 630287 327732 630685
rect 327732 630287 327742 630685
rect 327184 630276 327742 630287
rect 328002 630685 328560 630696
rect 328002 630664 328012 630685
rect 327924 630288 328012 630664
rect 328012 630288 328550 630685
rect 328550 630664 328560 630685
rect 328550 630288 328616 630664
rect 327924 630146 328616 630288
rect 328820 630685 329378 630696
rect 328820 630288 328830 630685
rect 328830 630288 329368 630685
rect 329368 630288 329378 630685
rect 328820 630276 329378 630288
rect 329638 630685 330196 630696
rect 329638 630288 329648 630685
rect 329648 630288 330186 630685
rect 330186 630288 330196 630685
rect 329638 630276 330196 630288
rect 330456 630685 331014 630696
rect 330456 630287 330466 630685
rect 330466 630287 331004 630685
rect 331004 630287 331014 630685
rect 330456 630276 331014 630287
rect 331274 630685 331832 630696
rect 331274 630288 331284 630685
rect 331284 630288 331822 630685
rect 331822 630288 331832 630685
rect 331274 630276 331832 630288
rect 322276 629476 322834 630034
rect 324730 629476 325288 630034
rect 327184 629476 327742 630034
rect 330456 629476 331014 630034
rect 332014 630685 332706 630696
rect 332014 630288 332102 630685
rect 332102 630288 332640 630685
rect 332640 630288 332706 630685
rect 332014 630004 332706 630288
rect 319400 628668 319600 628868
rect 319834 628668 320034 628868
rect 320268 628668 320468 628868
rect 320702 628668 320902 628868
rect 321136 628668 321336 628868
rect 321570 628668 321770 628868
rect 322004 628668 322204 628868
rect 322438 628668 322638 628868
rect 322872 628668 323072 628868
rect 323306 628668 323506 628868
rect 323740 628668 323940 628868
rect 324140 628668 324340 628868
rect 324540 628668 324740 628868
rect 324940 628668 325140 628868
rect 325340 628668 325540 628868
rect 325740 628668 325940 628868
rect 326140 628668 326340 628868
rect 326540 628668 326740 628868
rect 326940 628668 327140 628868
rect 327340 628668 327540 628868
rect 328940 628668 329140 628868
rect 329340 628668 329540 628868
rect 329740 628668 329940 628868
rect 330140 628668 330340 628868
rect 330540 628668 330740 628868
rect 330940 628668 331140 628868
rect 331340 628668 331540 628868
rect 331740 628668 331940 628868
rect 332140 628668 332340 628868
rect 319400 628234 319600 628434
rect 319834 628234 320034 628434
rect 320268 628234 320468 628434
rect 320702 628234 320902 628434
rect 321136 628234 321336 628434
rect 321570 628234 321770 628434
rect 322004 628234 322204 628434
rect 322438 628234 322638 628434
rect 322872 628234 323072 628434
rect 323306 628234 323506 628434
rect 323740 628234 323940 628434
rect 332832 630685 333524 630696
rect 332832 630288 332920 630685
rect 332920 630288 333458 630685
rect 333458 630288 333524 630685
rect 332832 630004 333524 630288
rect 319400 627800 319600 628000
rect 319834 627800 320034 628000
rect 320268 627800 320468 628000
rect 320702 627800 320902 628000
rect 321136 627800 321336 628000
rect 321570 627800 321770 628000
rect 322004 627800 322204 628000
rect 322438 627800 322638 628000
rect 322872 627800 323072 628000
rect 323306 627800 323506 628000
rect 323740 627800 323940 628000
rect 313820 626916 315808 627366
rect 312302 626196 312422 626610
rect 311846 625612 311966 625904
rect 297850 624496 297950 624596
rect 298074 624496 298174 624596
rect 298298 624496 298398 624596
rect 298522 624496 298622 624596
rect 298746 624496 298846 624596
rect 297850 624272 297950 624372
rect 298074 624272 298174 624372
rect 298298 624272 298398 624372
rect 298522 624272 298622 624372
rect 298746 624272 298846 624372
rect 297850 624048 297950 624148
rect 298074 624048 298174 624148
rect 298298 624048 298398 624148
rect 298522 624048 298622 624148
rect 298746 624048 298846 624148
rect 302972 624114 303032 624184
rect 303044 624114 303104 624184
rect 303116 624114 303176 624184
rect 303188 624114 303248 624184
rect 303260 624114 303320 624184
rect 303332 624114 303392 624184
rect 303404 624114 303464 624184
rect 303476 624114 303536 624184
rect 302972 624020 303032 624090
rect 303044 624020 303104 624090
rect 303116 624020 303176 624090
rect 303188 624020 303248 624090
rect 303260 624020 303320 624090
rect 303332 624020 303392 624090
rect 303404 624020 303464 624090
rect 303476 624020 303536 624090
rect 297850 623824 297950 623924
rect 298074 623824 298174 623924
rect 298298 623824 298398 623924
rect 298522 623824 298622 623924
rect 298746 623824 298846 623924
rect 297850 623600 297950 623700
rect 298074 623600 298174 623700
rect 298298 623600 298398 623700
rect 298522 623600 298622 623700
rect 298746 623600 298846 623700
rect 297850 623376 297950 623476
rect 298074 623376 298174 623476
rect 298298 623376 298398 623476
rect 298522 623376 298622 623476
rect 298746 623376 298846 623476
rect 297850 623152 297950 623252
rect 298074 623152 298174 623252
rect 298298 623152 298398 623252
rect 298522 623152 298622 623252
rect 298746 623152 298846 623252
rect 297850 622928 297950 623028
rect 298074 622928 298174 623028
rect 298298 622928 298398 623028
rect 298522 622928 298622 623028
rect 298746 622928 298846 623028
rect 297850 622704 297950 622804
rect 298074 622704 298174 622804
rect 298298 622704 298398 622804
rect 298522 622704 298622 622804
rect 298746 622704 298846 622804
rect 297850 622480 297950 622580
rect 298074 622480 298174 622580
rect 298298 622480 298398 622580
rect 298522 622480 298622 622580
rect 298746 622480 298846 622580
rect 297850 622256 297950 622356
rect 298074 622256 298174 622356
rect 298298 622256 298398 622356
rect 298522 622256 298622 622356
rect 298746 622256 298846 622356
rect 297850 622032 297950 622132
rect 298074 622032 298174 622132
rect 298298 622032 298398 622132
rect 298522 622032 298622 622132
rect 298746 622032 298846 622132
rect 297850 621808 297950 621908
rect 298074 621808 298174 621908
rect 298298 621808 298398 621908
rect 298522 621808 298622 621908
rect 298746 621808 298846 621908
rect 297850 621584 297950 621684
rect 298074 621584 298174 621684
rect 298298 621584 298398 621684
rect 298522 621584 298622 621684
rect 298746 621584 298846 621684
rect 297850 621360 297950 621460
rect 298074 621360 298174 621460
rect 298298 621360 298398 621460
rect 298522 621360 298622 621460
rect 298746 621360 298846 621460
rect 297850 621136 297950 621236
rect 298074 621136 298174 621236
rect 298298 621136 298398 621236
rect 298522 621136 298622 621236
rect 298746 621136 298846 621236
rect 297850 620912 297950 621012
rect 298074 620912 298174 621012
rect 298298 620912 298398 621012
rect 298522 620912 298622 621012
rect 298746 620912 298846 621012
rect 297850 620688 297950 620788
rect 298074 620688 298174 620788
rect 298298 620688 298398 620788
rect 298522 620688 298622 620788
rect 298746 620688 298846 620788
rect 297850 620464 297950 620564
rect 298074 620464 298174 620564
rect 298298 620464 298398 620564
rect 298522 620464 298622 620564
rect 298746 620464 298846 620564
rect 300840 620450 300892 620502
rect 297850 620240 297950 620340
rect 298074 620240 298174 620340
rect 298298 620240 298398 620340
rect 298522 620240 298622 620340
rect 298746 620240 298846 620340
rect 302674 620456 302726 620508
rect 303280 620450 303474 620508
rect 301758 620244 301810 620296
rect 297850 620016 297950 620116
rect 298074 620016 298174 620116
rect 298298 620016 298398 620116
rect 298522 620016 298622 620116
rect 298746 620016 298846 620116
rect 297850 619792 297950 619892
rect 298074 619792 298174 619892
rect 298298 619792 298398 619892
rect 298522 619792 298622 619892
rect 298746 619792 298846 619892
rect 297850 619568 297950 619668
rect 298074 619568 298174 619668
rect 298298 619568 298398 619668
rect 298522 619568 298622 619668
rect 298746 619568 298846 619668
rect 297850 619344 297950 619444
rect 298074 619344 298174 619444
rect 298298 619344 298398 619444
rect 298522 619344 298622 619444
rect 298746 619344 298846 619444
rect 297850 619120 297950 619220
rect 298074 619120 298174 619220
rect 298298 619120 298398 619220
rect 298522 619120 298622 619220
rect 298746 619120 298846 619220
rect 297850 618896 297950 618996
rect 298074 618896 298174 618996
rect 298298 618896 298398 618996
rect 298522 618896 298622 618996
rect 298746 618896 298846 618996
rect 297850 618672 297950 618772
rect 298074 618672 298174 618772
rect 298298 618672 298398 618772
rect 298522 618672 298622 618772
rect 298746 618672 298846 618772
rect 297850 618448 297950 618548
rect 298074 618448 298174 618548
rect 298298 618448 298398 618548
rect 298522 618448 298622 618548
rect 298746 618448 298846 618548
rect 297850 618224 297950 618324
rect 298074 618224 298174 618324
rect 298298 618224 298398 618324
rect 298522 618224 298622 618324
rect 298746 618224 298846 618324
rect 297850 618000 297950 618100
rect 298074 618000 298174 618100
rect 298298 618000 298398 618100
rect 298522 618000 298622 618100
rect 298746 618000 298846 618100
rect 302964 616954 303016 617058
rect 306640 622438 306784 622492
rect 306068 622298 306212 622352
rect 307784 622438 307928 622492
rect 307212 622298 307356 622352
rect 308928 622438 309072 622492
rect 308356 622298 308500 622352
rect 304436 619882 304488 620136
rect 304996 619882 305048 620136
rect 305556 619882 305608 620136
rect 306336 620182 306388 620286
rect 306908 620182 306960 620286
rect 306456 619882 306508 620136
rect 306034 619829 306242 619846
rect 306034 619795 306038 619829
rect 306038 619795 306222 619829
rect 306222 619795 306242 619829
rect 306034 619788 306242 619795
rect 306606 619829 306814 619842
rect 306606 619795 306610 619829
rect 306610 619795 306794 619829
rect 306794 619795 306814 619829
rect 306606 619784 306814 619795
rect 307480 620182 307532 620286
rect 308052 620182 308104 620286
rect 307600 619882 307652 620136
rect 307178 619829 307386 619846
rect 307178 619795 307182 619829
rect 307182 619795 307366 619829
rect 307366 619795 307386 619829
rect 307178 619788 307386 619795
rect 307750 619829 307958 619846
rect 307750 619795 307754 619829
rect 307754 619795 307938 619829
rect 307938 619795 307958 619829
rect 307750 619788 307958 619795
rect 308624 620182 308676 620286
rect 309196 620182 309248 620286
rect 308744 619882 308796 620136
rect 309544 619882 309596 620136
rect 308322 619829 308530 619846
rect 308322 619795 308326 619829
rect 308326 619795 308510 619829
rect 308510 619795 308530 619829
rect 308322 619788 308530 619795
rect 308894 619829 309102 619846
rect 308894 619795 308898 619829
rect 308898 619795 309082 619829
rect 309082 619795 309102 619829
rect 308894 619788 309102 619795
rect 310104 619882 310156 620136
rect 313820 626214 315808 626502
rect 316520 625614 318508 625902
rect 312302 622432 312422 622512
rect 311846 622292 311956 622372
rect 310664 619882 310716 620136
rect 312714 619882 313182 620136
rect 303586 616954 303638 617058
rect 304044 616954 304096 617058
rect 304620 616954 304672 617058
rect 305192 616954 305244 617058
rect 305764 616954 305816 617058
rect 306336 616954 306388 617058
rect 306908 616954 306960 617058
rect 307480 616954 307532 617058
rect 308052 616954 308104 617058
rect 308624 616954 308676 617058
rect 309196 616954 309248 617058
rect 309768 616954 309820 617058
rect 310340 616954 310392 617058
rect 310912 616954 310964 617058
rect 311022 616954 311074 617058
rect 311480 616954 311532 617058
rect 312092 616954 312144 617058
rect 312714 616894 313182 617042
rect 331490 627628 332424 628146
rect 327520 626916 329508 627366
rect 327520 626214 329508 626502
rect 324820 625614 326808 625902
rect 303280 616750 303474 616864
rect 304160 616754 304212 616858
rect 304732 616754 304784 616858
rect 305304 616754 305356 616858
rect 309308 616754 309360 616858
rect 309880 616754 309932 616858
rect 310452 616754 310504 616858
rect 314034 616908 314174 617028
rect 314494 616908 314634 617028
rect 314954 616908 315094 617028
rect 315414 616908 315554 617028
rect 315874 616908 316014 617028
rect 316334 616908 316474 617028
rect 316794 616908 316934 617028
rect 317254 616908 317394 617028
rect 317714 616908 317854 617028
rect 318174 616908 318314 617028
rect 319534 616908 319674 617028
rect 319994 616908 320134 617028
rect 320454 616908 320594 617028
rect 320914 616908 321054 617028
rect 321374 616908 321514 617028
rect 321834 616908 321974 617028
rect 322294 616908 322434 617028
rect 322754 616908 322894 617028
rect 323214 616908 323354 617028
rect 323674 616908 323814 617028
rect 325034 616908 325174 617028
rect 325494 616908 325634 617028
rect 325954 616908 326094 617028
rect 326414 616908 326554 617028
rect 326874 616908 327014 617028
rect 327334 616908 327474 617028
rect 327794 616908 327934 617028
rect 328254 616908 328394 617028
rect 328714 616908 328854 617028
rect 332832 626916 333524 627366
rect 333650 630685 334342 630696
rect 333650 630288 333738 630685
rect 333738 630288 334276 630685
rect 334276 630288 334342 630685
rect 333650 630004 334342 630288
rect 333652 625614 334342 625902
rect 332832 622886 333524 623578
rect 331488 617732 332424 618668
rect 337522 623506 338214 623578
rect 337522 623472 337608 623506
rect 337608 623472 337642 623506
rect 337642 623472 337708 623506
rect 337708 623472 337742 623506
rect 337742 623472 337808 623506
rect 337808 623472 337842 623506
rect 337842 623472 337908 623506
rect 337908 623472 337942 623506
rect 337942 623472 338008 623506
rect 338008 623472 338042 623506
rect 338042 623472 338108 623506
rect 338108 623472 338142 623506
rect 338142 623472 338214 623506
rect 337522 623406 338214 623472
rect 337522 623372 337608 623406
rect 337608 623372 337642 623406
rect 337642 623372 337708 623406
rect 337708 623372 337742 623406
rect 337742 623372 337808 623406
rect 337808 623372 337842 623406
rect 337842 623372 337908 623406
rect 337908 623372 337942 623406
rect 337942 623372 338008 623406
rect 338008 623372 338042 623406
rect 338042 623372 338108 623406
rect 338108 623372 338142 623406
rect 338142 623372 338214 623406
rect 337522 623306 338214 623372
rect 337522 623272 337608 623306
rect 337608 623272 337642 623306
rect 337642 623272 337708 623306
rect 337708 623272 337742 623306
rect 337742 623272 337808 623306
rect 337808 623272 337842 623306
rect 337842 623272 337908 623306
rect 337908 623272 337942 623306
rect 337942 623272 338008 623306
rect 338008 623272 338042 623306
rect 338042 623272 338108 623306
rect 338108 623272 338142 623306
rect 338142 623272 338214 623306
rect 337522 623206 338214 623272
rect 337522 623172 337608 623206
rect 337608 623172 337642 623206
rect 337642 623172 337708 623206
rect 337708 623172 337742 623206
rect 337742 623172 337808 623206
rect 337808 623172 337842 623206
rect 337842 623172 337908 623206
rect 337908 623172 337942 623206
rect 337942 623172 338008 623206
rect 338008 623172 338042 623206
rect 338042 623172 338108 623206
rect 338108 623172 338142 623206
rect 338142 623172 338214 623206
rect 337522 623106 338214 623172
rect 337522 623072 337608 623106
rect 337608 623072 337642 623106
rect 337642 623072 337708 623106
rect 337708 623072 337742 623106
rect 337742 623072 337808 623106
rect 337808 623072 337842 623106
rect 337842 623072 337908 623106
rect 337908 623072 337942 623106
rect 337942 623072 338008 623106
rect 338008 623072 338042 623106
rect 338042 623072 338108 623106
rect 338108 623072 338142 623106
rect 338142 623072 338214 623106
rect 337522 623006 338214 623072
rect 337522 622972 337608 623006
rect 337608 622972 337642 623006
rect 337642 622972 337708 623006
rect 337708 622972 337742 623006
rect 337742 622972 337808 623006
rect 337808 622972 337842 623006
rect 337842 622972 337908 623006
rect 337908 622972 337942 623006
rect 337942 622972 338008 623006
rect 338008 622972 338042 623006
rect 338042 622972 338108 623006
rect 338108 622972 338142 623006
rect 338142 622972 338214 623006
rect 337522 622886 338214 622972
rect 334946 618354 335628 618414
rect 334946 618320 335032 618354
rect 335032 618320 335066 618354
rect 335066 618320 335132 618354
rect 335132 618320 335166 618354
rect 335166 618320 335232 618354
rect 335232 618320 335266 618354
rect 335266 618320 335332 618354
rect 335332 618320 335366 618354
rect 335366 618320 335432 618354
rect 335432 618320 335466 618354
rect 335466 618320 335532 618354
rect 335532 618320 335566 618354
rect 335566 618320 335628 618354
rect 334946 618254 335628 618320
rect 334946 618220 335032 618254
rect 335032 618220 335066 618254
rect 335066 618220 335132 618254
rect 335132 618220 335166 618254
rect 335166 618220 335232 618254
rect 335232 618220 335266 618254
rect 335266 618220 335332 618254
rect 335332 618220 335366 618254
rect 335366 618220 335432 618254
rect 335432 618220 335466 618254
rect 335466 618220 335532 618254
rect 335532 618220 335566 618254
rect 335566 618220 335628 618254
rect 334946 618154 335628 618220
rect 334946 618120 335032 618154
rect 335032 618120 335066 618154
rect 335066 618120 335132 618154
rect 335132 618120 335166 618154
rect 335166 618120 335232 618154
rect 335232 618120 335266 618154
rect 335266 618120 335332 618154
rect 335332 618120 335366 618154
rect 335366 618120 335432 618154
rect 335432 618120 335466 618154
rect 335466 618120 335532 618154
rect 335532 618120 335566 618154
rect 335566 618120 335628 618154
rect 334946 618054 335628 618120
rect 334946 618020 335032 618054
rect 335032 618020 335066 618054
rect 335066 618020 335132 618054
rect 335132 618020 335166 618054
rect 335166 618020 335232 618054
rect 335232 618020 335266 618054
rect 335266 618020 335332 618054
rect 335332 618020 335366 618054
rect 335366 618020 335432 618054
rect 335432 618020 335466 618054
rect 335466 618020 335532 618054
rect 335532 618020 335566 618054
rect 335566 618020 335628 618054
rect 334946 617954 335628 618020
rect 334946 617920 335032 617954
rect 335032 617920 335066 617954
rect 335066 617920 335132 617954
rect 335132 617920 335166 617954
rect 335166 617920 335232 617954
rect 335232 617920 335266 617954
rect 335266 617920 335332 617954
rect 335332 617920 335366 617954
rect 335366 617920 335432 617954
rect 335432 617920 335466 617954
rect 335466 617920 335532 617954
rect 335532 617920 335566 617954
rect 335566 617920 335628 617954
rect 334946 617854 335628 617920
rect 334946 617820 335032 617854
rect 335032 617820 335066 617854
rect 335066 617820 335132 617854
rect 335132 617820 335166 617854
rect 335166 617820 335232 617854
rect 335232 617820 335266 617854
rect 335266 617820 335332 617854
rect 335332 617820 335366 617854
rect 335366 617820 335432 617854
rect 335432 617820 335466 617854
rect 335466 617820 335532 617854
rect 335532 617820 335566 617854
rect 335566 617820 335628 617854
rect 334946 617738 335628 617820
rect 336240 618354 336922 618422
rect 336240 618320 336320 618354
rect 336320 618320 336354 618354
rect 336354 618320 336420 618354
rect 336420 618320 336454 618354
rect 336454 618320 336520 618354
rect 336520 618320 336554 618354
rect 336554 618320 336620 618354
rect 336620 618320 336654 618354
rect 336654 618320 336720 618354
rect 336720 618320 336754 618354
rect 336754 618320 336820 618354
rect 336820 618320 336854 618354
rect 336854 618320 336922 618354
rect 336240 618254 336922 618320
rect 336240 618220 336320 618254
rect 336320 618220 336354 618254
rect 336354 618220 336420 618254
rect 336420 618220 336454 618254
rect 336454 618220 336520 618254
rect 336520 618220 336554 618254
rect 336554 618220 336620 618254
rect 336620 618220 336654 618254
rect 336654 618220 336720 618254
rect 336720 618220 336754 618254
rect 336754 618220 336820 618254
rect 336820 618220 336854 618254
rect 336854 618220 336922 618254
rect 336240 618154 336922 618220
rect 336240 618120 336320 618154
rect 336320 618120 336354 618154
rect 336354 618120 336420 618154
rect 336420 618120 336454 618154
rect 336454 618120 336520 618154
rect 336520 618120 336554 618154
rect 336554 618120 336620 618154
rect 336620 618120 336654 618154
rect 336654 618120 336720 618154
rect 336720 618120 336754 618154
rect 336754 618120 336820 618154
rect 336820 618120 336854 618154
rect 336854 618120 336922 618154
rect 336240 618054 336922 618120
rect 336240 618020 336320 618054
rect 336320 618020 336354 618054
rect 336354 618020 336420 618054
rect 336420 618020 336454 618054
rect 336454 618020 336520 618054
rect 336520 618020 336554 618054
rect 336554 618020 336620 618054
rect 336620 618020 336654 618054
rect 336654 618020 336720 618054
rect 336720 618020 336754 618054
rect 336754 618020 336820 618054
rect 336820 618020 336854 618054
rect 336854 618020 336922 618054
rect 336240 617954 336922 618020
rect 342130 624496 342230 624596
rect 342354 624496 342454 624596
rect 342578 624496 342678 624596
rect 342802 624496 342902 624596
rect 343026 624496 343126 624596
rect 342130 624272 342230 624372
rect 342354 624272 342454 624372
rect 342578 624272 342678 624372
rect 342802 624272 342902 624372
rect 343026 624272 343126 624372
rect 342130 624048 342230 624148
rect 342354 624048 342454 624148
rect 342578 624048 342678 624148
rect 342802 624048 342902 624148
rect 343026 624048 343126 624148
rect 342130 623824 342230 623924
rect 342354 623824 342454 623924
rect 342578 623824 342678 623924
rect 342802 623824 342902 623924
rect 343026 623824 343126 623924
rect 342130 623600 342230 623700
rect 342354 623600 342454 623700
rect 342578 623600 342678 623700
rect 342802 623600 342902 623700
rect 343026 623600 343126 623700
rect 342130 623376 342230 623476
rect 342354 623376 342454 623476
rect 342578 623376 342678 623476
rect 342802 623376 342902 623476
rect 343026 623376 343126 623476
rect 342130 623152 342230 623252
rect 342354 623152 342454 623252
rect 342578 623152 342678 623252
rect 342802 623152 342902 623252
rect 343026 623152 343126 623252
rect 342130 622928 342230 623028
rect 342354 622928 342454 623028
rect 342578 622928 342678 623028
rect 342802 622928 342902 623028
rect 343026 622928 343126 623028
rect 342130 622704 342230 622804
rect 342354 622704 342454 622804
rect 342578 622704 342678 622804
rect 342802 622704 342902 622804
rect 343026 622704 343126 622804
rect 342130 622480 342230 622580
rect 342354 622480 342454 622580
rect 342578 622480 342678 622580
rect 342802 622480 342902 622580
rect 343026 622480 343126 622580
rect 342130 622256 342230 622356
rect 342354 622256 342454 622356
rect 342578 622256 342678 622356
rect 342802 622256 342902 622356
rect 343026 622256 343126 622356
rect 342130 622032 342230 622132
rect 342354 622032 342454 622132
rect 342578 622032 342678 622132
rect 342802 622032 342902 622132
rect 343026 622032 343126 622132
rect 342130 621808 342230 621908
rect 342354 621808 342454 621908
rect 342578 621808 342678 621908
rect 342802 621808 342902 621908
rect 343026 621808 343126 621908
rect 342130 621584 342230 621684
rect 342354 621584 342454 621684
rect 342578 621584 342678 621684
rect 342802 621584 342902 621684
rect 343026 621584 343126 621684
rect 342130 621360 342230 621460
rect 342354 621360 342454 621460
rect 342578 621360 342678 621460
rect 342802 621360 342902 621460
rect 343026 621360 343126 621460
rect 342130 621136 342230 621236
rect 342354 621136 342454 621236
rect 342578 621136 342678 621236
rect 342802 621136 342902 621236
rect 343026 621136 343126 621236
rect 342130 620912 342230 621012
rect 342354 620912 342454 621012
rect 342578 620912 342678 621012
rect 342802 620912 342902 621012
rect 343026 620912 343126 621012
rect 342130 620688 342230 620788
rect 342354 620688 342454 620788
rect 342578 620688 342678 620788
rect 342802 620688 342902 620788
rect 343026 620688 343126 620788
rect 342130 620464 342230 620564
rect 342354 620464 342454 620564
rect 342578 620464 342678 620564
rect 342802 620464 342902 620564
rect 343026 620464 343126 620564
rect 342130 620240 342230 620340
rect 342354 620240 342454 620340
rect 342578 620240 342678 620340
rect 342802 620240 342902 620340
rect 343026 620240 343126 620340
rect 342130 620016 342230 620116
rect 342354 620016 342454 620116
rect 342578 620016 342678 620116
rect 342802 620016 342902 620116
rect 343026 620016 343126 620116
rect 342130 619792 342230 619892
rect 342354 619792 342454 619892
rect 342578 619792 342678 619892
rect 342802 619792 342902 619892
rect 343026 619792 343126 619892
rect 342130 619568 342230 619668
rect 342354 619568 342454 619668
rect 342578 619568 342678 619668
rect 342802 619568 342902 619668
rect 343026 619568 343126 619668
rect 342130 619344 342230 619444
rect 342354 619344 342454 619444
rect 342578 619344 342678 619444
rect 342802 619344 342902 619444
rect 343026 619344 343126 619444
rect 342130 619120 342230 619220
rect 342354 619120 342454 619220
rect 342578 619120 342678 619220
rect 342802 619120 342902 619220
rect 343026 619120 343126 619220
rect 342130 618896 342230 618996
rect 342354 618896 342454 618996
rect 342578 618896 342678 618996
rect 342802 618896 342902 618996
rect 343026 618896 343126 618996
rect 342130 618672 342230 618772
rect 342354 618672 342454 618772
rect 342578 618672 342678 618772
rect 342802 618672 342902 618772
rect 343026 618672 343126 618772
rect 342130 618448 342230 618548
rect 342354 618448 342454 618548
rect 342578 618448 342678 618548
rect 342802 618448 342902 618548
rect 343026 618448 343126 618548
rect 342130 618224 342230 618324
rect 342354 618224 342454 618324
rect 342578 618224 342678 618324
rect 342802 618224 342902 618324
rect 343026 618224 343126 618324
rect 342130 618000 342230 618100
rect 342354 618000 342454 618100
rect 342578 618000 342678 618100
rect 342802 618000 342902 618100
rect 343026 618000 343126 618100
rect 336240 617920 336320 617954
rect 336320 617920 336354 617954
rect 336354 617920 336420 617954
rect 336420 617920 336454 617954
rect 336454 617920 336520 617954
rect 336520 617920 336554 617954
rect 336554 617920 336620 617954
rect 336620 617920 336654 617954
rect 336654 617920 336720 617954
rect 336720 617920 336754 617954
rect 336754 617920 336820 617954
rect 336820 617920 336854 617954
rect 336854 617920 336922 617954
rect 336240 617854 336922 617920
rect 336240 617820 336320 617854
rect 336320 617820 336354 617854
rect 336354 617820 336420 617854
rect 336420 617820 336454 617854
rect 336454 617820 336520 617854
rect 336520 617820 336554 617854
rect 336554 617820 336620 617854
rect 336620 617820 336654 617854
rect 336654 617820 336720 617854
rect 336720 617820 336754 617854
rect 336754 617820 336820 617854
rect 336820 617820 336854 617854
rect 336854 617820 336922 617854
rect 336240 617746 336922 617820
rect 329174 616908 329314 617028
rect 314294 616748 314374 616828
rect 315214 616748 315294 616828
rect 316134 616748 316214 616828
rect 317054 616748 317134 616828
rect 317974 616748 318054 616828
rect 312804 616608 313204 616708
rect 319794 616748 319874 616828
rect 320714 616748 320794 616828
rect 321634 616748 321714 616828
rect 322554 616748 322634 616828
rect 323474 616748 323554 616828
rect 318714 616608 319114 616708
rect 325294 616748 325374 616828
rect 326214 616748 326294 616828
rect 327134 616748 327214 616828
rect 328054 616748 328134 616828
rect 328974 616748 329054 616828
rect 324214 616608 324614 616708
rect 330170 616606 330570 616706
rect 298876 615374 298976 615474
rect 299100 615374 299200 615474
rect 299324 615374 299424 615474
rect 299548 615374 299648 615474
rect 299772 615374 299872 615474
rect 299996 615374 300096 615474
rect 300220 615374 300320 615474
rect 300444 615374 300544 615474
rect 300668 615374 300768 615474
rect 300892 615374 300992 615474
rect 301116 615374 301216 615474
rect 301340 615374 301440 615474
rect 301564 615374 301664 615474
rect 301788 615374 301888 615474
rect 302012 615374 302112 615474
rect 302236 615374 302336 615474
rect 302460 615374 302560 615474
rect 302684 615374 302784 615474
rect 302908 615374 303008 615474
rect 303132 615374 303232 615474
rect 303356 615374 303456 615474
rect 303580 615374 303680 615474
rect 303804 615374 303904 615474
rect 304028 615374 304128 615474
rect 304252 615374 304352 615474
rect 304476 615374 304576 615474
rect 304700 615374 304800 615474
rect 304924 615374 305024 615474
rect 305148 615374 305248 615474
rect 305372 615374 305472 615474
rect 298876 615150 298976 615250
rect 299100 615150 299200 615250
rect 299324 615150 299424 615250
rect 299548 615150 299648 615250
rect 299772 615150 299872 615250
rect 299996 615150 300096 615250
rect 300220 615150 300320 615250
rect 300444 615150 300544 615250
rect 300668 615150 300768 615250
rect 300892 615150 300992 615250
rect 301116 615150 301216 615250
rect 301340 615150 301440 615250
rect 301564 615150 301664 615250
rect 301788 615150 301888 615250
rect 302012 615150 302112 615250
rect 302236 615150 302336 615250
rect 302460 615150 302560 615250
rect 302684 615150 302784 615250
rect 302908 615150 303008 615250
rect 303132 615150 303232 615250
rect 303356 615150 303456 615250
rect 303580 615150 303680 615250
rect 303804 615150 303904 615250
rect 304028 615150 304128 615250
rect 304252 615150 304352 615250
rect 304476 615150 304576 615250
rect 304700 615150 304800 615250
rect 304924 615150 305024 615250
rect 305148 615150 305248 615250
rect 305372 615150 305472 615250
rect 298876 614926 298976 615026
rect 299100 614926 299200 615026
rect 299324 614926 299424 615026
rect 299548 614926 299648 615026
rect 299772 614926 299872 615026
rect 299996 614926 300096 615026
rect 300220 614926 300320 615026
rect 300444 614926 300544 615026
rect 300668 614926 300768 615026
rect 300892 614926 300992 615026
rect 301116 614926 301216 615026
rect 301340 614926 301440 615026
rect 301564 614926 301664 615026
rect 301788 614926 301888 615026
rect 302012 614926 302112 615026
rect 302236 614926 302336 615026
rect 302460 614926 302560 615026
rect 302684 614926 302784 615026
rect 302908 614926 303008 615026
rect 303132 614926 303232 615026
rect 303356 614926 303456 615026
rect 303580 614926 303680 615026
rect 303804 614926 303904 615026
rect 304028 614926 304128 615026
rect 304252 614926 304352 615026
rect 304476 614926 304576 615026
rect 304700 614926 304800 615026
rect 304924 614926 305024 615026
rect 305148 614926 305248 615026
rect 305372 614926 305472 615026
rect 298876 614702 298976 614802
rect 299100 614702 299200 614802
rect 299324 614702 299424 614802
rect 299548 614702 299648 614802
rect 299772 614702 299872 614802
rect 299996 614702 300096 614802
rect 300220 614702 300320 614802
rect 300444 614702 300544 614802
rect 300668 614702 300768 614802
rect 300892 614702 300992 614802
rect 301116 614702 301216 614802
rect 301340 614702 301440 614802
rect 301564 614702 301664 614802
rect 301788 614702 301888 614802
rect 302012 614702 302112 614802
rect 302236 614702 302336 614802
rect 302460 614702 302560 614802
rect 302684 614702 302784 614802
rect 302908 614702 303008 614802
rect 303132 614702 303232 614802
rect 303356 614702 303456 614802
rect 303580 614702 303680 614802
rect 303804 614702 303904 614802
rect 304028 614702 304128 614802
rect 304252 614702 304352 614802
rect 304476 614702 304576 614802
rect 304700 614702 304800 614802
rect 304924 614702 305024 614802
rect 305148 614702 305248 614802
rect 305372 614702 305472 614802
rect 298876 614478 298976 614578
rect 299100 614478 299200 614578
rect 299324 614478 299424 614578
rect 299548 614478 299648 614578
rect 299772 614478 299872 614578
rect 299996 614478 300096 614578
rect 300220 614478 300320 614578
rect 300444 614478 300544 614578
rect 300668 614478 300768 614578
rect 300892 614478 300992 614578
rect 301116 614478 301216 614578
rect 301340 614478 301440 614578
rect 301564 614478 301664 614578
rect 301788 614478 301888 614578
rect 302012 614478 302112 614578
rect 302236 614478 302336 614578
rect 302460 614478 302560 614578
rect 302684 614478 302784 614578
rect 302908 614478 303008 614578
rect 303132 614478 303232 614578
rect 303356 614478 303456 614578
rect 303580 614478 303680 614578
rect 303804 614478 303904 614578
rect 304028 614478 304128 614578
rect 304252 614478 304352 614578
rect 304476 614478 304576 614578
rect 304700 614478 304800 614578
rect 304924 614478 305024 614578
rect 305148 614478 305248 614578
rect 305372 614478 305472 614578
rect 309346 615374 309446 615474
rect 309570 615374 309670 615474
rect 309794 615374 309894 615474
rect 310018 615374 310118 615474
rect 310242 615374 310342 615474
rect 310466 615374 310566 615474
rect 310690 615374 310790 615474
rect 310914 615374 311014 615474
rect 311138 615374 311238 615474
rect 311362 615374 311462 615474
rect 311586 615374 311686 615474
rect 311810 615374 311910 615474
rect 312034 615374 312134 615474
rect 312258 615374 312358 615474
rect 312482 615374 312582 615474
rect 312706 615374 312806 615474
rect 312930 615374 313030 615474
rect 313154 615374 313254 615474
rect 313378 615374 313478 615474
rect 313602 615374 313702 615474
rect 313826 615374 313926 615474
rect 314050 615374 314150 615474
rect 314274 615374 314374 615474
rect 314498 615374 314598 615474
rect 314722 615374 314822 615474
rect 314946 615374 315046 615474
rect 315170 615374 315270 615474
rect 315394 615374 315494 615474
rect 315618 615374 315718 615474
rect 315842 615374 315942 615474
rect 309346 615150 309446 615250
rect 309570 615150 309670 615250
rect 309794 615150 309894 615250
rect 310018 615150 310118 615250
rect 310242 615150 310342 615250
rect 310466 615150 310566 615250
rect 310690 615150 310790 615250
rect 310914 615150 311014 615250
rect 311138 615150 311238 615250
rect 311362 615150 311462 615250
rect 311586 615150 311686 615250
rect 311810 615150 311910 615250
rect 312034 615150 312134 615250
rect 312258 615150 312358 615250
rect 312482 615150 312582 615250
rect 312706 615150 312806 615250
rect 312930 615150 313030 615250
rect 313154 615150 313254 615250
rect 313378 615150 313478 615250
rect 313602 615150 313702 615250
rect 313826 615150 313926 615250
rect 314050 615150 314150 615250
rect 314274 615150 314374 615250
rect 314498 615150 314598 615250
rect 314722 615150 314822 615250
rect 314946 615150 315046 615250
rect 315170 615150 315270 615250
rect 315394 615150 315494 615250
rect 315618 615150 315718 615250
rect 315842 615150 315942 615250
rect 309346 614926 309446 615026
rect 309570 614926 309670 615026
rect 309794 614926 309894 615026
rect 310018 614926 310118 615026
rect 310242 614926 310342 615026
rect 310466 614926 310566 615026
rect 310690 614926 310790 615026
rect 310914 614926 311014 615026
rect 311138 614926 311238 615026
rect 311362 614926 311462 615026
rect 311586 614926 311686 615026
rect 311810 614926 311910 615026
rect 312034 614926 312134 615026
rect 312258 614926 312358 615026
rect 312482 614926 312582 615026
rect 312706 614926 312806 615026
rect 312930 614926 313030 615026
rect 313154 614926 313254 615026
rect 313378 614926 313478 615026
rect 313602 614926 313702 615026
rect 313826 614926 313926 615026
rect 314050 614926 314150 615026
rect 314274 614926 314374 615026
rect 314498 614926 314598 615026
rect 314722 614926 314822 615026
rect 314946 614926 315046 615026
rect 315170 614926 315270 615026
rect 315394 614926 315494 615026
rect 315618 614926 315718 615026
rect 315842 614926 315942 615026
rect 309346 614702 309446 614802
rect 309570 614702 309670 614802
rect 309794 614702 309894 614802
rect 310018 614702 310118 614802
rect 310242 614702 310342 614802
rect 310466 614702 310566 614802
rect 310690 614702 310790 614802
rect 310914 614702 311014 614802
rect 311138 614702 311238 614802
rect 311362 614702 311462 614802
rect 311586 614702 311686 614802
rect 311810 614702 311910 614802
rect 312034 614702 312134 614802
rect 312258 614702 312358 614802
rect 312482 614702 312582 614802
rect 312706 614702 312806 614802
rect 312930 614702 313030 614802
rect 313154 614702 313254 614802
rect 313378 614702 313478 614802
rect 313602 614702 313702 614802
rect 313826 614702 313926 614802
rect 314050 614702 314150 614802
rect 314274 614702 314374 614802
rect 314498 614702 314598 614802
rect 314722 614702 314822 614802
rect 314946 614702 315046 614802
rect 315170 614702 315270 614802
rect 315394 614702 315494 614802
rect 315618 614702 315718 614802
rect 315842 614702 315942 614802
rect 309346 614478 309446 614578
rect 309570 614478 309670 614578
rect 309794 614478 309894 614578
rect 310018 614478 310118 614578
rect 310242 614478 310342 614578
rect 310466 614478 310566 614578
rect 310690 614478 310790 614578
rect 310914 614478 311014 614578
rect 311138 614478 311238 614578
rect 311362 614478 311462 614578
rect 311586 614478 311686 614578
rect 311810 614478 311910 614578
rect 312034 614478 312134 614578
rect 312258 614478 312358 614578
rect 312482 614478 312582 614578
rect 312706 614478 312806 614578
rect 312930 614478 313030 614578
rect 313154 614478 313254 614578
rect 313378 614478 313478 614578
rect 313602 614478 313702 614578
rect 313826 614478 313926 614578
rect 314050 614478 314150 614578
rect 314274 614478 314374 614578
rect 314498 614478 314598 614578
rect 314722 614478 314822 614578
rect 314946 614478 315046 614578
rect 315170 614478 315270 614578
rect 315394 614478 315494 614578
rect 315618 614478 315718 614578
rect 315842 614478 315942 614578
rect 335616 615394 335716 615494
rect 335840 615394 335940 615494
rect 336064 615394 336164 615494
rect 336288 615394 336388 615494
rect 336512 615394 336612 615494
rect 336736 615394 336836 615494
rect 336960 615394 337060 615494
rect 337184 615394 337284 615494
rect 337408 615394 337508 615494
rect 337632 615394 337732 615494
rect 337856 615394 337956 615494
rect 338080 615394 338180 615494
rect 338304 615394 338404 615494
rect 338528 615394 338628 615494
rect 338752 615394 338852 615494
rect 338976 615394 339076 615494
rect 339200 615394 339300 615494
rect 339424 615394 339524 615494
rect 339648 615394 339748 615494
rect 339872 615394 339972 615494
rect 340096 615394 340196 615494
rect 340320 615394 340420 615494
rect 340544 615394 340644 615494
rect 340768 615394 340868 615494
rect 340992 615394 341092 615494
rect 341216 615394 341316 615494
rect 341440 615394 341540 615494
rect 341664 615394 341764 615494
rect 341888 615394 341988 615494
rect 342112 615394 342212 615494
rect 335616 615170 335716 615270
rect 335840 615170 335940 615270
rect 336064 615170 336164 615270
rect 336288 615170 336388 615270
rect 336512 615170 336612 615270
rect 336736 615170 336836 615270
rect 336960 615170 337060 615270
rect 337184 615170 337284 615270
rect 337408 615170 337508 615270
rect 337632 615170 337732 615270
rect 337856 615170 337956 615270
rect 338080 615170 338180 615270
rect 338304 615170 338404 615270
rect 338528 615170 338628 615270
rect 338752 615170 338852 615270
rect 338976 615170 339076 615270
rect 339200 615170 339300 615270
rect 339424 615170 339524 615270
rect 339648 615170 339748 615270
rect 339872 615170 339972 615270
rect 340096 615170 340196 615270
rect 340320 615170 340420 615270
rect 340544 615170 340644 615270
rect 340768 615170 340868 615270
rect 340992 615170 341092 615270
rect 341216 615170 341316 615270
rect 341440 615170 341540 615270
rect 341664 615170 341764 615270
rect 341888 615170 341988 615270
rect 342112 615170 342212 615270
rect 335616 614946 335716 615046
rect 335840 614946 335940 615046
rect 336064 614946 336164 615046
rect 336288 614946 336388 615046
rect 336512 614946 336612 615046
rect 336736 614946 336836 615046
rect 336960 614946 337060 615046
rect 337184 614946 337284 615046
rect 337408 614946 337508 615046
rect 337632 614946 337732 615046
rect 337856 614946 337956 615046
rect 338080 614946 338180 615046
rect 338304 614946 338404 615046
rect 338528 614946 338628 615046
rect 338752 614946 338852 615046
rect 338976 614946 339076 615046
rect 339200 614946 339300 615046
rect 339424 614946 339524 615046
rect 339648 614946 339748 615046
rect 339872 614946 339972 615046
rect 340096 614946 340196 615046
rect 340320 614946 340420 615046
rect 340544 614946 340644 615046
rect 340768 614946 340868 615046
rect 340992 614946 341092 615046
rect 341216 614946 341316 615046
rect 341440 614946 341540 615046
rect 341664 614946 341764 615046
rect 341888 614946 341988 615046
rect 342112 614946 342212 615046
rect 335616 614722 335716 614822
rect 335840 614722 335940 614822
rect 336064 614722 336164 614822
rect 336288 614722 336388 614822
rect 336512 614722 336612 614822
rect 336736 614722 336836 614822
rect 336960 614722 337060 614822
rect 337184 614722 337284 614822
rect 337408 614722 337508 614822
rect 337632 614722 337732 614822
rect 337856 614722 337956 614822
rect 338080 614722 338180 614822
rect 338304 614722 338404 614822
rect 338528 614722 338628 614822
rect 338752 614722 338852 614822
rect 338976 614722 339076 614822
rect 339200 614722 339300 614822
rect 339424 614722 339524 614822
rect 339648 614722 339748 614822
rect 339872 614722 339972 614822
rect 340096 614722 340196 614822
rect 340320 614722 340420 614822
rect 340544 614722 340644 614822
rect 340768 614722 340868 614822
rect 340992 614722 341092 614822
rect 341216 614722 341316 614822
rect 341440 614722 341540 614822
rect 341664 614722 341764 614822
rect 341888 614722 341988 614822
rect 342112 614722 342212 614822
rect 335616 614498 335716 614598
rect 335840 614498 335940 614598
rect 336064 614498 336164 614598
rect 336288 614498 336388 614598
rect 336512 614498 336612 614598
rect 336736 614498 336836 614598
rect 336960 614498 337060 614598
rect 337184 614498 337284 614598
rect 337408 614498 337508 614598
rect 337632 614498 337732 614598
rect 337856 614498 337956 614598
rect 338080 614498 338180 614598
rect 338304 614498 338404 614598
rect 338528 614498 338628 614598
rect 338752 614498 338852 614598
rect 338976 614498 339076 614598
rect 339200 614498 339300 614598
rect 339424 614498 339524 614598
rect 339648 614498 339748 614598
rect 339872 614498 339972 614598
rect 340096 614498 340196 614598
rect 340320 614498 340420 614598
rect 340544 614498 340644 614598
rect 340768 614498 340868 614598
rect 340992 614498 341092 614598
rect 341216 614498 341316 614598
rect 341440 614498 341540 614598
rect 341664 614498 341764 614598
rect 341888 614498 341988 614598
rect 342112 614498 342212 614598
<< metal2 >>
rect 298836 642694 305496 642724
rect 298836 642594 298876 642694
rect 298976 642594 299100 642694
rect 299200 642594 299324 642694
rect 299424 642594 299548 642694
rect 299648 642594 299772 642694
rect 299872 642594 299996 642694
rect 300096 642594 300220 642694
rect 300320 642594 300444 642694
rect 300544 642594 300668 642694
rect 300768 642594 300892 642694
rect 300992 642594 301116 642694
rect 301216 642594 301340 642694
rect 301440 642594 301564 642694
rect 301664 642594 301788 642694
rect 301888 642594 302012 642694
rect 302112 642594 302236 642694
rect 302336 642594 302460 642694
rect 302560 642594 302684 642694
rect 302784 642594 302908 642694
rect 303008 642594 303132 642694
rect 303232 642594 303356 642694
rect 303456 642594 303580 642694
rect 303680 642594 303804 642694
rect 303904 642594 304028 642694
rect 304128 642594 304252 642694
rect 304352 642594 304476 642694
rect 304576 642594 304700 642694
rect 304800 642594 304924 642694
rect 305024 642594 305148 642694
rect 305248 642594 305372 642694
rect 305472 642594 305496 642694
rect 298836 642470 305496 642594
rect 298836 642370 298876 642470
rect 298976 642370 299100 642470
rect 299200 642370 299324 642470
rect 299424 642370 299548 642470
rect 299648 642370 299772 642470
rect 299872 642370 299996 642470
rect 300096 642370 300220 642470
rect 300320 642370 300444 642470
rect 300544 642370 300668 642470
rect 300768 642370 300892 642470
rect 300992 642370 301116 642470
rect 301216 642370 301340 642470
rect 301440 642370 301564 642470
rect 301664 642370 301788 642470
rect 301888 642370 302012 642470
rect 302112 642370 302236 642470
rect 302336 642370 302460 642470
rect 302560 642370 302684 642470
rect 302784 642370 302908 642470
rect 303008 642370 303132 642470
rect 303232 642370 303356 642470
rect 303456 642370 303580 642470
rect 303680 642370 303804 642470
rect 303904 642370 304028 642470
rect 304128 642370 304252 642470
rect 304352 642370 304476 642470
rect 304576 642370 304700 642470
rect 304800 642370 304924 642470
rect 305024 642370 305148 642470
rect 305248 642370 305372 642470
rect 305472 642370 305496 642470
rect 298836 642246 305496 642370
rect 298836 642146 298876 642246
rect 298976 642146 299100 642246
rect 299200 642146 299324 642246
rect 299424 642146 299548 642246
rect 299648 642146 299772 642246
rect 299872 642146 299996 642246
rect 300096 642146 300220 642246
rect 300320 642146 300444 642246
rect 300544 642146 300668 642246
rect 300768 642146 300892 642246
rect 300992 642146 301116 642246
rect 301216 642146 301340 642246
rect 301440 642146 301564 642246
rect 301664 642146 301788 642246
rect 301888 642146 302012 642246
rect 302112 642146 302236 642246
rect 302336 642146 302460 642246
rect 302560 642146 302684 642246
rect 302784 642146 302908 642246
rect 303008 642146 303132 642246
rect 303232 642146 303356 642246
rect 303456 642146 303580 642246
rect 303680 642146 303804 642246
rect 303904 642146 304028 642246
rect 304128 642146 304252 642246
rect 304352 642146 304476 642246
rect 304576 642146 304700 642246
rect 304800 642146 304924 642246
rect 305024 642146 305148 642246
rect 305248 642146 305372 642246
rect 305472 642146 305496 642246
rect 298836 642022 305496 642146
rect 298836 641922 298876 642022
rect 298976 641922 299100 642022
rect 299200 641922 299324 642022
rect 299424 641922 299548 642022
rect 299648 641922 299772 642022
rect 299872 641922 299996 642022
rect 300096 641922 300220 642022
rect 300320 641922 300444 642022
rect 300544 641922 300668 642022
rect 300768 641922 300892 642022
rect 300992 641922 301116 642022
rect 301216 641922 301340 642022
rect 301440 641922 301564 642022
rect 301664 641922 301788 642022
rect 301888 641922 302012 642022
rect 302112 641922 302236 642022
rect 302336 641922 302460 642022
rect 302560 641922 302684 642022
rect 302784 641922 302908 642022
rect 303008 641922 303132 642022
rect 303232 641922 303356 642022
rect 303456 641922 303580 642022
rect 303680 641922 303804 642022
rect 303904 641922 304028 642022
rect 304128 641922 304252 642022
rect 304352 641922 304476 642022
rect 304576 641922 304700 642022
rect 304800 641922 304924 642022
rect 305024 641922 305148 642022
rect 305248 641922 305372 642022
rect 305472 641922 305496 642022
rect 298836 641798 305496 641922
rect 298836 641698 298876 641798
rect 298976 641698 299100 641798
rect 299200 641698 299324 641798
rect 299424 641698 299548 641798
rect 299648 641698 299772 641798
rect 299872 641698 299996 641798
rect 300096 641698 300220 641798
rect 300320 641698 300444 641798
rect 300544 641698 300668 641798
rect 300768 641698 300892 641798
rect 300992 641698 301116 641798
rect 301216 641698 301340 641798
rect 301440 641698 301564 641798
rect 301664 641698 301788 641798
rect 301888 641698 302012 641798
rect 302112 641698 302236 641798
rect 302336 641698 302460 641798
rect 302560 641698 302684 641798
rect 302784 641698 302908 641798
rect 303008 641698 303132 641798
rect 303232 641698 303356 641798
rect 303456 641698 303580 641798
rect 303680 641698 303804 641798
rect 303904 641698 304028 641798
rect 304128 641698 304252 641798
rect 304352 641698 304476 641798
rect 304576 641698 304700 641798
rect 304800 641698 304924 641798
rect 305024 641698 305148 641798
rect 305248 641698 305372 641798
rect 305472 641698 305496 641798
rect 298836 641664 305496 641698
rect 309306 642694 315966 642724
rect 309306 642594 309346 642694
rect 309446 642594 309570 642694
rect 309670 642594 309794 642694
rect 309894 642594 310018 642694
rect 310118 642594 310242 642694
rect 310342 642594 310466 642694
rect 310566 642594 310690 642694
rect 310790 642594 310914 642694
rect 311014 642594 311138 642694
rect 311238 642594 311362 642694
rect 311462 642594 311586 642694
rect 311686 642594 311810 642694
rect 311910 642594 312034 642694
rect 312134 642594 312258 642694
rect 312358 642594 312482 642694
rect 312582 642594 312706 642694
rect 312806 642594 312930 642694
rect 313030 642594 313154 642694
rect 313254 642594 313378 642694
rect 313478 642594 313602 642694
rect 313702 642594 313826 642694
rect 313926 642594 314050 642694
rect 314150 642594 314274 642694
rect 314374 642594 314498 642694
rect 314598 642594 314722 642694
rect 314822 642594 314946 642694
rect 315046 642594 315170 642694
rect 315270 642594 315394 642694
rect 315494 642594 315618 642694
rect 315718 642594 315842 642694
rect 315942 642594 315966 642694
rect 309306 642470 315966 642594
rect 309306 642370 309346 642470
rect 309446 642370 309570 642470
rect 309670 642370 309794 642470
rect 309894 642370 310018 642470
rect 310118 642370 310242 642470
rect 310342 642370 310466 642470
rect 310566 642370 310690 642470
rect 310790 642370 310914 642470
rect 311014 642370 311138 642470
rect 311238 642370 311362 642470
rect 311462 642370 311586 642470
rect 311686 642370 311810 642470
rect 311910 642370 312034 642470
rect 312134 642370 312258 642470
rect 312358 642370 312482 642470
rect 312582 642370 312706 642470
rect 312806 642370 312930 642470
rect 313030 642370 313154 642470
rect 313254 642370 313378 642470
rect 313478 642370 313602 642470
rect 313702 642370 313826 642470
rect 313926 642370 314050 642470
rect 314150 642370 314274 642470
rect 314374 642370 314498 642470
rect 314598 642370 314722 642470
rect 314822 642370 314946 642470
rect 315046 642370 315170 642470
rect 315270 642370 315394 642470
rect 315494 642370 315618 642470
rect 315718 642370 315842 642470
rect 315942 642370 315966 642470
rect 309306 642246 315966 642370
rect 309306 642146 309346 642246
rect 309446 642146 309570 642246
rect 309670 642146 309794 642246
rect 309894 642146 310018 642246
rect 310118 642146 310242 642246
rect 310342 642146 310466 642246
rect 310566 642146 310690 642246
rect 310790 642146 310914 642246
rect 311014 642146 311138 642246
rect 311238 642146 311362 642246
rect 311462 642146 311586 642246
rect 311686 642146 311810 642246
rect 311910 642146 312034 642246
rect 312134 642146 312258 642246
rect 312358 642146 312482 642246
rect 312582 642146 312706 642246
rect 312806 642146 312930 642246
rect 313030 642146 313154 642246
rect 313254 642146 313378 642246
rect 313478 642146 313602 642246
rect 313702 642146 313826 642246
rect 313926 642146 314050 642246
rect 314150 642146 314274 642246
rect 314374 642146 314498 642246
rect 314598 642146 314722 642246
rect 314822 642146 314946 642246
rect 315046 642146 315170 642246
rect 315270 642146 315394 642246
rect 315494 642146 315618 642246
rect 315718 642146 315842 642246
rect 315942 642146 315966 642246
rect 309306 642022 315966 642146
rect 309306 641922 309346 642022
rect 309446 641922 309570 642022
rect 309670 641922 309794 642022
rect 309894 641922 310018 642022
rect 310118 641922 310242 642022
rect 310342 641922 310466 642022
rect 310566 641922 310690 642022
rect 310790 641922 310914 642022
rect 311014 641922 311138 642022
rect 311238 641922 311362 642022
rect 311462 641922 311586 642022
rect 311686 641922 311810 642022
rect 311910 641922 312034 642022
rect 312134 641922 312258 642022
rect 312358 641922 312482 642022
rect 312582 641922 312706 642022
rect 312806 641922 312930 642022
rect 313030 641922 313154 642022
rect 313254 641922 313378 642022
rect 313478 641922 313602 642022
rect 313702 641922 313826 642022
rect 313926 641922 314050 642022
rect 314150 641922 314274 642022
rect 314374 641922 314498 642022
rect 314598 641922 314722 642022
rect 314822 641922 314946 642022
rect 315046 641922 315170 642022
rect 315270 641922 315394 642022
rect 315494 641922 315618 642022
rect 315718 641922 315842 642022
rect 315942 641922 315966 642022
rect 309306 641798 315966 641922
rect 309306 641698 309346 641798
rect 309446 641698 309570 641798
rect 309670 641698 309794 641798
rect 309894 641698 310018 641798
rect 310118 641698 310242 641798
rect 310342 641698 310466 641798
rect 310566 641698 310690 641798
rect 310790 641698 310914 641798
rect 311014 641698 311138 641798
rect 311238 641698 311362 641798
rect 311462 641698 311586 641798
rect 311686 641698 311810 641798
rect 311910 641698 312034 641798
rect 312134 641698 312258 641798
rect 312358 641698 312482 641798
rect 312582 641698 312706 641798
rect 312806 641698 312930 641798
rect 313030 641698 313154 641798
rect 313254 641698 313378 641798
rect 313478 641698 313602 641798
rect 313702 641698 313826 641798
rect 313926 641698 314050 641798
rect 314150 641698 314274 641798
rect 314374 641698 314498 641798
rect 314598 641698 314722 641798
rect 314822 641698 314946 641798
rect 315046 641698 315170 641798
rect 315270 641698 315394 641798
rect 315494 641698 315618 641798
rect 315718 641698 315842 641798
rect 315942 641698 315966 641798
rect 309306 641664 315966 641698
rect 335576 642714 342236 642744
rect 335576 642614 335616 642714
rect 335716 642614 335840 642714
rect 335940 642614 336064 642714
rect 336164 642614 336288 642714
rect 336388 642614 336512 642714
rect 336612 642614 336736 642714
rect 336836 642614 336960 642714
rect 337060 642614 337184 642714
rect 337284 642614 337408 642714
rect 337508 642614 337632 642714
rect 337732 642614 337856 642714
rect 337956 642614 338080 642714
rect 338180 642614 338304 642714
rect 338404 642614 338528 642714
rect 338628 642614 338752 642714
rect 338852 642614 338976 642714
rect 339076 642614 339200 642714
rect 339300 642614 339424 642714
rect 339524 642614 339648 642714
rect 339748 642614 339872 642714
rect 339972 642614 340096 642714
rect 340196 642614 340320 642714
rect 340420 642614 340544 642714
rect 340644 642614 340768 642714
rect 340868 642614 340992 642714
rect 341092 642614 341216 642714
rect 341316 642614 341440 642714
rect 341540 642614 341664 642714
rect 341764 642614 341888 642714
rect 341988 642614 342112 642714
rect 342212 642614 342236 642714
rect 335576 642490 342236 642614
rect 335576 642390 335616 642490
rect 335716 642390 335840 642490
rect 335940 642390 336064 642490
rect 336164 642390 336288 642490
rect 336388 642390 336512 642490
rect 336612 642390 336736 642490
rect 336836 642390 336960 642490
rect 337060 642390 337184 642490
rect 337284 642390 337408 642490
rect 337508 642390 337632 642490
rect 337732 642390 337856 642490
rect 337956 642390 338080 642490
rect 338180 642390 338304 642490
rect 338404 642390 338528 642490
rect 338628 642390 338752 642490
rect 338852 642390 338976 642490
rect 339076 642390 339200 642490
rect 339300 642390 339424 642490
rect 339524 642390 339648 642490
rect 339748 642390 339872 642490
rect 339972 642390 340096 642490
rect 340196 642390 340320 642490
rect 340420 642390 340544 642490
rect 340644 642390 340768 642490
rect 340868 642390 340992 642490
rect 341092 642390 341216 642490
rect 341316 642390 341440 642490
rect 341540 642390 341664 642490
rect 341764 642390 341888 642490
rect 341988 642390 342112 642490
rect 342212 642390 342236 642490
rect 335576 642266 342236 642390
rect 335576 642166 335616 642266
rect 335716 642166 335840 642266
rect 335940 642166 336064 642266
rect 336164 642166 336288 642266
rect 336388 642166 336512 642266
rect 336612 642166 336736 642266
rect 336836 642166 336960 642266
rect 337060 642166 337184 642266
rect 337284 642166 337408 642266
rect 337508 642166 337632 642266
rect 337732 642166 337856 642266
rect 337956 642166 338080 642266
rect 338180 642166 338304 642266
rect 338404 642166 338528 642266
rect 338628 642166 338752 642266
rect 338852 642166 338976 642266
rect 339076 642166 339200 642266
rect 339300 642166 339424 642266
rect 339524 642166 339648 642266
rect 339748 642166 339872 642266
rect 339972 642166 340096 642266
rect 340196 642166 340320 642266
rect 340420 642166 340544 642266
rect 340644 642166 340768 642266
rect 340868 642166 340992 642266
rect 341092 642166 341216 642266
rect 341316 642166 341440 642266
rect 341540 642166 341664 642266
rect 341764 642166 341888 642266
rect 341988 642166 342112 642266
rect 342212 642166 342236 642266
rect 335576 642042 342236 642166
rect 335576 641942 335616 642042
rect 335716 641942 335840 642042
rect 335940 641942 336064 642042
rect 336164 641942 336288 642042
rect 336388 641942 336512 642042
rect 336612 641942 336736 642042
rect 336836 641942 336960 642042
rect 337060 641942 337184 642042
rect 337284 641942 337408 642042
rect 337508 641942 337632 642042
rect 337732 641942 337856 642042
rect 337956 641942 338080 642042
rect 338180 641942 338304 642042
rect 338404 641942 338528 642042
rect 338628 641942 338752 642042
rect 338852 641942 338976 642042
rect 339076 641942 339200 642042
rect 339300 641942 339424 642042
rect 339524 641942 339648 642042
rect 339748 641942 339872 642042
rect 339972 641942 340096 642042
rect 340196 641942 340320 642042
rect 340420 641942 340544 642042
rect 340644 641942 340768 642042
rect 340868 641942 340992 642042
rect 341092 641942 341216 642042
rect 341316 641942 341440 642042
rect 341540 641942 341664 642042
rect 341764 641942 341888 642042
rect 341988 641942 342112 642042
rect 342212 641942 342236 642042
rect 335576 641818 342236 641942
rect 335576 641718 335616 641818
rect 335716 641718 335840 641818
rect 335940 641718 336064 641818
rect 336164 641718 336288 641818
rect 336388 641718 336512 641818
rect 336612 641718 336736 641818
rect 336836 641718 336960 641818
rect 337060 641718 337184 641818
rect 337284 641718 337408 641818
rect 337508 641718 337632 641818
rect 337732 641718 337856 641818
rect 337956 641718 338080 641818
rect 338180 641718 338304 641818
rect 338404 641718 338528 641818
rect 338628 641718 338752 641818
rect 338852 641718 338976 641818
rect 339076 641718 339200 641818
rect 339300 641718 339424 641818
rect 339524 641718 339648 641818
rect 339748 641718 339872 641818
rect 339972 641718 340096 641818
rect 340196 641718 340320 641818
rect 340420 641718 340544 641818
rect 340644 641718 340768 641818
rect 340868 641718 340992 641818
rect 341092 641718 341216 641818
rect 341316 641718 341440 641818
rect 341540 641718 341664 641818
rect 341764 641718 341888 641818
rect 341988 641718 342112 641818
rect 342212 641718 342236 641818
rect 335576 641684 342236 641718
rect 300643 640578 311917 640587
rect 300643 639740 300652 640578
rect 311908 639740 311917 640578
rect 300643 639731 311917 639740
rect 323918 639032 324488 639038
rect 323918 638474 323924 639032
rect 324482 638474 324488 639032
rect 317362 638232 317932 638238
rect 297820 637996 298880 638020
rect 297820 637896 297850 637996
rect 297950 637896 298074 637996
rect 298174 637896 298298 637996
rect 298398 637896 298522 637996
rect 298622 637896 298746 637996
rect 298846 637896 298880 637996
rect 297820 637772 298880 637896
rect 297820 637672 297850 637772
rect 297950 637672 298074 637772
rect 298174 637672 298298 637772
rect 298398 637672 298522 637772
rect 298622 637672 298746 637772
rect 298846 637672 298880 637772
rect 297820 637548 298880 637672
rect 297820 637448 297850 637548
rect 297950 637448 298074 637548
rect 298174 637448 298298 637548
rect 298398 637448 298522 637548
rect 298622 637448 298746 637548
rect 298846 637448 298880 637548
rect 297820 637324 298880 637448
rect 297820 637224 297850 637324
rect 297950 637224 298074 637324
rect 298174 637224 298298 637324
rect 298398 637224 298522 637324
rect 298622 637224 298746 637324
rect 298846 637224 298880 637324
rect 297820 637100 298880 637224
rect 297820 637000 297850 637100
rect 297950 637000 298074 637100
rect 298174 637000 298298 637100
rect 298398 637000 298522 637100
rect 298622 637000 298746 637100
rect 298846 637000 298880 637100
rect 317362 637674 317368 638232
rect 317926 637674 317932 638232
rect 317362 637494 317932 637674
rect 323088 638232 323658 638238
rect 323088 637674 323094 638232
rect 323652 637674 323658 638232
rect 317362 637074 317368 637494
rect 317926 637074 317932 637494
rect 317362 637068 317932 637074
rect 318180 637494 318750 637500
rect 318180 637074 318186 637494
rect 318744 637074 318750 637494
rect 297820 636876 298880 637000
rect 297820 636776 297850 636876
rect 297950 636776 298074 636876
rect 298174 636776 298298 636876
rect 298398 636776 298522 636876
rect 298622 636776 298746 636876
rect 298846 636776 298880 636876
rect 297820 636652 298880 636776
rect 297820 636552 297850 636652
rect 297950 636552 298074 636652
rect 298174 636552 298298 636652
rect 298398 636552 298522 636652
rect 298622 636552 298746 636652
rect 298846 636552 298880 636652
rect 297820 636428 298880 636552
rect 297820 636328 297850 636428
rect 297950 636328 298074 636428
rect 298174 636328 298298 636428
rect 298398 636328 298522 636428
rect 298622 636328 298746 636428
rect 298846 636328 298880 636428
rect 297820 636204 298880 636328
rect 318180 636770 318750 637074
rect 318180 636278 318186 636770
rect 318744 636278 318750 636770
rect 318180 636268 318750 636278
rect 322270 637432 322840 637438
rect 322270 637012 322276 637432
rect 322834 637012 322840 637432
rect 322270 636770 322840 637012
rect 323088 637432 323658 637674
rect 323918 637438 324488 638474
rect 325542 639032 326112 639038
rect 325542 638474 325548 639032
rect 326106 638474 326112 639032
rect 323088 637012 323094 637432
rect 323652 637012 323658 637432
rect 323088 637006 323658 637012
rect 323906 637432 324488 637438
rect 323906 637012 323912 637432
rect 324470 637024 324488 637432
rect 324724 637432 325294 637438
rect 324470 637012 324476 637024
rect 323906 637006 324476 637012
rect 324724 637012 324730 637432
rect 325288 637012 325294 637432
rect 322270 636212 322276 636770
rect 322834 636212 322840 636770
rect 322270 636206 322840 636212
rect 324724 636770 325294 637012
rect 325542 637432 326112 638474
rect 329632 639032 330202 639038
rect 329632 638474 329638 639032
rect 330196 638474 330202 639032
rect 325542 637012 325548 637432
rect 326106 637012 326112 637432
rect 325542 637006 326112 637012
rect 326360 638232 326930 638238
rect 326360 637674 326366 638232
rect 326924 637674 326930 638232
rect 326360 637432 326930 637674
rect 328814 638232 329384 638238
rect 328814 637674 328820 638232
rect 329378 637674 329384 638232
rect 326360 637012 326366 637432
rect 326924 637012 326930 637432
rect 326360 637006 326930 637012
rect 327178 637432 327748 637438
rect 327178 637012 327184 637432
rect 327742 637012 327748 637432
rect 324724 636212 324730 636770
rect 325288 636212 325294 636770
rect 324724 636206 325294 636212
rect 327178 636770 327748 637012
rect 327178 636212 327184 636770
rect 327742 636212 327748 636770
rect 327178 636206 327748 636212
rect 327996 637432 328566 637438
rect 327996 637012 328002 637432
rect 328560 637012 328566 637432
rect 297820 636104 297850 636204
rect 297950 636104 298074 636204
rect 298174 636104 298298 636204
rect 298398 636104 298522 636204
rect 298622 636104 298746 636204
rect 298846 636104 298880 636204
rect 297820 635980 298880 636104
rect 297820 635880 297850 635980
rect 297950 635880 298074 635980
rect 298174 635880 298298 635980
rect 298398 635880 298522 635980
rect 298622 635880 298746 635980
rect 298846 635880 298880 635980
rect 297820 635756 298880 635880
rect 297820 635656 297850 635756
rect 297950 635656 298074 635756
rect 298174 635656 298298 635756
rect 298398 635656 298522 635756
rect 298622 635656 298746 635756
rect 298846 635656 298880 635756
rect 297820 635532 298880 635656
rect 297820 635432 297850 635532
rect 297950 635432 298074 635532
rect 298174 635432 298298 635532
rect 298398 635432 298522 635532
rect 298622 635432 298746 635532
rect 298846 635432 298880 635532
rect 297820 635308 298880 635432
rect 297820 635208 297850 635308
rect 297950 635208 298074 635308
rect 298174 635208 298298 635308
rect 298398 635208 298522 635308
rect 298622 635208 298746 635308
rect 298846 635208 298880 635308
rect 297820 635084 298880 635208
rect 297820 634984 297850 635084
rect 297950 634984 298074 635084
rect 298174 634984 298298 635084
rect 298398 634984 298522 635084
rect 298622 634984 298746 635084
rect 298846 634984 298880 635084
rect 297820 634860 298880 634984
rect 297820 634760 297850 634860
rect 297950 634760 298074 634860
rect 298174 634760 298298 634860
rect 298398 634760 298522 634860
rect 298622 634760 298746 634860
rect 298846 634760 298880 634860
rect 297820 634636 298880 634760
rect 297820 634536 297850 634636
rect 297950 634536 298074 634636
rect 298174 634536 298298 634636
rect 298398 634536 298522 634636
rect 298622 634536 298746 634636
rect 298846 634536 298880 634636
rect 297820 634412 298880 634536
rect 297820 634312 297850 634412
rect 297950 634312 298074 634412
rect 298174 634312 298298 634412
rect 298398 634312 298522 634412
rect 298622 634312 298746 634412
rect 298846 634312 298880 634412
rect 297820 634188 298880 634312
rect 297820 634088 297850 634188
rect 297950 634088 298074 634188
rect 298174 634088 298298 634188
rect 298398 634088 298522 634188
rect 298622 634088 298746 634188
rect 298846 634088 298880 634188
rect 297820 633964 298880 634088
rect 327996 634576 328566 637012
rect 328814 637432 329384 637674
rect 328814 637012 328820 637432
rect 329378 637012 329384 637432
rect 328814 637006 329384 637012
rect 329632 637432 330202 638474
rect 332092 639032 332656 639038
rect 332650 638474 332656 639032
rect 332092 638468 332656 638474
rect 331268 638232 331838 638238
rect 331268 637674 331274 638232
rect 331832 637674 331838 638232
rect 329632 637012 329638 637432
rect 330196 637012 330202 637432
rect 329632 637006 330202 637012
rect 330450 637432 331020 637438
rect 330450 637012 330456 637432
rect 331014 637012 331020 637432
rect 330450 636770 331020 637012
rect 331268 637432 331838 637674
rect 331268 637012 331274 637432
rect 331832 637012 331838 637432
rect 331268 637006 331838 637012
rect 332086 637432 332656 638468
rect 333722 638232 334292 638238
rect 333722 637674 333728 638232
rect 334286 637674 334292 638232
rect 332086 637012 332092 637432
rect 332650 637012 332656 637432
rect 332086 637006 332656 637012
rect 332904 637432 333474 637438
rect 332904 637012 332910 637432
rect 333468 637012 333474 637432
rect 330450 636212 330456 636770
rect 331014 636212 331020 636770
rect 330450 636206 331020 636212
rect 332904 636770 333474 637012
rect 333722 637432 334292 637674
rect 333722 637012 333728 637432
rect 334286 637012 334292 637432
rect 333722 637006 334292 637012
rect 342100 637996 343160 638020
rect 342100 637896 342130 637996
rect 342230 637896 342354 637996
rect 342454 637896 342578 637996
rect 342678 637896 342802 637996
rect 342902 637896 343026 637996
rect 343126 637896 343160 637996
rect 342100 637772 343160 637896
rect 342100 637672 342130 637772
rect 342230 637672 342354 637772
rect 342454 637672 342578 637772
rect 342678 637672 342802 637772
rect 342902 637672 343026 637772
rect 343126 637672 343160 637772
rect 342100 637548 343160 637672
rect 342100 637448 342130 637548
rect 342230 637448 342354 637548
rect 342454 637448 342578 637548
rect 342678 637448 342802 637548
rect 342902 637448 343026 637548
rect 343126 637448 343160 637548
rect 342100 637324 343160 637448
rect 342100 637224 342130 637324
rect 342230 637224 342354 637324
rect 342454 637224 342578 637324
rect 342678 637224 342802 637324
rect 342902 637224 343026 637324
rect 343126 637224 343160 637324
rect 342100 637100 343160 637224
rect 332904 636212 332910 636770
rect 333468 636212 333474 636770
rect 332904 636206 333474 636212
rect 342100 637000 342130 637100
rect 342230 637000 342354 637100
rect 342454 637000 342578 637100
rect 342678 637000 342802 637100
rect 342902 637000 343026 637100
rect 343126 637000 343160 637100
rect 342100 636876 343160 637000
rect 342100 636776 342130 636876
rect 342230 636776 342354 636876
rect 342454 636776 342578 636876
rect 342678 636776 342802 636876
rect 342902 636776 343026 636876
rect 343126 636776 343160 636876
rect 342100 636652 343160 636776
rect 342100 636552 342130 636652
rect 342230 636552 342354 636652
rect 342454 636552 342578 636652
rect 342678 636552 342802 636652
rect 342902 636552 343026 636652
rect 343126 636552 343160 636652
rect 342100 636428 343160 636552
rect 342100 636328 342130 636428
rect 342230 636328 342354 636428
rect 342454 636328 342578 636428
rect 342678 636328 342802 636428
rect 342902 636328 343026 636428
rect 343126 636328 343160 636428
rect 342100 636204 343160 636328
rect 342100 636104 342130 636204
rect 342230 636104 342354 636204
rect 342454 636104 342578 636204
rect 342678 636104 342802 636204
rect 342902 636104 343026 636204
rect 343126 636104 343160 636204
rect 342100 635980 343160 636104
rect 342100 635880 342130 635980
rect 342230 635880 342354 635980
rect 342454 635880 342578 635980
rect 342678 635880 342802 635980
rect 342902 635880 343026 635980
rect 343126 635880 343160 635980
rect 342100 635756 343160 635880
rect 342100 635656 342130 635756
rect 342230 635656 342354 635756
rect 342454 635656 342578 635756
rect 342678 635656 342802 635756
rect 342902 635656 343026 635756
rect 343126 635656 343160 635756
rect 342100 635532 343160 635656
rect 342100 635432 342130 635532
rect 342230 635432 342354 635532
rect 342454 635432 342578 635532
rect 342678 635432 342802 635532
rect 342902 635432 343026 635532
rect 343126 635432 343160 635532
rect 342100 635308 343160 635432
rect 342100 635208 342130 635308
rect 342230 635208 342354 635308
rect 342454 635208 342578 635308
rect 342678 635208 342802 635308
rect 342902 635208 343026 635308
rect 343126 635208 343160 635308
rect 342100 635084 343160 635208
rect 342100 634984 342130 635084
rect 342230 634984 342354 635084
rect 342454 634984 342578 635084
rect 342678 634984 342802 635084
rect 342902 634984 343026 635084
rect 343126 634984 343160 635084
rect 342100 634860 343160 634984
rect 342100 634760 342130 634860
rect 342230 634760 342354 634860
rect 342454 634760 342578 634860
rect 342678 634760 342802 634860
rect 342902 634760 343026 634860
rect 343126 634760 343160 634860
rect 342100 634636 343160 634760
rect 327996 634006 334280 634576
rect 297820 633864 297850 633964
rect 297950 633864 298074 633964
rect 298174 633864 298298 633964
rect 298398 633864 298522 633964
rect 298622 633864 298746 633964
rect 298846 633864 298880 633964
rect 297820 633740 298880 633864
rect 297820 633640 297850 633740
rect 297950 633640 298074 633740
rect 298174 633640 298298 633740
rect 298398 633640 298522 633740
rect 298622 633640 298746 633740
rect 298846 633640 298880 633740
rect 297820 633516 298880 633640
rect 297820 633416 297850 633516
rect 297950 633416 298074 633516
rect 298174 633416 298298 633516
rect 298398 633416 298522 633516
rect 298622 633416 298746 633516
rect 298846 633416 298880 633516
rect 297820 633292 298880 633416
rect 297820 633192 297850 633292
rect 297950 633192 298074 633292
rect 298174 633192 298298 633292
rect 298398 633192 298522 633292
rect 298622 633192 298746 633292
rect 298846 633192 298880 633292
rect 297820 633068 298880 633192
rect 297820 632968 297850 633068
rect 297950 632968 298074 633068
rect 298174 632968 298298 633068
rect 298398 632968 298522 633068
rect 298622 632968 298746 633068
rect 298846 632968 298880 633068
rect 297820 632844 298880 632968
rect 297820 632744 297850 632844
rect 297950 632744 298074 632844
rect 298174 632744 298298 632844
rect 298398 632744 298522 632844
rect 298622 632744 298746 632844
rect 298846 632744 298880 632844
rect 297820 632620 298880 632744
rect 297820 632520 297850 632620
rect 297950 632520 298074 632620
rect 298174 632520 298298 632620
rect 298398 632520 298522 632620
rect 298622 632520 298746 632620
rect 298846 632520 298880 632620
rect 297820 632396 298880 632520
rect 297820 632296 297850 632396
rect 297950 632296 298074 632396
rect 298174 632296 298298 632396
rect 298398 632296 298522 632396
rect 298622 632296 298746 632396
rect 298846 632296 298880 632396
rect 297820 632172 298880 632296
rect 297820 632072 297850 632172
rect 297950 632072 298074 632172
rect 298174 632072 298298 632172
rect 298398 632072 298522 632172
rect 298622 632072 298746 632172
rect 298846 632072 298880 632172
rect 297820 631948 298880 632072
rect 297820 631848 297850 631948
rect 297950 631848 298074 631948
rect 298174 631848 298298 631948
rect 298398 631848 298522 631948
rect 298622 631848 298746 631948
rect 298846 631848 298880 631948
rect 297820 631724 298880 631848
rect 297820 631624 297850 631724
rect 297950 631624 298074 631724
rect 298174 631624 298298 631724
rect 298398 631624 298522 631724
rect 298622 631624 298746 631724
rect 298846 631624 298880 631724
rect 297820 631500 298880 631624
rect 297820 631400 297850 631500
rect 297950 631400 298074 631500
rect 298174 631400 298298 631500
rect 298398 631400 298522 631500
rect 298622 631400 298746 631500
rect 298846 631400 298880 631500
rect 297820 631360 298880 631400
rect 323088 632296 323658 632302
rect 323088 631738 323094 632296
rect 323652 631738 323658 632296
rect 322270 630696 322840 630702
rect 322270 630276 322276 630696
rect 322834 630276 322840 630696
rect 322270 630034 322840 630276
rect 323088 630696 323658 631738
rect 326360 632296 326930 632302
rect 326360 631738 326366 632296
rect 326924 631738 326930 632296
rect 323088 630276 323094 630696
rect 323652 630276 323658 630696
rect 323088 630270 323658 630276
rect 323906 631496 324476 631502
rect 323906 630938 323912 631496
rect 324470 630938 324476 631496
rect 323906 630696 324476 630938
rect 325542 631496 326112 631502
rect 325542 630938 325548 631496
rect 326106 630938 326112 631496
rect 323906 630276 323912 630696
rect 324470 630276 324476 630696
rect 323906 630270 324476 630276
rect 324724 630696 325294 630702
rect 324724 630276 324730 630696
rect 325288 630276 325294 630696
rect 322270 629476 322276 630034
rect 322834 629476 322840 630034
rect 324724 630034 325294 630276
rect 325542 630696 326112 630938
rect 325542 630276 325548 630696
rect 326106 630276 326112 630696
rect 325542 630270 326112 630276
rect 326360 630696 326930 631738
rect 328814 632296 329384 632302
rect 328814 631738 328820 632296
rect 329378 631738 329384 632296
rect 326360 630276 326366 630696
rect 326924 630276 326930 630696
rect 326360 630270 326930 630276
rect 327178 630696 327748 630702
rect 327178 630276 327184 630696
rect 327742 630276 327748 630696
rect 327996 630696 328566 630702
rect 327996 630664 328002 630696
rect 328560 630664 328566 630696
rect 328814 630696 329384 631738
rect 331268 632296 331838 632302
rect 331268 631738 331274 632296
rect 331832 631738 331838 632296
rect 324724 629476 324730 630034
rect 325288 629476 325294 630034
rect 327178 630034 327748 630276
rect 327178 629476 327184 630034
rect 327742 629476 327748 630034
rect 327918 630146 327924 630664
rect 328616 630146 328622 630664
rect 328814 630276 328820 630696
rect 329378 630276 329384 630696
rect 328814 630270 329384 630276
rect 329632 631496 330202 631502
rect 329632 630938 329638 631496
rect 330196 630938 330202 631496
rect 329632 630696 330202 630938
rect 329632 630276 329638 630696
rect 330196 630276 330202 630696
rect 329632 630270 330202 630276
rect 330450 630696 331020 630702
rect 330450 630276 330456 630696
rect 331014 630276 331020 630696
rect 322270 629470 322834 629476
rect 324724 629470 325288 629476
rect 327178 629470 327742 629476
rect 327918 629398 328622 630146
rect 330450 630034 331020 630276
rect 331268 630696 331838 631738
rect 333710 630702 334280 634006
rect 342100 634536 342130 634636
rect 342230 634536 342354 634636
rect 342454 634536 342578 634636
rect 342678 634536 342802 634636
rect 342902 634536 343026 634636
rect 343126 634536 343160 634636
rect 342100 634412 343160 634536
rect 342100 634312 342130 634412
rect 342230 634312 342354 634412
rect 342454 634312 342578 634412
rect 342678 634312 342802 634412
rect 342902 634312 343026 634412
rect 343126 634312 343160 634412
rect 342100 634188 343160 634312
rect 342100 634088 342130 634188
rect 342230 634088 342354 634188
rect 342454 634088 342578 634188
rect 342678 634088 342802 634188
rect 342902 634088 343026 634188
rect 343126 634088 343160 634188
rect 342100 633964 343160 634088
rect 342100 633864 342130 633964
rect 342230 633864 342354 633964
rect 342454 633864 342578 633964
rect 342678 633864 342802 633964
rect 342902 633864 343026 633964
rect 343126 633864 343160 633964
rect 342100 633740 343160 633864
rect 342100 633640 342130 633740
rect 342230 633640 342354 633740
rect 342454 633640 342578 633740
rect 342678 633640 342802 633740
rect 342902 633640 343026 633740
rect 343126 633640 343160 633740
rect 342100 633516 343160 633640
rect 342100 633416 342130 633516
rect 342230 633416 342354 633516
rect 342454 633416 342578 633516
rect 342678 633416 342802 633516
rect 342902 633416 343026 633516
rect 343126 633416 343160 633516
rect 342100 633292 343160 633416
rect 342100 633192 342130 633292
rect 342230 633192 342354 633292
rect 342454 633192 342578 633292
rect 342678 633192 342802 633292
rect 342902 633192 343026 633292
rect 343126 633192 343160 633292
rect 342100 633068 343160 633192
rect 342100 632968 342130 633068
rect 342230 632968 342354 633068
rect 342454 632968 342578 633068
rect 342678 632968 342802 633068
rect 342902 632968 343026 633068
rect 343126 632968 343160 633068
rect 342100 632844 343160 632968
rect 342100 632744 342130 632844
rect 342230 632744 342354 632844
rect 342454 632744 342578 632844
rect 342678 632744 342802 632844
rect 342902 632744 343026 632844
rect 343126 632744 343160 632844
rect 342100 632620 343160 632744
rect 342100 632520 342130 632620
rect 342230 632520 342354 632620
rect 342454 632520 342578 632620
rect 342678 632520 342802 632620
rect 342902 632520 343026 632620
rect 343126 632520 343160 632620
rect 342100 632396 343160 632520
rect 342100 632296 342130 632396
rect 342230 632296 342354 632396
rect 342454 632296 342578 632396
rect 342678 632296 342802 632396
rect 342902 632296 343026 632396
rect 343126 632296 343160 632396
rect 342100 632172 343160 632296
rect 342100 632072 342130 632172
rect 342230 632072 342354 632172
rect 342454 632072 342578 632172
rect 342678 632072 342802 632172
rect 342902 632072 343026 632172
rect 343126 632072 343160 632172
rect 342100 631948 343160 632072
rect 342100 631848 342130 631948
rect 342230 631848 342354 631948
rect 342454 631848 342578 631948
rect 342678 631848 342802 631948
rect 342902 631848 343026 631948
rect 343126 631848 343160 631948
rect 342100 631724 343160 631848
rect 342100 631624 342130 631724
rect 342230 631624 342354 631724
rect 342454 631624 342578 631724
rect 342678 631624 342802 631724
rect 342902 631624 343026 631724
rect 343126 631624 343160 631724
rect 342100 631500 343160 631624
rect 342100 631400 342130 631500
rect 342230 631400 342354 631500
rect 342454 631400 342578 631500
rect 342678 631400 342802 631500
rect 342902 631400 343026 631500
rect 343126 631400 343160 631500
rect 342100 631360 343160 631400
rect 331268 630276 331274 630696
rect 331832 630276 331838 630696
rect 331268 630270 331838 630276
rect 332008 630696 332712 630702
rect 330450 629476 330456 630034
rect 331014 629476 331020 630034
rect 332008 630004 332014 630696
rect 332706 630004 332712 630696
rect 332826 630696 333530 630702
rect 332826 630004 332832 630696
rect 333524 630004 333530 630696
rect 333644 630696 334348 630702
rect 333644 630004 333650 630696
rect 334342 630004 334348 630696
rect 332008 629998 332712 630004
rect 333644 629998 334348 630004
rect 330450 629470 331020 629476
rect 319383 628868 319617 628885
rect 319383 628668 319400 628868
rect 319600 628668 319617 628868
rect 319383 628651 319617 628668
rect 319817 628868 320051 628885
rect 319817 628668 319834 628868
rect 320034 628668 320051 628868
rect 319817 628651 320051 628668
rect 320251 628868 320485 628885
rect 320251 628668 320268 628868
rect 320468 628668 320485 628868
rect 320251 628651 320485 628668
rect 320685 628868 320919 628885
rect 320685 628668 320702 628868
rect 320902 628668 320919 628868
rect 320685 628651 320919 628668
rect 321119 628868 321353 628885
rect 321119 628668 321136 628868
rect 321336 628668 321353 628868
rect 321119 628651 321353 628668
rect 321553 628868 321787 628885
rect 321553 628668 321570 628868
rect 321770 628668 321787 628868
rect 321553 628651 321787 628668
rect 321987 628868 322221 628885
rect 321987 628668 322004 628868
rect 322204 628668 322221 628868
rect 321987 628651 322221 628668
rect 322421 628868 322655 628885
rect 322421 628668 322438 628868
rect 322638 628668 322655 628868
rect 322421 628651 322655 628668
rect 322855 628868 323089 628885
rect 322855 628668 322872 628868
rect 323072 628668 323089 628868
rect 322855 628651 323089 628668
rect 323289 628868 323523 628885
rect 323289 628668 323306 628868
rect 323506 628668 323523 628868
rect 323289 628651 323523 628668
rect 323723 628868 323957 628885
rect 323723 628668 323740 628868
rect 323940 628668 323957 628868
rect 323723 628651 323957 628668
rect 324123 628868 324357 628885
rect 324123 628668 324140 628868
rect 324340 628668 324357 628868
rect 324123 628651 324357 628668
rect 324523 628868 324757 628885
rect 324523 628668 324540 628868
rect 324740 628668 324757 628868
rect 324523 628651 324757 628668
rect 324923 628868 325157 628885
rect 324923 628668 324940 628868
rect 325140 628668 325157 628868
rect 324923 628651 325157 628668
rect 325323 628868 325557 628885
rect 325323 628668 325340 628868
rect 325540 628668 325557 628868
rect 325323 628651 325557 628668
rect 325723 628868 325957 628885
rect 325723 628668 325740 628868
rect 325940 628668 325957 628868
rect 325723 628651 325957 628668
rect 326123 628868 326357 628885
rect 326123 628668 326140 628868
rect 326340 628668 326357 628868
rect 326123 628651 326357 628668
rect 326523 628868 326757 628885
rect 326523 628668 326540 628868
rect 326740 628668 326757 628868
rect 326523 628651 326757 628668
rect 326923 628868 327157 628885
rect 326923 628668 326940 628868
rect 327140 628668 327157 628868
rect 326923 628651 327157 628668
rect 327323 628868 327557 628885
rect 327323 628668 327340 628868
rect 327540 628668 327557 628868
rect 327323 628651 327557 628668
rect 319383 628434 319617 628451
rect 319383 628234 319400 628434
rect 319600 628234 319617 628434
rect 319383 628217 319617 628234
rect 319817 628434 320051 628451
rect 319817 628234 319834 628434
rect 320034 628234 320051 628434
rect 319817 628217 320051 628234
rect 320251 628434 320485 628451
rect 320251 628234 320268 628434
rect 320468 628234 320485 628434
rect 320251 628217 320485 628234
rect 320685 628434 320919 628451
rect 320685 628234 320702 628434
rect 320902 628234 320919 628434
rect 320685 628217 320919 628234
rect 321119 628434 321353 628451
rect 321119 628234 321136 628434
rect 321336 628234 321353 628434
rect 321119 628217 321353 628234
rect 321553 628434 321787 628451
rect 321553 628234 321570 628434
rect 321770 628234 321787 628434
rect 321553 628217 321787 628234
rect 321987 628434 322221 628451
rect 321987 628234 322004 628434
rect 322204 628234 322221 628434
rect 321987 628217 322221 628234
rect 322421 628434 322655 628451
rect 322421 628234 322438 628434
rect 322638 628234 322655 628434
rect 322421 628217 322655 628234
rect 322855 628434 323089 628451
rect 322855 628234 322872 628434
rect 323072 628234 323089 628434
rect 322855 628217 323089 628234
rect 323289 628434 323523 628451
rect 323289 628234 323306 628434
rect 323506 628234 323523 628434
rect 323289 628217 323523 628234
rect 323723 628434 323957 628451
rect 323723 628234 323740 628434
rect 323940 628234 323957 628434
rect 323723 628217 323957 628234
rect 327918 628152 328620 629398
rect 328923 628868 329157 628885
rect 328923 628668 328940 628868
rect 329140 628668 329157 628868
rect 328923 628651 329157 628668
rect 329323 628868 329557 628885
rect 329323 628668 329340 628868
rect 329540 628668 329557 628868
rect 329323 628651 329557 628668
rect 329723 628868 329957 628885
rect 329723 628668 329740 628868
rect 329940 628668 329957 628868
rect 329723 628651 329957 628668
rect 330123 628868 330357 628885
rect 330123 628668 330140 628868
rect 330340 628668 330357 628868
rect 330123 628651 330357 628668
rect 330523 628868 330757 628885
rect 330523 628668 330540 628868
rect 330740 628668 330757 628868
rect 330523 628651 330757 628668
rect 330923 628868 331157 628885
rect 330923 628668 330940 628868
rect 331140 628668 331157 628868
rect 330923 628651 331157 628668
rect 331323 628868 331557 628885
rect 331323 628668 331340 628868
rect 331540 628668 331557 628868
rect 331323 628651 331557 628668
rect 331723 628868 331957 628885
rect 331723 628668 331740 628868
rect 331940 628668 331957 628868
rect 331723 628651 331957 628668
rect 332123 628868 332357 628885
rect 332123 628668 332140 628868
rect 332340 628668 332357 628868
rect 332123 628651 332357 628668
rect 327918 628146 332430 628152
rect 319383 628000 319617 628017
rect 319383 627800 319400 628000
rect 319600 627800 319617 628000
rect 319383 627783 319617 627800
rect 319817 628000 320051 628017
rect 319817 627800 319834 628000
rect 320034 627800 320051 628000
rect 319817 627783 320051 627800
rect 320251 628000 320485 628017
rect 320251 627800 320268 628000
rect 320468 627800 320485 628000
rect 320251 627783 320485 627800
rect 320685 628000 320919 628017
rect 320685 627800 320702 628000
rect 320902 627800 320919 628000
rect 320685 627783 320919 627800
rect 321119 628000 321353 628017
rect 321119 627800 321136 628000
rect 321336 627800 321353 628000
rect 321119 627783 321353 627800
rect 321553 628000 321787 628017
rect 321553 627800 321570 628000
rect 321770 627800 321787 628000
rect 321553 627783 321787 627800
rect 321987 628000 322221 628017
rect 321987 627800 322004 628000
rect 322204 627800 322221 628000
rect 321987 627783 322221 627800
rect 322421 628000 322655 628017
rect 322421 627800 322438 628000
rect 322638 627800 322655 628000
rect 322421 627783 322655 627800
rect 322855 628000 323089 628017
rect 322855 627800 322872 628000
rect 323072 627800 323089 628000
rect 322855 627783 323089 627800
rect 323289 628000 323523 628017
rect 323289 627800 323306 628000
rect 323506 627800 323523 628000
rect 323289 627783 323523 627800
rect 323723 628000 323957 628017
rect 323723 627800 323740 628000
rect 323940 627800 323957 628000
rect 323723 627783 323957 627800
rect 327918 627628 331490 628146
rect 332424 627628 332430 628146
rect 327918 627622 332430 627628
rect 312298 627366 333544 627374
rect 312298 627292 313820 627366
rect 315808 627292 327520 627366
rect 329508 627292 332832 627366
rect 312298 626616 312952 627292
rect 333524 626916 333544 627366
rect 312296 626610 312952 626616
rect 312296 626196 312302 626610
rect 312422 626308 312952 626610
rect 333274 626308 333544 626916
rect 312422 626214 313820 626308
rect 315808 626214 327520 626308
rect 329508 626214 333544 626308
rect 312422 626196 333544 626214
rect 312296 626192 333544 626196
rect 312296 626190 312428 626192
rect 302960 626030 303550 626090
rect 302960 625970 302980 626030
rect 303040 625970 303100 626030
rect 303160 625970 303220 626030
rect 303280 625970 303340 626030
rect 303400 625970 303460 626030
rect 303520 625970 303550 626030
rect 302960 625910 303550 625970
rect 302960 625850 302980 625910
rect 303040 625850 303100 625910
rect 303160 625850 303220 625910
rect 303280 625850 303340 625910
rect 303400 625850 303460 625910
rect 303520 625850 303550 625910
rect 297820 624596 298878 624606
rect 297820 624496 297850 624596
rect 297950 624496 298074 624596
rect 298174 624496 298298 624596
rect 298398 624496 298522 624596
rect 298622 624496 298746 624596
rect 298846 624496 298878 624596
rect 297820 624372 298878 624496
rect 297820 624272 297850 624372
rect 297950 624272 298074 624372
rect 298174 624272 298298 624372
rect 298398 624272 298522 624372
rect 298622 624272 298746 624372
rect 298846 624272 298878 624372
rect 297820 624148 298878 624272
rect 297820 624048 297850 624148
rect 297950 624048 298074 624148
rect 298174 624048 298298 624148
rect 298398 624048 298522 624148
rect 298622 624048 298746 624148
rect 298846 624048 298878 624148
rect 297820 623924 298878 624048
rect 302960 624184 303550 625850
rect 311840 625904 334348 625908
rect 311840 625612 311846 625904
rect 311966 625902 334348 625904
rect 311966 625614 316520 625902
rect 318508 625614 324820 625902
rect 326808 625614 333652 625902
rect 334342 625614 334348 625902
rect 311966 625612 334348 625614
rect 311840 625308 334348 625612
rect 302960 624114 302972 624184
rect 303032 624114 303044 624184
rect 303104 624114 303116 624184
rect 303176 624114 303188 624184
rect 303248 624114 303260 624184
rect 303320 624114 303332 624184
rect 303392 624114 303404 624184
rect 303464 624114 303476 624184
rect 303536 624114 303550 624184
rect 302960 624090 303550 624114
rect 302960 624020 302972 624090
rect 303032 624020 303044 624090
rect 303104 624020 303116 624090
rect 303176 624020 303188 624090
rect 303248 624020 303260 624090
rect 303320 624020 303332 624090
rect 303392 624020 303404 624090
rect 303464 624020 303476 624090
rect 303536 624020 303550 624090
rect 302960 624010 303550 624020
rect 342100 624596 343158 624606
rect 342100 624496 342130 624596
rect 342230 624496 342354 624596
rect 342454 624496 342578 624596
rect 342678 624496 342802 624596
rect 342902 624496 343026 624596
rect 343126 624496 343158 624596
rect 342100 624372 343158 624496
rect 342100 624272 342130 624372
rect 342230 624272 342354 624372
rect 342454 624272 342578 624372
rect 342678 624272 342802 624372
rect 342902 624272 343026 624372
rect 343126 624272 343158 624372
rect 342100 624148 343158 624272
rect 342100 624048 342130 624148
rect 342230 624048 342354 624148
rect 342454 624048 342578 624148
rect 342678 624048 342802 624148
rect 342902 624048 343026 624148
rect 343126 624048 343158 624148
rect 297820 623824 297850 623924
rect 297950 623824 298074 623924
rect 298174 623824 298298 623924
rect 298398 623824 298522 623924
rect 298622 623824 298746 623924
rect 298846 623824 298878 623924
rect 297820 623700 298878 623824
rect 297820 623600 297850 623700
rect 297950 623600 298074 623700
rect 298174 623600 298298 623700
rect 298398 623600 298522 623700
rect 298622 623600 298746 623700
rect 298846 623600 298878 623700
rect 297820 623476 298878 623600
rect 342100 623924 343158 624048
rect 342100 623824 342130 623924
rect 342230 623824 342354 623924
rect 342454 623824 342578 623924
rect 342678 623824 342802 623924
rect 342902 623824 343026 623924
rect 343126 623824 343158 623924
rect 342100 623700 343158 623824
rect 342100 623600 342130 623700
rect 342230 623600 342354 623700
rect 342454 623600 342578 623700
rect 342678 623600 342802 623700
rect 342902 623600 343026 623700
rect 343126 623600 343158 623700
rect 297820 623376 297850 623476
rect 297950 623376 298074 623476
rect 298174 623376 298298 623476
rect 298398 623376 298522 623476
rect 298622 623376 298746 623476
rect 298846 623376 298878 623476
rect 297820 623252 298878 623376
rect 297820 623152 297850 623252
rect 297950 623152 298074 623252
rect 298174 623152 298298 623252
rect 298398 623152 298522 623252
rect 298622 623152 298746 623252
rect 298846 623152 298878 623252
rect 297820 623028 298878 623152
rect 297820 622928 297850 623028
rect 297950 622928 298074 623028
rect 298174 622928 298298 623028
rect 298398 622928 298522 623028
rect 298622 622928 298746 623028
rect 298846 622928 298878 623028
rect 297820 622804 298878 622928
rect 332826 623578 338220 623584
rect 332826 622886 332832 623578
rect 333524 622886 337522 623578
rect 338214 622886 338220 623578
rect 332826 622880 338220 622886
rect 342100 623476 343158 623600
rect 342100 623376 342130 623476
rect 342230 623376 342354 623476
rect 342454 623376 342578 623476
rect 342678 623376 342802 623476
rect 342902 623376 343026 623476
rect 343126 623376 343158 623476
rect 342100 623252 343158 623376
rect 342100 623152 342130 623252
rect 342230 623152 342354 623252
rect 342454 623152 342578 623252
rect 342678 623152 342802 623252
rect 342902 623152 343026 623252
rect 343126 623152 343158 623252
rect 342100 623028 343158 623152
rect 342100 622928 342130 623028
rect 342230 622928 342354 623028
rect 342454 622928 342578 623028
rect 342678 622928 342802 623028
rect 342902 622928 343026 623028
rect 343126 622928 343158 623028
rect 297820 622704 297850 622804
rect 297950 622704 298074 622804
rect 298174 622704 298298 622804
rect 298398 622704 298522 622804
rect 298622 622704 298746 622804
rect 298846 622704 298878 622804
rect 297820 622580 298878 622704
rect 297820 622480 297850 622580
rect 297950 622480 298074 622580
rect 298174 622480 298298 622580
rect 298398 622480 298522 622580
rect 298622 622480 298746 622580
rect 298846 622480 298878 622580
rect 342100 622804 343158 622928
rect 342100 622704 342130 622804
rect 342230 622704 342354 622804
rect 342454 622704 342578 622804
rect 342678 622704 342802 622804
rect 342902 622704 343026 622804
rect 343126 622704 343158 622804
rect 342100 622580 343158 622704
rect 297820 622356 298878 622480
rect 306620 622492 312302 622512
rect 306620 622438 306640 622492
rect 306784 622438 307784 622492
rect 307928 622438 308928 622492
rect 309072 622438 312302 622492
rect 306620 622432 312302 622438
rect 312422 622432 312428 622512
rect 342100 622480 342130 622580
rect 342230 622480 342354 622580
rect 342454 622480 342578 622580
rect 342678 622480 342802 622580
rect 342902 622480 343026 622580
rect 343126 622480 343158 622580
rect 297820 622256 297850 622356
rect 297950 622256 298074 622356
rect 298174 622256 298298 622356
rect 298398 622256 298522 622356
rect 298622 622256 298746 622356
rect 298846 622256 298878 622356
rect 306048 622352 311846 622372
rect 306048 622298 306068 622352
rect 306212 622298 307212 622352
rect 307356 622298 308356 622352
rect 308500 622298 311846 622352
rect 306048 622292 311846 622298
rect 311956 622292 311962 622372
rect 342100 622356 343158 622480
rect 297820 622132 298878 622256
rect 297820 622032 297850 622132
rect 297950 622032 298074 622132
rect 298174 622032 298298 622132
rect 298398 622032 298522 622132
rect 298622 622032 298746 622132
rect 298846 622032 298878 622132
rect 297820 621908 298878 622032
rect 297820 621808 297850 621908
rect 297950 621808 298074 621908
rect 298174 621808 298298 621908
rect 298398 621808 298522 621908
rect 298622 621808 298746 621908
rect 298846 621808 298878 621908
rect 297820 621684 298878 621808
rect 297820 621584 297850 621684
rect 297950 621584 298074 621684
rect 298174 621584 298298 621684
rect 298398 621584 298522 621684
rect 298622 621584 298746 621684
rect 298846 621584 298878 621684
rect 297820 621460 298878 621584
rect 297820 621360 297850 621460
rect 297950 621360 298074 621460
rect 298174 621360 298298 621460
rect 298398 621360 298522 621460
rect 298622 621360 298746 621460
rect 298846 621360 298878 621460
rect 297820 621236 298878 621360
rect 297820 621136 297850 621236
rect 297950 621136 298074 621236
rect 298174 621136 298298 621236
rect 298398 621136 298522 621236
rect 298622 621136 298746 621236
rect 298846 621136 298878 621236
rect 297820 621012 298878 621136
rect 297820 620912 297850 621012
rect 297950 620912 298074 621012
rect 298174 620912 298298 621012
rect 298398 620912 298522 621012
rect 298622 620912 298746 621012
rect 298846 620912 298878 621012
rect 297820 620788 298878 620912
rect 297820 620688 297850 620788
rect 297950 620688 298074 620788
rect 298174 620688 298298 620788
rect 298398 620688 298522 620788
rect 298622 620688 298746 620788
rect 298846 620688 298878 620788
rect 297820 620564 298878 620688
rect 297820 620464 297850 620564
rect 297950 620464 298074 620564
rect 298174 620464 298298 620564
rect 298398 620464 298522 620564
rect 298622 620464 298746 620564
rect 298846 620464 298878 620564
rect 342100 622256 342130 622356
rect 342230 622256 342354 622356
rect 342454 622256 342578 622356
rect 342678 622256 342802 622356
rect 342902 622256 343026 622356
rect 343126 622256 343158 622356
rect 342100 622132 343158 622256
rect 342100 622032 342130 622132
rect 342230 622032 342354 622132
rect 342454 622032 342578 622132
rect 342678 622032 342802 622132
rect 342902 622032 343026 622132
rect 343126 622032 343158 622132
rect 342100 621908 343158 622032
rect 342100 621808 342130 621908
rect 342230 621808 342354 621908
rect 342454 621808 342578 621908
rect 342678 621808 342802 621908
rect 342902 621808 343026 621908
rect 343126 621808 343158 621908
rect 342100 621684 343158 621808
rect 342100 621584 342130 621684
rect 342230 621584 342354 621684
rect 342454 621584 342578 621684
rect 342678 621584 342802 621684
rect 342902 621584 343026 621684
rect 343126 621584 343158 621684
rect 342100 621460 343158 621584
rect 342100 621360 342130 621460
rect 342230 621360 342354 621460
rect 342454 621360 342578 621460
rect 342678 621360 342802 621460
rect 342902 621360 343026 621460
rect 343126 621360 343158 621460
rect 342100 621236 343158 621360
rect 342100 621136 342130 621236
rect 342230 621136 342354 621236
rect 342454 621136 342578 621236
rect 342678 621136 342802 621236
rect 342902 621136 343026 621236
rect 343126 621136 343158 621236
rect 342100 621012 343158 621136
rect 342100 620912 342130 621012
rect 342230 620912 342354 621012
rect 342454 620912 342578 621012
rect 342678 620912 342802 621012
rect 342902 620912 343026 621012
rect 343126 620912 343158 621012
rect 342100 620788 343158 620912
rect 342100 620688 342130 620788
rect 342230 620688 342354 620788
rect 342454 620688 342578 620788
rect 342678 620688 342802 620788
rect 342902 620688 343026 620788
rect 343126 620688 343158 620788
rect 342100 620564 343158 620688
rect 297820 620340 298878 620464
rect 300834 620508 303480 620514
rect 300834 620502 302674 620508
rect 300834 620450 300840 620502
rect 300892 620456 302674 620502
rect 302726 620456 303280 620508
rect 300892 620450 303280 620456
rect 303474 620450 303480 620508
rect 300834 620444 303480 620450
rect 342100 620464 342130 620564
rect 342230 620464 342354 620564
rect 342454 620464 342578 620564
rect 342678 620464 342802 620564
rect 342902 620464 343026 620564
rect 343126 620464 343158 620564
rect 297820 620240 297850 620340
rect 297950 620240 298074 620340
rect 298174 620240 298298 620340
rect 298398 620240 298522 620340
rect 298622 620240 298746 620340
rect 298846 620240 298878 620340
rect 342100 620340 343158 620464
rect 297820 620116 298878 620240
rect 300887 620296 309258 620304
rect 300887 620244 301758 620296
rect 301810 620286 309258 620296
rect 301810 620244 306336 620286
rect 300887 620182 306336 620244
rect 306388 620182 306908 620286
rect 306960 620182 307480 620286
rect 307532 620182 308052 620286
rect 308104 620182 308624 620286
rect 308676 620182 309196 620286
rect 309248 620182 309258 620286
rect 300887 620170 309258 620182
rect 342100 620240 342130 620340
rect 342230 620240 342354 620340
rect 342454 620240 342578 620340
rect 342678 620240 342802 620340
rect 342902 620240 343026 620340
rect 343126 620240 343158 620340
rect 297820 620016 297850 620116
rect 297950 620016 298074 620116
rect 298174 620016 298298 620116
rect 298398 620016 298522 620116
rect 298622 620016 298746 620116
rect 298846 620016 298878 620116
rect 297820 619892 298878 620016
rect 297820 619792 297850 619892
rect 297950 619792 298074 619892
rect 298174 619792 298298 619892
rect 298398 619792 298522 619892
rect 298622 619792 298746 619892
rect 298846 619792 298878 619892
rect 303584 620136 313188 620142
rect 303584 620135 304436 620136
rect 303584 619883 303604 620135
rect 304204 619883 304436 620135
rect 303584 619882 304436 619883
rect 304488 619882 304996 620136
rect 305048 619882 305556 620136
rect 305608 619882 306456 620136
rect 306508 619882 307600 620136
rect 307652 619882 308744 620136
rect 308796 619882 309544 620136
rect 309596 619882 310104 620136
rect 310156 619882 310664 620136
rect 310716 620135 312714 620136
rect 310716 619883 312095 620135
rect 312695 619883 312714 620135
rect 310716 619882 312714 619883
rect 313182 619882 313188 620136
rect 303584 619876 313188 619882
rect 342100 620116 343158 620240
rect 342100 620016 342130 620116
rect 342230 620016 342354 620116
rect 342454 620016 342578 620116
rect 342678 620016 342802 620116
rect 342902 620016 343026 620116
rect 343126 620016 343158 620116
rect 342100 619892 343158 620016
rect 297820 619668 298878 619792
rect 306028 619846 309108 619848
rect 306028 619788 306034 619846
rect 306242 619842 307178 619846
rect 306242 619788 306606 619842
rect 306028 619784 306606 619788
rect 306814 619788 307178 619842
rect 307386 619788 307750 619846
rect 307958 619788 308322 619846
rect 308530 619788 308894 619846
rect 309102 619788 309108 619846
rect 306814 619784 309108 619788
rect 306028 619782 309108 619784
rect 342100 619792 342130 619892
rect 342230 619792 342354 619892
rect 342454 619792 342578 619892
rect 342678 619792 342802 619892
rect 342902 619792 343026 619892
rect 343126 619792 343158 619892
rect 306028 619778 307074 619782
rect 297820 619568 297850 619668
rect 297950 619568 298074 619668
rect 298174 619568 298298 619668
rect 298398 619568 298522 619668
rect 298622 619568 298746 619668
rect 298846 619568 298878 619668
rect 297820 619444 298878 619568
rect 297820 619344 297850 619444
rect 297950 619344 298074 619444
rect 298174 619344 298298 619444
rect 298398 619344 298522 619444
rect 298622 619344 298746 619444
rect 298846 619344 298878 619444
rect 297820 619220 298878 619344
rect 297820 619120 297850 619220
rect 297950 619120 298074 619220
rect 298174 619120 298298 619220
rect 298398 619120 298522 619220
rect 298622 619120 298746 619220
rect 298846 619120 298878 619220
rect 297820 618996 298878 619120
rect 297820 618896 297850 618996
rect 297950 618896 298074 618996
rect 298174 618896 298298 618996
rect 298398 618896 298522 618996
rect 298622 618896 298746 618996
rect 298846 618896 298878 618996
rect 297820 618772 298878 618896
rect 297820 618672 297850 618772
rect 297950 618672 298074 618772
rect 298174 618672 298298 618772
rect 298398 618672 298522 618772
rect 298622 618672 298746 618772
rect 298846 618672 298878 618772
rect 342100 619668 343158 619792
rect 342100 619568 342130 619668
rect 342230 619568 342354 619668
rect 342454 619568 342578 619668
rect 342678 619568 342802 619668
rect 342902 619568 343026 619668
rect 343126 619568 343158 619668
rect 342100 619444 343158 619568
rect 342100 619344 342130 619444
rect 342230 619344 342354 619444
rect 342454 619344 342578 619444
rect 342678 619344 342802 619444
rect 342902 619344 343026 619444
rect 343126 619344 343158 619444
rect 342100 619220 343158 619344
rect 342100 619120 342130 619220
rect 342230 619120 342354 619220
rect 342454 619120 342578 619220
rect 342678 619120 342802 619220
rect 342902 619120 343026 619220
rect 343126 619120 343158 619220
rect 342100 618996 343158 619120
rect 342100 618896 342130 618996
rect 342230 618896 342354 618996
rect 342454 618896 342578 618996
rect 342678 618896 342802 618996
rect 342902 618896 343026 618996
rect 343126 618896 343158 618996
rect 342100 618772 343158 618896
rect 297820 618548 298878 618672
rect 297820 618448 297850 618548
rect 297950 618448 298074 618548
rect 298174 618448 298298 618548
rect 298398 618448 298522 618548
rect 298622 618448 298746 618548
rect 298846 618448 298878 618548
rect 297820 618324 298878 618448
rect 297820 618224 297850 618324
rect 297950 618224 298074 618324
rect 298174 618224 298298 618324
rect 298398 618224 298522 618324
rect 298622 618224 298746 618324
rect 298846 618224 298878 618324
rect 297820 618100 298878 618224
rect 297820 618000 297850 618100
rect 297950 618000 298074 618100
rect 298174 618000 298298 618100
rect 298398 618000 298522 618100
rect 298622 618000 298746 618100
rect 298846 618000 298878 618100
rect 297820 617980 298878 618000
rect 331482 618668 336972 618674
rect 331482 617732 331488 618668
rect 332424 618422 336972 618668
rect 332424 618414 336240 618422
rect 332424 617738 334946 618414
rect 335628 617746 336240 618414
rect 336922 617746 336972 618422
rect 342100 618672 342130 618772
rect 342230 618672 342354 618772
rect 342454 618672 342578 618772
rect 342678 618672 342802 618772
rect 342902 618672 343026 618772
rect 343126 618672 343158 618772
rect 342100 618548 343158 618672
rect 342100 618448 342130 618548
rect 342230 618448 342354 618548
rect 342454 618448 342578 618548
rect 342678 618448 342802 618548
rect 342902 618448 343026 618548
rect 343126 618448 343158 618548
rect 342100 618324 343158 618448
rect 342100 618224 342130 618324
rect 342230 618224 342354 618324
rect 342454 618224 342578 618324
rect 342678 618224 342802 618324
rect 342902 618224 343026 618324
rect 343126 618224 343158 618324
rect 342100 618100 343158 618224
rect 342100 618000 342130 618100
rect 342230 618000 342354 618100
rect 342454 618000 342578 618100
rect 342678 618000 342802 618100
rect 342902 618000 343026 618100
rect 343126 618000 343158 618100
rect 342100 617980 343158 618000
rect 335628 617738 336972 617746
rect 332424 617732 336972 617738
rect 331482 617726 336972 617732
rect 302936 617062 312202 617068
rect 302936 616948 302946 617062
rect 312192 616948 312202 617062
rect 302936 616944 312202 616948
rect 312708 617042 329334 617048
rect 312708 616894 312714 617042
rect 313182 617028 329334 617042
rect 313182 616908 314034 617028
rect 314174 616908 314494 617028
rect 314634 616908 314954 617028
rect 315094 616908 315414 617028
rect 315554 616908 315874 617028
rect 316014 616908 316334 617028
rect 316474 616908 316794 617028
rect 316934 616908 317254 617028
rect 317394 616908 317714 617028
rect 317854 616908 318174 617028
rect 318314 616908 319534 617028
rect 319674 616908 319994 617028
rect 320134 616908 320454 617028
rect 320594 616908 320914 617028
rect 321054 616908 321374 617028
rect 321514 616908 321834 617028
rect 321974 616908 322294 617028
rect 322434 616908 322754 617028
rect 322894 616908 323214 617028
rect 323354 616908 323674 617028
rect 323814 616908 325034 617028
rect 325174 616908 325494 617028
rect 325634 616908 325954 617028
rect 326094 616908 326414 617028
rect 326554 616908 326874 617028
rect 327014 616908 327334 617028
rect 327474 616908 327794 617028
rect 327934 616908 328254 617028
rect 328394 616908 328714 617028
rect 328854 616908 329174 617028
rect 329314 616908 329334 617028
rect 313182 616894 329334 616908
rect 312708 616888 329334 616894
rect 303274 616868 303480 616870
rect 303274 616864 310514 616868
rect 303274 616750 303280 616864
rect 303474 616858 310514 616864
rect 303474 616754 304160 616858
rect 304212 616754 304732 616858
rect 304784 616754 305304 616858
rect 305356 616754 309308 616858
rect 309360 616754 309880 616858
rect 309932 616754 310452 616858
rect 310504 616754 310514 616858
rect 314274 616840 314394 616848
rect 315194 616840 315314 616848
rect 316114 616840 316234 616848
rect 317034 616840 317154 616848
rect 317954 616840 318074 616848
rect 319774 616840 319894 616848
rect 320694 616840 320814 616848
rect 321614 616840 321734 616848
rect 322534 616840 322654 616848
rect 323454 616840 323574 616848
rect 325274 616840 325394 616848
rect 326194 616840 326314 616848
rect 327114 616840 327234 616848
rect 328034 616840 328154 616848
rect 328954 616840 329074 616848
rect 303474 616750 310514 616754
rect 303274 616744 310514 616750
rect 312700 616830 330658 616840
rect 312700 616512 312710 616830
rect 330648 616806 330658 616830
rect 330648 616512 330670 616806
rect 312700 616506 330670 616512
rect 312700 616504 330658 616506
rect 298836 615474 305496 615504
rect 298836 615374 298876 615474
rect 298976 615374 299100 615474
rect 299200 615374 299324 615474
rect 299424 615374 299548 615474
rect 299648 615374 299772 615474
rect 299872 615374 299996 615474
rect 300096 615374 300220 615474
rect 300320 615374 300444 615474
rect 300544 615374 300668 615474
rect 300768 615374 300892 615474
rect 300992 615374 301116 615474
rect 301216 615374 301340 615474
rect 301440 615374 301564 615474
rect 301664 615374 301788 615474
rect 301888 615374 302012 615474
rect 302112 615374 302236 615474
rect 302336 615374 302460 615474
rect 302560 615374 302684 615474
rect 302784 615374 302908 615474
rect 303008 615374 303132 615474
rect 303232 615374 303356 615474
rect 303456 615374 303580 615474
rect 303680 615374 303804 615474
rect 303904 615374 304028 615474
rect 304128 615374 304252 615474
rect 304352 615374 304476 615474
rect 304576 615374 304700 615474
rect 304800 615374 304924 615474
rect 305024 615374 305148 615474
rect 305248 615374 305372 615474
rect 305472 615374 305496 615474
rect 298836 615250 305496 615374
rect 298836 615150 298876 615250
rect 298976 615150 299100 615250
rect 299200 615150 299324 615250
rect 299424 615150 299548 615250
rect 299648 615150 299772 615250
rect 299872 615150 299996 615250
rect 300096 615150 300220 615250
rect 300320 615150 300444 615250
rect 300544 615150 300668 615250
rect 300768 615150 300892 615250
rect 300992 615150 301116 615250
rect 301216 615150 301340 615250
rect 301440 615150 301564 615250
rect 301664 615150 301788 615250
rect 301888 615150 302012 615250
rect 302112 615150 302236 615250
rect 302336 615150 302460 615250
rect 302560 615150 302684 615250
rect 302784 615150 302908 615250
rect 303008 615150 303132 615250
rect 303232 615150 303356 615250
rect 303456 615150 303580 615250
rect 303680 615150 303804 615250
rect 303904 615150 304028 615250
rect 304128 615150 304252 615250
rect 304352 615150 304476 615250
rect 304576 615150 304700 615250
rect 304800 615150 304924 615250
rect 305024 615150 305148 615250
rect 305248 615150 305372 615250
rect 305472 615150 305496 615250
rect 298836 615026 305496 615150
rect 298836 614926 298876 615026
rect 298976 614926 299100 615026
rect 299200 614926 299324 615026
rect 299424 614926 299548 615026
rect 299648 614926 299772 615026
rect 299872 614926 299996 615026
rect 300096 614926 300220 615026
rect 300320 614926 300444 615026
rect 300544 614926 300668 615026
rect 300768 614926 300892 615026
rect 300992 614926 301116 615026
rect 301216 614926 301340 615026
rect 301440 614926 301564 615026
rect 301664 614926 301788 615026
rect 301888 614926 302012 615026
rect 302112 614926 302236 615026
rect 302336 614926 302460 615026
rect 302560 614926 302684 615026
rect 302784 614926 302908 615026
rect 303008 614926 303132 615026
rect 303232 614926 303356 615026
rect 303456 614926 303580 615026
rect 303680 614926 303804 615026
rect 303904 614926 304028 615026
rect 304128 614926 304252 615026
rect 304352 614926 304476 615026
rect 304576 614926 304700 615026
rect 304800 614926 304924 615026
rect 305024 614926 305148 615026
rect 305248 614926 305372 615026
rect 305472 614926 305496 615026
rect 298836 614802 305496 614926
rect 298836 614702 298876 614802
rect 298976 614702 299100 614802
rect 299200 614702 299324 614802
rect 299424 614702 299548 614802
rect 299648 614702 299772 614802
rect 299872 614702 299996 614802
rect 300096 614702 300220 614802
rect 300320 614702 300444 614802
rect 300544 614702 300668 614802
rect 300768 614702 300892 614802
rect 300992 614702 301116 614802
rect 301216 614702 301340 614802
rect 301440 614702 301564 614802
rect 301664 614702 301788 614802
rect 301888 614702 302012 614802
rect 302112 614702 302236 614802
rect 302336 614702 302460 614802
rect 302560 614702 302684 614802
rect 302784 614702 302908 614802
rect 303008 614702 303132 614802
rect 303232 614702 303356 614802
rect 303456 614702 303580 614802
rect 303680 614702 303804 614802
rect 303904 614702 304028 614802
rect 304128 614702 304252 614802
rect 304352 614702 304476 614802
rect 304576 614702 304700 614802
rect 304800 614702 304924 614802
rect 305024 614702 305148 614802
rect 305248 614702 305372 614802
rect 305472 614702 305496 614802
rect 298836 614578 305496 614702
rect 298836 614478 298876 614578
rect 298976 614478 299100 614578
rect 299200 614478 299324 614578
rect 299424 614478 299548 614578
rect 299648 614478 299772 614578
rect 299872 614478 299996 614578
rect 300096 614478 300220 614578
rect 300320 614478 300444 614578
rect 300544 614478 300668 614578
rect 300768 614478 300892 614578
rect 300992 614478 301116 614578
rect 301216 614478 301340 614578
rect 301440 614478 301564 614578
rect 301664 614478 301788 614578
rect 301888 614478 302012 614578
rect 302112 614478 302236 614578
rect 302336 614478 302460 614578
rect 302560 614478 302684 614578
rect 302784 614478 302908 614578
rect 303008 614478 303132 614578
rect 303232 614478 303356 614578
rect 303456 614478 303580 614578
rect 303680 614478 303804 614578
rect 303904 614478 304028 614578
rect 304128 614478 304252 614578
rect 304352 614478 304476 614578
rect 304576 614478 304700 614578
rect 304800 614478 304924 614578
rect 305024 614478 305148 614578
rect 305248 614478 305372 614578
rect 305472 614478 305496 614578
rect 298836 614444 305496 614478
rect 309306 615474 315966 615504
rect 309306 615374 309346 615474
rect 309446 615374 309570 615474
rect 309670 615374 309794 615474
rect 309894 615374 310018 615474
rect 310118 615374 310242 615474
rect 310342 615374 310466 615474
rect 310566 615374 310690 615474
rect 310790 615374 310914 615474
rect 311014 615374 311138 615474
rect 311238 615374 311362 615474
rect 311462 615374 311586 615474
rect 311686 615374 311810 615474
rect 311910 615374 312034 615474
rect 312134 615374 312258 615474
rect 312358 615374 312482 615474
rect 312582 615374 312706 615474
rect 312806 615374 312930 615474
rect 313030 615374 313154 615474
rect 313254 615374 313378 615474
rect 313478 615374 313602 615474
rect 313702 615374 313826 615474
rect 313926 615374 314050 615474
rect 314150 615374 314274 615474
rect 314374 615374 314498 615474
rect 314598 615374 314722 615474
rect 314822 615374 314946 615474
rect 315046 615374 315170 615474
rect 315270 615374 315394 615474
rect 315494 615374 315618 615474
rect 315718 615374 315842 615474
rect 315942 615374 315966 615474
rect 309306 615250 315966 615374
rect 309306 615150 309346 615250
rect 309446 615150 309570 615250
rect 309670 615150 309794 615250
rect 309894 615150 310018 615250
rect 310118 615150 310242 615250
rect 310342 615150 310466 615250
rect 310566 615150 310690 615250
rect 310790 615150 310914 615250
rect 311014 615150 311138 615250
rect 311238 615150 311362 615250
rect 311462 615150 311586 615250
rect 311686 615150 311810 615250
rect 311910 615150 312034 615250
rect 312134 615150 312258 615250
rect 312358 615150 312482 615250
rect 312582 615150 312706 615250
rect 312806 615150 312930 615250
rect 313030 615150 313154 615250
rect 313254 615150 313378 615250
rect 313478 615150 313602 615250
rect 313702 615150 313826 615250
rect 313926 615150 314050 615250
rect 314150 615150 314274 615250
rect 314374 615150 314498 615250
rect 314598 615150 314722 615250
rect 314822 615150 314946 615250
rect 315046 615150 315170 615250
rect 315270 615150 315394 615250
rect 315494 615150 315618 615250
rect 315718 615150 315842 615250
rect 315942 615150 315966 615250
rect 309306 615026 315966 615150
rect 309306 614926 309346 615026
rect 309446 614926 309570 615026
rect 309670 614926 309794 615026
rect 309894 614926 310018 615026
rect 310118 614926 310242 615026
rect 310342 614926 310466 615026
rect 310566 614926 310690 615026
rect 310790 614926 310914 615026
rect 311014 614926 311138 615026
rect 311238 614926 311362 615026
rect 311462 614926 311586 615026
rect 311686 614926 311810 615026
rect 311910 614926 312034 615026
rect 312134 614926 312258 615026
rect 312358 614926 312482 615026
rect 312582 614926 312706 615026
rect 312806 614926 312930 615026
rect 313030 614926 313154 615026
rect 313254 614926 313378 615026
rect 313478 614926 313602 615026
rect 313702 614926 313826 615026
rect 313926 614926 314050 615026
rect 314150 614926 314274 615026
rect 314374 614926 314498 615026
rect 314598 614926 314722 615026
rect 314822 614926 314946 615026
rect 315046 614926 315170 615026
rect 315270 614926 315394 615026
rect 315494 614926 315618 615026
rect 315718 614926 315842 615026
rect 315942 614926 315966 615026
rect 309306 614802 315966 614926
rect 309306 614702 309346 614802
rect 309446 614702 309570 614802
rect 309670 614702 309794 614802
rect 309894 614702 310018 614802
rect 310118 614702 310242 614802
rect 310342 614702 310466 614802
rect 310566 614702 310690 614802
rect 310790 614702 310914 614802
rect 311014 614702 311138 614802
rect 311238 614702 311362 614802
rect 311462 614702 311586 614802
rect 311686 614702 311810 614802
rect 311910 614702 312034 614802
rect 312134 614702 312258 614802
rect 312358 614702 312482 614802
rect 312582 614702 312706 614802
rect 312806 614702 312930 614802
rect 313030 614702 313154 614802
rect 313254 614702 313378 614802
rect 313478 614702 313602 614802
rect 313702 614702 313826 614802
rect 313926 614702 314050 614802
rect 314150 614702 314274 614802
rect 314374 614702 314498 614802
rect 314598 614702 314722 614802
rect 314822 614702 314946 614802
rect 315046 614702 315170 614802
rect 315270 614702 315394 614802
rect 315494 614702 315618 614802
rect 315718 614702 315842 614802
rect 315942 614702 315966 614802
rect 309306 614578 315966 614702
rect 309306 614478 309346 614578
rect 309446 614478 309570 614578
rect 309670 614478 309794 614578
rect 309894 614478 310018 614578
rect 310118 614478 310242 614578
rect 310342 614478 310466 614578
rect 310566 614478 310690 614578
rect 310790 614478 310914 614578
rect 311014 614478 311138 614578
rect 311238 614478 311362 614578
rect 311462 614478 311586 614578
rect 311686 614478 311810 614578
rect 311910 614478 312034 614578
rect 312134 614478 312258 614578
rect 312358 614478 312482 614578
rect 312582 614478 312706 614578
rect 312806 614478 312930 614578
rect 313030 614478 313154 614578
rect 313254 614478 313378 614578
rect 313478 614478 313602 614578
rect 313702 614478 313826 614578
rect 313926 614478 314050 614578
rect 314150 614478 314274 614578
rect 314374 614478 314498 614578
rect 314598 614478 314722 614578
rect 314822 614478 314946 614578
rect 315046 614478 315170 614578
rect 315270 614478 315394 614578
rect 315494 614478 315618 614578
rect 315718 614478 315842 614578
rect 315942 614478 315966 614578
rect 309306 614444 315966 614478
rect 335576 615494 342236 615524
rect 335576 615394 335616 615494
rect 335716 615394 335840 615494
rect 335940 615394 336064 615494
rect 336164 615394 336288 615494
rect 336388 615394 336512 615494
rect 336612 615394 336736 615494
rect 336836 615394 336960 615494
rect 337060 615394 337184 615494
rect 337284 615394 337408 615494
rect 337508 615394 337632 615494
rect 337732 615394 337856 615494
rect 337956 615394 338080 615494
rect 338180 615394 338304 615494
rect 338404 615394 338528 615494
rect 338628 615394 338752 615494
rect 338852 615394 338976 615494
rect 339076 615394 339200 615494
rect 339300 615394 339424 615494
rect 339524 615394 339648 615494
rect 339748 615394 339872 615494
rect 339972 615394 340096 615494
rect 340196 615394 340320 615494
rect 340420 615394 340544 615494
rect 340644 615394 340768 615494
rect 340868 615394 340992 615494
rect 341092 615394 341216 615494
rect 341316 615394 341440 615494
rect 341540 615394 341664 615494
rect 341764 615394 341888 615494
rect 341988 615394 342112 615494
rect 342212 615394 342236 615494
rect 335576 615270 342236 615394
rect 335576 615170 335616 615270
rect 335716 615170 335840 615270
rect 335940 615170 336064 615270
rect 336164 615170 336288 615270
rect 336388 615170 336512 615270
rect 336612 615170 336736 615270
rect 336836 615170 336960 615270
rect 337060 615170 337184 615270
rect 337284 615170 337408 615270
rect 337508 615170 337632 615270
rect 337732 615170 337856 615270
rect 337956 615170 338080 615270
rect 338180 615170 338304 615270
rect 338404 615170 338528 615270
rect 338628 615170 338752 615270
rect 338852 615170 338976 615270
rect 339076 615170 339200 615270
rect 339300 615170 339424 615270
rect 339524 615170 339648 615270
rect 339748 615170 339872 615270
rect 339972 615170 340096 615270
rect 340196 615170 340320 615270
rect 340420 615170 340544 615270
rect 340644 615170 340768 615270
rect 340868 615170 340992 615270
rect 341092 615170 341216 615270
rect 341316 615170 341440 615270
rect 341540 615170 341664 615270
rect 341764 615170 341888 615270
rect 341988 615170 342112 615270
rect 342212 615170 342236 615270
rect 335576 615046 342236 615170
rect 335576 614946 335616 615046
rect 335716 614946 335840 615046
rect 335940 614946 336064 615046
rect 336164 614946 336288 615046
rect 336388 614946 336512 615046
rect 336612 614946 336736 615046
rect 336836 614946 336960 615046
rect 337060 614946 337184 615046
rect 337284 614946 337408 615046
rect 337508 614946 337632 615046
rect 337732 614946 337856 615046
rect 337956 614946 338080 615046
rect 338180 614946 338304 615046
rect 338404 614946 338528 615046
rect 338628 614946 338752 615046
rect 338852 614946 338976 615046
rect 339076 614946 339200 615046
rect 339300 614946 339424 615046
rect 339524 614946 339648 615046
rect 339748 614946 339872 615046
rect 339972 614946 340096 615046
rect 340196 614946 340320 615046
rect 340420 614946 340544 615046
rect 340644 614946 340768 615046
rect 340868 614946 340992 615046
rect 341092 614946 341216 615046
rect 341316 614946 341440 615046
rect 341540 614946 341664 615046
rect 341764 614946 341888 615046
rect 341988 614946 342112 615046
rect 342212 614946 342236 615046
rect 335576 614822 342236 614946
rect 335576 614722 335616 614822
rect 335716 614722 335840 614822
rect 335940 614722 336064 614822
rect 336164 614722 336288 614822
rect 336388 614722 336512 614822
rect 336612 614722 336736 614822
rect 336836 614722 336960 614822
rect 337060 614722 337184 614822
rect 337284 614722 337408 614822
rect 337508 614722 337632 614822
rect 337732 614722 337856 614822
rect 337956 614722 338080 614822
rect 338180 614722 338304 614822
rect 338404 614722 338528 614822
rect 338628 614722 338752 614822
rect 338852 614722 338976 614822
rect 339076 614722 339200 614822
rect 339300 614722 339424 614822
rect 339524 614722 339648 614822
rect 339748 614722 339872 614822
rect 339972 614722 340096 614822
rect 340196 614722 340320 614822
rect 340420 614722 340544 614822
rect 340644 614722 340768 614822
rect 340868 614722 340992 614822
rect 341092 614722 341216 614822
rect 341316 614722 341440 614822
rect 341540 614722 341664 614822
rect 341764 614722 341888 614822
rect 341988 614722 342112 614822
rect 342212 614722 342236 614822
rect 335576 614598 342236 614722
rect 335576 614498 335616 614598
rect 335716 614498 335840 614598
rect 335940 614498 336064 614598
rect 336164 614498 336288 614598
rect 336388 614498 336512 614598
rect 336612 614498 336736 614598
rect 336836 614498 336960 614598
rect 337060 614498 337184 614598
rect 337284 614498 337408 614598
rect 337508 614498 337632 614598
rect 337732 614498 337856 614598
rect 337956 614498 338080 614598
rect 338180 614498 338304 614598
rect 338404 614498 338528 614598
rect 338628 614498 338752 614598
rect 338852 614498 338976 614598
rect 339076 614498 339200 614598
rect 339300 614498 339424 614598
rect 339524 614498 339648 614598
rect 339748 614498 339872 614598
rect 339972 614498 340096 614598
rect 340196 614498 340320 614598
rect 340420 614498 340544 614598
rect 340644 614498 340768 614598
rect 340868 614498 340992 614598
rect 341092 614498 341216 614598
rect 341316 614498 341440 614598
rect 341540 614498 341664 614598
rect 341764 614498 341888 614598
rect 341988 614498 342112 614598
rect 342212 614498 342236 614598
rect 335576 614464 342236 614498
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 298876 642594 298976 642694
rect 299100 642594 299200 642694
rect 299324 642594 299424 642694
rect 299548 642594 299648 642694
rect 299772 642594 299872 642694
rect 299996 642594 300096 642694
rect 300220 642594 300320 642694
rect 300444 642594 300544 642694
rect 300668 642594 300768 642694
rect 300892 642594 300992 642694
rect 301116 642594 301216 642694
rect 301340 642594 301440 642694
rect 301564 642594 301664 642694
rect 301788 642594 301888 642694
rect 302012 642594 302112 642694
rect 302236 642594 302336 642694
rect 302460 642594 302560 642694
rect 302684 642594 302784 642694
rect 302908 642594 303008 642694
rect 303132 642594 303232 642694
rect 303356 642594 303456 642694
rect 303580 642594 303680 642694
rect 303804 642594 303904 642694
rect 304028 642594 304128 642694
rect 304252 642594 304352 642694
rect 304476 642594 304576 642694
rect 304700 642594 304800 642694
rect 304924 642594 305024 642694
rect 305148 642594 305248 642694
rect 305372 642594 305472 642694
rect 298876 642370 298976 642470
rect 299100 642370 299200 642470
rect 299324 642370 299424 642470
rect 299548 642370 299648 642470
rect 299772 642370 299872 642470
rect 299996 642370 300096 642470
rect 300220 642370 300320 642470
rect 300444 642370 300544 642470
rect 300668 642370 300768 642470
rect 300892 642370 300992 642470
rect 301116 642370 301216 642470
rect 301340 642370 301440 642470
rect 301564 642370 301664 642470
rect 301788 642370 301888 642470
rect 302012 642370 302112 642470
rect 302236 642370 302336 642470
rect 302460 642370 302560 642470
rect 302684 642370 302784 642470
rect 302908 642370 303008 642470
rect 303132 642370 303232 642470
rect 303356 642370 303456 642470
rect 303580 642370 303680 642470
rect 303804 642370 303904 642470
rect 304028 642370 304128 642470
rect 304252 642370 304352 642470
rect 304476 642370 304576 642470
rect 304700 642370 304800 642470
rect 304924 642370 305024 642470
rect 305148 642370 305248 642470
rect 305372 642370 305472 642470
rect 298876 642146 298976 642246
rect 299100 642146 299200 642246
rect 299324 642146 299424 642246
rect 299548 642146 299648 642246
rect 299772 642146 299872 642246
rect 299996 642146 300096 642246
rect 300220 642146 300320 642246
rect 300444 642146 300544 642246
rect 300668 642146 300768 642246
rect 300892 642146 300992 642246
rect 301116 642146 301216 642246
rect 301340 642146 301440 642246
rect 301564 642146 301664 642246
rect 301788 642146 301888 642246
rect 302012 642146 302112 642246
rect 302236 642146 302336 642246
rect 302460 642146 302560 642246
rect 302684 642146 302784 642246
rect 302908 642146 303008 642246
rect 303132 642146 303232 642246
rect 303356 642146 303456 642246
rect 303580 642146 303680 642246
rect 303804 642146 303904 642246
rect 304028 642146 304128 642246
rect 304252 642146 304352 642246
rect 304476 642146 304576 642246
rect 304700 642146 304800 642246
rect 304924 642146 305024 642246
rect 305148 642146 305248 642246
rect 305372 642146 305472 642246
rect 298876 641922 298976 642022
rect 299100 641922 299200 642022
rect 299324 641922 299424 642022
rect 299548 641922 299648 642022
rect 299772 641922 299872 642022
rect 299996 641922 300096 642022
rect 300220 641922 300320 642022
rect 300444 641922 300544 642022
rect 300668 641922 300768 642022
rect 300892 641922 300992 642022
rect 301116 641922 301216 642022
rect 301340 641922 301440 642022
rect 301564 641922 301664 642022
rect 301788 641922 301888 642022
rect 302012 641922 302112 642022
rect 302236 641922 302336 642022
rect 302460 641922 302560 642022
rect 302684 641922 302784 642022
rect 302908 641922 303008 642022
rect 303132 641922 303232 642022
rect 303356 641922 303456 642022
rect 303580 641922 303680 642022
rect 303804 641922 303904 642022
rect 304028 641922 304128 642022
rect 304252 641922 304352 642022
rect 304476 641922 304576 642022
rect 304700 641922 304800 642022
rect 304924 641922 305024 642022
rect 305148 641922 305248 642022
rect 305372 641922 305472 642022
rect 298876 641698 298976 641798
rect 299100 641698 299200 641798
rect 299324 641698 299424 641798
rect 299548 641698 299648 641798
rect 299772 641698 299872 641798
rect 299996 641698 300096 641798
rect 300220 641698 300320 641798
rect 300444 641698 300544 641798
rect 300668 641698 300768 641798
rect 300892 641698 300992 641798
rect 301116 641698 301216 641798
rect 301340 641698 301440 641798
rect 301564 641698 301664 641798
rect 301788 641698 301888 641798
rect 302012 641698 302112 641798
rect 302236 641698 302336 641798
rect 302460 641698 302560 641798
rect 302684 641698 302784 641798
rect 302908 641698 303008 641798
rect 303132 641698 303232 641798
rect 303356 641698 303456 641798
rect 303580 641698 303680 641798
rect 303804 641698 303904 641798
rect 304028 641698 304128 641798
rect 304252 641698 304352 641798
rect 304476 641698 304576 641798
rect 304700 641698 304800 641798
rect 304924 641698 305024 641798
rect 305148 641698 305248 641798
rect 305372 641698 305472 641798
rect 309346 642594 309446 642694
rect 309570 642594 309670 642694
rect 309794 642594 309894 642694
rect 310018 642594 310118 642694
rect 310242 642594 310342 642694
rect 310466 642594 310566 642694
rect 310690 642594 310790 642694
rect 310914 642594 311014 642694
rect 311138 642594 311238 642694
rect 311362 642594 311462 642694
rect 311586 642594 311686 642694
rect 311810 642594 311910 642694
rect 312034 642594 312134 642694
rect 312258 642594 312358 642694
rect 312482 642594 312582 642694
rect 312706 642594 312806 642694
rect 312930 642594 313030 642694
rect 313154 642594 313254 642694
rect 313378 642594 313478 642694
rect 313602 642594 313702 642694
rect 313826 642594 313926 642694
rect 314050 642594 314150 642694
rect 314274 642594 314374 642694
rect 314498 642594 314598 642694
rect 314722 642594 314822 642694
rect 314946 642594 315046 642694
rect 315170 642594 315270 642694
rect 315394 642594 315494 642694
rect 315618 642594 315718 642694
rect 315842 642594 315942 642694
rect 309346 642370 309446 642470
rect 309570 642370 309670 642470
rect 309794 642370 309894 642470
rect 310018 642370 310118 642470
rect 310242 642370 310342 642470
rect 310466 642370 310566 642470
rect 310690 642370 310790 642470
rect 310914 642370 311014 642470
rect 311138 642370 311238 642470
rect 311362 642370 311462 642470
rect 311586 642370 311686 642470
rect 311810 642370 311910 642470
rect 312034 642370 312134 642470
rect 312258 642370 312358 642470
rect 312482 642370 312582 642470
rect 312706 642370 312806 642470
rect 312930 642370 313030 642470
rect 313154 642370 313254 642470
rect 313378 642370 313478 642470
rect 313602 642370 313702 642470
rect 313826 642370 313926 642470
rect 314050 642370 314150 642470
rect 314274 642370 314374 642470
rect 314498 642370 314598 642470
rect 314722 642370 314822 642470
rect 314946 642370 315046 642470
rect 315170 642370 315270 642470
rect 315394 642370 315494 642470
rect 315618 642370 315718 642470
rect 315842 642370 315942 642470
rect 309346 642146 309446 642246
rect 309570 642146 309670 642246
rect 309794 642146 309894 642246
rect 310018 642146 310118 642246
rect 310242 642146 310342 642246
rect 310466 642146 310566 642246
rect 310690 642146 310790 642246
rect 310914 642146 311014 642246
rect 311138 642146 311238 642246
rect 311362 642146 311462 642246
rect 311586 642146 311686 642246
rect 311810 642146 311910 642246
rect 312034 642146 312134 642246
rect 312258 642146 312358 642246
rect 312482 642146 312582 642246
rect 312706 642146 312806 642246
rect 312930 642146 313030 642246
rect 313154 642146 313254 642246
rect 313378 642146 313478 642246
rect 313602 642146 313702 642246
rect 313826 642146 313926 642246
rect 314050 642146 314150 642246
rect 314274 642146 314374 642246
rect 314498 642146 314598 642246
rect 314722 642146 314822 642246
rect 314946 642146 315046 642246
rect 315170 642146 315270 642246
rect 315394 642146 315494 642246
rect 315618 642146 315718 642246
rect 315842 642146 315942 642246
rect 309346 641922 309446 642022
rect 309570 641922 309670 642022
rect 309794 641922 309894 642022
rect 310018 641922 310118 642022
rect 310242 641922 310342 642022
rect 310466 641922 310566 642022
rect 310690 641922 310790 642022
rect 310914 641922 311014 642022
rect 311138 641922 311238 642022
rect 311362 641922 311462 642022
rect 311586 641922 311686 642022
rect 311810 641922 311910 642022
rect 312034 641922 312134 642022
rect 312258 641922 312358 642022
rect 312482 641922 312582 642022
rect 312706 641922 312806 642022
rect 312930 641922 313030 642022
rect 313154 641922 313254 642022
rect 313378 641922 313478 642022
rect 313602 641922 313702 642022
rect 313826 641922 313926 642022
rect 314050 641922 314150 642022
rect 314274 641922 314374 642022
rect 314498 641922 314598 642022
rect 314722 641922 314822 642022
rect 314946 641922 315046 642022
rect 315170 641922 315270 642022
rect 315394 641922 315494 642022
rect 315618 641922 315718 642022
rect 315842 641922 315942 642022
rect 309346 641698 309446 641798
rect 309570 641698 309670 641798
rect 309794 641698 309894 641798
rect 310018 641698 310118 641798
rect 310242 641698 310342 641798
rect 310466 641698 310566 641798
rect 310690 641698 310790 641798
rect 310914 641698 311014 641798
rect 311138 641698 311238 641798
rect 311362 641698 311462 641798
rect 311586 641698 311686 641798
rect 311810 641698 311910 641798
rect 312034 641698 312134 641798
rect 312258 641698 312358 641798
rect 312482 641698 312582 641798
rect 312706 641698 312806 641798
rect 312930 641698 313030 641798
rect 313154 641698 313254 641798
rect 313378 641698 313478 641798
rect 313602 641698 313702 641798
rect 313826 641698 313926 641798
rect 314050 641698 314150 641798
rect 314274 641698 314374 641798
rect 314498 641698 314598 641798
rect 314722 641698 314822 641798
rect 314946 641698 315046 641798
rect 315170 641698 315270 641798
rect 315394 641698 315494 641798
rect 315618 641698 315718 641798
rect 315842 641698 315942 641798
rect 335616 642614 335716 642714
rect 335840 642614 335940 642714
rect 336064 642614 336164 642714
rect 336288 642614 336388 642714
rect 336512 642614 336612 642714
rect 336736 642614 336836 642714
rect 336960 642614 337060 642714
rect 337184 642614 337284 642714
rect 337408 642614 337508 642714
rect 337632 642614 337732 642714
rect 337856 642614 337956 642714
rect 338080 642614 338180 642714
rect 338304 642614 338404 642714
rect 338528 642614 338628 642714
rect 338752 642614 338852 642714
rect 338976 642614 339076 642714
rect 339200 642614 339300 642714
rect 339424 642614 339524 642714
rect 339648 642614 339748 642714
rect 339872 642614 339972 642714
rect 340096 642614 340196 642714
rect 340320 642614 340420 642714
rect 340544 642614 340644 642714
rect 340768 642614 340868 642714
rect 340992 642614 341092 642714
rect 341216 642614 341316 642714
rect 341440 642614 341540 642714
rect 341664 642614 341764 642714
rect 341888 642614 341988 642714
rect 342112 642614 342212 642714
rect 335616 642390 335716 642490
rect 335840 642390 335940 642490
rect 336064 642390 336164 642490
rect 336288 642390 336388 642490
rect 336512 642390 336612 642490
rect 336736 642390 336836 642490
rect 336960 642390 337060 642490
rect 337184 642390 337284 642490
rect 337408 642390 337508 642490
rect 337632 642390 337732 642490
rect 337856 642390 337956 642490
rect 338080 642390 338180 642490
rect 338304 642390 338404 642490
rect 338528 642390 338628 642490
rect 338752 642390 338852 642490
rect 338976 642390 339076 642490
rect 339200 642390 339300 642490
rect 339424 642390 339524 642490
rect 339648 642390 339748 642490
rect 339872 642390 339972 642490
rect 340096 642390 340196 642490
rect 340320 642390 340420 642490
rect 340544 642390 340644 642490
rect 340768 642390 340868 642490
rect 340992 642390 341092 642490
rect 341216 642390 341316 642490
rect 341440 642390 341540 642490
rect 341664 642390 341764 642490
rect 341888 642390 341988 642490
rect 342112 642390 342212 642490
rect 335616 642166 335716 642266
rect 335840 642166 335940 642266
rect 336064 642166 336164 642266
rect 336288 642166 336388 642266
rect 336512 642166 336612 642266
rect 336736 642166 336836 642266
rect 336960 642166 337060 642266
rect 337184 642166 337284 642266
rect 337408 642166 337508 642266
rect 337632 642166 337732 642266
rect 337856 642166 337956 642266
rect 338080 642166 338180 642266
rect 338304 642166 338404 642266
rect 338528 642166 338628 642266
rect 338752 642166 338852 642266
rect 338976 642166 339076 642266
rect 339200 642166 339300 642266
rect 339424 642166 339524 642266
rect 339648 642166 339748 642266
rect 339872 642166 339972 642266
rect 340096 642166 340196 642266
rect 340320 642166 340420 642266
rect 340544 642166 340644 642266
rect 340768 642166 340868 642266
rect 340992 642166 341092 642266
rect 341216 642166 341316 642266
rect 341440 642166 341540 642266
rect 341664 642166 341764 642266
rect 341888 642166 341988 642266
rect 342112 642166 342212 642266
rect 335616 641942 335716 642042
rect 335840 641942 335940 642042
rect 336064 641942 336164 642042
rect 336288 641942 336388 642042
rect 336512 641942 336612 642042
rect 336736 641942 336836 642042
rect 336960 641942 337060 642042
rect 337184 641942 337284 642042
rect 337408 641942 337508 642042
rect 337632 641942 337732 642042
rect 337856 641942 337956 642042
rect 338080 641942 338180 642042
rect 338304 641942 338404 642042
rect 338528 641942 338628 642042
rect 338752 641942 338852 642042
rect 338976 641942 339076 642042
rect 339200 641942 339300 642042
rect 339424 641942 339524 642042
rect 339648 641942 339748 642042
rect 339872 641942 339972 642042
rect 340096 641942 340196 642042
rect 340320 641942 340420 642042
rect 340544 641942 340644 642042
rect 340768 641942 340868 642042
rect 340992 641942 341092 642042
rect 341216 641942 341316 642042
rect 341440 641942 341540 642042
rect 341664 641942 341764 642042
rect 341888 641942 341988 642042
rect 342112 641942 342212 642042
rect 335616 641718 335716 641818
rect 335840 641718 335940 641818
rect 336064 641718 336164 641818
rect 336288 641718 336388 641818
rect 336512 641718 336612 641818
rect 336736 641718 336836 641818
rect 336960 641718 337060 641818
rect 337184 641718 337284 641818
rect 337408 641718 337508 641818
rect 337632 641718 337732 641818
rect 337856 641718 337956 641818
rect 338080 641718 338180 641818
rect 338304 641718 338404 641818
rect 338528 641718 338628 641818
rect 338752 641718 338852 641818
rect 338976 641718 339076 641818
rect 339200 641718 339300 641818
rect 339424 641718 339524 641818
rect 339648 641718 339748 641818
rect 339872 641718 339972 641818
rect 340096 641718 340196 641818
rect 340320 641718 340420 641818
rect 340544 641718 340644 641818
rect 340768 641718 340868 641818
rect 340992 641718 341092 641818
rect 341216 641718 341316 641818
rect 341440 641718 341540 641818
rect 341664 641718 341764 641818
rect 341888 641718 341988 641818
rect 342112 641718 342212 641818
rect 300652 640572 311908 640578
rect 300652 639746 300658 640572
rect 300658 639746 311902 640572
rect 311902 639746 311908 640572
rect 300652 639740 311908 639746
rect 297850 637896 297950 637996
rect 298074 637896 298174 637996
rect 298298 637896 298398 637996
rect 298522 637896 298622 637996
rect 298746 637896 298846 637996
rect 297850 637672 297950 637772
rect 298074 637672 298174 637772
rect 298298 637672 298398 637772
rect 298522 637672 298622 637772
rect 298746 637672 298846 637772
rect 297850 637448 297950 637548
rect 298074 637448 298174 637548
rect 298298 637448 298398 637548
rect 298522 637448 298622 637548
rect 298746 637448 298846 637548
rect 297850 637224 297950 637324
rect 298074 637224 298174 637324
rect 298298 637224 298398 637324
rect 298522 637224 298622 637324
rect 298746 637224 298846 637324
rect 297850 637000 297950 637100
rect 298074 637000 298174 637100
rect 298298 637000 298398 637100
rect 298522 637000 298622 637100
rect 298746 637000 298846 637100
rect 297850 636776 297950 636876
rect 298074 636776 298174 636876
rect 298298 636776 298398 636876
rect 298522 636776 298622 636876
rect 298746 636776 298846 636876
rect 297850 636552 297950 636652
rect 298074 636552 298174 636652
rect 298298 636552 298398 636652
rect 298522 636552 298622 636652
rect 298746 636552 298846 636652
rect 297850 636328 297950 636428
rect 298074 636328 298174 636428
rect 298298 636328 298398 636428
rect 298522 636328 298622 636428
rect 298746 636328 298846 636428
rect 297850 636104 297950 636204
rect 298074 636104 298174 636204
rect 298298 636104 298398 636204
rect 298522 636104 298622 636204
rect 298746 636104 298846 636204
rect 297850 635880 297950 635980
rect 298074 635880 298174 635980
rect 298298 635880 298398 635980
rect 298522 635880 298622 635980
rect 298746 635880 298846 635980
rect 297850 635656 297950 635756
rect 298074 635656 298174 635756
rect 298298 635656 298398 635756
rect 298522 635656 298622 635756
rect 298746 635656 298846 635756
rect 297850 635432 297950 635532
rect 298074 635432 298174 635532
rect 298298 635432 298398 635532
rect 298522 635432 298622 635532
rect 298746 635432 298846 635532
rect 297850 635208 297950 635308
rect 298074 635208 298174 635308
rect 298298 635208 298398 635308
rect 298522 635208 298622 635308
rect 298746 635208 298846 635308
rect 297850 634984 297950 635084
rect 298074 634984 298174 635084
rect 298298 634984 298398 635084
rect 298522 634984 298622 635084
rect 298746 634984 298846 635084
rect 297850 634760 297950 634860
rect 298074 634760 298174 634860
rect 298298 634760 298398 634860
rect 298522 634760 298622 634860
rect 298746 634760 298846 634860
rect 297850 634536 297950 634636
rect 298074 634536 298174 634636
rect 298298 634536 298398 634636
rect 298522 634536 298622 634636
rect 298746 634536 298846 634636
rect 297850 634312 297950 634412
rect 298074 634312 298174 634412
rect 298298 634312 298398 634412
rect 298522 634312 298622 634412
rect 298746 634312 298846 634412
rect 297850 634088 297950 634188
rect 298074 634088 298174 634188
rect 298298 634088 298398 634188
rect 298522 634088 298622 634188
rect 298746 634088 298846 634188
rect 342130 637896 342230 637996
rect 342354 637896 342454 637996
rect 342578 637896 342678 637996
rect 342802 637896 342902 637996
rect 343026 637896 343126 637996
rect 342130 637672 342230 637772
rect 342354 637672 342454 637772
rect 342578 637672 342678 637772
rect 342802 637672 342902 637772
rect 343026 637672 343126 637772
rect 342130 637448 342230 637548
rect 342354 637448 342454 637548
rect 342578 637448 342678 637548
rect 342802 637448 342902 637548
rect 343026 637448 343126 637548
rect 342130 637224 342230 637324
rect 342354 637224 342454 637324
rect 342578 637224 342678 637324
rect 342802 637224 342902 637324
rect 343026 637224 343126 637324
rect 342130 637000 342230 637100
rect 342354 637000 342454 637100
rect 342578 637000 342678 637100
rect 342802 637000 342902 637100
rect 343026 637000 343126 637100
rect 342130 636776 342230 636876
rect 342354 636776 342454 636876
rect 342578 636776 342678 636876
rect 342802 636776 342902 636876
rect 343026 636776 343126 636876
rect 342130 636552 342230 636652
rect 342354 636552 342454 636652
rect 342578 636552 342678 636652
rect 342802 636552 342902 636652
rect 343026 636552 343126 636652
rect 342130 636328 342230 636428
rect 342354 636328 342454 636428
rect 342578 636328 342678 636428
rect 342802 636328 342902 636428
rect 343026 636328 343126 636428
rect 342130 636104 342230 636204
rect 342354 636104 342454 636204
rect 342578 636104 342678 636204
rect 342802 636104 342902 636204
rect 343026 636104 343126 636204
rect 342130 635880 342230 635980
rect 342354 635880 342454 635980
rect 342578 635880 342678 635980
rect 342802 635880 342902 635980
rect 343026 635880 343126 635980
rect 342130 635656 342230 635756
rect 342354 635656 342454 635756
rect 342578 635656 342678 635756
rect 342802 635656 342902 635756
rect 343026 635656 343126 635756
rect 342130 635432 342230 635532
rect 342354 635432 342454 635532
rect 342578 635432 342678 635532
rect 342802 635432 342902 635532
rect 343026 635432 343126 635532
rect 342130 635208 342230 635308
rect 342354 635208 342454 635308
rect 342578 635208 342678 635308
rect 342802 635208 342902 635308
rect 343026 635208 343126 635308
rect 342130 634984 342230 635084
rect 342354 634984 342454 635084
rect 342578 634984 342678 635084
rect 342802 634984 342902 635084
rect 343026 634984 343126 635084
rect 342130 634760 342230 634860
rect 342354 634760 342454 634860
rect 342578 634760 342678 634860
rect 342802 634760 342902 634860
rect 343026 634760 343126 634860
rect 297850 633864 297950 633964
rect 298074 633864 298174 633964
rect 298298 633864 298398 633964
rect 298522 633864 298622 633964
rect 298746 633864 298846 633964
rect 297850 633640 297950 633740
rect 298074 633640 298174 633740
rect 298298 633640 298398 633740
rect 298522 633640 298622 633740
rect 298746 633640 298846 633740
rect 297850 633416 297950 633516
rect 298074 633416 298174 633516
rect 298298 633416 298398 633516
rect 298522 633416 298622 633516
rect 298746 633416 298846 633516
rect 297850 633192 297950 633292
rect 298074 633192 298174 633292
rect 298298 633192 298398 633292
rect 298522 633192 298622 633292
rect 298746 633192 298846 633292
rect 297850 632968 297950 633068
rect 298074 632968 298174 633068
rect 298298 632968 298398 633068
rect 298522 632968 298622 633068
rect 298746 632968 298846 633068
rect 297850 632744 297950 632844
rect 298074 632744 298174 632844
rect 298298 632744 298398 632844
rect 298522 632744 298622 632844
rect 298746 632744 298846 632844
rect 297850 632520 297950 632620
rect 298074 632520 298174 632620
rect 298298 632520 298398 632620
rect 298522 632520 298622 632620
rect 298746 632520 298846 632620
rect 297850 632296 297950 632396
rect 298074 632296 298174 632396
rect 298298 632296 298398 632396
rect 298522 632296 298622 632396
rect 298746 632296 298846 632396
rect 297850 632072 297950 632172
rect 298074 632072 298174 632172
rect 298298 632072 298398 632172
rect 298522 632072 298622 632172
rect 298746 632072 298846 632172
rect 297850 631848 297950 631948
rect 298074 631848 298174 631948
rect 298298 631848 298398 631948
rect 298522 631848 298622 631948
rect 298746 631848 298846 631948
rect 297850 631624 297950 631724
rect 298074 631624 298174 631724
rect 298298 631624 298398 631724
rect 298522 631624 298622 631724
rect 298746 631624 298846 631724
rect 297850 631400 297950 631500
rect 298074 631400 298174 631500
rect 298298 631400 298398 631500
rect 298522 631400 298622 631500
rect 298746 631400 298846 631500
rect 342130 634536 342230 634636
rect 342354 634536 342454 634636
rect 342578 634536 342678 634636
rect 342802 634536 342902 634636
rect 343026 634536 343126 634636
rect 342130 634312 342230 634412
rect 342354 634312 342454 634412
rect 342578 634312 342678 634412
rect 342802 634312 342902 634412
rect 343026 634312 343126 634412
rect 342130 634088 342230 634188
rect 342354 634088 342454 634188
rect 342578 634088 342678 634188
rect 342802 634088 342902 634188
rect 343026 634088 343126 634188
rect 342130 633864 342230 633964
rect 342354 633864 342454 633964
rect 342578 633864 342678 633964
rect 342802 633864 342902 633964
rect 343026 633864 343126 633964
rect 342130 633640 342230 633740
rect 342354 633640 342454 633740
rect 342578 633640 342678 633740
rect 342802 633640 342902 633740
rect 343026 633640 343126 633740
rect 342130 633416 342230 633516
rect 342354 633416 342454 633516
rect 342578 633416 342678 633516
rect 342802 633416 342902 633516
rect 343026 633416 343126 633516
rect 342130 633192 342230 633292
rect 342354 633192 342454 633292
rect 342578 633192 342678 633292
rect 342802 633192 342902 633292
rect 343026 633192 343126 633292
rect 342130 632968 342230 633068
rect 342354 632968 342454 633068
rect 342578 632968 342678 633068
rect 342802 632968 342902 633068
rect 343026 632968 343126 633068
rect 342130 632744 342230 632844
rect 342354 632744 342454 632844
rect 342578 632744 342678 632844
rect 342802 632744 342902 632844
rect 343026 632744 343126 632844
rect 342130 632520 342230 632620
rect 342354 632520 342454 632620
rect 342578 632520 342678 632620
rect 342802 632520 342902 632620
rect 343026 632520 343126 632620
rect 342130 632296 342230 632396
rect 342354 632296 342454 632396
rect 342578 632296 342678 632396
rect 342802 632296 342902 632396
rect 343026 632296 343126 632396
rect 342130 632072 342230 632172
rect 342354 632072 342454 632172
rect 342578 632072 342678 632172
rect 342802 632072 342902 632172
rect 343026 632072 343126 632172
rect 342130 631848 342230 631948
rect 342354 631848 342454 631948
rect 342578 631848 342678 631948
rect 342802 631848 342902 631948
rect 343026 631848 343126 631948
rect 342130 631624 342230 631724
rect 342354 631624 342454 631724
rect 342578 631624 342678 631724
rect 342802 631624 342902 631724
rect 343026 631624 343126 631724
rect 342130 631400 342230 631500
rect 342354 631400 342454 631500
rect 342578 631400 342678 631500
rect 342802 631400 342902 631500
rect 343026 631400 343126 631500
rect 319400 628668 319600 628868
rect 319834 628668 320034 628868
rect 320268 628668 320468 628868
rect 320702 628668 320902 628868
rect 321136 628668 321336 628868
rect 321570 628668 321770 628868
rect 322004 628668 322204 628868
rect 322438 628668 322638 628868
rect 322872 628668 323072 628868
rect 323306 628668 323506 628868
rect 323740 628668 323940 628868
rect 324140 628668 324340 628868
rect 324540 628668 324740 628868
rect 324940 628668 325140 628868
rect 325340 628668 325540 628868
rect 325740 628668 325940 628868
rect 326140 628668 326340 628868
rect 326540 628668 326740 628868
rect 326940 628668 327140 628868
rect 327340 628668 327540 628868
rect 319400 628234 319600 628434
rect 319834 628234 320034 628434
rect 320268 628234 320468 628434
rect 320702 628234 320902 628434
rect 321136 628234 321336 628434
rect 321570 628234 321770 628434
rect 322004 628234 322204 628434
rect 322438 628234 322638 628434
rect 322872 628234 323072 628434
rect 323306 628234 323506 628434
rect 323740 628234 323940 628434
rect 328940 628668 329140 628868
rect 329340 628668 329540 628868
rect 329740 628668 329940 628868
rect 330140 628668 330340 628868
rect 330540 628668 330740 628868
rect 330940 628668 331140 628868
rect 331340 628668 331540 628868
rect 331740 628668 331940 628868
rect 332140 628668 332340 628868
rect 319400 627800 319600 628000
rect 319834 627800 320034 628000
rect 320268 627800 320468 628000
rect 320702 627800 320902 628000
rect 321136 627800 321336 628000
rect 321570 627800 321770 628000
rect 322004 627800 322204 628000
rect 322438 627800 322638 628000
rect 322872 627800 323072 628000
rect 323306 627800 323506 628000
rect 323740 627800 323940 628000
rect 312952 626916 313820 627292
rect 313820 626916 315808 627292
rect 315808 626916 327520 627292
rect 327520 626916 329508 627292
rect 329508 626916 332832 627292
rect 332832 626916 333274 627292
rect 312952 626502 333274 626916
rect 312952 626308 313820 626502
rect 313820 626308 315808 626502
rect 315808 626308 327520 626502
rect 327520 626308 329508 626502
rect 329508 626308 333274 626502
rect 302980 625970 303040 626030
rect 303100 625970 303160 626030
rect 303220 625970 303280 626030
rect 303340 625970 303400 626030
rect 303460 625970 303520 626030
rect 302980 625850 303040 625910
rect 303100 625850 303160 625910
rect 303220 625850 303280 625910
rect 303340 625850 303400 625910
rect 303460 625850 303520 625910
rect 297850 624496 297950 624596
rect 298074 624496 298174 624596
rect 298298 624496 298398 624596
rect 298522 624496 298622 624596
rect 298746 624496 298846 624596
rect 297850 624272 297950 624372
rect 298074 624272 298174 624372
rect 298298 624272 298398 624372
rect 298522 624272 298622 624372
rect 298746 624272 298846 624372
rect 297850 624048 297950 624148
rect 298074 624048 298174 624148
rect 298298 624048 298398 624148
rect 298522 624048 298622 624148
rect 298746 624048 298846 624148
rect 342130 624496 342230 624596
rect 342354 624496 342454 624596
rect 342578 624496 342678 624596
rect 342802 624496 342902 624596
rect 343026 624496 343126 624596
rect 342130 624272 342230 624372
rect 342354 624272 342454 624372
rect 342578 624272 342678 624372
rect 342802 624272 342902 624372
rect 343026 624272 343126 624372
rect 342130 624048 342230 624148
rect 342354 624048 342454 624148
rect 342578 624048 342678 624148
rect 342802 624048 342902 624148
rect 343026 624048 343126 624148
rect 297850 623824 297950 623924
rect 298074 623824 298174 623924
rect 298298 623824 298398 623924
rect 298522 623824 298622 623924
rect 298746 623824 298846 623924
rect 297850 623600 297950 623700
rect 298074 623600 298174 623700
rect 298298 623600 298398 623700
rect 298522 623600 298622 623700
rect 298746 623600 298846 623700
rect 342130 623824 342230 623924
rect 342354 623824 342454 623924
rect 342578 623824 342678 623924
rect 342802 623824 342902 623924
rect 343026 623824 343126 623924
rect 342130 623600 342230 623700
rect 342354 623600 342454 623700
rect 342578 623600 342678 623700
rect 342802 623600 342902 623700
rect 343026 623600 343126 623700
rect 297850 623376 297950 623476
rect 298074 623376 298174 623476
rect 298298 623376 298398 623476
rect 298522 623376 298622 623476
rect 298746 623376 298846 623476
rect 297850 623152 297950 623252
rect 298074 623152 298174 623252
rect 298298 623152 298398 623252
rect 298522 623152 298622 623252
rect 298746 623152 298846 623252
rect 297850 622928 297950 623028
rect 298074 622928 298174 623028
rect 298298 622928 298398 623028
rect 298522 622928 298622 623028
rect 298746 622928 298846 623028
rect 342130 623376 342230 623476
rect 342354 623376 342454 623476
rect 342578 623376 342678 623476
rect 342802 623376 342902 623476
rect 343026 623376 343126 623476
rect 342130 623152 342230 623252
rect 342354 623152 342454 623252
rect 342578 623152 342678 623252
rect 342802 623152 342902 623252
rect 343026 623152 343126 623252
rect 342130 622928 342230 623028
rect 342354 622928 342454 623028
rect 342578 622928 342678 623028
rect 342802 622928 342902 623028
rect 343026 622928 343126 623028
rect 297850 622704 297950 622804
rect 298074 622704 298174 622804
rect 298298 622704 298398 622804
rect 298522 622704 298622 622804
rect 298746 622704 298846 622804
rect 297850 622480 297950 622580
rect 298074 622480 298174 622580
rect 298298 622480 298398 622580
rect 298522 622480 298622 622580
rect 298746 622480 298846 622580
rect 342130 622704 342230 622804
rect 342354 622704 342454 622804
rect 342578 622704 342678 622804
rect 342802 622704 342902 622804
rect 343026 622704 343126 622804
rect 342130 622480 342230 622580
rect 342354 622480 342454 622580
rect 342578 622480 342678 622580
rect 342802 622480 342902 622580
rect 343026 622480 343126 622580
rect 297850 622256 297950 622356
rect 298074 622256 298174 622356
rect 298298 622256 298398 622356
rect 298522 622256 298622 622356
rect 298746 622256 298846 622356
rect 297850 622032 297950 622132
rect 298074 622032 298174 622132
rect 298298 622032 298398 622132
rect 298522 622032 298622 622132
rect 298746 622032 298846 622132
rect 297850 621808 297950 621908
rect 298074 621808 298174 621908
rect 298298 621808 298398 621908
rect 298522 621808 298622 621908
rect 298746 621808 298846 621908
rect 297850 621584 297950 621684
rect 298074 621584 298174 621684
rect 298298 621584 298398 621684
rect 298522 621584 298622 621684
rect 298746 621584 298846 621684
rect 297850 621360 297950 621460
rect 298074 621360 298174 621460
rect 298298 621360 298398 621460
rect 298522 621360 298622 621460
rect 298746 621360 298846 621460
rect 297850 621136 297950 621236
rect 298074 621136 298174 621236
rect 298298 621136 298398 621236
rect 298522 621136 298622 621236
rect 298746 621136 298846 621236
rect 297850 620912 297950 621012
rect 298074 620912 298174 621012
rect 298298 620912 298398 621012
rect 298522 620912 298622 621012
rect 298746 620912 298846 621012
rect 297850 620688 297950 620788
rect 298074 620688 298174 620788
rect 298298 620688 298398 620788
rect 298522 620688 298622 620788
rect 298746 620688 298846 620788
rect 297850 620464 297950 620564
rect 298074 620464 298174 620564
rect 298298 620464 298398 620564
rect 298522 620464 298622 620564
rect 298746 620464 298846 620564
rect 342130 622256 342230 622356
rect 342354 622256 342454 622356
rect 342578 622256 342678 622356
rect 342802 622256 342902 622356
rect 343026 622256 343126 622356
rect 342130 622032 342230 622132
rect 342354 622032 342454 622132
rect 342578 622032 342678 622132
rect 342802 622032 342902 622132
rect 343026 622032 343126 622132
rect 342130 621808 342230 621908
rect 342354 621808 342454 621908
rect 342578 621808 342678 621908
rect 342802 621808 342902 621908
rect 343026 621808 343126 621908
rect 342130 621584 342230 621684
rect 342354 621584 342454 621684
rect 342578 621584 342678 621684
rect 342802 621584 342902 621684
rect 343026 621584 343126 621684
rect 342130 621360 342230 621460
rect 342354 621360 342454 621460
rect 342578 621360 342678 621460
rect 342802 621360 342902 621460
rect 343026 621360 343126 621460
rect 342130 621136 342230 621236
rect 342354 621136 342454 621236
rect 342578 621136 342678 621236
rect 342802 621136 342902 621236
rect 343026 621136 343126 621236
rect 342130 620912 342230 621012
rect 342354 620912 342454 621012
rect 342578 620912 342678 621012
rect 342802 620912 342902 621012
rect 343026 620912 343126 621012
rect 342130 620688 342230 620788
rect 342354 620688 342454 620788
rect 342578 620688 342678 620788
rect 342802 620688 342902 620788
rect 343026 620688 343126 620788
rect 342130 620464 342230 620564
rect 342354 620464 342454 620564
rect 342578 620464 342678 620564
rect 342802 620464 342902 620564
rect 343026 620464 343126 620564
rect 297850 620240 297950 620340
rect 298074 620240 298174 620340
rect 298298 620240 298398 620340
rect 298522 620240 298622 620340
rect 298746 620240 298846 620340
rect 342130 620240 342230 620340
rect 342354 620240 342454 620340
rect 342578 620240 342678 620340
rect 342802 620240 342902 620340
rect 343026 620240 343126 620340
rect 297850 620016 297950 620116
rect 298074 620016 298174 620116
rect 298298 620016 298398 620116
rect 298522 620016 298622 620116
rect 298746 620016 298846 620116
rect 297850 619792 297950 619892
rect 298074 619792 298174 619892
rect 298298 619792 298398 619892
rect 298522 619792 298622 619892
rect 298746 619792 298846 619892
rect 303604 619883 304204 620135
rect 312095 619883 312695 620135
rect 342130 620016 342230 620116
rect 342354 620016 342454 620116
rect 342578 620016 342678 620116
rect 342802 620016 342902 620116
rect 343026 620016 343126 620116
rect 342130 619792 342230 619892
rect 342354 619792 342454 619892
rect 342578 619792 342678 619892
rect 342802 619792 342902 619892
rect 343026 619792 343126 619892
rect 297850 619568 297950 619668
rect 298074 619568 298174 619668
rect 298298 619568 298398 619668
rect 298522 619568 298622 619668
rect 298746 619568 298846 619668
rect 297850 619344 297950 619444
rect 298074 619344 298174 619444
rect 298298 619344 298398 619444
rect 298522 619344 298622 619444
rect 298746 619344 298846 619444
rect 297850 619120 297950 619220
rect 298074 619120 298174 619220
rect 298298 619120 298398 619220
rect 298522 619120 298622 619220
rect 298746 619120 298846 619220
rect 297850 618896 297950 618996
rect 298074 618896 298174 618996
rect 298298 618896 298398 618996
rect 298522 618896 298622 618996
rect 298746 618896 298846 618996
rect 297850 618672 297950 618772
rect 298074 618672 298174 618772
rect 298298 618672 298398 618772
rect 298522 618672 298622 618772
rect 298746 618672 298846 618772
rect 342130 619568 342230 619668
rect 342354 619568 342454 619668
rect 342578 619568 342678 619668
rect 342802 619568 342902 619668
rect 343026 619568 343126 619668
rect 342130 619344 342230 619444
rect 342354 619344 342454 619444
rect 342578 619344 342678 619444
rect 342802 619344 342902 619444
rect 343026 619344 343126 619444
rect 342130 619120 342230 619220
rect 342354 619120 342454 619220
rect 342578 619120 342678 619220
rect 342802 619120 342902 619220
rect 343026 619120 343126 619220
rect 342130 618896 342230 618996
rect 342354 618896 342454 618996
rect 342578 618896 342678 618996
rect 342802 618896 342902 618996
rect 343026 618896 343126 618996
rect 297850 618448 297950 618548
rect 298074 618448 298174 618548
rect 298298 618448 298398 618548
rect 298522 618448 298622 618548
rect 298746 618448 298846 618548
rect 297850 618224 297950 618324
rect 298074 618224 298174 618324
rect 298298 618224 298398 618324
rect 298522 618224 298622 618324
rect 298746 618224 298846 618324
rect 297850 618000 297950 618100
rect 298074 618000 298174 618100
rect 298298 618000 298398 618100
rect 298522 618000 298622 618100
rect 298746 618000 298846 618100
rect 342130 618672 342230 618772
rect 342354 618672 342454 618772
rect 342578 618672 342678 618772
rect 342802 618672 342902 618772
rect 343026 618672 343126 618772
rect 342130 618448 342230 618548
rect 342354 618448 342454 618548
rect 342578 618448 342678 618548
rect 342802 618448 342902 618548
rect 343026 618448 343126 618548
rect 342130 618224 342230 618324
rect 342354 618224 342454 618324
rect 342578 618224 342678 618324
rect 342802 618224 342902 618324
rect 343026 618224 343126 618324
rect 342130 618000 342230 618100
rect 342354 618000 342454 618100
rect 342578 618000 342678 618100
rect 342802 618000 342902 618100
rect 343026 618000 343126 618100
rect 302946 617058 312192 617062
rect 302946 616954 302964 617058
rect 302964 616954 303016 617058
rect 303016 616954 303586 617058
rect 303586 616954 303638 617058
rect 303638 616954 304044 617058
rect 304044 616954 304096 617058
rect 304096 616954 304620 617058
rect 304620 616954 304672 617058
rect 304672 616954 305192 617058
rect 305192 616954 305244 617058
rect 305244 616954 305764 617058
rect 305764 616954 305816 617058
rect 305816 616954 306336 617058
rect 306336 616954 306388 617058
rect 306388 616954 306908 617058
rect 306908 616954 306960 617058
rect 306960 616954 307480 617058
rect 307480 616954 307532 617058
rect 307532 616954 308052 617058
rect 308052 616954 308104 617058
rect 308104 616954 308624 617058
rect 308624 616954 308676 617058
rect 308676 616954 309196 617058
rect 309196 616954 309248 617058
rect 309248 616954 309768 617058
rect 309768 616954 309820 617058
rect 309820 616954 310340 617058
rect 310340 616954 310392 617058
rect 310392 616954 310912 617058
rect 310912 616954 310964 617058
rect 310964 616954 311022 617058
rect 311022 616954 311074 617058
rect 311074 616954 311480 617058
rect 311480 616954 311532 617058
rect 311532 616954 312092 617058
rect 312092 616954 312144 617058
rect 312144 616954 312192 617058
rect 302946 616948 312192 616954
rect 312710 616828 330648 616830
rect 312710 616748 314294 616828
rect 314294 616748 314374 616828
rect 314374 616748 315214 616828
rect 315214 616748 315294 616828
rect 315294 616748 316134 616828
rect 316134 616748 316214 616828
rect 316214 616748 317054 616828
rect 317054 616748 317134 616828
rect 317134 616748 317974 616828
rect 317974 616748 318054 616828
rect 318054 616748 319794 616828
rect 319794 616748 319874 616828
rect 319874 616748 320714 616828
rect 320714 616748 320794 616828
rect 320794 616748 321634 616828
rect 321634 616748 321714 616828
rect 321714 616748 322554 616828
rect 322554 616748 322634 616828
rect 322634 616748 323474 616828
rect 323474 616748 323554 616828
rect 323554 616748 325294 616828
rect 325294 616748 325374 616828
rect 325374 616748 326214 616828
rect 326214 616748 326294 616828
rect 326294 616748 327134 616828
rect 327134 616748 327214 616828
rect 327214 616748 328054 616828
rect 328054 616748 328134 616828
rect 328134 616748 328974 616828
rect 328974 616748 329054 616828
rect 329054 616748 330648 616828
rect 312710 616708 330648 616748
rect 312710 616608 312804 616708
rect 312804 616608 313204 616708
rect 313204 616608 318714 616708
rect 318714 616608 319114 616708
rect 319114 616608 324214 616708
rect 324214 616608 324614 616708
rect 324614 616706 330648 616708
rect 324614 616608 330170 616706
rect 312710 616606 330170 616608
rect 330170 616606 330570 616706
rect 330570 616606 330648 616706
rect 312710 616512 330648 616606
rect 298876 615374 298976 615474
rect 299100 615374 299200 615474
rect 299324 615374 299424 615474
rect 299548 615374 299648 615474
rect 299772 615374 299872 615474
rect 299996 615374 300096 615474
rect 300220 615374 300320 615474
rect 300444 615374 300544 615474
rect 300668 615374 300768 615474
rect 300892 615374 300992 615474
rect 301116 615374 301216 615474
rect 301340 615374 301440 615474
rect 301564 615374 301664 615474
rect 301788 615374 301888 615474
rect 302012 615374 302112 615474
rect 302236 615374 302336 615474
rect 302460 615374 302560 615474
rect 302684 615374 302784 615474
rect 302908 615374 303008 615474
rect 303132 615374 303232 615474
rect 303356 615374 303456 615474
rect 303580 615374 303680 615474
rect 303804 615374 303904 615474
rect 304028 615374 304128 615474
rect 304252 615374 304352 615474
rect 304476 615374 304576 615474
rect 304700 615374 304800 615474
rect 304924 615374 305024 615474
rect 305148 615374 305248 615474
rect 305372 615374 305472 615474
rect 298876 615150 298976 615250
rect 299100 615150 299200 615250
rect 299324 615150 299424 615250
rect 299548 615150 299648 615250
rect 299772 615150 299872 615250
rect 299996 615150 300096 615250
rect 300220 615150 300320 615250
rect 300444 615150 300544 615250
rect 300668 615150 300768 615250
rect 300892 615150 300992 615250
rect 301116 615150 301216 615250
rect 301340 615150 301440 615250
rect 301564 615150 301664 615250
rect 301788 615150 301888 615250
rect 302012 615150 302112 615250
rect 302236 615150 302336 615250
rect 302460 615150 302560 615250
rect 302684 615150 302784 615250
rect 302908 615150 303008 615250
rect 303132 615150 303232 615250
rect 303356 615150 303456 615250
rect 303580 615150 303680 615250
rect 303804 615150 303904 615250
rect 304028 615150 304128 615250
rect 304252 615150 304352 615250
rect 304476 615150 304576 615250
rect 304700 615150 304800 615250
rect 304924 615150 305024 615250
rect 305148 615150 305248 615250
rect 305372 615150 305472 615250
rect 298876 614926 298976 615026
rect 299100 614926 299200 615026
rect 299324 614926 299424 615026
rect 299548 614926 299648 615026
rect 299772 614926 299872 615026
rect 299996 614926 300096 615026
rect 300220 614926 300320 615026
rect 300444 614926 300544 615026
rect 300668 614926 300768 615026
rect 300892 614926 300992 615026
rect 301116 614926 301216 615026
rect 301340 614926 301440 615026
rect 301564 614926 301664 615026
rect 301788 614926 301888 615026
rect 302012 614926 302112 615026
rect 302236 614926 302336 615026
rect 302460 614926 302560 615026
rect 302684 614926 302784 615026
rect 302908 614926 303008 615026
rect 303132 614926 303232 615026
rect 303356 614926 303456 615026
rect 303580 614926 303680 615026
rect 303804 614926 303904 615026
rect 304028 614926 304128 615026
rect 304252 614926 304352 615026
rect 304476 614926 304576 615026
rect 304700 614926 304800 615026
rect 304924 614926 305024 615026
rect 305148 614926 305248 615026
rect 305372 614926 305472 615026
rect 298876 614702 298976 614802
rect 299100 614702 299200 614802
rect 299324 614702 299424 614802
rect 299548 614702 299648 614802
rect 299772 614702 299872 614802
rect 299996 614702 300096 614802
rect 300220 614702 300320 614802
rect 300444 614702 300544 614802
rect 300668 614702 300768 614802
rect 300892 614702 300992 614802
rect 301116 614702 301216 614802
rect 301340 614702 301440 614802
rect 301564 614702 301664 614802
rect 301788 614702 301888 614802
rect 302012 614702 302112 614802
rect 302236 614702 302336 614802
rect 302460 614702 302560 614802
rect 302684 614702 302784 614802
rect 302908 614702 303008 614802
rect 303132 614702 303232 614802
rect 303356 614702 303456 614802
rect 303580 614702 303680 614802
rect 303804 614702 303904 614802
rect 304028 614702 304128 614802
rect 304252 614702 304352 614802
rect 304476 614702 304576 614802
rect 304700 614702 304800 614802
rect 304924 614702 305024 614802
rect 305148 614702 305248 614802
rect 305372 614702 305472 614802
rect 298876 614478 298976 614578
rect 299100 614478 299200 614578
rect 299324 614478 299424 614578
rect 299548 614478 299648 614578
rect 299772 614478 299872 614578
rect 299996 614478 300096 614578
rect 300220 614478 300320 614578
rect 300444 614478 300544 614578
rect 300668 614478 300768 614578
rect 300892 614478 300992 614578
rect 301116 614478 301216 614578
rect 301340 614478 301440 614578
rect 301564 614478 301664 614578
rect 301788 614478 301888 614578
rect 302012 614478 302112 614578
rect 302236 614478 302336 614578
rect 302460 614478 302560 614578
rect 302684 614478 302784 614578
rect 302908 614478 303008 614578
rect 303132 614478 303232 614578
rect 303356 614478 303456 614578
rect 303580 614478 303680 614578
rect 303804 614478 303904 614578
rect 304028 614478 304128 614578
rect 304252 614478 304352 614578
rect 304476 614478 304576 614578
rect 304700 614478 304800 614578
rect 304924 614478 305024 614578
rect 305148 614478 305248 614578
rect 305372 614478 305472 614578
rect 309346 615374 309446 615474
rect 309570 615374 309670 615474
rect 309794 615374 309894 615474
rect 310018 615374 310118 615474
rect 310242 615374 310342 615474
rect 310466 615374 310566 615474
rect 310690 615374 310790 615474
rect 310914 615374 311014 615474
rect 311138 615374 311238 615474
rect 311362 615374 311462 615474
rect 311586 615374 311686 615474
rect 311810 615374 311910 615474
rect 312034 615374 312134 615474
rect 312258 615374 312358 615474
rect 312482 615374 312582 615474
rect 312706 615374 312806 615474
rect 312930 615374 313030 615474
rect 313154 615374 313254 615474
rect 313378 615374 313478 615474
rect 313602 615374 313702 615474
rect 313826 615374 313926 615474
rect 314050 615374 314150 615474
rect 314274 615374 314374 615474
rect 314498 615374 314598 615474
rect 314722 615374 314822 615474
rect 314946 615374 315046 615474
rect 315170 615374 315270 615474
rect 315394 615374 315494 615474
rect 315618 615374 315718 615474
rect 315842 615374 315942 615474
rect 309346 615150 309446 615250
rect 309570 615150 309670 615250
rect 309794 615150 309894 615250
rect 310018 615150 310118 615250
rect 310242 615150 310342 615250
rect 310466 615150 310566 615250
rect 310690 615150 310790 615250
rect 310914 615150 311014 615250
rect 311138 615150 311238 615250
rect 311362 615150 311462 615250
rect 311586 615150 311686 615250
rect 311810 615150 311910 615250
rect 312034 615150 312134 615250
rect 312258 615150 312358 615250
rect 312482 615150 312582 615250
rect 312706 615150 312806 615250
rect 312930 615150 313030 615250
rect 313154 615150 313254 615250
rect 313378 615150 313478 615250
rect 313602 615150 313702 615250
rect 313826 615150 313926 615250
rect 314050 615150 314150 615250
rect 314274 615150 314374 615250
rect 314498 615150 314598 615250
rect 314722 615150 314822 615250
rect 314946 615150 315046 615250
rect 315170 615150 315270 615250
rect 315394 615150 315494 615250
rect 315618 615150 315718 615250
rect 315842 615150 315942 615250
rect 309346 614926 309446 615026
rect 309570 614926 309670 615026
rect 309794 614926 309894 615026
rect 310018 614926 310118 615026
rect 310242 614926 310342 615026
rect 310466 614926 310566 615026
rect 310690 614926 310790 615026
rect 310914 614926 311014 615026
rect 311138 614926 311238 615026
rect 311362 614926 311462 615026
rect 311586 614926 311686 615026
rect 311810 614926 311910 615026
rect 312034 614926 312134 615026
rect 312258 614926 312358 615026
rect 312482 614926 312582 615026
rect 312706 614926 312806 615026
rect 312930 614926 313030 615026
rect 313154 614926 313254 615026
rect 313378 614926 313478 615026
rect 313602 614926 313702 615026
rect 313826 614926 313926 615026
rect 314050 614926 314150 615026
rect 314274 614926 314374 615026
rect 314498 614926 314598 615026
rect 314722 614926 314822 615026
rect 314946 614926 315046 615026
rect 315170 614926 315270 615026
rect 315394 614926 315494 615026
rect 315618 614926 315718 615026
rect 315842 614926 315942 615026
rect 309346 614702 309446 614802
rect 309570 614702 309670 614802
rect 309794 614702 309894 614802
rect 310018 614702 310118 614802
rect 310242 614702 310342 614802
rect 310466 614702 310566 614802
rect 310690 614702 310790 614802
rect 310914 614702 311014 614802
rect 311138 614702 311238 614802
rect 311362 614702 311462 614802
rect 311586 614702 311686 614802
rect 311810 614702 311910 614802
rect 312034 614702 312134 614802
rect 312258 614702 312358 614802
rect 312482 614702 312582 614802
rect 312706 614702 312806 614802
rect 312930 614702 313030 614802
rect 313154 614702 313254 614802
rect 313378 614702 313478 614802
rect 313602 614702 313702 614802
rect 313826 614702 313926 614802
rect 314050 614702 314150 614802
rect 314274 614702 314374 614802
rect 314498 614702 314598 614802
rect 314722 614702 314822 614802
rect 314946 614702 315046 614802
rect 315170 614702 315270 614802
rect 315394 614702 315494 614802
rect 315618 614702 315718 614802
rect 315842 614702 315942 614802
rect 309346 614478 309446 614578
rect 309570 614478 309670 614578
rect 309794 614478 309894 614578
rect 310018 614478 310118 614578
rect 310242 614478 310342 614578
rect 310466 614478 310566 614578
rect 310690 614478 310790 614578
rect 310914 614478 311014 614578
rect 311138 614478 311238 614578
rect 311362 614478 311462 614578
rect 311586 614478 311686 614578
rect 311810 614478 311910 614578
rect 312034 614478 312134 614578
rect 312258 614478 312358 614578
rect 312482 614478 312582 614578
rect 312706 614478 312806 614578
rect 312930 614478 313030 614578
rect 313154 614478 313254 614578
rect 313378 614478 313478 614578
rect 313602 614478 313702 614578
rect 313826 614478 313926 614578
rect 314050 614478 314150 614578
rect 314274 614478 314374 614578
rect 314498 614478 314598 614578
rect 314722 614478 314822 614578
rect 314946 614478 315046 614578
rect 315170 614478 315270 614578
rect 315394 614478 315494 614578
rect 315618 614478 315718 614578
rect 315842 614478 315942 614578
rect 335616 615394 335716 615494
rect 335840 615394 335940 615494
rect 336064 615394 336164 615494
rect 336288 615394 336388 615494
rect 336512 615394 336612 615494
rect 336736 615394 336836 615494
rect 336960 615394 337060 615494
rect 337184 615394 337284 615494
rect 337408 615394 337508 615494
rect 337632 615394 337732 615494
rect 337856 615394 337956 615494
rect 338080 615394 338180 615494
rect 338304 615394 338404 615494
rect 338528 615394 338628 615494
rect 338752 615394 338852 615494
rect 338976 615394 339076 615494
rect 339200 615394 339300 615494
rect 339424 615394 339524 615494
rect 339648 615394 339748 615494
rect 339872 615394 339972 615494
rect 340096 615394 340196 615494
rect 340320 615394 340420 615494
rect 340544 615394 340644 615494
rect 340768 615394 340868 615494
rect 340992 615394 341092 615494
rect 341216 615394 341316 615494
rect 341440 615394 341540 615494
rect 341664 615394 341764 615494
rect 341888 615394 341988 615494
rect 342112 615394 342212 615494
rect 335616 615170 335716 615270
rect 335840 615170 335940 615270
rect 336064 615170 336164 615270
rect 336288 615170 336388 615270
rect 336512 615170 336612 615270
rect 336736 615170 336836 615270
rect 336960 615170 337060 615270
rect 337184 615170 337284 615270
rect 337408 615170 337508 615270
rect 337632 615170 337732 615270
rect 337856 615170 337956 615270
rect 338080 615170 338180 615270
rect 338304 615170 338404 615270
rect 338528 615170 338628 615270
rect 338752 615170 338852 615270
rect 338976 615170 339076 615270
rect 339200 615170 339300 615270
rect 339424 615170 339524 615270
rect 339648 615170 339748 615270
rect 339872 615170 339972 615270
rect 340096 615170 340196 615270
rect 340320 615170 340420 615270
rect 340544 615170 340644 615270
rect 340768 615170 340868 615270
rect 340992 615170 341092 615270
rect 341216 615170 341316 615270
rect 341440 615170 341540 615270
rect 341664 615170 341764 615270
rect 341888 615170 341988 615270
rect 342112 615170 342212 615270
rect 335616 614946 335716 615046
rect 335840 614946 335940 615046
rect 336064 614946 336164 615046
rect 336288 614946 336388 615046
rect 336512 614946 336612 615046
rect 336736 614946 336836 615046
rect 336960 614946 337060 615046
rect 337184 614946 337284 615046
rect 337408 614946 337508 615046
rect 337632 614946 337732 615046
rect 337856 614946 337956 615046
rect 338080 614946 338180 615046
rect 338304 614946 338404 615046
rect 338528 614946 338628 615046
rect 338752 614946 338852 615046
rect 338976 614946 339076 615046
rect 339200 614946 339300 615046
rect 339424 614946 339524 615046
rect 339648 614946 339748 615046
rect 339872 614946 339972 615046
rect 340096 614946 340196 615046
rect 340320 614946 340420 615046
rect 340544 614946 340644 615046
rect 340768 614946 340868 615046
rect 340992 614946 341092 615046
rect 341216 614946 341316 615046
rect 341440 614946 341540 615046
rect 341664 614946 341764 615046
rect 341888 614946 341988 615046
rect 342112 614946 342212 615046
rect 335616 614722 335716 614822
rect 335840 614722 335940 614822
rect 336064 614722 336164 614822
rect 336288 614722 336388 614822
rect 336512 614722 336612 614822
rect 336736 614722 336836 614822
rect 336960 614722 337060 614822
rect 337184 614722 337284 614822
rect 337408 614722 337508 614822
rect 337632 614722 337732 614822
rect 337856 614722 337956 614822
rect 338080 614722 338180 614822
rect 338304 614722 338404 614822
rect 338528 614722 338628 614822
rect 338752 614722 338852 614822
rect 338976 614722 339076 614822
rect 339200 614722 339300 614822
rect 339424 614722 339524 614822
rect 339648 614722 339748 614822
rect 339872 614722 339972 614822
rect 340096 614722 340196 614822
rect 340320 614722 340420 614822
rect 340544 614722 340644 614822
rect 340768 614722 340868 614822
rect 340992 614722 341092 614822
rect 341216 614722 341316 614822
rect 341440 614722 341540 614822
rect 341664 614722 341764 614822
rect 341888 614722 341988 614822
rect 342112 614722 342212 614822
rect 335616 614498 335716 614598
rect 335840 614498 335940 614598
rect 336064 614498 336164 614598
rect 336288 614498 336388 614598
rect 336512 614498 336612 614598
rect 336736 614498 336836 614598
rect 336960 614498 337060 614598
rect 337184 614498 337284 614598
rect 337408 614498 337508 614598
rect 337632 614498 337732 614598
rect 337856 614498 337956 614598
rect 338080 614498 338180 614598
rect 338304 614498 338404 614598
rect 338528 614498 338628 614598
rect 338752 614498 338852 614598
rect 338976 614498 339076 614598
rect 339200 614498 339300 614598
rect 339424 614498 339524 614598
rect 339648 614498 339748 614598
rect 339872 614498 339972 614598
rect 340096 614498 340196 614598
rect 340320 614498 340420 614598
rect 340544 614498 340644 614598
rect 340768 614498 340868 614598
rect 340992 614498 341092 614598
rect 341216 614498 341316 614598
rect 341440 614498 341540 614598
rect 341664 614498 341764 614598
rect 341888 614498 341988 614598
rect 342112 614498 342212 614598
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 690577 173094 704800
rect -800 680242 1700 685242
rect 170894 684353 170922 690577
rect 173066 684353 173094 690577
rect 170894 683764 173094 684353
rect 173394 690577 175594 704800
rect 175894 702300 180894 704800
rect 173394 684353 173422 690577
rect 175566 684353 175594 690577
rect 173394 683764 175594 684353
rect -800 643842 1660 648642
rect -800 633842 1660 638642
rect 217294 626176 222294 704800
rect 222594 690610 224794 704800
rect 222594 684386 222622 690610
rect 224766 684386 224794 690610
rect 222594 683913 224794 684386
rect 225094 694292 227294 704800
rect 227594 694292 232594 704800
rect 225094 692092 232594 694292
rect 225094 683913 227294 692092
rect 217294 626112 217344 626176
rect 217408 626112 217472 626176
rect 217536 626112 217600 626176
rect 217664 626112 217728 626176
rect 217792 626112 217856 626176
rect 217920 626112 217984 626176
rect 218048 626112 218112 626176
rect 218176 626112 218240 626176
rect 218304 626112 218368 626176
rect 218432 626112 218496 626176
rect 218560 626112 218624 626176
rect 218688 626112 218752 626176
rect 218816 626112 218880 626176
rect 218944 626112 219008 626176
rect 219072 626112 219136 626176
rect 219200 626112 219264 626176
rect 219328 626112 219392 626176
rect 219456 626112 219520 626176
rect 219584 626112 219648 626176
rect 219712 626112 219776 626176
rect 219840 626112 219904 626176
rect 219968 626112 220032 626176
rect 220096 626112 220160 626176
rect 220224 626112 220288 626176
rect 220352 626112 220416 626176
rect 220480 626112 220544 626176
rect 220608 626112 220672 626176
rect 220736 626112 220800 626176
rect 220864 626112 220928 626176
rect 220992 626112 221056 626176
rect 221120 626112 221184 626176
rect 221248 626112 221312 626176
rect 221376 626112 221440 626176
rect 221504 626112 221568 626176
rect 221632 626112 221696 626176
rect 221760 626112 221824 626176
rect 221888 626112 221952 626176
rect 222016 626112 222080 626176
rect 222144 626112 222294 626176
rect 217294 626048 222294 626112
rect 217294 625984 217344 626048
rect 217408 625984 217472 626048
rect 217536 625984 217600 626048
rect 217664 625984 217728 626048
rect 217792 625984 217856 626048
rect 217920 625984 217984 626048
rect 218048 625984 218112 626048
rect 218176 625984 218240 626048
rect 218304 625984 218368 626048
rect 218432 625984 218496 626048
rect 218560 625984 218624 626048
rect 218688 625984 218752 626048
rect 218816 625984 218880 626048
rect 218944 625984 219008 626048
rect 219072 625984 219136 626048
rect 219200 625984 219264 626048
rect 219328 625984 219392 626048
rect 219456 625984 219520 626048
rect 219584 625984 219648 626048
rect 219712 625984 219776 626048
rect 219840 625984 219904 626048
rect 219968 625984 220032 626048
rect 220096 625984 220160 626048
rect 220224 625984 220288 626048
rect 220352 625984 220416 626048
rect 220480 625984 220544 626048
rect 220608 625984 220672 626048
rect 220736 625984 220800 626048
rect 220864 625984 220928 626048
rect 220992 625984 221056 626048
rect 221120 625984 221184 626048
rect 221248 625984 221312 626048
rect 221376 625984 221440 626048
rect 221504 625984 221568 626048
rect 221632 625984 221696 626048
rect 221760 625984 221824 626048
rect 221888 625984 221952 626048
rect 222016 625984 222080 626048
rect 222144 625984 222294 626048
rect 217294 625920 222294 625984
rect 217294 625856 217344 625920
rect 217408 625856 217472 625920
rect 217536 625856 217600 625920
rect 217664 625856 217728 625920
rect 217792 625856 217856 625920
rect 217920 625856 217984 625920
rect 218048 625856 218112 625920
rect 218176 625856 218240 625920
rect 218304 625856 218368 625920
rect 218432 625856 218496 625920
rect 218560 625856 218624 625920
rect 218688 625856 218752 625920
rect 218816 625856 218880 625920
rect 218944 625856 219008 625920
rect 219072 625856 219136 625920
rect 219200 625856 219264 625920
rect 219328 625856 219392 625920
rect 219456 625856 219520 625920
rect 219584 625856 219648 625920
rect 219712 625856 219776 625920
rect 219840 625856 219904 625920
rect 219968 625856 220032 625920
rect 220096 625856 220160 625920
rect 220224 625856 220288 625920
rect 220352 625856 220416 625920
rect 220480 625856 220544 625920
rect 220608 625856 220672 625920
rect 220736 625856 220800 625920
rect 220864 625856 220928 625920
rect 220992 625856 221056 625920
rect 221120 625856 221184 625920
rect 221248 625856 221312 625920
rect 221376 625856 221440 625920
rect 221504 625856 221568 625920
rect 221632 625856 221696 625920
rect 221760 625856 221824 625920
rect 221888 625856 221952 625920
rect 222016 625856 222080 625920
rect 222144 625856 222294 625920
rect 217294 625792 222294 625856
rect 217294 625728 217344 625792
rect 217408 625728 217472 625792
rect 217536 625728 217600 625792
rect 217664 625728 217728 625792
rect 217792 625728 217856 625792
rect 217920 625728 217984 625792
rect 218048 625728 218112 625792
rect 218176 625728 218240 625792
rect 218304 625728 218368 625792
rect 218432 625728 218496 625792
rect 218560 625728 218624 625792
rect 218688 625728 218752 625792
rect 218816 625728 218880 625792
rect 218944 625728 219008 625792
rect 219072 625728 219136 625792
rect 219200 625728 219264 625792
rect 219328 625728 219392 625792
rect 219456 625728 219520 625792
rect 219584 625728 219648 625792
rect 219712 625728 219776 625792
rect 219840 625728 219904 625792
rect 219968 625728 220032 625792
rect 220096 625728 220160 625792
rect 220224 625728 220288 625792
rect 220352 625728 220416 625792
rect 220480 625728 220544 625792
rect 220608 625728 220672 625792
rect 220736 625728 220800 625792
rect 220864 625728 220928 625792
rect 220992 625728 221056 625792
rect 221120 625728 221184 625792
rect 221248 625728 221312 625792
rect 221376 625728 221440 625792
rect 221504 625728 221568 625792
rect 221632 625728 221696 625792
rect 221760 625728 221824 625792
rect 221888 625728 221952 625792
rect 222016 625728 222080 625792
rect 222144 625728 222294 625792
rect 217294 625700 222294 625728
rect 227594 626176 232594 692092
rect 227594 626112 227640 626176
rect 227704 626112 227768 626176
rect 227832 626112 227896 626176
rect 227960 626112 228024 626176
rect 228088 626112 228152 626176
rect 228216 626112 228280 626176
rect 228344 626112 228408 626176
rect 228472 626112 228536 626176
rect 228600 626112 228664 626176
rect 228728 626112 228792 626176
rect 228856 626112 228920 626176
rect 228984 626112 229048 626176
rect 229112 626112 229176 626176
rect 229240 626112 229304 626176
rect 229368 626112 229432 626176
rect 229496 626112 229560 626176
rect 229624 626112 229688 626176
rect 229752 626112 229816 626176
rect 229880 626112 229944 626176
rect 230008 626112 230072 626176
rect 230136 626112 230200 626176
rect 230264 626112 230328 626176
rect 230392 626112 230456 626176
rect 230520 626112 230584 626176
rect 230648 626112 230712 626176
rect 230776 626112 230840 626176
rect 230904 626112 230968 626176
rect 231032 626112 231096 626176
rect 231160 626112 231224 626176
rect 231288 626112 231352 626176
rect 231416 626112 231480 626176
rect 231544 626112 231608 626176
rect 231672 626112 231736 626176
rect 231800 626112 231864 626176
rect 231928 626112 231992 626176
rect 232056 626112 232120 626176
rect 232184 626112 232248 626176
rect 232312 626112 232376 626176
rect 232440 626112 232594 626176
rect 227594 626048 232594 626112
rect 227594 625984 227640 626048
rect 227704 625984 227768 626048
rect 227832 625984 227896 626048
rect 227960 625984 228024 626048
rect 228088 625984 228152 626048
rect 228216 625984 228280 626048
rect 228344 625984 228408 626048
rect 228472 625984 228536 626048
rect 228600 625984 228664 626048
rect 228728 625984 228792 626048
rect 228856 625984 228920 626048
rect 228984 625984 229048 626048
rect 229112 625984 229176 626048
rect 229240 625984 229304 626048
rect 229368 625984 229432 626048
rect 229496 625984 229560 626048
rect 229624 625984 229688 626048
rect 229752 625984 229816 626048
rect 229880 625984 229944 626048
rect 230008 625984 230072 626048
rect 230136 625984 230200 626048
rect 230264 625984 230328 626048
rect 230392 625984 230456 626048
rect 230520 625984 230584 626048
rect 230648 625984 230712 626048
rect 230776 625984 230840 626048
rect 230904 625984 230968 626048
rect 231032 625984 231096 626048
rect 231160 625984 231224 626048
rect 231288 625984 231352 626048
rect 231416 625984 231480 626048
rect 231544 625984 231608 626048
rect 231672 625984 231736 626048
rect 231800 625984 231864 626048
rect 231928 625984 231992 626048
rect 232056 625984 232120 626048
rect 232184 625984 232248 626048
rect 232312 625984 232376 626048
rect 232440 625984 232594 626048
rect 227594 625920 232594 625984
rect 227594 625856 227640 625920
rect 227704 625856 227768 625920
rect 227832 625856 227896 625920
rect 227960 625856 228024 625920
rect 228088 625856 228152 625920
rect 228216 625856 228280 625920
rect 228344 625856 228408 625920
rect 228472 625856 228536 625920
rect 228600 625856 228664 625920
rect 228728 625856 228792 625920
rect 228856 625856 228920 625920
rect 228984 625856 229048 625920
rect 229112 625856 229176 625920
rect 229240 625856 229304 625920
rect 229368 625856 229432 625920
rect 229496 625856 229560 625920
rect 229624 625856 229688 625920
rect 229752 625856 229816 625920
rect 229880 625856 229944 625920
rect 230008 625856 230072 625920
rect 230136 625856 230200 625920
rect 230264 625856 230328 625920
rect 230392 625856 230456 625920
rect 230520 625856 230584 625920
rect 230648 625856 230712 625920
rect 230776 625856 230840 625920
rect 230904 625856 230968 625920
rect 231032 625856 231096 625920
rect 231160 625856 231224 625920
rect 231288 625856 231352 625920
rect 231416 625856 231480 625920
rect 231544 625856 231608 625920
rect 231672 625856 231736 625920
rect 231800 625856 231864 625920
rect 231928 625856 231992 625920
rect 232056 625856 232120 625920
rect 232184 625856 232248 625920
rect 232312 625856 232376 625920
rect 232440 625856 232594 625920
rect 227594 625792 232594 625856
rect 227594 625728 227640 625792
rect 227704 625728 227768 625792
rect 227832 625728 227896 625792
rect 227960 625728 228024 625792
rect 228088 625728 228152 625792
rect 228216 625728 228280 625792
rect 228344 625728 228408 625792
rect 228472 625728 228536 625792
rect 228600 625728 228664 625792
rect 228728 625728 228792 625792
rect 228856 625728 228920 625792
rect 228984 625728 229048 625792
rect 229112 625728 229176 625792
rect 229240 625728 229304 625792
rect 229368 625728 229432 625792
rect 229496 625728 229560 625792
rect 229624 625728 229688 625792
rect 229752 625728 229816 625792
rect 229880 625728 229944 625792
rect 230008 625728 230072 625792
rect 230136 625728 230200 625792
rect 230264 625728 230328 625792
rect 230392 625728 230456 625792
rect 230520 625728 230584 625792
rect 230648 625728 230712 625792
rect 230776 625728 230840 625792
rect 230904 625728 230968 625792
rect 231032 625728 231096 625792
rect 231160 625728 231224 625792
rect 231288 625728 231352 625792
rect 231416 625728 231480 625792
rect 231544 625728 231608 625792
rect 231672 625728 231736 625792
rect 231800 625728 231864 625792
rect 231928 625728 231992 625792
rect 232056 625728 232120 625792
rect 232184 625728 232248 625792
rect 232312 625728 232376 625792
rect 232440 625728 232594 625792
rect 227594 625700 232594 625728
rect 288920 690084 295576 690584
rect 288920 684340 289800 690084
rect 294584 684340 295576 690084
rect 288920 650584 295576 684340
rect 318994 683600 323994 704800
rect 324294 690593 326494 704800
rect 326794 694292 328994 704800
rect 329294 694292 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 326794 692092 334294 694292
rect 324294 684369 324322 690593
rect 326466 684369 326494 690593
rect 324294 684038 326494 684369
rect 329294 683600 334294 692092
rect 510594 690560 515394 704800
rect 510594 684336 510602 690560
rect 515386 684336 515394 690560
rect 288920 644840 289920 650584
rect 294704 644840 295576 650584
rect 288920 637184 295576 644840
rect 298820 650584 315980 651400
rect 298820 644840 298920 650584
rect 303704 644840 304920 650584
rect 309704 644840 310920 650584
rect 315704 644840 315980 650584
rect 318994 650200 334400 683600
rect 510594 651406 515394 684336
rect 298820 642694 315980 644840
rect 298820 642594 298876 642694
rect 298976 642594 299100 642694
rect 299200 642594 299324 642694
rect 299424 642594 299548 642694
rect 299648 642594 299772 642694
rect 299872 642594 299996 642694
rect 300096 642594 300220 642694
rect 300320 642594 300444 642694
rect 300544 642594 300668 642694
rect 300768 642594 300892 642694
rect 300992 642594 301116 642694
rect 301216 642594 301340 642694
rect 301440 642594 301564 642694
rect 301664 642594 301788 642694
rect 301888 642594 302012 642694
rect 302112 642594 302236 642694
rect 302336 642594 302460 642694
rect 302560 642594 302684 642694
rect 302784 642594 302908 642694
rect 303008 642594 303132 642694
rect 303232 642594 303356 642694
rect 303456 642594 303580 642694
rect 303680 642594 303804 642694
rect 303904 642594 304028 642694
rect 304128 642594 304252 642694
rect 304352 642594 304476 642694
rect 304576 642594 304700 642694
rect 304800 642594 304924 642694
rect 305024 642594 305148 642694
rect 305248 642594 305372 642694
rect 305472 642594 309346 642694
rect 309446 642594 309570 642694
rect 309670 642594 309794 642694
rect 309894 642594 310018 642694
rect 310118 642594 310242 642694
rect 310342 642594 310466 642694
rect 310566 642594 310690 642694
rect 310790 642594 310914 642694
rect 311014 642594 311138 642694
rect 311238 642594 311362 642694
rect 311462 642594 311586 642694
rect 311686 642594 311810 642694
rect 311910 642594 312034 642694
rect 312134 642594 312258 642694
rect 312358 642594 312482 642694
rect 312582 642594 312706 642694
rect 312806 642594 312930 642694
rect 313030 642594 313154 642694
rect 313254 642594 313378 642694
rect 313478 642594 313602 642694
rect 313702 642594 313826 642694
rect 313926 642594 314050 642694
rect 314150 642594 314274 642694
rect 314374 642594 314498 642694
rect 314598 642594 314722 642694
rect 314822 642594 314946 642694
rect 315046 642594 315170 642694
rect 315270 642594 315394 642694
rect 315494 642594 315618 642694
rect 315718 642594 315842 642694
rect 315942 642594 315980 642694
rect 298820 642470 315980 642594
rect 298820 642370 298876 642470
rect 298976 642370 299100 642470
rect 299200 642370 299324 642470
rect 299424 642370 299548 642470
rect 299648 642370 299772 642470
rect 299872 642370 299996 642470
rect 300096 642370 300220 642470
rect 300320 642370 300444 642470
rect 300544 642370 300668 642470
rect 300768 642370 300892 642470
rect 300992 642370 301116 642470
rect 301216 642370 301340 642470
rect 301440 642370 301564 642470
rect 301664 642370 301788 642470
rect 301888 642370 302012 642470
rect 302112 642370 302236 642470
rect 302336 642370 302460 642470
rect 302560 642370 302684 642470
rect 302784 642370 302908 642470
rect 303008 642370 303132 642470
rect 303232 642370 303356 642470
rect 303456 642370 303580 642470
rect 303680 642370 303804 642470
rect 303904 642370 304028 642470
rect 304128 642370 304252 642470
rect 304352 642370 304476 642470
rect 304576 642370 304700 642470
rect 304800 642370 304924 642470
rect 305024 642370 305148 642470
rect 305248 642370 305372 642470
rect 305472 642370 309346 642470
rect 309446 642370 309570 642470
rect 309670 642370 309794 642470
rect 309894 642370 310018 642470
rect 310118 642370 310242 642470
rect 310342 642370 310466 642470
rect 310566 642370 310690 642470
rect 310790 642370 310914 642470
rect 311014 642370 311138 642470
rect 311238 642370 311362 642470
rect 311462 642370 311586 642470
rect 311686 642370 311810 642470
rect 311910 642370 312034 642470
rect 312134 642370 312258 642470
rect 312358 642370 312482 642470
rect 312582 642370 312706 642470
rect 312806 642370 312930 642470
rect 313030 642370 313154 642470
rect 313254 642370 313378 642470
rect 313478 642370 313602 642470
rect 313702 642370 313826 642470
rect 313926 642370 314050 642470
rect 314150 642370 314274 642470
rect 314374 642370 314498 642470
rect 314598 642370 314722 642470
rect 314822 642370 314946 642470
rect 315046 642370 315170 642470
rect 315270 642370 315394 642470
rect 315494 642370 315618 642470
rect 315718 642370 315842 642470
rect 315942 642370 315980 642470
rect 298820 642246 315980 642370
rect 298820 642146 298876 642246
rect 298976 642146 299100 642246
rect 299200 642146 299324 642246
rect 299424 642146 299548 642246
rect 299648 642146 299772 642246
rect 299872 642146 299996 642246
rect 300096 642146 300220 642246
rect 300320 642146 300444 642246
rect 300544 642146 300668 642246
rect 300768 642146 300892 642246
rect 300992 642146 301116 642246
rect 301216 642146 301340 642246
rect 301440 642146 301564 642246
rect 301664 642146 301788 642246
rect 301888 642146 302012 642246
rect 302112 642146 302236 642246
rect 302336 642146 302460 642246
rect 302560 642146 302684 642246
rect 302784 642146 302908 642246
rect 303008 642146 303132 642246
rect 303232 642146 303356 642246
rect 303456 642146 303580 642246
rect 303680 642146 303804 642246
rect 303904 642146 304028 642246
rect 304128 642146 304252 642246
rect 304352 642146 304476 642246
rect 304576 642146 304700 642246
rect 304800 642146 304924 642246
rect 305024 642146 305148 642246
rect 305248 642146 305372 642246
rect 305472 642146 309346 642246
rect 309446 642146 309570 642246
rect 309670 642146 309794 642246
rect 309894 642146 310018 642246
rect 310118 642146 310242 642246
rect 310342 642146 310466 642246
rect 310566 642146 310690 642246
rect 310790 642146 310914 642246
rect 311014 642146 311138 642246
rect 311238 642146 311362 642246
rect 311462 642146 311586 642246
rect 311686 642146 311810 642246
rect 311910 642146 312034 642246
rect 312134 642146 312258 642246
rect 312358 642146 312482 642246
rect 312582 642146 312706 642246
rect 312806 642146 312930 642246
rect 313030 642146 313154 642246
rect 313254 642146 313378 642246
rect 313478 642146 313602 642246
rect 313702 642146 313826 642246
rect 313926 642146 314050 642246
rect 314150 642146 314274 642246
rect 314374 642146 314498 642246
rect 314598 642146 314722 642246
rect 314822 642146 314946 642246
rect 315046 642146 315170 642246
rect 315270 642146 315394 642246
rect 315494 642146 315618 642246
rect 315718 642146 315842 642246
rect 315942 642146 315980 642246
rect 298820 642022 315980 642146
rect 298820 641922 298876 642022
rect 298976 641922 299100 642022
rect 299200 641922 299324 642022
rect 299424 641922 299548 642022
rect 299648 641922 299772 642022
rect 299872 641922 299996 642022
rect 300096 641922 300220 642022
rect 300320 641922 300444 642022
rect 300544 641922 300668 642022
rect 300768 641922 300892 642022
rect 300992 641922 301116 642022
rect 301216 641922 301340 642022
rect 301440 641922 301564 642022
rect 301664 641922 301788 642022
rect 301888 641922 302012 642022
rect 302112 641922 302236 642022
rect 302336 641922 302460 642022
rect 302560 641922 302684 642022
rect 302784 641922 302908 642022
rect 303008 641922 303132 642022
rect 303232 641922 303356 642022
rect 303456 641922 303580 642022
rect 303680 641922 303804 642022
rect 303904 641922 304028 642022
rect 304128 641922 304252 642022
rect 304352 641922 304476 642022
rect 304576 641922 304700 642022
rect 304800 641922 304924 642022
rect 305024 641922 305148 642022
rect 305248 641922 305372 642022
rect 305472 641922 309346 642022
rect 309446 641922 309570 642022
rect 309670 641922 309794 642022
rect 309894 641922 310018 642022
rect 310118 641922 310242 642022
rect 310342 641922 310466 642022
rect 310566 641922 310690 642022
rect 310790 641922 310914 642022
rect 311014 641922 311138 642022
rect 311238 641922 311362 642022
rect 311462 641922 311586 642022
rect 311686 641922 311810 642022
rect 311910 641922 312034 642022
rect 312134 641922 312258 642022
rect 312358 641922 312482 642022
rect 312582 641922 312706 642022
rect 312806 641922 312930 642022
rect 313030 641922 313154 642022
rect 313254 641922 313378 642022
rect 313478 641922 313602 642022
rect 313702 641922 313826 642022
rect 313926 641922 314050 642022
rect 314150 641922 314274 642022
rect 314374 641922 314498 642022
rect 314598 641922 314722 642022
rect 314822 641922 314946 642022
rect 315046 641922 315170 642022
rect 315270 641922 315394 642022
rect 315494 641922 315618 642022
rect 315718 641922 315842 642022
rect 315942 641922 315980 642022
rect 298820 641798 315980 641922
rect 298820 641698 298876 641798
rect 298976 641698 299100 641798
rect 299200 641698 299324 641798
rect 299424 641698 299548 641798
rect 299648 641698 299772 641798
rect 299872 641698 299996 641798
rect 300096 641698 300220 641798
rect 300320 641698 300444 641798
rect 300544 641698 300668 641798
rect 300768 641698 300892 641798
rect 300992 641698 301116 641798
rect 301216 641698 301340 641798
rect 301440 641698 301564 641798
rect 301664 641698 301788 641798
rect 301888 641698 302012 641798
rect 302112 641698 302236 641798
rect 302336 641698 302460 641798
rect 302560 641698 302684 641798
rect 302784 641698 302908 641798
rect 303008 641698 303132 641798
rect 303232 641698 303356 641798
rect 303456 641698 303580 641798
rect 303680 641698 303804 641798
rect 303904 641698 304028 641798
rect 304128 641698 304252 641798
rect 304352 641698 304476 641798
rect 304576 641698 304700 641798
rect 304800 641698 304924 641798
rect 305024 641698 305148 641798
rect 305248 641698 305372 641798
rect 305472 641698 309346 641798
rect 309446 641698 309570 641798
rect 309670 641698 309794 641798
rect 309894 641698 310018 641798
rect 310118 641698 310242 641798
rect 310342 641698 310466 641798
rect 310566 641698 310690 641798
rect 310790 641698 310914 641798
rect 311014 641698 311138 641798
rect 311238 641698 311362 641798
rect 311462 641698 311586 641798
rect 311686 641698 311810 641798
rect 311910 641698 312034 641798
rect 312134 641698 312258 641798
rect 312358 641698 312482 641798
rect 312582 641698 312706 641798
rect 312806 641698 312930 641798
rect 313030 641698 313154 641798
rect 313254 641698 313378 641798
rect 313478 641698 313602 641798
rect 313702 641698 313826 641798
rect 313926 641698 314050 641798
rect 314150 641698 314274 641798
rect 314374 641698 314498 641798
rect 314598 641698 314722 641798
rect 314822 641698 314946 641798
rect 315046 641698 315170 641798
rect 315270 641698 315394 641798
rect 315494 641698 315618 641798
rect 315718 641698 315842 641798
rect 315942 641698 315980 641798
rect 298820 641660 315980 641698
rect 300637 640587 311923 640593
rect 300637 639731 300643 640587
rect 311917 639731 311923 640587
rect 300637 639725 311923 639731
rect 288920 631440 289920 637184
rect 294704 631440 295576 637184
rect 288920 623784 295576 631440
rect 297820 637996 298880 638020
rect 297820 637896 297850 637996
rect 297950 637896 298074 637996
rect 298174 637896 298298 637996
rect 298398 637896 298522 637996
rect 298622 637896 298746 637996
rect 298846 637896 298880 637996
rect 297820 637772 298880 637896
rect 297820 637672 297850 637772
rect 297950 637672 298074 637772
rect 298174 637672 298298 637772
rect 298398 637672 298522 637772
rect 298622 637672 298746 637772
rect 298846 637672 298880 637772
rect 297820 637548 298880 637672
rect 297820 637448 297850 637548
rect 297950 637448 298074 637548
rect 298174 637448 298298 637548
rect 298398 637448 298522 637548
rect 298622 637448 298746 637548
rect 298846 637448 298880 637548
rect 297820 637324 298880 637448
rect 297820 637224 297850 637324
rect 297950 637224 298074 637324
rect 298174 637224 298298 637324
rect 298398 637224 298522 637324
rect 298622 637224 298746 637324
rect 298846 637224 298880 637324
rect 297820 637100 298880 637224
rect 297820 637000 297850 637100
rect 297950 637000 298074 637100
rect 298174 637000 298298 637100
rect 298398 637000 298522 637100
rect 298622 637000 298746 637100
rect 298846 637000 298880 637100
rect 297820 636876 298880 637000
rect 297820 636776 297850 636876
rect 297950 636776 298074 636876
rect 298174 636776 298298 636876
rect 298398 636776 298522 636876
rect 298622 636776 298746 636876
rect 298846 636776 298880 636876
rect 297820 636652 298880 636776
rect 297820 636552 297850 636652
rect 297950 636552 298074 636652
rect 298174 636552 298298 636652
rect 298398 636552 298522 636652
rect 298622 636552 298746 636652
rect 298846 636552 298880 636652
rect 297820 636428 298880 636552
rect 297820 636328 297850 636428
rect 297950 636328 298074 636428
rect 298174 636328 298298 636428
rect 298398 636328 298522 636428
rect 298622 636328 298746 636428
rect 298846 636328 298880 636428
rect 297820 636204 298880 636328
rect 297820 636104 297850 636204
rect 297950 636104 298074 636204
rect 298174 636104 298298 636204
rect 298398 636104 298522 636204
rect 298622 636104 298746 636204
rect 298846 636104 298880 636204
rect 297820 635980 298880 636104
rect 297820 635880 297850 635980
rect 297950 635880 298074 635980
rect 298174 635880 298298 635980
rect 298398 635880 298522 635980
rect 298622 635880 298746 635980
rect 298846 635880 298880 635980
rect 297820 635756 298880 635880
rect 297820 635656 297850 635756
rect 297950 635656 298074 635756
rect 298174 635656 298298 635756
rect 298398 635656 298522 635756
rect 298622 635656 298746 635756
rect 298846 635656 298880 635756
rect 297820 635532 298880 635656
rect 297820 635432 297850 635532
rect 297950 635432 298074 635532
rect 298174 635432 298298 635532
rect 298398 635432 298522 635532
rect 298622 635432 298746 635532
rect 298846 635432 298880 635532
rect 297820 635308 298880 635432
rect 297820 635208 297850 635308
rect 297950 635208 298074 635308
rect 298174 635208 298298 635308
rect 298398 635208 298522 635308
rect 298622 635208 298746 635308
rect 298846 635208 298880 635308
rect 297820 635084 298880 635208
rect 297820 634984 297850 635084
rect 297950 634984 298074 635084
rect 298174 634984 298298 635084
rect 298398 634984 298522 635084
rect 298622 634984 298746 635084
rect 298846 634984 298880 635084
rect 297820 634860 298880 634984
rect 297820 634760 297850 634860
rect 297950 634760 298074 634860
rect 298174 634760 298298 634860
rect 298398 634760 298522 634860
rect 298622 634760 298746 634860
rect 298846 634760 298880 634860
rect 297820 634636 298880 634760
rect 297820 634536 297850 634636
rect 297950 634536 298074 634636
rect 298174 634536 298298 634636
rect 298398 634536 298522 634636
rect 298622 634536 298746 634636
rect 298846 634536 298880 634636
rect 297820 634412 298880 634536
rect 297820 634312 297850 634412
rect 297950 634312 298074 634412
rect 298174 634312 298298 634412
rect 298398 634312 298522 634412
rect 298622 634312 298746 634412
rect 298846 634312 298880 634412
rect 297820 634188 298880 634312
rect 297820 634088 297850 634188
rect 297950 634088 298074 634188
rect 298174 634088 298298 634188
rect 298398 634088 298522 634188
rect 298622 634088 298746 634188
rect 298846 634088 298880 634188
rect 297820 633964 298880 634088
rect 297820 633864 297850 633964
rect 297950 633864 298074 633964
rect 298174 633864 298298 633964
rect 298398 633864 298522 633964
rect 298622 633864 298746 633964
rect 298846 633864 298880 633964
rect 297820 633740 298880 633864
rect 297820 633640 297850 633740
rect 297950 633640 298074 633740
rect 298174 633640 298298 633740
rect 298398 633640 298522 633740
rect 298622 633640 298746 633740
rect 298846 633640 298880 633740
rect 297820 633516 298880 633640
rect 297820 633416 297850 633516
rect 297950 633416 298074 633516
rect 298174 633416 298298 633516
rect 298398 633416 298522 633516
rect 298622 633416 298746 633516
rect 298846 633416 298880 633516
rect 297820 633292 298880 633416
rect 297820 633192 297850 633292
rect 297950 633192 298074 633292
rect 298174 633192 298298 633292
rect 298398 633192 298522 633292
rect 298622 633192 298746 633292
rect 298846 633192 298880 633292
rect 297820 633068 298880 633192
rect 297820 632968 297850 633068
rect 297950 632968 298074 633068
rect 298174 632968 298298 633068
rect 298398 632968 298522 633068
rect 298622 632968 298746 633068
rect 298846 632968 298880 633068
rect 297820 632844 298880 632968
rect 297820 632744 297850 632844
rect 297950 632744 298074 632844
rect 298174 632744 298298 632844
rect 298398 632744 298522 632844
rect 298622 632744 298746 632844
rect 298846 632744 298880 632844
rect 297820 632620 298880 632744
rect 297820 632520 297850 632620
rect 297950 632520 298074 632620
rect 298174 632520 298298 632620
rect 298398 632520 298522 632620
rect 298622 632520 298746 632620
rect 298846 632520 298880 632620
rect 297820 632396 298880 632520
rect 297820 632296 297850 632396
rect 297950 632296 298074 632396
rect 298174 632296 298298 632396
rect 298398 632296 298522 632396
rect 298622 632296 298746 632396
rect 298846 632296 298880 632396
rect 297820 632172 298880 632296
rect 297820 632072 297850 632172
rect 297950 632072 298074 632172
rect 298174 632072 298298 632172
rect 298398 632072 298522 632172
rect 298622 632072 298746 632172
rect 298846 632072 298880 632172
rect 297820 631948 298880 632072
rect 297820 631848 297850 631948
rect 297950 631848 298074 631948
rect 298174 631848 298298 631948
rect 298398 631848 298522 631948
rect 298622 631848 298746 631948
rect 298846 631848 298880 631948
rect 297820 631724 298880 631848
rect 297820 631624 297850 631724
rect 297950 631624 298074 631724
rect 298174 631624 298298 631724
rect 298398 631624 298522 631724
rect 298622 631624 298746 631724
rect 298846 631624 298880 631724
rect 297820 631500 298880 631624
rect 297820 631400 297850 631500
rect 297950 631400 298074 631500
rect 298174 631400 298298 631500
rect 298398 631400 298522 631500
rect 298622 631400 298746 631500
rect 298846 631400 298880 631500
rect 297820 631360 298880 631400
rect 304316 632144 311486 632172
rect 304316 631600 304931 632144
rect 304995 631600 305650 632144
rect 305714 631600 306369 632144
rect 306433 631600 307088 632144
rect 307152 631600 307807 632144
rect 307871 631600 308526 632144
rect 308590 631600 309245 632144
rect 309309 631600 309964 632144
rect 310028 631600 310683 632144
rect 310747 631600 311402 632144
rect 311466 631600 311486 632144
rect 304316 631444 311486 631600
rect 304316 630900 304931 631444
rect 304995 630900 305650 631444
rect 305714 630900 306369 631444
rect 306433 630900 307088 631444
rect 307152 630900 307807 631444
rect 307871 630900 308526 631444
rect 308590 630900 309245 631444
rect 309309 630900 309964 631444
rect 310028 630900 310683 631444
rect 310747 630900 311402 631444
rect 311466 630900 311486 631444
rect 304316 630744 311486 630900
rect 304316 630200 304931 630744
rect 304995 630200 305650 630744
rect 305714 630200 306369 630744
rect 306433 630200 307088 630744
rect 307152 630200 307807 630744
rect 307871 630200 308526 630744
rect 308590 630200 309245 630744
rect 309309 630200 309964 630744
rect 310028 630200 310683 630744
rect 310747 630200 311402 630744
rect 311466 630200 311486 630744
rect 304316 630044 311486 630200
rect 304316 629500 304931 630044
rect 304995 629500 305650 630044
rect 305714 629500 306369 630044
rect 306433 629500 307088 630044
rect 307152 629500 307807 630044
rect 307871 629500 308526 630044
rect 308590 629500 309245 630044
rect 309309 629500 309964 630044
rect 310028 629500 310683 630044
rect 310747 629500 311402 630044
rect 311466 629500 311486 630044
rect 304316 629344 311486 629500
rect 304316 628800 304931 629344
rect 304995 628800 305650 629344
rect 305714 628800 306369 629344
rect 306433 628800 307088 629344
rect 307152 628800 307807 629344
rect 307871 628800 308526 629344
rect 308590 628800 309245 629344
rect 309309 628800 309964 629344
rect 310028 628800 310683 629344
rect 310747 628800 311402 629344
rect 311466 628800 311486 629344
rect 304316 628644 311486 628800
rect 304316 628100 304931 628644
rect 304995 628100 305650 628644
rect 305714 628100 306369 628644
rect 306433 628100 307088 628644
rect 307152 628100 307807 628644
rect 307871 628100 308526 628644
rect 308590 628100 309245 628644
rect 309309 628100 309964 628644
rect 310028 628100 310683 628644
rect 310747 628100 311402 628644
rect 311466 628100 311486 628644
rect 304316 627944 311486 628100
rect 304316 627400 304931 627944
rect 304995 627400 305650 627944
rect 305714 627400 306369 627944
rect 306433 627400 307088 627944
rect 307152 627400 307807 627944
rect 307871 627400 308526 627944
rect 308590 627400 309245 627944
rect 309309 627400 309964 627944
rect 310028 627400 310683 627944
rect 310747 627400 311402 627944
rect 311466 627400 311486 627944
rect 319000 628868 334400 650200
rect 335580 650904 342400 651380
rect 335580 645160 336480 650904
rect 341264 645160 342400 650904
rect 335580 642744 342400 645160
rect 510602 650961 515394 651406
rect 515386 645217 515394 650961
rect 510602 644744 515394 645217
rect 335576 642714 342400 642744
rect 335576 642614 335616 642714
rect 335716 642614 335840 642714
rect 335940 642614 336064 642714
rect 336164 642614 336288 642714
rect 336388 642614 336512 642714
rect 336612 642614 336736 642714
rect 336836 642614 336960 642714
rect 337060 642614 337184 642714
rect 337284 642614 337408 642714
rect 337508 642614 337632 642714
rect 337732 642614 337856 642714
rect 337956 642614 338080 642714
rect 338180 642614 338304 642714
rect 338404 642614 338528 642714
rect 338628 642614 338752 642714
rect 338852 642614 338976 642714
rect 339076 642614 339200 642714
rect 339300 642614 339424 642714
rect 339524 642614 339648 642714
rect 339748 642614 339872 642714
rect 339972 642614 340096 642714
rect 340196 642614 340320 642714
rect 340420 642614 340544 642714
rect 340644 642614 340768 642714
rect 340868 642614 340992 642714
rect 341092 642614 341216 642714
rect 341316 642614 341440 642714
rect 341540 642614 341664 642714
rect 341764 642614 341888 642714
rect 341988 642614 342112 642714
rect 342212 642614 342400 642714
rect 335576 642490 342400 642614
rect 335576 642390 335616 642490
rect 335716 642390 335840 642490
rect 335940 642390 336064 642490
rect 336164 642390 336288 642490
rect 336388 642390 336512 642490
rect 336612 642390 336736 642490
rect 336836 642390 336960 642490
rect 337060 642390 337184 642490
rect 337284 642390 337408 642490
rect 337508 642390 337632 642490
rect 337732 642390 337856 642490
rect 337956 642390 338080 642490
rect 338180 642390 338304 642490
rect 338404 642390 338528 642490
rect 338628 642390 338752 642490
rect 338852 642390 338976 642490
rect 339076 642390 339200 642490
rect 339300 642390 339424 642490
rect 339524 642390 339648 642490
rect 339748 642390 339872 642490
rect 339972 642390 340096 642490
rect 340196 642390 340320 642490
rect 340420 642390 340544 642490
rect 340644 642390 340768 642490
rect 340868 642390 340992 642490
rect 341092 642390 341216 642490
rect 341316 642390 341440 642490
rect 341540 642390 341664 642490
rect 341764 642390 341888 642490
rect 341988 642390 342112 642490
rect 342212 642390 342400 642490
rect 335576 642266 342400 642390
rect 335576 642166 335616 642266
rect 335716 642166 335840 642266
rect 335940 642166 336064 642266
rect 336164 642166 336288 642266
rect 336388 642166 336512 642266
rect 336612 642166 336736 642266
rect 336836 642166 336960 642266
rect 337060 642166 337184 642266
rect 337284 642166 337408 642266
rect 337508 642166 337632 642266
rect 337732 642166 337856 642266
rect 337956 642166 338080 642266
rect 338180 642166 338304 642266
rect 338404 642166 338528 642266
rect 338628 642166 338752 642266
rect 338852 642166 338976 642266
rect 339076 642166 339200 642266
rect 339300 642166 339424 642266
rect 339524 642166 339648 642266
rect 339748 642166 339872 642266
rect 339972 642166 340096 642266
rect 340196 642166 340320 642266
rect 340420 642166 340544 642266
rect 340644 642166 340768 642266
rect 340868 642166 340992 642266
rect 341092 642166 341216 642266
rect 341316 642166 341440 642266
rect 341540 642166 341664 642266
rect 341764 642166 341888 642266
rect 341988 642166 342112 642266
rect 342212 642166 342400 642266
rect 335576 642042 342400 642166
rect 335576 641942 335616 642042
rect 335716 641942 335840 642042
rect 335940 641942 336064 642042
rect 336164 641942 336288 642042
rect 336388 641942 336512 642042
rect 336612 641942 336736 642042
rect 336836 641942 336960 642042
rect 337060 641942 337184 642042
rect 337284 641942 337408 642042
rect 337508 641942 337632 642042
rect 337732 641942 337856 642042
rect 337956 641942 338080 642042
rect 338180 641942 338304 642042
rect 338404 641942 338528 642042
rect 338628 641942 338752 642042
rect 338852 641942 338976 642042
rect 339076 641942 339200 642042
rect 339300 641942 339424 642042
rect 339524 641942 339648 642042
rect 339748 641942 339872 642042
rect 339972 641942 340096 642042
rect 340196 641942 340320 642042
rect 340420 641942 340544 642042
rect 340644 641942 340768 642042
rect 340868 641942 340992 642042
rect 341092 641942 341216 642042
rect 341316 641942 341440 642042
rect 341540 641942 341664 642042
rect 341764 641942 341888 642042
rect 341988 641942 342112 642042
rect 342212 641942 342400 642042
rect 335576 641818 342400 641942
rect 335576 641718 335616 641818
rect 335716 641718 335840 641818
rect 335940 641718 336064 641818
rect 336164 641718 336288 641818
rect 336388 641718 336512 641818
rect 336612 641718 336736 641818
rect 336836 641718 336960 641818
rect 337060 641718 337184 641818
rect 337284 641718 337408 641818
rect 337508 641718 337632 641818
rect 337732 641718 337856 641818
rect 337956 641718 338080 641818
rect 338180 641718 338304 641818
rect 338404 641718 338528 641818
rect 338628 641718 338752 641818
rect 338852 641718 338976 641818
rect 339076 641718 339200 641818
rect 339300 641718 339424 641818
rect 339524 641718 339648 641818
rect 339748 641718 339872 641818
rect 339972 641718 340096 641818
rect 340196 641718 340320 641818
rect 340420 641718 340544 641818
rect 340644 641718 340768 641818
rect 340868 641718 340992 641818
rect 341092 641718 341216 641818
rect 341316 641718 341440 641818
rect 341540 641718 341664 641818
rect 341764 641718 341888 641818
rect 341988 641718 342112 641818
rect 342212 641718 342400 641818
rect 335576 641684 342400 641718
rect 335580 641660 342400 641684
rect 342100 637996 343160 638020
rect 342100 637896 342130 637996
rect 342230 637896 342354 637996
rect 342454 637896 342578 637996
rect 342678 637896 342802 637996
rect 342902 637896 343026 637996
rect 343126 637896 343160 637996
rect 342100 637772 343160 637896
rect 342100 637672 342130 637772
rect 342230 637672 342354 637772
rect 342454 637672 342578 637772
rect 342678 637672 342802 637772
rect 342902 637672 343026 637772
rect 343126 637672 343160 637772
rect 342100 637548 343160 637672
rect 342100 637448 342130 637548
rect 342230 637448 342354 637548
rect 342454 637448 342578 637548
rect 342678 637448 342802 637548
rect 342902 637448 343026 637548
rect 343126 637448 343160 637548
rect 342100 637324 343160 637448
rect 342100 637224 342130 637324
rect 342230 637224 342354 637324
rect 342454 637224 342578 637324
rect 342678 637224 342802 637324
rect 342902 637224 343026 637324
rect 343126 637224 343160 637324
rect 342100 637100 343160 637224
rect 342100 637000 342130 637100
rect 342230 637000 342354 637100
rect 342454 637000 342578 637100
rect 342678 637000 342802 637100
rect 342902 637000 343026 637100
rect 343126 637000 343160 637100
rect 342100 636876 343160 637000
rect 342100 636776 342130 636876
rect 342230 636776 342354 636876
rect 342454 636776 342578 636876
rect 342678 636776 342802 636876
rect 342902 636776 343026 636876
rect 343126 636776 343160 636876
rect 342100 636652 343160 636776
rect 342100 636552 342130 636652
rect 342230 636552 342354 636652
rect 342454 636552 342578 636652
rect 342678 636552 342802 636652
rect 342902 636552 343026 636652
rect 343126 636552 343160 636652
rect 342100 636428 343160 636552
rect 342100 636328 342130 636428
rect 342230 636328 342354 636428
rect 342454 636328 342578 636428
rect 342678 636328 342802 636428
rect 342902 636328 343026 636428
rect 343126 636328 343160 636428
rect 342100 636204 343160 636328
rect 342100 636104 342130 636204
rect 342230 636104 342354 636204
rect 342454 636104 342578 636204
rect 342678 636104 342802 636204
rect 342902 636104 343026 636204
rect 343126 636104 343160 636204
rect 342100 635980 343160 636104
rect 342100 635880 342130 635980
rect 342230 635880 342354 635980
rect 342454 635880 342578 635980
rect 342678 635880 342802 635980
rect 342902 635880 343026 635980
rect 343126 635880 343160 635980
rect 342100 635756 343160 635880
rect 342100 635656 342130 635756
rect 342230 635656 342354 635756
rect 342454 635656 342578 635756
rect 342678 635656 342802 635756
rect 342902 635656 343026 635756
rect 343126 635656 343160 635756
rect 342100 635532 343160 635656
rect 342100 635432 342130 635532
rect 342230 635432 342354 635532
rect 342454 635432 342578 635532
rect 342678 635432 342802 635532
rect 342902 635432 343026 635532
rect 343126 635432 343160 635532
rect 342100 635308 343160 635432
rect 342100 635208 342130 635308
rect 342230 635208 342354 635308
rect 342454 635208 342578 635308
rect 342678 635208 342802 635308
rect 342902 635208 343026 635308
rect 343126 635208 343160 635308
rect 342100 635084 343160 635208
rect 342100 634984 342130 635084
rect 342230 634984 342354 635084
rect 342454 634984 342578 635084
rect 342678 634984 342802 635084
rect 342902 634984 343026 635084
rect 343126 634984 343160 635084
rect 342100 634860 343160 634984
rect 342100 634760 342130 634860
rect 342230 634760 342354 634860
rect 342454 634760 342578 634860
rect 342678 634760 342802 634860
rect 342902 634760 343026 634860
rect 343126 634760 343160 634860
rect 342100 634636 343160 634760
rect 342100 634536 342130 634636
rect 342230 634536 342354 634636
rect 342454 634536 342578 634636
rect 342678 634536 342802 634636
rect 342902 634536 343026 634636
rect 343126 634536 343160 634636
rect 342100 634412 343160 634536
rect 342100 634312 342130 634412
rect 342230 634312 342354 634412
rect 342454 634312 342578 634412
rect 342678 634312 342802 634412
rect 342902 634312 343026 634412
rect 343126 634312 343160 634412
rect 342100 634188 343160 634312
rect 342100 634088 342130 634188
rect 342230 634088 342354 634188
rect 342454 634088 342578 634188
rect 342678 634088 342802 634188
rect 342902 634088 343026 634188
rect 343126 634088 343160 634188
rect 342100 633964 343160 634088
rect 342100 633864 342130 633964
rect 342230 633864 342354 633964
rect 342454 633864 342578 633964
rect 342678 633864 342802 633964
rect 342902 633864 343026 633964
rect 343126 633864 343160 633964
rect 342100 633740 343160 633864
rect 342100 633640 342130 633740
rect 342230 633640 342354 633740
rect 342454 633640 342578 633740
rect 342678 633640 342802 633740
rect 342902 633640 343026 633740
rect 343126 633640 343160 633740
rect 342100 633516 343160 633640
rect 342100 633416 342130 633516
rect 342230 633416 342354 633516
rect 342454 633416 342578 633516
rect 342678 633416 342802 633516
rect 342902 633416 343026 633516
rect 343126 633416 343160 633516
rect 342100 633292 343160 633416
rect 342100 633192 342130 633292
rect 342230 633192 342354 633292
rect 342454 633192 342578 633292
rect 342678 633192 342802 633292
rect 342902 633192 343026 633292
rect 343126 633192 343160 633292
rect 342100 633068 343160 633192
rect 342100 632968 342130 633068
rect 342230 632968 342354 633068
rect 342454 632968 342578 633068
rect 342678 632968 342802 633068
rect 342902 632968 343026 633068
rect 343126 632968 343160 633068
rect 342100 632844 343160 632968
rect 342100 632744 342130 632844
rect 342230 632744 342354 632844
rect 342454 632744 342578 632844
rect 342678 632744 342802 632844
rect 342902 632744 343026 632844
rect 343126 632744 343160 632844
rect 342100 632620 343160 632744
rect 342100 632520 342130 632620
rect 342230 632520 342354 632620
rect 342454 632520 342578 632620
rect 342678 632520 342802 632620
rect 342902 632520 343026 632620
rect 343126 632520 343160 632620
rect 342100 632396 343160 632520
rect 342100 632296 342130 632396
rect 342230 632296 342354 632396
rect 342454 632296 342578 632396
rect 342678 632296 342802 632396
rect 342902 632296 343026 632396
rect 343126 632296 343160 632396
rect 342100 632172 343160 632296
rect 342100 632072 342130 632172
rect 342230 632072 342354 632172
rect 342454 632072 342578 632172
rect 342678 632072 342802 632172
rect 342902 632072 343026 632172
rect 343126 632072 343160 632172
rect 342100 631948 343160 632072
rect 342100 631848 342130 631948
rect 342230 631848 342354 631948
rect 342454 631848 342578 631948
rect 342678 631848 342802 631948
rect 342902 631848 343026 631948
rect 343126 631848 343160 631948
rect 342100 631724 343160 631848
rect 342100 631624 342130 631724
rect 342230 631624 342354 631724
rect 342454 631624 342578 631724
rect 342678 631624 342802 631724
rect 342902 631624 343026 631724
rect 343126 631624 343160 631724
rect 342100 631500 343160 631624
rect 342100 631400 342130 631500
rect 342230 631400 342354 631500
rect 342454 631400 342578 631500
rect 342678 631400 342802 631500
rect 342902 631400 343026 631500
rect 343126 631400 343160 631500
rect 342100 631360 343160 631400
rect 510594 637561 515394 644744
rect 510594 631817 510602 637561
rect 515386 631817 515394 637561
rect 319000 628668 319400 628868
rect 319600 628668 319834 628868
rect 320034 628668 320268 628868
rect 320468 628668 320702 628868
rect 320902 628668 321136 628868
rect 321336 628668 321570 628868
rect 321770 628668 322004 628868
rect 322204 628668 322438 628868
rect 322638 628668 322872 628868
rect 323072 628668 323306 628868
rect 323506 628668 323740 628868
rect 323940 628668 324140 628868
rect 324340 628668 324540 628868
rect 324740 628668 324940 628868
rect 325140 628668 325340 628868
rect 325540 628668 325740 628868
rect 325940 628668 326140 628868
rect 326340 628668 326540 628868
rect 326740 628668 326940 628868
rect 327140 628668 327340 628868
rect 327540 628668 328940 628868
rect 329140 628668 329340 628868
rect 329540 628668 329740 628868
rect 329940 628668 330140 628868
rect 330340 628668 330540 628868
rect 330740 628668 330940 628868
rect 331140 628668 331340 628868
rect 331540 628668 331740 628868
rect 331940 628668 332140 628868
rect 332340 628668 334400 628868
rect 319000 628434 334400 628668
rect 319000 628234 319400 628434
rect 319600 628234 319834 628434
rect 320034 628234 320268 628434
rect 320468 628234 320702 628434
rect 320902 628234 321136 628434
rect 321336 628234 321570 628434
rect 321770 628234 322004 628434
rect 322204 628234 322438 628434
rect 322638 628234 322872 628434
rect 323072 628234 323306 628434
rect 323506 628234 323740 628434
rect 323940 628234 334400 628434
rect 319000 628000 334400 628234
rect 319000 627800 319400 628000
rect 319600 627800 319834 628000
rect 320034 627800 320268 628000
rect 320468 627800 320702 628000
rect 320902 627800 321136 628000
rect 321336 627800 321570 628000
rect 321770 627800 322004 628000
rect 322204 627800 322438 628000
rect 322638 627800 322872 628000
rect 323072 627800 323306 628000
rect 323506 627800 323740 628000
rect 323940 627800 334400 628000
rect 319000 627600 334400 627800
rect 304316 627244 311486 627400
rect 304316 626700 304931 627244
rect 304995 626700 305650 627244
rect 305714 626700 306369 627244
rect 306433 626700 307088 627244
rect 307152 626700 307807 627244
rect 307871 626700 308526 627244
rect 308590 626700 309245 627244
rect 309309 626700 309964 627244
rect 310028 626700 310683 627244
rect 310747 626700 311402 627244
rect 311466 626700 311486 627244
rect 304316 626544 311486 626700
rect 297792 626176 303552 626240
rect 297792 626112 297856 626176
rect 297920 626112 297984 626176
rect 298048 626112 298112 626176
rect 298176 626112 298240 626176
rect 298304 626112 298368 626176
rect 298432 626112 298496 626176
rect 298560 626112 298624 626176
rect 298688 626112 298752 626176
rect 298816 626112 298880 626176
rect 298944 626112 303552 626176
rect 297792 626048 303552 626112
rect 297792 625984 297856 626048
rect 297920 625984 297984 626048
rect 298048 625984 298112 626048
rect 298176 625984 298240 626048
rect 298304 625984 298368 626048
rect 298432 625984 298496 626048
rect 298560 625984 298624 626048
rect 298688 625984 298752 626048
rect 298816 625984 298880 626048
rect 298944 626030 303552 626048
rect 298944 625984 302980 626030
rect 297792 625970 302980 625984
rect 303040 625970 303100 626030
rect 303160 625970 303220 626030
rect 303280 625970 303340 626030
rect 303400 625970 303460 626030
rect 303520 625970 303552 626030
rect 297792 625920 303552 625970
rect 297792 625856 297856 625920
rect 297920 625856 297984 625920
rect 298048 625856 298112 625920
rect 298176 625856 298240 625920
rect 298304 625856 298368 625920
rect 298432 625856 298496 625920
rect 298560 625856 298624 625920
rect 298688 625856 298752 625920
rect 298816 625856 298880 625920
rect 298944 625910 303552 625920
rect 298944 625856 302980 625910
rect 297792 625850 302980 625856
rect 303040 625850 303100 625910
rect 303160 625850 303220 625910
rect 303280 625850 303340 625910
rect 303400 625850 303460 625910
rect 303520 625850 303552 625910
rect 297792 625792 303552 625850
rect 297792 625728 297856 625792
rect 297920 625728 297984 625792
rect 298048 625728 298112 625792
rect 298176 625728 298240 625792
rect 298304 625728 298368 625792
rect 298432 625728 298496 625792
rect 298560 625728 298624 625792
rect 298688 625728 298752 625792
rect 298816 625728 298880 625792
rect 298944 625728 303552 625792
rect 297792 625664 303552 625728
rect 304316 626000 304931 626544
rect 304995 626000 305650 626544
rect 305714 626000 306369 626544
rect 306433 626000 307088 626544
rect 307152 626000 307807 626544
rect 307871 626000 308526 626544
rect 308590 626000 309245 626544
rect 309309 626000 309964 626544
rect 310028 626000 310683 626544
rect 310747 626000 311402 626544
rect 311466 626000 311486 626544
rect 312947 627292 333279 627297
rect 312947 626308 312952 627292
rect 333274 626308 333279 627292
rect 312947 626303 333279 626308
rect 304316 625844 311486 626000
rect 304316 625300 304931 625844
rect 304995 625300 305650 625844
rect 305714 625300 306369 625844
rect 306433 625300 307088 625844
rect 307152 625300 307807 625844
rect 307871 625300 308526 625844
rect 308590 625300 309245 625844
rect 309309 625300 309964 625844
rect 310028 625300 310683 625844
rect 310747 625300 311402 625844
rect 311466 625300 311486 625844
rect 297820 624600 298878 624606
rect 288920 618040 289920 623784
rect 294704 618040 295576 623784
rect 288920 610764 295576 618040
rect 297720 624596 298880 624600
rect 297720 624496 297850 624596
rect 297950 624496 298074 624596
rect 298174 624496 298298 624596
rect 298398 624496 298522 624596
rect 298622 624496 298746 624596
rect 298846 624496 298880 624596
rect 297720 624372 298880 624496
rect 297720 624272 297850 624372
rect 297950 624272 298074 624372
rect 298174 624272 298298 624372
rect 298398 624272 298522 624372
rect 298622 624272 298746 624372
rect 298846 624272 298880 624372
rect 297720 624148 298880 624272
rect 297720 624048 297850 624148
rect 297950 624048 298074 624148
rect 298174 624048 298298 624148
rect 298398 624048 298522 624148
rect 298622 624048 298746 624148
rect 298846 624048 298880 624148
rect 297720 623924 298880 624048
rect 297720 623824 297850 623924
rect 297950 623824 298074 623924
rect 298174 623824 298298 623924
rect 298398 623824 298522 623924
rect 298622 623824 298746 623924
rect 298846 623824 298880 623924
rect 297720 623700 298880 623824
rect 297720 623600 297850 623700
rect 297950 623600 298074 623700
rect 298174 623600 298298 623700
rect 298398 623600 298522 623700
rect 298622 623600 298746 623700
rect 298846 623600 298880 623700
rect 297720 623476 298880 623600
rect 297720 623376 297850 623476
rect 297950 623376 298074 623476
rect 298174 623376 298298 623476
rect 298398 623376 298522 623476
rect 298622 623376 298746 623476
rect 298846 623376 298880 623476
rect 297720 623252 298880 623376
rect 297720 623152 297850 623252
rect 297950 623152 298074 623252
rect 298174 623152 298298 623252
rect 298398 623152 298522 623252
rect 298622 623152 298746 623252
rect 298846 623152 298880 623252
rect 297720 623028 298880 623152
rect 297720 622928 297850 623028
rect 297950 622928 298074 623028
rect 298174 622928 298298 623028
rect 298398 622928 298522 623028
rect 298622 622928 298746 623028
rect 298846 622928 298880 623028
rect 297720 622804 298880 622928
rect 297720 622704 297850 622804
rect 297950 622704 298074 622804
rect 298174 622704 298298 622804
rect 298398 622704 298522 622804
rect 298622 622704 298746 622804
rect 298846 622704 298880 622804
rect 297720 622580 298880 622704
rect 297720 622480 297850 622580
rect 297950 622480 298074 622580
rect 298174 622480 298298 622580
rect 298398 622480 298522 622580
rect 298622 622480 298746 622580
rect 298846 622480 298880 622580
rect 297720 622356 298880 622480
rect 297720 622256 297850 622356
rect 297950 622256 298074 622356
rect 298174 622256 298298 622356
rect 298398 622256 298522 622356
rect 298622 622256 298746 622356
rect 298846 622256 298880 622356
rect 297720 622132 298880 622256
rect 297720 622032 297850 622132
rect 297950 622032 298074 622132
rect 298174 622032 298298 622132
rect 298398 622032 298522 622132
rect 298622 622032 298746 622132
rect 298846 622032 298880 622132
rect 297720 621908 298880 622032
rect 297720 621808 297850 621908
rect 297950 621808 298074 621908
rect 298174 621808 298298 621908
rect 298398 621808 298522 621908
rect 298622 621808 298746 621908
rect 298846 621808 298880 621908
rect 297720 621684 298880 621808
rect 297720 621584 297850 621684
rect 297950 621584 298074 621684
rect 298174 621584 298298 621684
rect 298398 621584 298522 621684
rect 298622 621584 298746 621684
rect 298846 621584 298880 621684
rect 297720 621460 298880 621584
rect 297720 621360 297850 621460
rect 297950 621360 298074 621460
rect 298174 621360 298298 621460
rect 298398 621360 298522 621460
rect 298622 621360 298746 621460
rect 298846 621360 298880 621460
rect 297720 621236 298880 621360
rect 297720 621136 297850 621236
rect 297950 621136 298074 621236
rect 298174 621136 298298 621236
rect 298398 621136 298522 621236
rect 298622 621136 298746 621236
rect 298846 621136 298880 621236
rect 297720 621012 298880 621136
rect 297720 620912 297850 621012
rect 297950 620912 298074 621012
rect 298174 620912 298298 621012
rect 298398 620912 298522 621012
rect 298622 620912 298746 621012
rect 298846 620912 298880 621012
rect 297720 620788 298880 620912
rect 297720 620688 297850 620788
rect 297950 620688 298074 620788
rect 298174 620688 298298 620788
rect 298398 620688 298522 620788
rect 298622 620688 298746 620788
rect 298846 620688 298880 620788
rect 297720 620564 298880 620688
rect 297720 620464 297850 620564
rect 297950 620464 298074 620564
rect 298174 620464 298298 620564
rect 298398 620464 298522 620564
rect 298622 620464 298746 620564
rect 298846 620464 298880 620564
rect 297720 620340 298880 620464
rect 297720 620240 297850 620340
rect 297950 620240 298074 620340
rect 298174 620240 298298 620340
rect 298398 620240 298522 620340
rect 298622 620240 298746 620340
rect 298846 620240 298880 620340
rect 297720 620116 298880 620240
rect 297720 620016 297850 620116
rect 297950 620016 298074 620116
rect 298174 620016 298298 620116
rect 298398 620016 298522 620116
rect 298622 620016 298746 620116
rect 298846 620016 298880 620116
rect 297720 619892 298880 620016
rect 297720 619792 297850 619892
rect 297950 619792 298074 619892
rect 298174 619792 298298 619892
rect 298398 619792 298522 619892
rect 298622 619792 298746 619892
rect 298846 619792 298880 619892
rect 303584 620149 304224 620155
rect 303584 619869 303590 620149
rect 304218 619869 304224 620149
rect 303584 619863 304224 619869
rect 297720 619668 298880 619792
rect 297720 619568 297850 619668
rect 297950 619568 298074 619668
rect 298174 619568 298298 619668
rect 298398 619568 298522 619668
rect 298622 619568 298746 619668
rect 298846 619568 298880 619668
rect 297720 619444 298880 619568
rect 297720 619344 297850 619444
rect 297950 619344 298074 619444
rect 298174 619344 298298 619444
rect 298398 619344 298522 619444
rect 298622 619344 298746 619444
rect 298846 619344 298880 619444
rect 297720 619220 298880 619344
rect 297720 619120 297850 619220
rect 297950 619120 298074 619220
rect 298174 619120 298298 619220
rect 298398 619120 298522 619220
rect 298622 619120 298746 619220
rect 298846 619120 298880 619220
rect 297720 618996 298880 619120
rect 297720 618896 297850 618996
rect 297950 618896 298074 618996
rect 298174 618896 298298 618996
rect 298398 618896 298522 618996
rect 298622 618896 298746 618996
rect 298846 618896 298880 618996
rect 297720 618772 298880 618896
rect 297720 618672 297850 618772
rect 297950 618672 298074 618772
rect 298174 618672 298298 618772
rect 298398 618672 298522 618772
rect 298622 618672 298746 618772
rect 298846 618672 298880 618772
rect 297720 618548 298880 618672
rect 297720 618448 297850 618548
rect 297950 618448 298074 618548
rect 298174 618448 298298 618548
rect 298398 618448 298522 618548
rect 298622 618448 298746 618548
rect 298846 618448 298880 618548
rect 297720 618324 298880 618448
rect 297720 618224 297850 618324
rect 297950 618224 298074 618324
rect 298174 618224 298298 618324
rect 298398 618224 298522 618324
rect 298622 618224 298746 618324
rect 298846 618224 298880 618324
rect 297720 618100 298880 618224
rect 297720 618000 297850 618100
rect 297950 618000 298074 618100
rect 298174 618000 298298 618100
rect 298398 618000 298522 618100
rect 298622 618000 298746 618100
rect 298846 618000 298880 618100
rect 297720 617944 298880 618000
rect 304316 617068 311486 625300
rect 510594 624606 515394 631817
rect 342100 624600 343186 624606
rect 342000 624596 343186 624600
rect 342000 624496 342130 624596
rect 342230 624496 342354 624596
rect 342454 624496 342578 624596
rect 342678 624496 342802 624596
rect 342902 624496 343026 624596
rect 343126 624496 343186 624596
rect 342000 624372 343186 624496
rect 342000 624272 342130 624372
rect 342230 624272 342354 624372
rect 342454 624272 342578 624372
rect 342678 624272 342802 624372
rect 342902 624272 343026 624372
rect 343126 624272 343186 624372
rect 342000 624148 343186 624272
rect 342000 624048 342130 624148
rect 342230 624048 342354 624148
rect 342454 624048 342578 624148
rect 342678 624048 342802 624148
rect 342902 624048 343026 624148
rect 343126 624048 343186 624148
rect 342000 623924 343186 624048
rect 342000 623824 342130 623924
rect 342230 623824 342354 623924
rect 342454 623824 342578 623924
rect 342678 623824 342802 623924
rect 342902 623824 343026 623924
rect 343126 623824 343186 623924
rect 342000 623700 343186 623824
rect 342000 623600 342130 623700
rect 342230 623600 342354 623700
rect 342454 623600 342578 623700
rect 342678 623600 342802 623700
rect 342902 623600 343026 623700
rect 343126 623600 343186 623700
rect 342000 623476 343186 623600
rect 342000 623376 342130 623476
rect 342230 623376 342354 623476
rect 342454 623376 342578 623476
rect 342678 623376 342802 623476
rect 342902 623376 343026 623476
rect 343126 623376 343186 623476
rect 342000 623252 343186 623376
rect 342000 623152 342130 623252
rect 342230 623152 342354 623252
rect 342454 623152 342578 623252
rect 342678 623152 342802 623252
rect 342902 623152 343026 623252
rect 343126 623152 343186 623252
rect 342000 623028 343186 623152
rect 342000 622928 342130 623028
rect 342230 622928 342354 623028
rect 342454 622928 342578 623028
rect 342678 622928 342802 623028
rect 342902 622928 343026 623028
rect 343126 622928 343186 623028
rect 342000 622804 343186 622928
rect 342000 622704 342130 622804
rect 342230 622704 342354 622804
rect 342454 622704 342578 622804
rect 342678 622704 342802 622804
rect 342902 622704 343026 622804
rect 343126 622704 343186 622804
rect 342000 622580 343186 622704
rect 342000 622480 342130 622580
rect 342230 622480 342354 622580
rect 342454 622480 342578 622580
rect 342678 622480 342802 622580
rect 342902 622480 343026 622580
rect 343126 622480 343186 622580
rect 342000 622356 343186 622480
rect 342000 622256 342130 622356
rect 342230 622256 342354 622356
rect 342454 622256 342578 622356
rect 342678 622256 342802 622356
rect 342902 622256 343026 622356
rect 343126 622256 343186 622356
rect 342000 622132 343186 622256
rect 342000 622032 342130 622132
rect 342230 622032 342354 622132
rect 342454 622032 342578 622132
rect 342678 622032 342802 622132
rect 342902 622032 343026 622132
rect 343126 622032 343186 622132
rect 342000 621908 343186 622032
rect 342000 621808 342130 621908
rect 342230 621808 342354 621908
rect 342454 621808 342578 621908
rect 342678 621808 342802 621908
rect 342902 621808 343026 621908
rect 343126 621808 343186 621908
rect 342000 621684 343186 621808
rect 342000 621584 342130 621684
rect 342230 621584 342354 621684
rect 342454 621584 342578 621684
rect 342678 621584 342802 621684
rect 342902 621584 343026 621684
rect 343126 621584 343186 621684
rect 342000 621460 343186 621584
rect 342000 621360 342130 621460
rect 342230 621360 342354 621460
rect 342454 621360 342578 621460
rect 342678 621360 342802 621460
rect 342902 621360 343026 621460
rect 343126 621360 343186 621460
rect 342000 621236 343186 621360
rect 342000 621136 342130 621236
rect 342230 621136 342354 621236
rect 342454 621136 342578 621236
rect 342678 621136 342802 621236
rect 342902 621136 343026 621236
rect 343126 621136 343186 621236
rect 342000 621012 343186 621136
rect 342000 620912 342130 621012
rect 342230 620912 342354 621012
rect 342454 620912 342578 621012
rect 342678 620912 342802 621012
rect 342902 620912 343026 621012
rect 343126 620912 343186 621012
rect 342000 620788 343186 620912
rect 342000 620688 342130 620788
rect 342230 620688 342354 620788
rect 342454 620688 342578 620788
rect 342678 620688 342802 620788
rect 342902 620688 343026 620788
rect 343126 620688 343186 620788
rect 342000 620564 343186 620688
rect 342000 620464 342130 620564
rect 342230 620464 342354 620564
rect 342454 620464 342578 620564
rect 342678 620464 342802 620564
rect 342902 620464 343026 620564
rect 343126 620464 343186 620564
rect 342000 620340 343186 620464
rect 342000 620240 342130 620340
rect 342230 620240 342354 620340
rect 342454 620240 342578 620340
rect 342678 620240 342802 620340
rect 342902 620240 343026 620340
rect 343126 620240 343186 620340
rect 312075 620149 312715 620155
rect 312075 619869 312081 620149
rect 312709 619869 312715 620149
rect 312075 619863 312715 619869
rect 342000 620116 343186 620240
rect 342000 620016 342130 620116
rect 342230 620016 342354 620116
rect 342454 620016 342578 620116
rect 342678 620016 342802 620116
rect 342902 620016 343026 620116
rect 343126 620016 343186 620116
rect 342000 619892 343186 620016
rect 342000 619792 342130 619892
rect 342230 619792 342354 619892
rect 342454 619792 342578 619892
rect 342678 619792 342802 619892
rect 342902 619792 343026 619892
rect 343126 619792 343186 619892
rect 342000 619668 343186 619792
rect 342000 619568 342130 619668
rect 342230 619568 342354 619668
rect 342454 619568 342578 619668
rect 342678 619568 342802 619668
rect 342902 619568 343026 619668
rect 343126 619568 343186 619668
rect 342000 619444 343186 619568
rect 342000 619344 342130 619444
rect 342230 619344 342354 619444
rect 342454 619344 342578 619444
rect 342678 619344 342802 619444
rect 342902 619344 343026 619444
rect 343126 619344 343186 619444
rect 342000 619220 343186 619344
rect 342000 619120 342130 619220
rect 342230 619120 342354 619220
rect 342454 619120 342578 619220
rect 342678 619120 342802 619220
rect 342902 619120 343026 619220
rect 343126 619120 343186 619220
rect 342000 618996 343186 619120
rect 342000 618896 342130 618996
rect 342230 618896 342354 618996
rect 342454 618896 342578 618996
rect 342678 618896 342802 618996
rect 342902 618896 343026 618996
rect 343126 618896 343186 618996
rect 342000 618772 343186 618896
rect 342000 618672 342130 618772
rect 342230 618672 342354 618772
rect 342454 618672 342578 618772
rect 342678 618672 342802 618772
rect 342902 618672 343026 618772
rect 343126 618672 343186 618772
rect 342000 618548 343186 618672
rect 342000 618448 342130 618548
rect 342230 618448 342354 618548
rect 342454 618448 342578 618548
rect 342678 618448 342802 618548
rect 342902 618448 343026 618548
rect 343126 618448 343186 618548
rect 342000 618324 343186 618448
rect 342000 618224 342130 618324
rect 342230 618224 342354 618324
rect 342454 618224 342578 618324
rect 342678 618224 342802 618324
rect 342902 618224 343026 618324
rect 343126 618224 343186 618324
rect 342000 618100 343186 618224
rect 342000 618000 342130 618100
rect 342230 618000 342354 618100
rect 342454 618000 342578 618100
rect 342678 618000 342802 618100
rect 342902 618000 343026 618100
rect 343126 618000 343186 618100
rect 342000 617944 343186 618000
rect 510602 624161 515394 624606
rect 515386 618417 515394 624161
rect 510602 617944 515394 618417
rect 302938 617062 330669 617068
rect 302938 616948 302946 617062
rect 312192 616948 330669 617062
rect 301938 616846 330669 616948
rect 301938 616840 330670 616846
rect 301938 616830 330680 616840
rect 301938 616512 312710 616830
rect 330648 616512 330680 616830
rect 301938 616506 330680 616512
rect 304316 616472 311486 616506
rect 288920 605020 289920 610764
rect 294704 605020 295576 610764
rect 288920 604520 295576 605020
rect 298820 615474 315960 615520
rect 298820 615374 298876 615474
rect 298976 615374 299100 615474
rect 299200 615374 299324 615474
rect 299424 615374 299548 615474
rect 299648 615374 299772 615474
rect 299872 615374 299996 615474
rect 300096 615374 300220 615474
rect 300320 615374 300444 615474
rect 300544 615374 300668 615474
rect 300768 615374 300892 615474
rect 300992 615374 301116 615474
rect 301216 615374 301340 615474
rect 301440 615374 301564 615474
rect 301664 615374 301788 615474
rect 301888 615374 302012 615474
rect 302112 615374 302236 615474
rect 302336 615374 302460 615474
rect 302560 615374 302684 615474
rect 302784 615374 302908 615474
rect 303008 615374 303132 615474
rect 303232 615374 303356 615474
rect 303456 615374 303580 615474
rect 303680 615374 303804 615474
rect 303904 615374 304028 615474
rect 304128 615374 304252 615474
rect 304352 615374 304476 615474
rect 304576 615374 304700 615474
rect 304800 615374 304924 615474
rect 305024 615374 305148 615474
rect 305248 615374 305372 615474
rect 305472 615374 309346 615474
rect 309446 615374 309570 615474
rect 309670 615374 309794 615474
rect 309894 615374 310018 615474
rect 310118 615374 310242 615474
rect 310342 615374 310466 615474
rect 310566 615374 310690 615474
rect 310790 615374 310914 615474
rect 311014 615374 311138 615474
rect 311238 615374 311362 615474
rect 311462 615374 311586 615474
rect 311686 615374 311810 615474
rect 311910 615374 312034 615474
rect 312134 615374 312258 615474
rect 312358 615374 312482 615474
rect 312582 615374 312706 615474
rect 312806 615374 312930 615474
rect 313030 615374 313154 615474
rect 313254 615374 313378 615474
rect 313478 615374 313602 615474
rect 313702 615374 313826 615474
rect 313926 615374 314050 615474
rect 314150 615374 314274 615474
rect 314374 615374 314498 615474
rect 314598 615374 314722 615474
rect 314822 615374 314946 615474
rect 315046 615374 315170 615474
rect 315270 615374 315394 615474
rect 315494 615374 315618 615474
rect 315718 615374 315842 615474
rect 315942 615374 315960 615474
rect 298820 615250 315960 615374
rect 298820 615150 298876 615250
rect 298976 615150 299100 615250
rect 299200 615150 299324 615250
rect 299424 615150 299548 615250
rect 299648 615150 299772 615250
rect 299872 615150 299996 615250
rect 300096 615150 300220 615250
rect 300320 615150 300444 615250
rect 300544 615150 300668 615250
rect 300768 615150 300892 615250
rect 300992 615150 301116 615250
rect 301216 615150 301340 615250
rect 301440 615150 301564 615250
rect 301664 615150 301788 615250
rect 301888 615150 302012 615250
rect 302112 615150 302236 615250
rect 302336 615150 302460 615250
rect 302560 615150 302684 615250
rect 302784 615150 302908 615250
rect 303008 615150 303132 615250
rect 303232 615150 303356 615250
rect 303456 615150 303580 615250
rect 303680 615150 303804 615250
rect 303904 615150 304028 615250
rect 304128 615150 304252 615250
rect 304352 615150 304476 615250
rect 304576 615150 304700 615250
rect 304800 615150 304924 615250
rect 305024 615150 305148 615250
rect 305248 615150 305372 615250
rect 305472 615150 309346 615250
rect 309446 615150 309570 615250
rect 309670 615150 309794 615250
rect 309894 615150 310018 615250
rect 310118 615150 310242 615250
rect 310342 615150 310466 615250
rect 310566 615150 310690 615250
rect 310790 615150 310914 615250
rect 311014 615150 311138 615250
rect 311238 615150 311362 615250
rect 311462 615150 311586 615250
rect 311686 615150 311810 615250
rect 311910 615150 312034 615250
rect 312134 615150 312258 615250
rect 312358 615150 312482 615250
rect 312582 615150 312706 615250
rect 312806 615150 312930 615250
rect 313030 615150 313154 615250
rect 313254 615150 313378 615250
rect 313478 615150 313602 615250
rect 313702 615150 313826 615250
rect 313926 615150 314050 615250
rect 314150 615150 314274 615250
rect 314374 615150 314498 615250
rect 314598 615150 314722 615250
rect 314822 615150 314946 615250
rect 315046 615150 315170 615250
rect 315270 615150 315394 615250
rect 315494 615150 315618 615250
rect 315718 615150 315842 615250
rect 315942 615150 315960 615250
rect 298820 615026 315960 615150
rect 298820 614926 298876 615026
rect 298976 614926 299100 615026
rect 299200 614926 299324 615026
rect 299424 614926 299548 615026
rect 299648 614926 299772 615026
rect 299872 614926 299996 615026
rect 300096 614926 300220 615026
rect 300320 614926 300444 615026
rect 300544 614926 300668 615026
rect 300768 614926 300892 615026
rect 300992 614926 301116 615026
rect 301216 614926 301340 615026
rect 301440 614926 301564 615026
rect 301664 614926 301788 615026
rect 301888 614926 302012 615026
rect 302112 614926 302236 615026
rect 302336 614926 302460 615026
rect 302560 614926 302684 615026
rect 302784 614926 302908 615026
rect 303008 614926 303132 615026
rect 303232 614926 303356 615026
rect 303456 614926 303580 615026
rect 303680 614926 303804 615026
rect 303904 614926 304028 615026
rect 304128 614926 304252 615026
rect 304352 614926 304476 615026
rect 304576 614926 304700 615026
rect 304800 614926 304924 615026
rect 305024 614926 305148 615026
rect 305248 614926 305372 615026
rect 305472 614926 309346 615026
rect 309446 614926 309570 615026
rect 309670 614926 309794 615026
rect 309894 614926 310018 615026
rect 310118 614926 310242 615026
rect 310342 614926 310466 615026
rect 310566 614926 310690 615026
rect 310790 614926 310914 615026
rect 311014 614926 311138 615026
rect 311238 614926 311362 615026
rect 311462 614926 311586 615026
rect 311686 614926 311810 615026
rect 311910 614926 312034 615026
rect 312134 614926 312258 615026
rect 312358 614926 312482 615026
rect 312582 614926 312706 615026
rect 312806 614926 312930 615026
rect 313030 614926 313154 615026
rect 313254 614926 313378 615026
rect 313478 614926 313602 615026
rect 313702 614926 313826 615026
rect 313926 614926 314050 615026
rect 314150 614926 314274 615026
rect 314374 614926 314498 615026
rect 314598 614926 314722 615026
rect 314822 614926 314946 615026
rect 315046 614926 315170 615026
rect 315270 614926 315394 615026
rect 315494 614926 315618 615026
rect 315718 614926 315842 615026
rect 315942 614926 315960 615026
rect 298820 614802 315960 614926
rect 298820 614702 298876 614802
rect 298976 614702 299100 614802
rect 299200 614702 299324 614802
rect 299424 614702 299548 614802
rect 299648 614702 299772 614802
rect 299872 614702 299996 614802
rect 300096 614702 300220 614802
rect 300320 614702 300444 614802
rect 300544 614702 300668 614802
rect 300768 614702 300892 614802
rect 300992 614702 301116 614802
rect 301216 614702 301340 614802
rect 301440 614702 301564 614802
rect 301664 614702 301788 614802
rect 301888 614702 302012 614802
rect 302112 614702 302236 614802
rect 302336 614702 302460 614802
rect 302560 614702 302684 614802
rect 302784 614702 302908 614802
rect 303008 614702 303132 614802
rect 303232 614702 303356 614802
rect 303456 614702 303580 614802
rect 303680 614702 303804 614802
rect 303904 614702 304028 614802
rect 304128 614702 304252 614802
rect 304352 614702 304476 614802
rect 304576 614702 304700 614802
rect 304800 614702 304924 614802
rect 305024 614702 305148 614802
rect 305248 614702 305372 614802
rect 305472 614702 309346 614802
rect 309446 614702 309570 614802
rect 309670 614702 309794 614802
rect 309894 614702 310018 614802
rect 310118 614702 310242 614802
rect 310342 614702 310466 614802
rect 310566 614702 310690 614802
rect 310790 614702 310914 614802
rect 311014 614702 311138 614802
rect 311238 614702 311362 614802
rect 311462 614702 311586 614802
rect 311686 614702 311810 614802
rect 311910 614702 312034 614802
rect 312134 614702 312258 614802
rect 312358 614702 312482 614802
rect 312582 614702 312706 614802
rect 312806 614702 312930 614802
rect 313030 614702 313154 614802
rect 313254 614702 313378 614802
rect 313478 614702 313602 614802
rect 313702 614702 313826 614802
rect 313926 614702 314050 614802
rect 314150 614702 314274 614802
rect 314374 614702 314498 614802
rect 314598 614702 314722 614802
rect 314822 614702 314946 614802
rect 315046 614702 315170 614802
rect 315270 614702 315394 614802
rect 315494 614702 315618 614802
rect 315718 614702 315842 614802
rect 315942 614702 315960 614802
rect 298820 614578 315960 614702
rect 298820 614478 298876 614578
rect 298976 614478 299100 614578
rect 299200 614478 299324 614578
rect 299424 614478 299548 614578
rect 299648 614478 299772 614578
rect 299872 614478 299996 614578
rect 300096 614478 300220 614578
rect 300320 614478 300444 614578
rect 300544 614478 300668 614578
rect 300768 614478 300892 614578
rect 300992 614478 301116 614578
rect 301216 614478 301340 614578
rect 301440 614478 301564 614578
rect 301664 614478 301788 614578
rect 301888 614478 302012 614578
rect 302112 614478 302236 614578
rect 302336 614478 302460 614578
rect 302560 614478 302684 614578
rect 302784 614478 302908 614578
rect 303008 614478 303132 614578
rect 303232 614478 303356 614578
rect 303456 614478 303580 614578
rect 303680 614478 303804 614578
rect 303904 614478 304028 614578
rect 304128 614478 304252 614578
rect 304352 614478 304476 614578
rect 304576 614478 304700 614578
rect 304800 614478 304924 614578
rect 305024 614478 305148 614578
rect 305248 614478 305372 614578
rect 305472 614478 309346 614578
rect 309446 614478 309570 614578
rect 309670 614478 309794 614578
rect 309894 614478 310018 614578
rect 310118 614478 310242 614578
rect 310342 614478 310466 614578
rect 310566 614478 310690 614578
rect 310790 614478 310914 614578
rect 311014 614478 311138 614578
rect 311238 614478 311362 614578
rect 311462 614478 311586 614578
rect 311686 614478 311810 614578
rect 311910 614478 312034 614578
rect 312134 614478 312258 614578
rect 312358 614478 312482 614578
rect 312582 614478 312706 614578
rect 312806 614478 312930 614578
rect 313030 614478 313154 614578
rect 313254 614478 313378 614578
rect 313478 614478 313602 614578
rect 313702 614478 313826 614578
rect 313926 614478 314050 614578
rect 314150 614478 314274 614578
rect 314374 614478 314498 614578
rect 314598 614478 314722 614578
rect 314822 614478 314946 614578
rect 315046 614478 315170 614578
rect 315270 614478 315394 614578
rect 315494 614478 315618 614578
rect 315718 614478 315842 614578
rect 315942 614478 315960 614578
rect 298820 613100 315960 614478
rect 298820 611080 315980 613100
rect 298820 605336 298920 611080
rect 303704 605336 304920 611080
rect 309704 605336 310920 611080
rect 315704 605336 315980 611080
rect 298820 604520 315980 605336
rect 316960 597324 330680 616506
rect 335560 615494 342400 615540
rect 335560 615394 335616 615494
rect 335716 615394 335840 615494
rect 335940 615394 336064 615494
rect 336164 615394 336288 615494
rect 336388 615394 336512 615494
rect 336612 615394 336736 615494
rect 336836 615394 336960 615494
rect 337060 615394 337184 615494
rect 337284 615394 337408 615494
rect 337508 615394 337632 615494
rect 337732 615394 337856 615494
rect 337956 615394 338080 615494
rect 338180 615394 338304 615494
rect 338404 615394 338528 615494
rect 338628 615394 338752 615494
rect 338852 615394 338976 615494
rect 339076 615394 339200 615494
rect 339300 615394 339424 615494
rect 339524 615394 339648 615494
rect 339748 615394 339872 615494
rect 339972 615394 340096 615494
rect 340196 615394 340320 615494
rect 340420 615394 340544 615494
rect 340644 615394 340768 615494
rect 340868 615394 340992 615494
rect 341092 615394 341216 615494
rect 341316 615394 341440 615494
rect 341540 615394 341664 615494
rect 341764 615394 341888 615494
rect 341988 615394 342112 615494
rect 342212 615394 342400 615494
rect 335560 615270 342400 615394
rect 335560 615170 335616 615270
rect 335716 615170 335840 615270
rect 335940 615170 336064 615270
rect 336164 615170 336288 615270
rect 336388 615170 336512 615270
rect 336612 615170 336736 615270
rect 336836 615170 336960 615270
rect 337060 615170 337184 615270
rect 337284 615170 337408 615270
rect 337508 615170 337632 615270
rect 337732 615170 337856 615270
rect 337956 615170 338080 615270
rect 338180 615170 338304 615270
rect 338404 615170 338528 615270
rect 338628 615170 338752 615270
rect 338852 615170 338976 615270
rect 339076 615170 339200 615270
rect 339300 615170 339424 615270
rect 339524 615170 339648 615270
rect 339748 615170 339872 615270
rect 339972 615170 340096 615270
rect 340196 615170 340320 615270
rect 340420 615170 340544 615270
rect 340644 615170 340768 615270
rect 340868 615170 340992 615270
rect 341092 615170 341216 615270
rect 341316 615170 341440 615270
rect 341540 615170 341664 615270
rect 341764 615170 341888 615270
rect 341988 615170 342112 615270
rect 342212 615170 342400 615270
rect 335560 615046 342400 615170
rect 335560 614946 335616 615046
rect 335716 614946 335840 615046
rect 335940 614946 336064 615046
rect 336164 614946 336288 615046
rect 336388 614946 336512 615046
rect 336612 614946 336736 615046
rect 336836 614946 336960 615046
rect 337060 614946 337184 615046
rect 337284 614946 337408 615046
rect 337508 614946 337632 615046
rect 337732 614946 337856 615046
rect 337956 614946 338080 615046
rect 338180 614946 338304 615046
rect 338404 614946 338528 615046
rect 338628 614946 338752 615046
rect 338852 614946 338976 615046
rect 339076 614946 339200 615046
rect 339300 614946 339424 615046
rect 339524 614946 339648 615046
rect 339748 614946 339872 615046
rect 339972 614946 340096 615046
rect 340196 614946 340320 615046
rect 340420 614946 340544 615046
rect 340644 614946 340768 615046
rect 340868 614946 340992 615046
rect 341092 614946 341216 615046
rect 341316 614946 341440 615046
rect 341540 614946 341664 615046
rect 341764 614946 341888 615046
rect 341988 614946 342112 615046
rect 342212 614946 342400 615046
rect 335560 614822 342400 614946
rect 335560 614722 335616 614822
rect 335716 614722 335840 614822
rect 335940 614722 336064 614822
rect 336164 614722 336288 614822
rect 336388 614722 336512 614822
rect 336612 614722 336736 614822
rect 336836 614722 336960 614822
rect 337060 614722 337184 614822
rect 337284 614722 337408 614822
rect 337508 614722 337632 614822
rect 337732 614722 337856 614822
rect 337956 614722 338080 614822
rect 338180 614722 338304 614822
rect 338404 614722 338528 614822
rect 338628 614722 338752 614822
rect 338852 614722 338976 614822
rect 339076 614722 339200 614822
rect 339300 614722 339424 614822
rect 339524 614722 339648 614822
rect 339748 614722 339872 614822
rect 339972 614722 340096 614822
rect 340196 614722 340320 614822
rect 340420 614722 340544 614822
rect 340644 614722 340768 614822
rect 340868 614722 340992 614822
rect 341092 614722 341216 614822
rect 341316 614722 341440 614822
rect 341540 614722 341664 614822
rect 341764 614722 341888 614822
rect 341988 614722 342112 614822
rect 342212 614722 342400 614822
rect 335560 614598 342400 614722
rect 335560 614498 335616 614598
rect 335716 614498 335840 614598
rect 335940 614498 336064 614598
rect 336164 614498 336288 614598
rect 336388 614498 336512 614598
rect 336612 614498 336736 614598
rect 336836 614498 336960 614598
rect 337060 614498 337184 614598
rect 337284 614498 337408 614598
rect 337508 614498 337632 614598
rect 337732 614498 337856 614598
rect 337956 614498 338080 614598
rect 338180 614498 338304 614598
rect 338404 614498 338528 614598
rect 338628 614498 338752 614598
rect 338852 614498 338976 614598
rect 339076 614498 339200 614598
rect 339300 614498 339424 614598
rect 339524 614498 339648 614598
rect 339748 614498 339872 614598
rect 339972 614498 340096 614598
rect 340196 614498 340320 614598
rect 340420 614498 340544 614598
rect 340644 614498 340768 614598
rect 340868 614498 340992 614598
rect 341092 614498 341216 614598
rect 341316 614498 341440 614598
rect 341540 614498 341664 614598
rect 341764 614498 341888 614598
rect 341988 614498 342112 614598
rect 342212 614498 342400 614598
rect 335560 614464 342400 614498
rect 335580 611084 342400 614464
rect 510594 611200 515394 617944
rect 335580 605340 336480 611084
rect 341264 605340 342400 611084
rect 335580 604720 342400 605340
rect 510602 610761 515394 611200
rect 515386 605017 515394 610761
rect 510602 604544 515394 605017
rect 520594 690560 525394 704800
rect 566594 702300 571594 704800
rect 520594 684336 520602 690560
rect 525386 684336 525394 690560
rect 520594 650961 525394 684336
rect 582300 677984 584800 682984
rect 520594 645217 520602 650961
rect 525386 645217 525394 650961
rect 520594 637561 525394 645217
rect 560050 644576 584800 644584
rect 560050 639792 560582 644576
rect 566726 639792 584800 644576
rect 560050 639784 584800 639792
rect 520594 631817 520602 637561
rect 525386 631817 525394 637561
rect 520594 624161 525394 631817
rect 560050 634576 584800 634584
rect 560050 629792 560582 634576
rect 566726 629792 584800 634576
rect 560050 629784 584800 629792
rect 520594 618417 520602 624161
rect 525386 618417 525394 624161
rect 520594 610761 525394 618417
rect 520594 605017 520602 610761
rect 525386 605017 525394 610761
rect 520594 604544 525394 605017
rect 316960 591580 317480 597324
rect 322264 591580 325480 597324
rect 330264 591580 330680 597324
rect 316960 591080 330680 591580
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 339960 511642 340072 571500
rect -800 511530 340072 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect 340967 463692 341079 571500
rect -800 463580 341079 463692
rect -800 462486 17711 462510
rect -800 462422 13897 462486
rect 13961 462422 13977 462486
rect 14041 462422 14057 462486
rect 14121 462422 14137 462486
rect 14201 462422 14217 462486
rect 14281 462422 14297 462486
rect 14361 462422 14377 462486
rect 14441 462422 14457 462486
rect 14521 462422 14537 462486
rect 14601 462422 14617 462486
rect 14681 462422 14697 462486
rect 14761 462422 14777 462486
rect 14841 462422 14857 462486
rect 14921 462422 14937 462486
rect 15001 462422 15017 462486
rect 15081 462422 15097 462486
rect 15161 462422 15177 462486
rect 15241 462422 15257 462486
rect 15321 462422 15337 462486
rect 15401 462422 15417 462486
rect 15481 462422 15497 462486
rect 15561 462422 15577 462486
rect 15641 462422 15657 462486
rect 15721 462422 15737 462486
rect 15801 462422 15817 462486
rect 15881 462422 15897 462486
rect 15961 462422 15977 462486
rect 16041 462422 16057 462486
rect 16121 462422 16137 462486
rect 16201 462422 16217 462486
rect 16281 462422 16297 462486
rect 16361 462422 16377 462486
rect 16441 462422 16457 462486
rect 16521 462422 16537 462486
rect 16601 462422 16617 462486
rect 16681 462422 16697 462486
rect 16761 462422 16777 462486
rect 16841 462422 16857 462486
rect 16921 462422 16937 462486
rect 17001 462422 17017 462486
rect 17081 462422 17097 462486
rect 17161 462422 17177 462486
rect 17241 462422 17257 462486
rect 17321 462422 17337 462486
rect 17401 462422 17417 462486
rect 17481 462422 17497 462486
rect 17561 462422 17711 462486
rect -800 462398 17711 462422
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect 341738 420470 341850 571500
rect -800 420358 341850 420470
rect -800 419264 17694 419288
rect -800 419200 13911 419264
rect 13975 419200 13991 419264
rect 14055 419200 14071 419264
rect 14135 419200 14151 419264
rect 14215 419200 14231 419264
rect 14295 419200 14311 419264
rect 14375 419200 14391 419264
rect 14455 419200 14471 419264
rect 14535 419200 14551 419264
rect 14615 419200 14631 419264
rect 14695 419200 14711 419264
rect 14775 419200 14791 419264
rect 14855 419200 14871 419264
rect 14935 419200 14951 419264
rect 15015 419200 15031 419264
rect 15095 419200 15111 419264
rect 15175 419200 15191 419264
rect 15255 419200 15271 419264
rect 15335 419200 15351 419264
rect 15415 419200 15431 419264
rect 15495 419200 15511 419264
rect 15575 419200 15591 419264
rect 15655 419200 15671 419264
rect 15735 419200 15751 419264
rect 15815 419200 15831 419264
rect 15895 419200 15911 419264
rect 15975 419200 15991 419264
rect 16055 419200 16071 419264
rect 16135 419200 16151 419264
rect 16215 419200 16231 419264
rect 16295 419200 16311 419264
rect 16375 419200 16391 419264
rect 16455 419200 16471 419264
rect 16535 419200 16551 419264
rect 16615 419200 16631 419264
rect 16695 419200 16711 419264
rect 16775 419200 16791 419264
rect 16855 419200 16871 419264
rect 16935 419200 16951 419264
rect 17015 419200 17031 419264
rect 17095 419200 17111 419264
rect 17175 419200 17191 419264
rect 17255 419200 17271 419264
rect 17335 419200 17351 419264
rect 17415 419200 17431 419264
rect 17495 419200 17511 419264
rect 17575 419200 17694 419264
rect -800 419176 17694 419200
rect 533497 405408 533609 573580
rect 537376 454558 537488 573580
rect 539494 498980 539606 573580
rect 555452 555354 584800 555362
rect 555452 550570 556255 555354
rect 562319 550570 584800 555354
rect 555452 550562 584800 550570
rect 555452 545354 584800 545362
rect 555452 540570 556255 545354
rect 562319 540570 584800 545354
rect 555452 540562 584800 540570
rect 573371 500138 584800 500162
rect 573371 500074 573553 500138
rect 573617 500074 573633 500138
rect 573697 500074 573713 500138
rect 573777 500074 573793 500138
rect 573857 500074 573873 500138
rect 573937 500074 573953 500138
rect 574017 500074 574033 500138
rect 574097 500074 574113 500138
rect 574177 500074 574193 500138
rect 574257 500074 574273 500138
rect 574337 500074 574353 500138
rect 574417 500074 574433 500138
rect 574497 500074 574513 500138
rect 574577 500074 574593 500138
rect 574657 500074 574673 500138
rect 574737 500074 574753 500138
rect 574817 500074 574833 500138
rect 574897 500074 574913 500138
rect 574977 500074 574993 500138
rect 575057 500074 575073 500138
rect 575137 500074 575153 500138
rect 575217 500074 575233 500138
rect 575297 500074 575313 500138
rect 575377 500074 575393 500138
rect 575457 500074 575473 500138
rect 575537 500074 575553 500138
rect 575617 500074 575633 500138
rect 575697 500074 575713 500138
rect 575777 500074 575793 500138
rect 575857 500074 575873 500138
rect 575937 500074 575953 500138
rect 576017 500074 576033 500138
rect 576097 500074 576113 500138
rect 576177 500074 576193 500138
rect 576257 500074 576273 500138
rect 576337 500074 576353 500138
rect 576417 500074 576433 500138
rect 576497 500074 576513 500138
rect 576577 500074 576593 500138
rect 576657 500074 576673 500138
rect 576737 500074 584800 500138
rect 573371 500050 584800 500074
rect 539494 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 573405 455716 584800 455740
rect 573405 455652 573591 455716
rect 573655 455652 573671 455716
rect 573735 455652 573751 455716
rect 573815 455652 573831 455716
rect 573895 455652 573911 455716
rect 573975 455652 573991 455716
rect 574055 455652 574071 455716
rect 574135 455652 574151 455716
rect 574215 455652 574231 455716
rect 574295 455652 574311 455716
rect 574375 455652 574391 455716
rect 574455 455652 574471 455716
rect 574535 455652 574551 455716
rect 574615 455652 574631 455716
rect 574695 455652 574711 455716
rect 574775 455652 574791 455716
rect 574855 455652 574871 455716
rect 574935 455652 574951 455716
rect 575015 455652 575031 455716
rect 575095 455652 575111 455716
rect 575175 455652 575191 455716
rect 575255 455652 575271 455716
rect 575335 455652 575351 455716
rect 575415 455652 575431 455716
rect 575495 455652 575511 455716
rect 575575 455652 575591 455716
rect 575655 455652 575671 455716
rect 575735 455652 575751 455716
rect 575815 455652 575831 455716
rect 575895 455652 575911 455716
rect 575975 455652 575991 455716
rect 576055 455652 576071 455716
rect 576135 455652 576151 455716
rect 576215 455652 576231 455716
rect 576295 455652 576311 455716
rect 576375 455652 576391 455716
rect 576455 455652 576471 455716
rect 576535 455652 576551 455716
rect 576615 455652 576631 455716
rect 576695 455652 584800 455716
rect 573405 455628 584800 455652
rect 537376 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 533497 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 13406 196222 584800 196230
rect 13406 191438 13997 196222
rect 17421 191438 573605 196222
rect 576629 191438 584800 196222
rect 13406 191430 584800 191438
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 170922 684353 173066 690577
rect 173422 684353 175566 690577
rect 222622 684386 224766 690610
rect 217344 626112 217408 626176
rect 217472 626112 217536 626176
rect 217600 626112 217664 626176
rect 217728 626112 217792 626176
rect 217856 626112 217920 626176
rect 217984 626112 218048 626176
rect 218112 626112 218176 626176
rect 218240 626112 218304 626176
rect 218368 626112 218432 626176
rect 218496 626112 218560 626176
rect 218624 626112 218688 626176
rect 218752 626112 218816 626176
rect 218880 626112 218944 626176
rect 219008 626112 219072 626176
rect 219136 626112 219200 626176
rect 219264 626112 219328 626176
rect 219392 626112 219456 626176
rect 219520 626112 219584 626176
rect 219648 626112 219712 626176
rect 219776 626112 219840 626176
rect 219904 626112 219968 626176
rect 220032 626112 220096 626176
rect 220160 626112 220224 626176
rect 220288 626112 220352 626176
rect 220416 626112 220480 626176
rect 220544 626112 220608 626176
rect 220672 626112 220736 626176
rect 220800 626112 220864 626176
rect 220928 626112 220992 626176
rect 221056 626112 221120 626176
rect 221184 626112 221248 626176
rect 221312 626112 221376 626176
rect 221440 626112 221504 626176
rect 221568 626112 221632 626176
rect 221696 626112 221760 626176
rect 221824 626112 221888 626176
rect 221952 626112 222016 626176
rect 222080 626112 222144 626176
rect 217344 625984 217408 626048
rect 217472 625984 217536 626048
rect 217600 625984 217664 626048
rect 217728 625984 217792 626048
rect 217856 625984 217920 626048
rect 217984 625984 218048 626048
rect 218112 625984 218176 626048
rect 218240 625984 218304 626048
rect 218368 625984 218432 626048
rect 218496 625984 218560 626048
rect 218624 625984 218688 626048
rect 218752 625984 218816 626048
rect 218880 625984 218944 626048
rect 219008 625984 219072 626048
rect 219136 625984 219200 626048
rect 219264 625984 219328 626048
rect 219392 625984 219456 626048
rect 219520 625984 219584 626048
rect 219648 625984 219712 626048
rect 219776 625984 219840 626048
rect 219904 625984 219968 626048
rect 220032 625984 220096 626048
rect 220160 625984 220224 626048
rect 220288 625984 220352 626048
rect 220416 625984 220480 626048
rect 220544 625984 220608 626048
rect 220672 625984 220736 626048
rect 220800 625984 220864 626048
rect 220928 625984 220992 626048
rect 221056 625984 221120 626048
rect 221184 625984 221248 626048
rect 221312 625984 221376 626048
rect 221440 625984 221504 626048
rect 221568 625984 221632 626048
rect 221696 625984 221760 626048
rect 221824 625984 221888 626048
rect 221952 625984 222016 626048
rect 222080 625984 222144 626048
rect 217344 625856 217408 625920
rect 217472 625856 217536 625920
rect 217600 625856 217664 625920
rect 217728 625856 217792 625920
rect 217856 625856 217920 625920
rect 217984 625856 218048 625920
rect 218112 625856 218176 625920
rect 218240 625856 218304 625920
rect 218368 625856 218432 625920
rect 218496 625856 218560 625920
rect 218624 625856 218688 625920
rect 218752 625856 218816 625920
rect 218880 625856 218944 625920
rect 219008 625856 219072 625920
rect 219136 625856 219200 625920
rect 219264 625856 219328 625920
rect 219392 625856 219456 625920
rect 219520 625856 219584 625920
rect 219648 625856 219712 625920
rect 219776 625856 219840 625920
rect 219904 625856 219968 625920
rect 220032 625856 220096 625920
rect 220160 625856 220224 625920
rect 220288 625856 220352 625920
rect 220416 625856 220480 625920
rect 220544 625856 220608 625920
rect 220672 625856 220736 625920
rect 220800 625856 220864 625920
rect 220928 625856 220992 625920
rect 221056 625856 221120 625920
rect 221184 625856 221248 625920
rect 221312 625856 221376 625920
rect 221440 625856 221504 625920
rect 221568 625856 221632 625920
rect 221696 625856 221760 625920
rect 221824 625856 221888 625920
rect 221952 625856 222016 625920
rect 222080 625856 222144 625920
rect 217344 625728 217408 625792
rect 217472 625728 217536 625792
rect 217600 625728 217664 625792
rect 217728 625728 217792 625792
rect 217856 625728 217920 625792
rect 217984 625728 218048 625792
rect 218112 625728 218176 625792
rect 218240 625728 218304 625792
rect 218368 625728 218432 625792
rect 218496 625728 218560 625792
rect 218624 625728 218688 625792
rect 218752 625728 218816 625792
rect 218880 625728 218944 625792
rect 219008 625728 219072 625792
rect 219136 625728 219200 625792
rect 219264 625728 219328 625792
rect 219392 625728 219456 625792
rect 219520 625728 219584 625792
rect 219648 625728 219712 625792
rect 219776 625728 219840 625792
rect 219904 625728 219968 625792
rect 220032 625728 220096 625792
rect 220160 625728 220224 625792
rect 220288 625728 220352 625792
rect 220416 625728 220480 625792
rect 220544 625728 220608 625792
rect 220672 625728 220736 625792
rect 220800 625728 220864 625792
rect 220928 625728 220992 625792
rect 221056 625728 221120 625792
rect 221184 625728 221248 625792
rect 221312 625728 221376 625792
rect 221440 625728 221504 625792
rect 221568 625728 221632 625792
rect 221696 625728 221760 625792
rect 221824 625728 221888 625792
rect 221952 625728 222016 625792
rect 222080 625728 222144 625792
rect 227640 626112 227704 626176
rect 227768 626112 227832 626176
rect 227896 626112 227960 626176
rect 228024 626112 228088 626176
rect 228152 626112 228216 626176
rect 228280 626112 228344 626176
rect 228408 626112 228472 626176
rect 228536 626112 228600 626176
rect 228664 626112 228728 626176
rect 228792 626112 228856 626176
rect 228920 626112 228984 626176
rect 229048 626112 229112 626176
rect 229176 626112 229240 626176
rect 229304 626112 229368 626176
rect 229432 626112 229496 626176
rect 229560 626112 229624 626176
rect 229688 626112 229752 626176
rect 229816 626112 229880 626176
rect 229944 626112 230008 626176
rect 230072 626112 230136 626176
rect 230200 626112 230264 626176
rect 230328 626112 230392 626176
rect 230456 626112 230520 626176
rect 230584 626112 230648 626176
rect 230712 626112 230776 626176
rect 230840 626112 230904 626176
rect 230968 626112 231032 626176
rect 231096 626112 231160 626176
rect 231224 626112 231288 626176
rect 231352 626112 231416 626176
rect 231480 626112 231544 626176
rect 231608 626112 231672 626176
rect 231736 626112 231800 626176
rect 231864 626112 231928 626176
rect 231992 626112 232056 626176
rect 232120 626112 232184 626176
rect 232248 626112 232312 626176
rect 232376 626112 232440 626176
rect 227640 625984 227704 626048
rect 227768 625984 227832 626048
rect 227896 625984 227960 626048
rect 228024 625984 228088 626048
rect 228152 625984 228216 626048
rect 228280 625984 228344 626048
rect 228408 625984 228472 626048
rect 228536 625984 228600 626048
rect 228664 625984 228728 626048
rect 228792 625984 228856 626048
rect 228920 625984 228984 626048
rect 229048 625984 229112 626048
rect 229176 625984 229240 626048
rect 229304 625984 229368 626048
rect 229432 625984 229496 626048
rect 229560 625984 229624 626048
rect 229688 625984 229752 626048
rect 229816 625984 229880 626048
rect 229944 625984 230008 626048
rect 230072 625984 230136 626048
rect 230200 625984 230264 626048
rect 230328 625984 230392 626048
rect 230456 625984 230520 626048
rect 230584 625984 230648 626048
rect 230712 625984 230776 626048
rect 230840 625984 230904 626048
rect 230968 625984 231032 626048
rect 231096 625984 231160 626048
rect 231224 625984 231288 626048
rect 231352 625984 231416 626048
rect 231480 625984 231544 626048
rect 231608 625984 231672 626048
rect 231736 625984 231800 626048
rect 231864 625984 231928 626048
rect 231992 625984 232056 626048
rect 232120 625984 232184 626048
rect 232248 625984 232312 626048
rect 232376 625984 232440 626048
rect 227640 625856 227704 625920
rect 227768 625856 227832 625920
rect 227896 625856 227960 625920
rect 228024 625856 228088 625920
rect 228152 625856 228216 625920
rect 228280 625856 228344 625920
rect 228408 625856 228472 625920
rect 228536 625856 228600 625920
rect 228664 625856 228728 625920
rect 228792 625856 228856 625920
rect 228920 625856 228984 625920
rect 229048 625856 229112 625920
rect 229176 625856 229240 625920
rect 229304 625856 229368 625920
rect 229432 625856 229496 625920
rect 229560 625856 229624 625920
rect 229688 625856 229752 625920
rect 229816 625856 229880 625920
rect 229944 625856 230008 625920
rect 230072 625856 230136 625920
rect 230200 625856 230264 625920
rect 230328 625856 230392 625920
rect 230456 625856 230520 625920
rect 230584 625856 230648 625920
rect 230712 625856 230776 625920
rect 230840 625856 230904 625920
rect 230968 625856 231032 625920
rect 231096 625856 231160 625920
rect 231224 625856 231288 625920
rect 231352 625856 231416 625920
rect 231480 625856 231544 625920
rect 231608 625856 231672 625920
rect 231736 625856 231800 625920
rect 231864 625856 231928 625920
rect 231992 625856 232056 625920
rect 232120 625856 232184 625920
rect 232248 625856 232312 625920
rect 232376 625856 232440 625920
rect 227640 625728 227704 625792
rect 227768 625728 227832 625792
rect 227896 625728 227960 625792
rect 228024 625728 228088 625792
rect 228152 625728 228216 625792
rect 228280 625728 228344 625792
rect 228408 625728 228472 625792
rect 228536 625728 228600 625792
rect 228664 625728 228728 625792
rect 228792 625728 228856 625792
rect 228920 625728 228984 625792
rect 229048 625728 229112 625792
rect 229176 625728 229240 625792
rect 229304 625728 229368 625792
rect 229432 625728 229496 625792
rect 229560 625728 229624 625792
rect 229688 625728 229752 625792
rect 229816 625728 229880 625792
rect 229944 625728 230008 625792
rect 230072 625728 230136 625792
rect 230200 625728 230264 625792
rect 230328 625728 230392 625792
rect 230456 625728 230520 625792
rect 230584 625728 230648 625792
rect 230712 625728 230776 625792
rect 230840 625728 230904 625792
rect 230968 625728 231032 625792
rect 231096 625728 231160 625792
rect 231224 625728 231288 625792
rect 231352 625728 231416 625792
rect 231480 625728 231544 625792
rect 231608 625728 231672 625792
rect 231736 625728 231800 625792
rect 231864 625728 231928 625792
rect 231992 625728 232056 625792
rect 232120 625728 232184 625792
rect 232248 625728 232312 625792
rect 232376 625728 232440 625792
rect 289800 684340 294584 690084
rect 324322 684369 326466 690593
rect 510602 684336 515386 690560
rect 289920 644840 294704 650584
rect 298920 644840 303704 650584
rect 304920 644840 309704 650584
rect 310920 644840 315704 650584
rect 298876 642594 298976 642694
rect 299100 642594 299200 642694
rect 299324 642594 299424 642694
rect 299548 642594 299648 642694
rect 299772 642594 299872 642694
rect 299996 642594 300096 642694
rect 300220 642594 300320 642694
rect 300444 642594 300544 642694
rect 300668 642594 300768 642694
rect 300892 642594 300992 642694
rect 301116 642594 301216 642694
rect 301340 642594 301440 642694
rect 301564 642594 301664 642694
rect 301788 642594 301888 642694
rect 302012 642594 302112 642694
rect 302236 642594 302336 642694
rect 302460 642594 302560 642694
rect 302684 642594 302784 642694
rect 302908 642594 303008 642694
rect 303132 642594 303232 642694
rect 303356 642594 303456 642694
rect 303580 642594 303680 642694
rect 303804 642594 303904 642694
rect 304028 642594 304128 642694
rect 304252 642594 304352 642694
rect 304476 642594 304576 642694
rect 304700 642594 304800 642694
rect 304924 642594 305024 642694
rect 305148 642594 305248 642694
rect 305372 642594 305472 642694
rect 309346 642594 309446 642694
rect 309570 642594 309670 642694
rect 309794 642594 309894 642694
rect 310018 642594 310118 642694
rect 310242 642594 310342 642694
rect 310466 642594 310566 642694
rect 310690 642594 310790 642694
rect 310914 642594 311014 642694
rect 311138 642594 311238 642694
rect 311362 642594 311462 642694
rect 311586 642594 311686 642694
rect 311810 642594 311910 642694
rect 312034 642594 312134 642694
rect 312258 642594 312358 642694
rect 312482 642594 312582 642694
rect 312706 642594 312806 642694
rect 312930 642594 313030 642694
rect 313154 642594 313254 642694
rect 313378 642594 313478 642694
rect 313602 642594 313702 642694
rect 313826 642594 313926 642694
rect 314050 642594 314150 642694
rect 314274 642594 314374 642694
rect 314498 642594 314598 642694
rect 314722 642594 314822 642694
rect 314946 642594 315046 642694
rect 315170 642594 315270 642694
rect 315394 642594 315494 642694
rect 315618 642594 315718 642694
rect 315842 642594 315942 642694
rect 298876 642370 298976 642470
rect 299100 642370 299200 642470
rect 299324 642370 299424 642470
rect 299548 642370 299648 642470
rect 299772 642370 299872 642470
rect 299996 642370 300096 642470
rect 300220 642370 300320 642470
rect 300444 642370 300544 642470
rect 300668 642370 300768 642470
rect 300892 642370 300992 642470
rect 301116 642370 301216 642470
rect 301340 642370 301440 642470
rect 301564 642370 301664 642470
rect 301788 642370 301888 642470
rect 302012 642370 302112 642470
rect 302236 642370 302336 642470
rect 302460 642370 302560 642470
rect 302684 642370 302784 642470
rect 302908 642370 303008 642470
rect 303132 642370 303232 642470
rect 303356 642370 303456 642470
rect 303580 642370 303680 642470
rect 303804 642370 303904 642470
rect 304028 642370 304128 642470
rect 304252 642370 304352 642470
rect 304476 642370 304576 642470
rect 304700 642370 304800 642470
rect 304924 642370 305024 642470
rect 305148 642370 305248 642470
rect 305372 642370 305472 642470
rect 309346 642370 309446 642470
rect 309570 642370 309670 642470
rect 309794 642370 309894 642470
rect 310018 642370 310118 642470
rect 310242 642370 310342 642470
rect 310466 642370 310566 642470
rect 310690 642370 310790 642470
rect 310914 642370 311014 642470
rect 311138 642370 311238 642470
rect 311362 642370 311462 642470
rect 311586 642370 311686 642470
rect 311810 642370 311910 642470
rect 312034 642370 312134 642470
rect 312258 642370 312358 642470
rect 312482 642370 312582 642470
rect 312706 642370 312806 642470
rect 312930 642370 313030 642470
rect 313154 642370 313254 642470
rect 313378 642370 313478 642470
rect 313602 642370 313702 642470
rect 313826 642370 313926 642470
rect 314050 642370 314150 642470
rect 314274 642370 314374 642470
rect 314498 642370 314598 642470
rect 314722 642370 314822 642470
rect 314946 642370 315046 642470
rect 315170 642370 315270 642470
rect 315394 642370 315494 642470
rect 315618 642370 315718 642470
rect 315842 642370 315942 642470
rect 298876 642146 298976 642246
rect 299100 642146 299200 642246
rect 299324 642146 299424 642246
rect 299548 642146 299648 642246
rect 299772 642146 299872 642246
rect 299996 642146 300096 642246
rect 300220 642146 300320 642246
rect 300444 642146 300544 642246
rect 300668 642146 300768 642246
rect 300892 642146 300992 642246
rect 301116 642146 301216 642246
rect 301340 642146 301440 642246
rect 301564 642146 301664 642246
rect 301788 642146 301888 642246
rect 302012 642146 302112 642246
rect 302236 642146 302336 642246
rect 302460 642146 302560 642246
rect 302684 642146 302784 642246
rect 302908 642146 303008 642246
rect 303132 642146 303232 642246
rect 303356 642146 303456 642246
rect 303580 642146 303680 642246
rect 303804 642146 303904 642246
rect 304028 642146 304128 642246
rect 304252 642146 304352 642246
rect 304476 642146 304576 642246
rect 304700 642146 304800 642246
rect 304924 642146 305024 642246
rect 305148 642146 305248 642246
rect 305372 642146 305472 642246
rect 309346 642146 309446 642246
rect 309570 642146 309670 642246
rect 309794 642146 309894 642246
rect 310018 642146 310118 642246
rect 310242 642146 310342 642246
rect 310466 642146 310566 642246
rect 310690 642146 310790 642246
rect 310914 642146 311014 642246
rect 311138 642146 311238 642246
rect 311362 642146 311462 642246
rect 311586 642146 311686 642246
rect 311810 642146 311910 642246
rect 312034 642146 312134 642246
rect 312258 642146 312358 642246
rect 312482 642146 312582 642246
rect 312706 642146 312806 642246
rect 312930 642146 313030 642246
rect 313154 642146 313254 642246
rect 313378 642146 313478 642246
rect 313602 642146 313702 642246
rect 313826 642146 313926 642246
rect 314050 642146 314150 642246
rect 314274 642146 314374 642246
rect 314498 642146 314598 642246
rect 314722 642146 314822 642246
rect 314946 642146 315046 642246
rect 315170 642146 315270 642246
rect 315394 642146 315494 642246
rect 315618 642146 315718 642246
rect 315842 642146 315942 642246
rect 298876 641922 298976 642022
rect 299100 641922 299200 642022
rect 299324 641922 299424 642022
rect 299548 641922 299648 642022
rect 299772 641922 299872 642022
rect 299996 641922 300096 642022
rect 300220 641922 300320 642022
rect 300444 641922 300544 642022
rect 300668 641922 300768 642022
rect 300892 641922 300992 642022
rect 301116 641922 301216 642022
rect 301340 641922 301440 642022
rect 301564 641922 301664 642022
rect 301788 641922 301888 642022
rect 302012 641922 302112 642022
rect 302236 641922 302336 642022
rect 302460 641922 302560 642022
rect 302684 641922 302784 642022
rect 302908 641922 303008 642022
rect 303132 641922 303232 642022
rect 303356 641922 303456 642022
rect 303580 641922 303680 642022
rect 303804 641922 303904 642022
rect 304028 641922 304128 642022
rect 304252 641922 304352 642022
rect 304476 641922 304576 642022
rect 304700 641922 304800 642022
rect 304924 641922 305024 642022
rect 305148 641922 305248 642022
rect 305372 641922 305472 642022
rect 309346 641922 309446 642022
rect 309570 641922 309670 642022
rect 309794 641922 309894 642022
rect 310018 641922 310118 642022
rect 310242 641922 310342 642022
rect 310466 641922 310566 642022
rect 310690 641922 310790 642022
rect 310914 641922 311014 642022
rect 311138 641922 311238 642022
rect 311362 641922 311462 642022
rect 311586 641922 311686 642022
rect 311810 641922 311910 642022
rect 312034 641922 312134 642022
rect 312258 641922 312358 642022
rect 312482 641922 312582 642022
rect 312706 641922 312806 642022
rect 312930 641922 313030 642022
rect 313154 641922 313254 642022
rect 313378 641922 313478 642022
rect 313602 641922 313702 642022
rect 313826 641922 313926 642022
rect 314050 641922 314150 642022
rect 314274 641922 314374 642022
rect 314498 641922 314598 642022
rect 314722 641922 314822 642022
rect 314946 641922 315046 642022
rect 315170 641922 315270 642022
rect 315394 641922 315494 642022
rect 315618 641922 315718 642022
rect 315842 641922 315942 642022
rect 298876 641698 298976 641798
rect 299100 641698 299200 641798
rect 299324 641698 299424 641798
rect 299548 641698 299648 641798
rect 299772 641698 299872 641798
rect 299996 641698 300096 641798
rect 300220 641698 300320 641798
rect 300444 641698 300544 641798
rect 300668 641698 300768 641798
rect 300892 641698 300992 641798
rect 301116 641698 301216 641798
rect 301340 641698 301440 641798
rect 301564 641698 301664 641798
rect 301788 641698 301888 641798
rect 302012 641698 302112 641798
rect 302236 641698 302336 641798
rect 302460 641698 302560 641798
rect 302684 641698 302784 641798
rect 302908 641698 303008 641798
rect 303132 641698 303232 641798
rect 303356 641698 303456 641798
rect 303580 641698 303680 641798
rect 303804 641698 303904 641798
rect 304028 641698 304128 641798
rect 304252 641698 304352 641798
rect 304476 641698 304576 641798
rect 304700 641698 304800 641798
rect 304924 641698 305024 641798
rect 305148 641698 305248 641798
rect 305372 641698 305472 641798
rect 309346 641698 309446 641798
rect 309570 641698 309670 641798
rect 309794 641698 309894 641798
rect 310018 641698 310118 641798
rect 310242 641698 310342 641798
rect 310466 641698 310566 641798
rect 310690 641698 310790 641798
rect 310914 641698 311014 641798
rect 311138 641698 311238 641798
rect 311362 641698 311462 641798
rect 311586 641698 311686 641798
rect 311810 641698 311910 641798
rect 312034 641698 312134 641798
rect 312258 641698 312358 641798
rect 312482 641698 312582 641798
rect 312706 641698 312806 641798
rect 312930 641698 313030 641798
rect 313154 641698 313254 641798
rect 313378 641698 313478 641798
rect 313602 641698 313702 641798
rect 313826 641698 313926 641798
rect 314050 641698 314150 641798
rect 314274 641698 314374 641798
rect 314498 641698 314598 641798
rect 314722 641698 314822 641798
rect 314946 641698 315046 641798
rect 315170 641698 315270 641798
rect 315394 641698 315494 641798
rect 315618 641698 315718 641798
rect 315842 641698 315942 641798
rect 300643 640578 311917 640587
rect 300643 639740 300652 640578
rect 300652 639740 311908 640578
rect 311908 639740 311917 640578
rect 300643 639731 311917 639740
rect 289920 631440 294704 637184
rect 297850 637896 297950 637996
rect 298074 637896 298174 637996
rect 298298 637896 298398 637996
rect 298522 637896 298622 637996
rect 298746 637896 298846 637996
rect 297850 637672 297950 637772
rect 298074 637672 298174 637772
rect 298298 637672 298398 637772
rect 298522 637672 298622 637772
rect 298746 637672 298846 637772
rect 297850 637448 297950 637548
rect 298074 637448 298174 637548
rect 298298 637448 298398 637548
rect 298522 637448 298622 637548
rect 298746 637448 298846 637548
rect 297850 637224 297950 637324
rect 298074 637224 298174 637324
rect 298298 637224 298398 637324
rect 298522 637224 298622 637324
rect 298746 637224 298846 637324
rect 297850 637000 297950 637100
rect 298074 637000 298174 637100
rect 298298 637000 298398 637100
rect 298522 637000 298622 637100
rect 298746 637000 298846 637100
rect 297850 636776 297950 636876
rect 298074 636776 298174 636876
rect 298298 636776 298398 636876
rect 298522 636776 298622 636876
rect 298746 636776 298846 636876
rect 297850 636552 297950 636652
rect 298074 636552 298174 636652
rect 298298 636552 298398 636652
rect 298522 636552 298622 636652
rect 298746 636552 298846 636652
rect 297850 636328 297950 636428
rect 298074 636328 298174 636428
rect 298298 636328 298398 636428
rect 298522 636328 298622 636428
rect 298746 636328 298846 636428
rect 297850 636104 297950 636204
rect 298074 636104 298174 636204
rect 298298 636104 298398 636204
rect 298522 636104 298622 636204
rect 298746 636104 298846 636204
rect 297850 635880 297950 635980
rect 298074 635880 298174 635980
rect 298298 635880 298398 635980
rect 298522 635880 298622 635980
rect 298746 635880 298846 635980
rect 297850 635656 297950 635756
rect 298074 635656 298174 635756
rect 298298 635656 298398 635756
rect 298522 635656 298622 635756
rect 298746 635656 298846 635756
rect 297850 635432 297950 635532
rect 298074 635432 298174 635532
rect 298298 635432 298398 635532
rect 298522 635432 298622 635532
rect 298746 635432 298846 635532
rect 297850 635208 297950 635308
rect 298074 635208 298174 635308
rect 298298 635208 298398 635308
rect 298522 635208 298622 635308
rect 298746 635208 298846 635308
rect 297850 634984 297950 635084
rect 298074 634984 298174 635084
rect 298298 634984 298398 635084
rect 298522 634984 298622 635084
rect 298746 634984 298846 635084
rect 297850 634760 297950 634860
rect 298074 634760 298174 634860
rect 298298 634760 298398 634860
rect 298522 634760 298622 634860
rect 298746 634760 298846 634860
rect 297850 634536 297950 634636
rect 298074 634536 298174 634636
rect 298298 634536 298398 634636
rect 298522 634536 298622 634636
rect 298746 634536 298846 634636
rect 297850 634312 297950 634412
rect 298074 634312 298174 634412
rect 298298 634312 298398 634412
rect 298522 634312 298622 634412
rect 298746 634312 298846 634412
rect 297850 634088 297950 634188
rect 298074 634088 298174 634188
rect 298298 634088 298398 634188
rect 298522 634088 298622 634188
rect 298746 634088 298846 634188
rect 297850 633864 297950 633964
rect 298074 633864 298174 633964
rect 298298 633864 298398 633964
rect 298522 633864 298622 633964
rect 298746 633864 298846 633964
rect 297850 633640 297950 633740
rect 298074 633640 298174 633740
rect 298298 633640 298398 633740
rect 298522 633640 298622 633740
rect 298746 633640 298846 633740
rect 297850 633416 297950 633516
rect 298074 633416 298174 633516
rect 298298 633416 298398 633516
rect 298522 633416 298622 633516
rect 298746 633416 298846 633516
rect 297850 633192 297950 633292
rect 298074 633192 298174 633292
rect 298298 633192 298398 633292
rect 298522 633192 298622 633292
rect 298746 633192 298846 633292
rect 297850 632968 297950 633068
rect 298074 632968 298174 633068
rect 298298 632968 298398 633068
rect 298522 632968 298622 633068
rect 298746 632968 298846 633068
rect 297850 632744 297950 632844
rect 298074 632744 298174 632844
rect 298298 632744 298398 632844
rect 298522 632744 298622 632844
rect 298746 632744 298846 632844
rect 297850 632520 297950 632620
rect 298074 632520 298174 632620
rect 298298 632520 298398 632620
rect 298522 632520 298622 632620
rect 298746 632520 298846 632620
rect 297850 632296 297950 632396
rect 298074 632296 298174 632396
rect 298298 632296 298398 632396
rect 298522 632296 298622 632396
rect 298746 632296 298846 632396
rect 297850 632072 297950 632172
rect 298074 632072 298174 632172
rect 298298 632072 298398 632172
rect 298522 632072 298622 632172
rect 298746 632072 298846 632172
rect 297850 631848 297950 631948
rect 298074 631848 298174 631948
rect 298298 631848 298398 631948
rect 298522 631848 298622 631948
rect 298746 631848 298846 631948
rect 297850 631624 297950 631724
rect 298074 631624 298174 631724
rect 298298 631624 298398 631724
rect 298522 631624 298622 631724
rect 298746 631624 298846 631724
rect 297850 631400 297950 631500
rect 298074 631400 298174 631500
rect 298298 631400 298398 631500
rect 298522 631400 298622 631500
rect 298746 631400 298846 631500
rect 304931 631600 304995 632144
rect 305650 631600 305714 632144
rect 306369 631600 306433 632144
rect 307088 631600 307152 632144
rect 307807 631600 307871 632144
rect 308526 631600 308590 632144
rect 309245 631600 309309 632144
rect 309964 631600 310028 632144
rect 310683 631600 310747 632144
rect 311402 631600 311466 632144
rect 304931 630900 304995 631444
rect 305650 630900 305714 631444
rect 306369 630900 306433 631444
rect 307088 630900 307152 631444
rect 307807 630900 307871 631444
rect 308526 630900 308590 631444
rect 309245 630900 309309 631444
rect 309964 630900 310028 631444
rect 310683 630900 310747 631444
rect 311402 630900 311466 631444
rect 304931 630200 304995 630744
rect 305650 630200 305714 630744
rect 306369 630200 306433 630744
rect 307088 630200 307152 630744
rect 307807 630200 307871 630744
rect 308526 630200 308590 630744
rect 309245 630200 309309 630744
rect 309964 630200 310028 630744
rect 310683 630200 310747 630744
rect 311402 630200 311466 630744
rect 304931 629500 304995 630044
rect 305650 629500 305714 630044
rect 306369 629500 306433 630044
rect 307088 629500 307152 630044
rect 307807 629500 307871 630044
rect 308526 629500 308590 630044
rect 309245 629500 309309 630044
rect 309964 629500 310028 630044
rect 310683 629500 310747 630044
rect 311402 629500 311466 630044
rect 304931 628800 304995 629344
rect 305650 628800 305714 629344
rect 306369 628800 306433 629344
rect 307088 628800 307152 629344
rect 307807 628800 307871 629344
rect 308526 628800 308590 629344
rect 309245 628800 309309 629344
rect 309964 628800 310028 629344
rect 310683 628800 310747 629344
rect 311402 628800 311466 629344
rect 304931 628100 304995 628644
rect 305650 628100 305714 628644
rect 306369 628100 306433 628644
rect 307088 628100 307152 628644
rect 307807 628100 307871 628644
rect 308526 628100 308590 628644
rect 309245 628100 309309 628644
rect 309964 628100 310028 628644
rect 310683 628100 310747 628644
rect 311402 628100 311466 628644
rect 304931 627400 304995 627944
rect 305650 627400 305714 627944
rect 306369 627400 306433 627944
rect 307088 627400 307152 627944
rect 307807 627400 307871 627944
rect 308526 627400 308590 627944
rect 309245 627400 309309 627944
rect 309964 627400 310028 627944
rect 310683 627400 310747 627944
rect 311402 627400 311466 627944
rect 336480 645160 341264 650904
rect 510602 645217 515386 650961
rect 335616 642614 335716 642714
rect 335840 642614 335940 642714
rect 336064 642614 336164 642714
rect 336288 642614 336388 642714
rect 336512 642614 336612 642714
rect 336736 642614 336836 642714
rect 336960 642614 337060 642714
rect 337184 642614 337284 642714
rect 337408 642614 337508 642714
rect 337632 642614 337732 642714
rect 337856 642614 337956 642714
rect 338080 642614 338180 642714
rect 338304 642614 338404 642714
rect 338528 642614 338628 642714
rect 338752 642614 338852 642714
rect 338976 642614 339076 642714
rect 339200 642614 339300 642714
rect 339424 642614 339524 642714
rect 339648 642614 339748 642714
rect 339872 642614 339972 642714
rect 340096 642614 340196 642714
rect 340320 642614 340420 642714
rect 340544 642614 340644 642714
rect 340768 642614 340868 642714
rect 340992 642614 341092 642714
rect 341216 642614 341316 642714
rect 341440 642614 341540 642714
rect 341664 642614 341764 642714
rect 341888 642614 341988 642714
rect 342112 642614 342212 642714
rect 335616 642390 335716 642490
rect 335840 642390 335940 642490
rect 336064 642390 336164 642490
rect 336288 642390 336388 642490
rect 336512 642390 336612 642490
rect 336736 642390 336836 642490
rect 336960 642390 337060 642490
rect 337184 642390 337284 642490
rect 337408 642390 337508 642490
rect 337632 642390 337732 642490
rect 337856 642390 337956 642490
rect 338080 642390 338180 642490
rect 338304 642390 338404 642490
rect 338528 642390 338628 642490
rect 338752 642390 338852 642490
rect 338976 642390 339076 642490
rect 339200 642390 339300 642490
rect 339424 642390 339524 642490
rect 339648 642390 339748 642490
rect 339872 642390 339972 642490
rect 340096 642390 340196 642490
rect 340320 642390 340420 642490
rect 340544 642390 340644 642490
rect 340768 642390 340868 642490
rect 340992 642390 341092 642490
rect 341216 642390 341316 642490
rect 341440 642390 341540 642490
rect 341664 642390 341764 642490
rect 341888 642390 341988 642490
rect 342112 642390 342212 642490
rect 335616 642166 335716 642266
rect 335840 642166 335940 642266
rect 336064 642166 336164 642266
rect 336288 642166 336388 642266
rect 336512 642166 336612 642266
rect 336736 642166 336836 642266
rect 336960 642166 337060 642266
rect 337184 642166 337284 642266
rect 337408 642166 337508 642266
rect 337632 642166 337732 642266
rect 337856 642166 337956 642266
rect 338080 642166 338180 642266
rect 338304 642166 338404 642266
rect 338528 642166 338628 642266
rect 338752 642166 338852 642266
rect 338976 642166 339076 642266
rect 339200 642166 339300 642266
rect 339424 642166 339524 642266
rect 339648 642166 339748 642266
rect 339872 642166 339972 642266
rect 340096 642166 340196 642266
rect 340320 642166 340420 642266
rect 340544 642166 340644 642266
rect 340768 642166 340868 642266
rect 340992 642166 341092 642266
rect 341216 642166 341316 642266
rect 341440 642166 341540 642266
rect 341664 642166 341764 642266
rect 341888 642166 341988 642266
rect 342112 642166 342212 642266
rect 335616 641942 335716 642042
rect 335840 641942 335940 642042
rect 336064 641942 336164 642042
rect 336288 641942 336388 642042
rect 336512 641942 336612 642042
rect 336736 641942 336836 642042
rect 336960 641942 337060 642042
rect 337184 641942 337284 642042
rect 337408 641942 337508 642042
rect 337632 641942 337732 642042
rect 337856 641942 337956 642042
rect 338080 641942 338180 642042
rect 338304 641942 338404 642042
rect 338528 641942 338628 642042
rect 338752 641942 338852 642042
rect 338976 641942 339076 642042
rect 339200 641942 339300 642042
rect 339424 641942 339524 642042
rect 339648 641942 339748 642042
rect 339872 641942 339972 642042
rect 340096 641942 340196 642042
rect 340320 641942 340420 642042
rect 340544 641942 340644 642042
rect 340768 641942 340868 642042
rect 340992 641942 341092 642042
rect 341216 641942 341316 642042
rect 341440 641942 341540 642042
rect 341664 641942 341764 642042
rect 341888 641942 341988 642042
rect 342112 641942 342212 642042
rect 335616 641718 335716 641818
rect 335840 641718 335940 641818
rect 336064 641718 336164 641818
rect 336288 641718 336388 641818
rect 336512 641718 336612 641818
rect 336736 641718 336836 641818
rect 336960 641718 337060 641818
rect 337184 641718 337284 641818
rect 337408 641718 337508 641818
rect 337632 641718 337732 641818
rect 337856 641718 337956 641818
rect 338080 641718 338180 641818
rect 338304 641718 338404 641818
rect 338528 641718 338628 641818
rect 338752 641718 338852 641818
rect 338976 641718 339076 641818
rect 339200 641718 339300 641818
rect 339424 641718 339524 641818
rect 339648 641718 339748 641818
rect 339872 641718 339972 641818
rect 340096 641718 340196 641818
rect 340320 641718 340420 641818
rect 340544 641718 340644 641818
rect 340768 641718 340868 641818
rect 340992 641718 341092 641818
rect 341216 641718 341316 641818
rect 341440 641718 341540 641818
rect 341664 641718 341764 641818
rect 341888 641718 341988 641818
rect 342112 641718 342212 641818
rect 342130 637896 342230 637996
rect 342354 637896 342454 637996
rect 342578 637896 342678 637996
rect 342802 637896 342902 637996
rect 343026 637896 343126 637996
rect 342130 637672 342230 637772
rect 342354 637672 342454 637772
rect 342578 637672 342678 637772
rect 342802 637672 342902 637772
rect 343026 637672 343126 637772
rect 342130 637448 342230 637548
rect 342354 637448 342454 637548
rect 342578 637448 342678 637548
rect 342802 637448 342902 637548
rect 343026 637448 343126 637548
rect 342130 637224 342230 637324
rect 342354 637224 342454 637324
rect 342578 637224 342678 637324
rect 342802 637224 342902 637324
rect 343026 637224 343126 637324
rect 342130 637000 342230 637100
rect 342354 637000 342454 637100
rect 342578 637000 342678 637100
rect 342802 637000 342902 637100
rect 343026 637000 343126 637100
rect 342130 636776 342230 636876
rect 342354 636776 342454 636876
rect 342578 636776 342678 636876
rect 342802 636776 342902 636876
rect 343026 636776 343126 636876
rect 342130 636552 342230 636652
rect 342354 636552 342454 636652
rect 342578 636552 342678 636652
rect 342802 636552 342902 636652
rect 343026 636552 343126 636652
rect 342130 636328 342230 636428
rect 342354 636328 342454 636428
rect 342578 636328 342678 636428
rect 342802 636328 342902 636428
rect 343026 636328 343126 636428
rect 342130 636104 342230 636204
rect 342354 636104 342454 636204
rect 342578 636104 342678 636204
rect 342802 636104 342902 636204
rect 343026 636104 343126 636204
rect 342130 635880 342230 635980
rect 342354 635880 342454 635980
rect 342578 635880 342678 635980
rect 342802 635880 342902 635980
rect 343026 635880 343126 635980
rect 342130 635656 342230 635756
rect 342354 635656 342454 635756
rect 342578 635656 342678 635756
rect 342802 635656 342902 635756
rect 343026 635656 343126 635756
rect 342130 635432 342230 635532
rect 342354 635432 342454 635532
rect 342578 635432 342678 635532
rect 342802 635432 342902 635532
rect 343026 635432 343126 635532
rect 342130 635208 342230 635308
rect 342354 635208 342454 635308
rect 342578 635208 342678 635308
rect 342802 635208 342902 635308
rect 343026 635208 343126 635308
rect 342130 634984 342230 635084
rect 342354 634984 342454 635084
rect 342578 634984 342678 635084
rect 342802 634984 342902 635084
rect 343026 634984 343126 635084
rect 342130 634760 342230 634860
rect 342354 634760 342454 634860
rect 342578 634760 342678 634860
rect 342802 634760 342902 634860
rect 343026 634760 343126 634860
rect 342130 634536 342230 634636
rect 342354 634536 342454 634636
rect 342578 634536 342678 634636
rect 342802 634536 342902 634636
rect 343026 634536 343126 634636
rect 342130 634312 342230 634412
rect 342354 634312 342454 634412
rect 342578 634312 342678 634412
rect 342802 634312 342902 634412
rect 343026 634312 343126 634412
rect 342130 634088 342230 634188
rect 342354 634088 342454 634188
rect 342578 634088 342678 634188
rect 342802 634088 342902 634188
rect 343026 634088 343126 634188
rect 342130 633864 342230 633964
rect 342354 633864 342454 633964
rect 342578 633864 342678 633964
rect 342802 633864 342902 633964
rect 343026 633864 343126 633964
rect 342130 633640 342230 633740
rect 342354 633640 342454 633740
rect 342578 633640 342678 633740
rect 342802 633640 342902 633740
rect 343026 633640 343126 633740
rect 342130 633416 342230 633516
rect 342354 633416 342454 633516
rect 342578 633416 342678 633516
rect 342802 633416 342902 633516
rect 343026 633416 343126 633516
rect 342130 633192 342230 633292
rect 342354 633192 342454 633292
rect 342578 633192 342678 633292
rect 342802 633192 342902 633292
rect 343026 633192 343126 633292
rect 342130 632968 342230 633068
rect 342354 632968 342454 633068
rect 342578 632968 342678 633068
rect 342802 632968 342902 633068
rect 343026 632968 343126 633068
rect 342130 632744 342230 632844
rect 342354 632744 342454 632844
rect 342578 632744 342678 632844
rect 342802 632744 342902 632844
rect 343026 632744 343126 632844
rect 342130 632520 342230 632620
rect 342354 632520 342454 632620
rect 342578 632520 342678 632620
rect 342802 632520 342902 632620
rect 343026 632520 343126 632620
rect 342130 632296 342230 632396
rect 342354 632296 342454 632396
rect 342578 632296 342678 632396
rect 342802 632296 342902 632396
rect 343026 632296 343126 632396
rect 342130 632072 342230 632172
rect 342354 632072 342454 632172
rect 342578 632072 342678 632172
rect 342802 632072 342902 632172
rect 343026 632072 343126 632172
rect 342130 631848 342230 631948
rect 342354 631848 342454 631948
rect 342578 631848 342678 631948
rect 342802 631848 342902 631948
rect 343026 631848 343126 631948
rect 342130 631624 342230 631724
rect 342354 631624 342454 631724
rect 342578 631624 342678 631724
rect 342802 631624 342902 631724
rect 343026 631624 343126 631724
rect 342130 631400 342230 631500
rect 342354 631400 342454 631500
rect 342578 631400 342678 631500
rect 342802 631400 342902 631500
rect 343026 631400 343126 631500
rect 510602 631817 515386 637561
rect 319400 628668 319600 628868
rect 319834 628668 320034 628868
rect 320268 628668 320468 628868
rect 320702 628668 320902 628868
rect 321136 628668 321336 628868
rect 321570 628668 321770 628868
rect 322004 628668 322204 628868
rect 322438 628668 322638 628868
rect 322872 628668 323072 628868
rect 323306 628668 323506 628868
rect 323740 628668 323940 628868
rect 324140 628668 324340 628868
rect 324540 628668 324740 628868
rect 324940 628668 325140 628868
rect 325340 628668 325540 628868
rect 325740 628668 325940 628868
rect 326140 628668 326340 628868
rect 326540 628668 326740 628868
rect 326940 628668 327140 628868
rect 327340 628668 327540 628868
rect 328940 628668 329140 628868
rect 329340 628668 329540 628868
rect 329740 628668 329940 628868
rect 330140 628668 330340 628868
rect 330540 628668 330740 628868
rect 330940 628668 331140 628868
rect 331340 628668 331540 628868
rect 331740 628668 331940 628868
rect 332140 628668 332340 628868
rect 319400 628234 319600 628434
rect 319834 628234 320034 628434
rect 320268 628234 320468 628434
rect 320702 628234 320902 628434
rect 321136 628234 321336 628434
rect 321570 628234 321770 628434
rect 322004 628234 322204 628434
rect 322438 628234 322638 628434
rect 322872 628234 323072 628434
rect 323306 628234 323506 628434
rect 323740 628234 323940 628434
rect 319400 627800 319600 628000
rect 319834 627800 320034 628000
rect 320268 627800 320468 628000
rect 320702 627800 320902 628000
rect 321136 627800 321336 628000
rect 321570 627800 321770 628000
rect 322004 627800 322204 628000
rect 322438 627800 322638 628000
rect 322872 627800 323072 628000
rect 323306 627800 323506 628000
rect 323740 627800 323940 628000
rect 304931 626700 304995 627244
rect 305650 626700 305714 627244
rect 306369 626700 306433 627244
rect 307088 626700 307152 627244
rect 307807 626700 307871 627244
rect 308526 626700 308590 627244
rect 309245 626700 309309 627244
rect 309964 626700 310028 627244
rect 310683 626700 310747 627244
rect 311402 626700 311466 627244
rect 297856 626112 297920 626176
rect 297984 626112 298048 626176
rect 298112 626112 298176 626176
rect 298240 626112 298304 626176
rect 298368 626112 298432 626176
rect 298496 626112 298560 626176
rect 298624 626112 298688 626176
rect 298752 626112 298816 626176
rect 298880 626112 298944 626176
rect 297856 625984 297920 626048
rect 297984 625984 298048 626048
rect 298112 625984 298176 626048
rect 298240 625984 298304 626048
rect 298368 625984 298432 626048
rect 298496 625984 298560 626048
rect 298624 625984 298688 626048
rect 298752 625984 298816 626048
rect 298880 625984 298944 626048
rect 297856 625856 297920 625920
rect 297984 625856 298048 625920
rect 298112 625856 298176 625920
rect 298240 625856 298304 625920
rect 298368 625856 298432 625920
rect 298496 625856 298560 625920
rect 298624 625856 298688 625920
rect 298752 625856 298816 625920
rect 298880 625856 298944 625920
rect 297856 625728 297920 625792
rect 297984 625728 298048 625792
rect 298112 625728 298176 625792
rect 298240 625728 298304 625792
rect 298368 625728 298432 625792
rect 298496 625728 298560 625792
rect 298624 625728 298688 625792
rect 298752 625728 298816 625792
rect 298880 625728 298944 625792
rect 304931 626000 304995 626544
rect 305650 626000 305714 626544
rect 306369 626000 306433 626544
rect 307088 626000 307152 626544
rect 307807 626000 307871 626544
rect 308526 626000 308590 626544
rect 309245 626000 309309 626544
rect 309964 626000 310028 626544
rect 310683 626000 310747 626544
rect 311402 626000 311466 626544
rect 312958 626314 333268 627286
rect 304931 625300 304995 625844
rect 305650 625300 305714 625844
rect 306369 625300 306433 625844
rect 307088 625300 307152 625844
rect 307807 625300 307871 625844
rect 308526 625300 308590 625844
rect 309245 625300 309309 625844
rect 309964 625300 310028 625844
rect 310683 625300 310747 625844
rect 311402 625300 311466 625844
rect 289920 618040 294704 623784
rect 297850 624496 297950 624596
rect 298074 624496 298174 624596
rect 298298 624496 298398 624596
rect 298522 624496 298622 624596
rect 298746 624496 298846 624596
rect 297850 624272 297950 624372
rect 298074 624272 298174 624372
rect 298298 624272 298398 624372
rect 298522 624272 298622 624372
rect 298746 624272 298846 624372
rect 297850 624048 297950 624148
rect 298074 624048 298174 624148
rect 298298 624048 298398 624148
rect 298522 624048 298622 624148
rect 298746 624048 298846 624148
rect 297850 623824 297950 623924
rect 298074 623824 298174 623924
rect 298298 623824 298398 623924
rect 298522 623824 298622 623924
rect 298746 623824 298846 623924
rect 297850 623600 297950 623700
rect 298074 623600 298174 623700
rect 298298 623600 298398 623700
rect 298522 623600 298622 623700
rect 298746 623600 298846 623700
rect 297850 623376 297950 623476
rect 298074 623376 298174 623476
rect 298298 623376 298398 623476
rect 298522 623376 298622 623476
rect 298746 623376 298846 623476
rect 297850 623152 297950 623252
rect 298074 623152 298174 623252
rect 298298 623152 298398 623252
rect 298522 623152 298622 623252
rect 298746 623152 298846 623252
rect 297850 622928 297950 623028
rect 298074 622928 298174 623028
rect 298298 622928 298398 623028
rect 298522 622928 298622 623028
rect 298746 622928 298846 623028
rect 297850 622704 297950 622804
rect 298074 622704 298174 622804
rect 298298 622704 298398 622804
rect 298522 622704 298622 622804
rect 298746 622704 298846 622804
rect 297850 622480 297950 622580
rect 298074 622480 298174 622580
rect 298298 622480 298398 622580
rect 298522 622480 298622 622580
rect 298746 622480 298846 622580
rect 297850 622256 297950 622356
rect 298074 622256 298174 622356
rect 298298 622256 298398 622356
rect 298522 622256 298622 622356
rect 298746 622256 298846 622356
rect 297850 622032 297950 622132
rect 298074 622032 298174 622132
rect 298298 622032 298398 622132
rect 298522 622032 298622 622132
rect 298746 622032 298846 622132
rect 297850 621808 297950 621908
rect 298074 621808 298174 621908
rect 298298 621808 298398 621908
rect 298522 621808 298622 621908
rect 298746 621808 298846 621908
rect 297850 621584 297950 621684
rect 298074 621584 298174 621684
rect 298298 621584 298398 621684
rect 298522 621584 298622 621684
rect 298746 621584 298846 621684
rect 297850 621360 297950 621460
rect 298074 621360 298174 621460
rect 298298 621360 298398 621460
rect 298522 621360 298622 621460
rect 298746 621360 298846 621460
rect 297850 621136 297950 621236
rect 298074 621136 298174 621236
rect 298298 621136 298398 621236
rect 298522 621136 298622 621236
rect 298746 621136 298846 621236
rect 297850 620912 297950 621012
rect 298074 620912 298174 621012
rect 298298 620912 298398 621012
rect 298522 620912 298622 621012
rect 298746 620912 298846 621012
rect 297850 620688 297950 620788
rect 298074 620688 298174 620788
rect 298298 620688 298398 620788
rect 298522 620688 298622 620788
rect 298746 620688 298846 620788
rect 297850 620464 297950 620564
rect 298074 620464 298174 620564
rect 298298 620464 298398 620564
rect 298522 620464 298622 620564
rect 298746 620464 298846 620564
rect 297850 620240 297950 620340
rect 298074 620240 298174 620340
rect 298298 620240 298398 620340
rect 298522 620240 298622 620340
rect 298746 620240 298846 620340
rect 297850 620016 297950 620116
rect 298074 620016 298174 620116
rect 298298 620016 298398 620116
rect 298522 620016 298622 620116
rect 298746 620016 298846 620116
rect 297850 619792 297950 619892
rect 298074 619792 298174 619892
rect 298298 619792 298398 619892
rect 298522 619792 298622 619892
rect 298746 619792 298846 619892
rect 303590 620135 304218 620149
rect 303590 619883 303604 620135
rect 303604 619883 304204 620135
rect 304204 619883 304218 620135
rect 303590 619869 304218 619883
rect 297850 619568 297950 619668
rect 298074 619568 298174 619668
rect 298298 619568 298398 619668
rect 298522 619568 298622 619668
rect 298746 619568 298846 619668
rect 297850 619344 297950 619444
rect 298074 619344 298174 619444
rect 298298 619344 298398 619444
rect 298522 619344 298622 619444
rect 298746 619344 298846 619444
rect 297850 619120 297950 619220
rect 298074 619120 298174 619220
rect 298298 619120 298398 619220
rect 298522 619120 298622 619220
rect 298746 619120 298846 619220
rect 297850 618896 297950 618996
rect 298074 618896 298174 618996
rect 298298 618896 298398 618996
rect 298522 618896 298622 618996
rect 298746 618896 298846 618996
rect 297850 618672 297950 618772
rect 298074 618672 298174 618772
rect 298298 618672 298398 618772
rect 298522 618672 298622 618772
rect 298746 618672 298846 618772
rect 297850 618448 297950 618548
rect 298074 618448 298174 618548
rect 298298 618448 298398 618548
rect 298522 618448 298622 618548
rect 298746 618448 298846 618548
rect 297850 618224 297950 618324
rect 298074 618224 298174 618324
rect 298298 618224 298398 618324
rect 298522 618224 298622 618324
rect 298746 618224 298846 618324
rect 297850 618000 297950 618100
rect 298074 618000 298174 618100
rect 298298 618000 298398 618100
rect 298522 618000 298622 618100
rect 298746 618000 298846 618100
rect 342130 624496 342230 624596
rect 342354 624496 342454 624596
rect 342578 624496 342678 624596
rect 342802 624496 342902 624596
rect 343026 624496 343126 624596
rect 342130 624272 342230 624372
rect 342354 624272 342454 624372
rect 342578 624272 342678 624372
rect 342802 624272 342902 624372
rect 343026 624272 343126 624372
rect 342130 624048 342230 624148
rect 342354 624048 342454 624148
rect 342578 624048 342678 624148
rect 342802 624048 342902 624148
rect 343026 624048 343126 624148
rect 342130 623824 342230 623924
rect 342354 623824 342454 623924
rect 342578 623824 342678 623924
rect 342802 623824 342902 623924
rect 343026 623824 343126 623924
rect 342130 623600 342230 623700
rect 342354 623600 342454 623700
rect 342578 623600 342678 623700
rect 342802 623600 342902 623700
rect 343026 623600 343126 623700
rect 342130 623376 342230 623476
rect 342354 623376 342454 623476
rect 342578 623376 342678 623476
rect 342802 623376 342902 623476
rect 343026 623376 343126 623476
rect 342130 623152 342230 623252
rect 342354 623152 342454 623252
rect 342578 623152 342678 623252
rect 342802 623152 342902 623252
rect 343026 623152 343126 623252
rect 342130 622928 342230 623028
rect 342354 622928 342454 623028
rect 342578 622928 342678 623028
rect 342802 622928 342902 623028
rect 343026 622928 343126 623028
rect 342130 622704 342230 622804
rect 342354 622704 342454 622804
rect 342578 622704 342678 622804
rect 342802 622704 342902 622804
rect 343026 622704 343126 622804
rect 342130 622480 342230 622580
rect 342354 622480 342454 622580
rect 342578 622480 342678 622580
rect 342802 622480 342902 622580
rect 343026 622480 343126 622580
rect 342130 622256 342230 622356
rect 342354 622256 342454 622356
rect 342578 622256 342678 622356
rect 342802 622256 342902 622356
rect 343026 622256 343126 622356
rect 342130 622032 342230 622132
rect 342354 622032 342454 622132
rect 342578 622032 342678 622132
rect 342802 622032 342902 622132
rect 343026 622032 343126 622132
rect 342130 621808 342230 621908
rect 342354 621808 342454 621908
rect 342578 621808 342678 621908
rect 342802 621808 342902 621908
rect 343026 621808 343126 621908
rect 342130 621584 342230 621684
rect 342354 621584 342454 621684
rect 342578 621584 342678 621684
rect 342802 621584 342902 621684
rect 343026 621584 343126 621684
rect 342130 621360 342230 621460
rect 342354 621360 342454 621460
rect 342578 621360 342678 621460
rect 342802 621360 342902 621460
rect 343026 621360 343126 621460
rect 342130 621136 342230 621236
rect 342354 621136 342454 621236
rect 342578 621136 342678 621236
rect 342802 621136 342902 621236
rect 343026 621136 343126 621236
rect 342130 620912 342230 621012
rect 342354 620912 342454 621012
rect 342578 620912 342678 621012
rect 342802 620912 342902 621012
rect 343026 620912 343126 621012
rect 342130 620688 342230 620788
rect 342354 620688 342454 620788
rect 342578 620688 342678 620788
rect 342802 620688 342902 620788
rect 343026 620688 343126 620788
rect 342130 620464 342230 620564
rect 342354 620464 342454 620564
rect 342578 620464 342678 620564
rect 342802 620464 342902 620564
rect 343026 620464 343126 620564
rect 342130 620240 342230 620340
rect 342354 620240 342454 620340
rect 342578 620240 342678 620340
rect 342802 620240 342902 620340
rect 343026 620240 343126 620340
rect 312081 620135 312709 620149
rect 312081 619883 312095 620135
rect 312095 619883 312695 620135
rect 312695 619883 312709 620135
rect 312081 619869 312709 619883
rect 342130 620016 342230 620116
rect 342354 620016 342454 620116
rect 342578 620016 342678 620116
rect 342802 620016 342902 620116
rect 343026 620016 343126 620116
rect 342130 619792 342230 619892
rect 342354 619792 342454 619892
rect 342578 619792 342678 619892
rect 342802 619792 342902 619892
rect 343026 619792 343126 619892
rect 342130 619568 342230 619668
rect 342354 619568 342454 619668
rect 342578 619568 342678 619668
rect 342802 619568 342902 619668
rect 343026 619568 343126 619668
rect 342130 619344 342230 619444
rect 342354 619344 342454 619444
rect 342578 619344 342678 619444
rect 342802 619344 342902 619444
rect 343026 619344 343126 619444
rect 342130 619120 342230 619220
rect 342354 619120 342454 619220
rect 342578 619120 342678 619220
rect 342802 619120 342902 619220
rect 343026 619120 343126 619220
rect 342130 618896 342230 618996
rect 342354 618896 342454 618996
rect 342578 618896 342678 618996
rect 342802 618896 342902 618996
rect 343026 618896 343126 618996
rect 342130 618672 342230 618772
rect 342354 618672 342454 618772
rect 342578 618672 342678 618772
rect 342802 618672 342902 618772
rect 343026 618672 343126 618772
rect 342130 618448 342230 618548
rect 342354 618448 342454 618548
rect 342578 618448 342678 618548
rect 342802 618448 342902 618548
rect 343026 618448 343126 618548
rect 342130 618224 342230 618324
rect 342354 618224 342454 618324
rect 342578 618224 342678 618324
rect 342802 618224 342902 618324
rect 343026 618224 343126 618324
rect 342130 618000 342230 618100
rect 342354 618000 342454 618100
rect 342578 618000 342678 618100
rect 342802 618000 342902 618100
rect 343026 618000 343126 618100
rect 510602 618417 515386 624161
rect 289920 605020 294704 610764
rect 298876 615374 298976 615474
rect 299100 615374 299200 615474
rect 299324 615374 299424 615474
rect 299548 615374 299648 615474
rect 299772 615374 299872 615474
rect 299996 615374 300096 615474
rect 300220 615374 300320 615474
rect 300444 615374 300544 615474
rect 300668 615374 300768 615474
rect 300892 615374 300992 615474
rect 301116 615374 301216 615474
rect 301340 615374 301440 615474
rect 301564 615374 301664 615474
rect 301788 615374 301888 615474
rect 302012 615374 302112 615474
rect 302236 615374 302336 615474
rect 302460 615374 302560 615474
rect 302684 615374 302784 615474
rect 302908 615374 303008 615474
rect 303132 615374 303232 615474
rect 303356 615374 303456 615474
rect 303580 615374 303680 615474
rect 303804 615374 303904 615474
rect 304028 615374 304128 615474
rect 304252 615374 304352 615474
rect 304476 615374 304576 615474
rect 304700 615374 304800 615474
rect 304924 615374 305024 615474
rect 305148 615374 305248 615474
rect 305372 615374 305472 615474
rect 309346 615374 309446 615474
rect 309570 615374 309670 615474
rect 309794 615374 309894 615474
rect 310018 615374 310118 615474
rect 310242 615374 310342 615474
rect 310466 615374 310566 615474
rect 310690 615374 310790 615474
rect 310914 615374 311014 615474
rect 311138 615374 311238 615474
rect 311362 615374 311462 615474
rect 311586 615374 311686 615474
rect 311810 615374 311910 615474
rect 312034 615374 312134 615474
rect 312258 615374 312358 615474
rect 312482 615374 312582 615474
rect 312706 615374 312806 615474
rect 312930 615374 313030 615474
rect 313154 615374 313254 615474
rect 313378 615374 313478 615474
rect 313602 615374 313702 615474
rect 313826 615374 313926 615474
rect 314050 615374 314150 615474
rect 314274 615374 314374 615474
rect 314498 615374 314598 615474
rect 314722 615374 314822 615474
rect 314946 615374 315046 615474
rect 315170 615374 315270 615474
rect 315394 615374 315494 615474
rect 315618 615374 315718 615474
rect 315842 615374 315942 615474
rect 298876 615150 298976 615250
rect 299100 615150 299200 615250
rect 299324 615150 299424 615250
rect 299548 615150 299648 615250
rect 299772 615150 299872 615250
rect 299996 615150 300096 615250
rect 300220 615150 300320 615250
rect 300444 615150 300544 615250
rect 300668 615150 300768 615250
rect 300892 615150 300992 615250
rect 301116 615150 301216 615250
rect 301340 615150 301440 615250
rect 301564 615150 301664 615250
rect 301788 615150 301888 615250
rect 302012 615150 302112 615250
rect 302236 615150 302336 615250
rect 302460 615150 302560 615250
rect 302684 615150 302784 615250
rect 302908 615150 303008 615250
rect 303132 615150 303232 615250
rect 303356 615150 303456 615250
rect 303580 615150 303680 615250
rect 303804 615150 303904 615250
rect 304028 615150 304128 615250
rect 304252 615150 304352 615250
rect 304476 615150 304576 615250
rect 304700 615150 304800 615250
rect 304924 615150 305024 615250
rect 305148 615150 305248 615250
rect 305372 615150 305472 615250
rect 309346 615150 309446 615250
rect 309570 615150 309670 615250
rect 309794 615150 309894 615250
rect 310018 615150 310118 615250
rect 310242 615150 310342 615250
rect 310466 615150 310566 615250
rect 310690 615150 310790 615250
rect 310914 615150 311014 615250
rect 311138 615150 311238 615250
rect 311362 615150 311462 615250
rect 311586 615150 311686 615250
rect 311810 615150 311910 615250
rect 312034 615150 312134 615250
rect 312258 615150 312358 615250
rect 312482 615150 312582 615250
rect 312706 615150 312806 615250
rect 312930 615150 313030 615250
rect 313154 615150 313254 615250
rect 313378 615150 313478 615250
rect 313602 615150 313702 615250
rect 313826 615150 313926 615250
rect 314050 615150 314150 615250
rect 314274 615150 314374 615250
rect 314498 615150 314598 615250
rect 314722 615150 314822 615250
rect 314946 615150 315046 615250
rect 315170 615150 315270 615250
rect 315394 615150 315494 615250
rect 315618 615150 315718 615250
rect 315842 615150 315942 615250
rect 298876 614926 298976 615026
rect 299100 614926 299200 615026
rect 299324 614926 299424 615026
rect 299548 614926 299648 615026
rect 299772 614926 299872 615026
rect 299996 614926 300096 615026
rect 300220 614926 300320 615026
rect 300444 614926 300544 615026
rect 300668 614926 300768 615026
rect 300892 614926 300992 615026
rect 301116 614926 301216 615026
rect 301340 614926 301440 615026
rect 301564 614926 301664 615026
rect 301788 614926 301888 615026
rect 302012 614926 302112 615026
rect 302236 614926 302336 615026
rect 302460 614926 302560 615026
rect 302684 614926 302784 615026
rect 302908 614926 303008 615026
rect 303132 614926 303232 615026
rect 303356 614926 303456 615026
rect 303580 614926 303680 615026
rect 303804 614926 303904 615026
rect 304028 614926 304128 615026
rect 304252 614926 304352 615026
rect 304476 614926 304576 615026
rect 304700 614926 304800 615026
rect 304924 614926 305024 615026
rect 305148 614926 305248 615026
rect 305372 614926 305472 615026
rect 309346 614926 309446 615026
rect 309570 614926 309670 615026
rect 309794 614926 309894 615026
rect 310018 614926 310118 615026
rect 310242 614926 310342 615026
rect 310466 614926 310566 615026
rect 310690 614926 310790 615026
rect 310914 614926 311014 615026
rect 311138 614926 311238 615026
rect 311362 614926 311462 615026
rect 311586 614926 311686 615026
rect 311810 614926 311910 615026
rect 312034 614926 312134 615026
rect 312258 614926 312358 615026
rect 312482 614926 312582 615026
rect 312706 614926 312806 615026
rect 312930 614926 313030 615026
rect 313154 614926 313254 615026
rect 313378 614926 313478 615026
rect 313602 614926 313702 615026
rect 313826 614926 313926 615026
rect 314050 614926 314150 615026
rect 314274 614926 314374 615026
rect 314498 614926 314598 615026
rect 314722 614926 314822 615026
rect 314946 614926 315046 615026
rect 315170 614926 315270 615026
rect 315394 614926 315494 615026
rect 315618 614926 315718 615026
rect 315842 614926 315942 615026
rect 298876 614702 298976 614802
rect 299100 614702 299200 614802
rect 299324 614702 299424 614802
rect 299548 614702 299648 614802
rect 299772 614702 299872 614802
rect 299996 614702 300096 614802
rect 300220 614702 300320 614802
rect 300444 614702 300544 614802
rect 300668 614702 300768 614802
rect 300892 614702 300992 614802
rect 301116 614702 301216 614802
rect 301340 614702 301440 614802
rect 301564 614702 301664 614802
rect 301788 614702 301888 614802
rect 302012 614702 302112 614802
rect 302236 614702 302336 614802
rect 302460 614702 302560 614802
rect 302684 614702 302784 614802
rect 302908 614702 303008 614802
rect 303132 614702 303232 614802
rect 303356 614702 303456 614802
rect 303580 614702 303680 614802
rect 303804 614702 303904 614802
rect 304028 614702 304128 614802
rect 304252 614702 304352 614802
rect 304476 614702 304576 614802
rect 304700 614702 304800 614802
rect 304924 614702 305024 614802
rect 305148 614702 305248 614802
rect 305372 614702 305472 614802
rect 309346 614702 309446 614802
rect 309570 614702 309670 614802
rect 309794 614702 309894 614802
rect 310018 614702 310118 614802
rect 310242 614702 310342 614802
rect 310466 614702 310566 614802
rect 310690 614702 310790 614802
rect 310914 614702 311014 614802
rect 311138 614702 311238 614802
rect 311362 614702 311462 614802
rect 311586 614702 311686 614802
rect 311810 614702 311910 614802
rect 312034 614702 312134 614802
rect 312258 614702 312358 614802
rect 312482 614702 312582 614802
rect 312706 614702 312806 614802
rect 312930 614702 313030 614802
rect 313154 614702 313254 614802
rect 313378 614702 313478 614802
rect 313602 614702 313702 614802
rect 313826 614702 313926 614802
rect 314050 614702 314150 614802
rect 314274 614702 314374 614802
rect 314498 614702 314598 614802
rect 314722 614702 314822 614802
rect 314946 614702 315046 614802
rect 315170 614702 315270 614802
rect 315394 614702 315494 614802
rect 315618 614702 315718 614802
rect 315842 614702 315942 614802
rect 298876 614478 298976 614578
rect 299100 614478 299200 614578
rect 299324 614478 299424 614578
rect 299548 614478 299648 614578
rect 299772 614478 299872 614578
rect 299996 614478 300096 614578
rect 300220 614478 300320 614578
rect 300444 614478 300544 614578
rect 300668 614478 300768 614578
rect 300892 614478 300992 614578
rect 301116 614478 301216 614578
rect 301340 614478 301440 614578
rect 301564 614478 301664 614578
rect 301788 614478 301888 614578
rect 302012 614478 302112 614578
rect 302236 614478 302336 614578
rect 302460 614478 302560 614578
rect 302684 614478 302784 614578
rect 302908 614478 303008 614578
rect 303132 614478 303232 614578
rect 303356 614478 303456 614578
rect 303580 614478 303680 614578
rect 303804 614478 303904 614578
rect 304028 614478 304128 614578
rect 304252 614478 304352 614578
rect 304476 614478 304576 614578
rect 304700 614478 304800 614578
rect 304924 614478 305024 614578
rect 305148 614478 305248 614578
rect 305372 614478 305472 614578
rect 309346 614478 309446 614578
rect 309570 614478 309670 614578
rect 309794 614478 309894 614578
rect 310018 614478 310118 614578
rect 310242 614478 310342 614578
rect 310466 614478 310566 614578
rect 310690 614478 310790 614578
rect 310914 614478 311014 614578
rect 311138 614478 311238 614578
rect 311362 614478 311462 614578
rect 311586 614478 311686 614578
rect 311810 614478 311910 614578
rect 312034 614478 312134 614578
rect 312258 614478 312358 614578
rect 312482 614478 312582 614578
rect 312706 614478 312806 614578
rect 312930 614478 313030 614578
rect 313154 614478 313254 614578
rect 313378 614478 313478 614578
rect 313602 614478 313702 614578
rect 313826 614478 313926 614578
rect 314050 614478 314150 614578
rect 314274 614478 314374 614578
rect 314498 614478 314598 614578
rect 314722 614478 314822 614578
rect 314946 614478 315046 614578
rect 315170 614478 315270 614578
rect 315394 614478 315494 614578
rect 315618 614478 315718 614578
rect 315842 614478 315942 614578
rect 298920 605336 303704 611080
rect 304920 605336 309704 611080
rect 310920 605336 315704 611080
rect 335616 615394 335716 615494
rect 335840 615394 335940 615494
rect 336064 615394 336164 615494
rect 336288 615394 336388 615494
rect 336512 615394 336612 615494
rect 336736 615394 336836 615494
rect 336960 615394 337060 615494
rect 337184 615394 337284 615494
rect 337408 615394 337508 615494
rect 337632 615394 337732 615494
rect 337856 615394 337956 615494
rect 338080 615394 338180 615494
rect 338304 615394 338404 615494
rect 338528 615394 338628 615494
rect 338752 615394 338852 615494
rect 338976 615394 339076 615494
rect 339200 615394 339300 615494
rect 339424 615394 339524 615494
rect 339648 615394 339748 615494
rect 339872 615394 339972 615494
rect 340096 615394 340196 615494
rect 340320 615394 340420 615494
rect 340544 615394 340644 615494
rect 340768 615394 340868 615494
rect 340992 615394 341092 615494
rect 341216 615394 341316 615494
rect 341440 615394 341540 615494
rect 341664 615394 341764 615494
rect 341888 615394 341988 615494
rect 342112 615394 342212 615494
rect 335616 615170 335716 615270
rect 335840 615170 335940 615270
rect 336064 615170 336164 615270
rect 336288 615170 336388 615270
rect 336512 615170 336612 615270
rect 336736 615170 336836 615270
rect 336960 615170 337060 615270
rect 337184 615170 337284 615270
rect 337408 615170 337508 615270
rect 337632 615170 337732 615270
rect 337856 615170 337956 615270
rect 338080 615170 338180 615270
rect 338304 615170 338404 615270
rect 338528 615170 338628 615270
rect 338752 615170 338852 615270
rect 338976 615170 339076 615270
rect 339200 615170 339300 615270
rect 339424 615170 339524 615270
rect 339648 615170 339748 615270
rect 339872 615170 339972 615270
rect 340096 615170 340196 615270
rect 340320 615170 340420 615270
rect 340544 615170 340644 615270
rect 340768 615170 340868 615270
rect 340992 615170 341092 615270
rect 341216 615170 341316 615270
rect 341440 615170 341540 615270
rect 341664 615170 341764 615270
rect 341888 615170 341988 615270
rect 342112 615170 342212 615270
rect 335616 614946 335716 615046
rect 335840 614946 335940 615046
rect 336064 614946 336164 615046
rect 336288 614946 336388 615046
rect 336512 614946 336612 615046
rect 336736 614946 336836 615046
rect 336960 614946 337060 615046
rect 337184 614946 337284 615046
rect 337408 614946 337508 615046
rect 337632 614946 337732 615046
rect 337856 614946 337956 615046
rect 338080 614946 338180 615046
rect 338304 614946 338404 615046
rect 338528 614946 338628 615046
rect 338752 614946 338852 615046
rect 338976 614946 339076 615046
rect 339200 614946 339300 615046
rect 339424 614946 339524 615046
rect 339648 614946 339748 615046
rect 339872 614946 339972 615046
rect 340096 614946 340196 615046
rect 340320 614946 340420 615046
rect 340544 614946 340644 615046
rect 340768 614946 340868 615046
rect 340992 614946 341092 615046
rect 341216 614946 341316 615046
rect 341440 614946 341540 615046
rect 341664 614946 341764 615046
rect 341888 614946 341988 615046
rect 342112 614946 342212 615046
rect 335616 614722 335716 614822
rect 335840 614722 335940 614822
rect 336064 614722 336164 614822
rect 336288 614722 336388 614822
rect 336512 614722 336612 614822
rect 336736 614722 336836 614822
rect 336960 614722 337060 614822
rect 337184 614722 337284 614822
rect 337408 614722 337508 614822
rect 337632 614722 337732 614822
rect 337856 614722 337956 614822
rect 338080 614722 338180 614822
rect 338304 614722 338404 614822
rect 338528 614722 338628 614822
rect 338752 614722 338852 614822
rect 338976 614722 339076 614822
rect 339200 614722 339300 614822
rect 339424 614722 339524 614822
rect 339648 614722 339748 614822
rect 339872 614722 339972 614822
rect 340096 614722 340196 614822
rect 340320 614722 340420 614822
rect 340544 614722 340644 614822
rect 340768 614722 340868 614822
rect 340992 614722 341092 614822
rect 341216 614722 341316 614822
rect 341440 614722 341540 614822
rect 341664 614722 341764 614822
rect 341888 614722 341988 614822
rect 342112 614722 342212 614822
rect 335616 614498 335716 614598
rect 335840 614498 335940 614598
rect 336064 614498 336164 614598
rect 336288 614498 336388 614598
rect 336512 614498 336612 614598
rect 336736 614498 336836 614598
rect 336960 614498 337060 614598
rect 337184 614498 337284 614598
rect 337408 614498 337508 614598
rect 337632 614498 337732 614598
rect 337856 614498 337956 614598
rect 338080 614498 338180 614598
rect 338304 614498 338404 614598
rect 338528 614498 338628 614598
rect 338752 614498 338852 614598
rect 338976 614498 339076 614598
rect 339200 614498 339300 614598
rect 339424 614498 339524 614598
rect 339648 614498 339748 614598
rect 339872 614498 339972 614598
rect 340096 614498 340196 614598
rect 340320 614498 340420 614598
rect 340544 614498 340644 614598
rect 340768 614498 340868 614598
rect 340992 614498 341092 614598
rect 341216 614498 341316 614598
rect 341440 614498 341540 614598
rect 341664 614498 341764 614598
rect 341888 614498 341988 614598
rect 342112 614498 342212 614598
rect 336480 605340 341264 611084
rect 510602 605017 515386 610761
rect 520602 684336 525386 690560
rect 520602 645217 525386 650961
rect 560582 639792 566726 644576
rect 520602 631817 525386 637561
rect 560582 629792 566726 634576
rect 520602 618417 525386 624161
rect 520602 605017 525386 610761
rect 317480 591580 322264 597324
rect 325480 591580 330264 597324
rect 13897 462422 13961 462486
rect 13977 462422 14041 462486
rect 14057 462422 14121 462486
rect 14137 462422 14201 462486
rect 14217 462422 14281 462486
rect 14297 462422 14361 462486
rect 14377 462422 14441 462486
rect 14457 462422 14521 462486
rect 14537 462422 14601 462486
rect 14617 462422 14681 462486
rect 14697 462422 14761 462486
rect 14777 462422 14841 462486
rect 14857 462422 14921 462486
rect 14937 462422 15001 462486
rect 15017 462422 15081 462486
rect 15097 462422 15161 462486
rect 15177 462422 15241 462486
rect 15257 462422 15321 462486
rect 15337 462422 15401 462486
rect 15417 462422 15481 462486
rect 15497 462422 15561 462486
rect 15577 462422 15641 462486
rect 15657 462422 15721 462486
rect 15737 462422 15801 462486
rect 15817 462422 15881 462486
rect 15897 462422 15961 462486
rect 15977 462422 16041 462486
rect 16057 462422 16121 462486
rect 16137 462422 16201 462486
rect 16217 462422 16281 462486
rect 16297 462422 16361 462486
rect 16377 462422 16441 462486
rect 16457 462422 16521 462486
rect 16537 462422 16601 462486
rect 16617 462422 16681 462486
rect 16697 462422 16761 462486
rect 16777 462422 16841 462486
rect 16857 462422 16921 462486
rect 16937 462422 17001 462486
rect 17017 462422 17081 462486
rect 17097 462422 17161 462486
rect 17177 462422 17241 462486
rect 17257 462422 17321 462486
rect 17337 462422 17401 462486
rect 17417 462422 17481 462486
rect 17497 462422 17561 462486
rect 13911 419200 13975 419264
rect 13991 419200 14055 419264
rect 14071 419200 14135 419264
rect 14151 419200 14215 419264
rect 14231 419200 14295 419264
rect 14311 419200 14375 419264
rect 14391 419200 14455 419264
rect 14471 419200 14535 419264
rect 14551 419200 14615 419264
rect 14631 419200 14695 419264
rect 14711 419200 14775 419264
rect 14791 419200 14855 419264
rect 14871 419200 14935 419264
rect 14951 419200 15015 419264
rect 15031 419200 15095 419264
rect 15111 419200 15175 419264
rect 15191 419200 15255 419264
rect 15271 419200 15335 419264
rect 15351 419200 15415 419264
rect 15431 419200 15495 419264
rect 15511 419200 15575 419264
rect 15591 419200 15655 419264
rect 15671 419200 15735 419264
rect 15751 419200 15815 419264
rect 15831 419200 15895 419264
rect 15911 419200 15975 419264
rect 15991 419200 16055 419264
rect 16071 419200 16135 419264
rect 16151 419200 16215 419264
rect 16231 419200 16295 419264
rect 16311 419200 16375 419264
rect 16391 419200 16455 419264
rect 16471 419200 16535 419264
rect 16551 419200 16615 419264
rect 16631 419200 16695 419264
rect 16711 419200 16775 419264
rect 16791 419200 16855 419264
rect 16871 419200 16935 419264
rect 16951 419200 17015 419264
rect 17031 419200 17095 419264
rect 17111 419200 17175 419264
rect 17191 419200 17255 419264
rect 17271 419200 17335 419264
rect 17351 419200 17415 419264
rect 17431 419200 17495 419264
rect 17511 419200 17575 419264
rect 556255 550570 562319 555354
rect 556255 540570 562319 545354
rect 573553 500074 573617 500138
rect 573633 500074 573697 500138
rect 573713 500074 573777 500138
rect 573793 500074 573857 500138
rect 573873 500074 573937 500138
rect 573953 500074 574017 500138
rect 574033 500074 574097 500138
rect 574113 500074 574177 500138
rect 574193 500074 574257 500138
rect 574273 500074 574337 500138
rect 574353 500074 574417 500138
rect 574433 500074 574497 500138
rect 574513 500074 574577 500138
rect 574593 500074 574657 500138
rect 574673 500074 574737 500138
rect 574753 500074 574817 500138
rect 574833 500074 574897 500138
rect 574913 500074 574977 500138
rect 574993 500074 575057 500138
rect 575073 500074 575137 500138
rect 575153 500074 575217 500138
rect 575233 500074 575297 500138
rect 575313 500074 575377 500138
rect 575393 500074 575457 500138
rect 575473 500074 575537 500138
rect 575553 500074 575617 500138
rect 575633 500074 575697 500138
rect 575713 500074 575777 500138
rect 575793 500074 575857 500138
rect 575873 500074 575937 500138
rect 575953 500074 576017 500138
rect 576033 500074 576097 500138
rect 576113 500074 576177 500138
rect 576193 500074 576257 500138
rect 576273 500074 576337 500138
rect 576353 500074 576417 500138
rect 576433 500074 576497 500138
rect 576513 500074 576577 500138
rect 576593 500074 576657 500138
rect 576673 500074 576737 500138
rect 573591 455652 573655 455716
rect 573671 455652 573735 455716
rect 573751 455652 573815 455716
rect 573831 455652 573895 455716
rect 573911 455652 573975 455716
rect 573991 455652 574055 455716
rect 574071 455652 574135 455716
rect 574151 455652 574215 455716
rect 574231 455652 574295 455716
rect 574311 455652 574375 455716
rect 574391 455652 574455 455716
rect 574471 455652 574535 455716
rect 574551 455652 574615 455716
rect 574631 455652 574695 455716
rect 574711 455652 574775 455716
rect 574791 455652 574855 455716
rect 574871 455652 574935 455716
rect 574951 455652 575015 455716
rect 575031 455652 575095 455716
rect 575111 455652 575175 455716
rect 575191 455652 575255 455716
rect 575271 455652 575335 455716
rect 575351 455652 575415 455716
rect 575431 455652 575495 455716
rect 575511 455652 575575 455716
rect 575591 455652 575655 455716
rect 575671 455652 575735 455716
rect 575751 455652 575815 455716
rect 575831 455652 575895 455716
rect 575911 455652 575975 455716
rect 575991 455652 576055 455716
rect 576071 455652 576135 455716
rect 576151 455652 576215 455716
rect 576231 455652 576295 455716
rect 576311 455652 576375 455716
rect 576391 455652 576455 455716
rect 576471 455652 576535 455716
rect 576551 455652 576615 455716
rect 576631 455652 576695 455716
rect 13997 191438 17421 196222
rect 573605 191438 576629 196222
<< mimcap >>
rect 304416 632032 304816 632072
rect 304416 631712 304456 632032
rect 304776 631712 304816 632032
rect 304416 631672 304816 631712
rect 305135 632032 305535 632072
rect 305135 631712 305175 632032
rect 305495 631712 305535 632032
rect 305135 631672 305535 631712
rect 305854 632032 306254 632072
rect 305854 631712 305894 632032
rect 306214 631712 306254 632032
rect 305854 631672 306254 631712
rect 306573 632032 306973 632072
rect 306573 631712 306613 632032
rect 306933 631712 306973 632032
rect 306573 631672 306973 631712
rect 307292 632032 307692 632072
rect 307292 631712 307332 632032
rect 307652 631712 307692 632032
rect 307292 631672 307692 631712
rect 308011 632032 308411 632072
rect 308011 631712 308051 632032
rect 308371 631712 308411 632032
rect 308011 631672 308411 631712
rect 308730 632032 309130 632072
rect 308730 631712 308770 632032
rect 309090 631712 309130 632032
rect 308730 631672 309130 631712
rect 309449 632032 309849 632072
rect 309449 631712 309489 632032
rect 309809 631712 309849 632032
rect 309449 631672 309849 631712
rect 310168 632032 310568 632072
rect 310168 631712 310208 632032
rect 310528 631712 310568 632032
rect 310168 631672 310568 631712
rect 310887 632032 311287 632072
rect 310887 631712 310927 632032
rect 311247 631712 311287 632032
rect 310887 631672 311287 631712
rect 304416 631332 304816 631372
rect 304416 631012 304456 631332
rect 304776 631012 304816 631332
rect 304416 630972 304816 631012
rect 305135 631332 305535 631372
rect 305135 631012 305175 631332
rect 305495 631012 305535 631332
rect 305135 630972 305535 631012
rect 305854 631332 306254 631372
rect 305854 631012 305894 631332
rect 306214 631012 306254 631332
rect 305854 630972 306254 631012
rect 306573 631332 306973 631372
rect 306573 631012 306613 631332
rect 306933 631012 306973 631332
rect 306573 630972 306973 631012
rect 307292 631332 307692 631372
rect 307292 631012 307332 631332
rect 307652 631012 307692 631332
rect 307292 630972 307692 631012
rect 308011 631332 308411 631372
rect 308011 631012 308051 631332
rect 308371 631012 308411 631332
rect 308011 630972 308411 631012
rect 308730 631332 309130 631372
rect 308730 631012 308770 631332
rect 309090 631012 309130 631332
rect 308730 630972 309130 631012
rect 309449 631332 309849 631372
rect 309449 631012 309489 631332
rect 309809 631012 309849 631332
rect 309449 630972 309849 631012
rect 310168 631332 310568 631372
rect 310168 631012 310208 631332
rect 310528 631012 310568 631332
rect 310168 630972 310568 631012
rect 310887 631332 311287 631372
rect 310887 631012 310927 631332
rect 311247 631012 311287 631332
rect 310887 630972 311287 631012
rect 304416 630632 304816 630672
rect 304416 630312 304456 630632
rect 304776 630312 304816 630632
rect 304416 630272 304816 630312
rect 305135 630632 305535 630672
rect 305135 630312 305175 630632
rect 305495 630312 305535 630632
rect 305135 630272 305535 630312
rect 305854 630632 306254 630672
rect 305854 630312 305894 630632
rect 306214 630312 306254 630632
rect 305854 630272 306254 630312
rect 306573 630632 306973 630672
rect 306573 630312 306613 630632
rect 306933 630312 306973 630632
rect 306573 630272 306973 630312
rect 307292 630632 307692 630672
rect 307292 630312 307332 630632
rect 307652 630312 307692 630632
rect 307292 630272 307692 630312
rect 308011 630632 308411 630672
rect 308011 630312 308051 630632
rect 308371 630312 308411 630632
rect 308011 630272 308411 630312
rect 308730 630632 309130 630672
rect 308730 630312 308770 630632
rect 309090 630312 309130 630632
rect 308730 630272 309130 630312
rect 309449 630632 309849 630672
rect 309449 630312 309489 630632
rect 309809 630312 309849 630632
rect 309449 630272 309849 630312
rect 310168 630632 310568 630672
rect 310168 630312 310208 630632
rect 310528 630312 310568 630632
rect 310168 630272 310568 630312
rect 310887 630632 311287 630672
rect 310887 630312 310927 630632
rect 311247 630312 311287 630632
rect 310887 630272 311287 630312
rect 304416 629932 304816 629972
rect 304416 629612 304456 629932
rect 304776 629612 304816 629932
rect 304416 629572 304816 629612
rect 305135 629932 305535 629972
rect 305135 629612 305175 629932
rect 305495 629612 305535 629932
rect 305135 629572 305535 629612
rect 305854 629932 306254 629972
rect 305854 629612 305894 629932
rect 306214 629612 306254 629932
rect 305854 629572 306254 629612
rect 306573 629932 306973 629972
rect 306573 629612 306613 629932
rect 306933 629612 306973 629932
rect 306573 629572 306973 629612
rect 307292 629932 307692 629972
rect 307292 629612 307332 629932
rect 307652 629612 307692 629932
rect 307292 629572 307692 629612
rect 308011 629932 308411 629972
rect 308011 629612 308051 629932
rect 308371 629612 308411 629932
rect 308011 629572 308411 629612
rect 308730 629932 309130 629972
rect 308730 629612 308770 629932
rect 309090 629612 309130 629932
rect 308730 629572 309130 629612
rect 309449 629932 309849 629972
rect 309449 629612 309489 629932
rect 309809 629612 309849 629932
rect 309449 629572 309849 629612
rect 310168 629932 310568 629972
rect 310168 629612 310208 629932
rect 310528 629612 310568 629932
rect 310168 629572 310568 629612
rect 310887 629932 311287 629972
rect 310887 629612 310927 629932
rect 311247 629612 311287 629932
rect 310887 629572 311287 629612
rect 304416 629232 304816 629272
rect 304416 628912 304456 629232
rect 304776 628912 304816 629232
rect 304416 628872 304816 628912
rect 305135 629232 305535 629272
rect 305135 628912 305175 629232
rect 305495 628912 305535 629232
rect 305135 628872 305535 628912
rect 305854 629232 306254 629272
rect 305854 628912 305894 629232
rect 306214 628912 306254 629232
rect 305854 628872 306254 628912
rect 306573 629232 306973 629272
rect 306573 628912 306613 629232
rect 306933 628912 306973 629232
rect 306573 628872 306973 628912
rect 307292 629232 307692 629272
rect 307292 628912 307332 629232
rect 307652 628912 307692 629232
rect 307292 628872 307692 628912
rect 308011 629232 308411 629272
rect 308011 628912 308051 629232
rect 308371 628912 308411 629232
rect 308011 628872 308411 628912
rect 308730 629232 309130 629272
rect 308730 628912 308770 629232
rect 309090 628912 309130 629232
rect 308730 628872 309130 628912
rect 309449 629232 309849 629272
rect 309449 628912 309489 629232
rect 309809 628912 309849 629232
rect 309449 628872 309849 628912
rect 310168 629232 310568 629272
rect 310168 628912 310208 629232
rect 310528 628912 310568 629232
rect 310168 628872 310568 628912
rect 310887 629232 311287 629272
rect 310887 628912 310927 629232
rect 311247 628912 311287 629232
rect 310887 628872 311287 628912
rect 304416 628532 304816 628572
rect 304416 628212 304456 628532
rect 304776 628212 304816 628532
rect 304416 628172 304816 628212
rect 305135 628532 305535 628572
rect 305135 628212 305175 628532
rect 305495 628212 305535 628532
rect 305135 628172 305535 628212
rect 305854 628532 306254 628572
rect 305854 628212 305894 628532
rect 306214 628212 306254 628532
rect 305854 628172 306254 628212
rect 306573 628532 306973 628572
rect 306573 628212 306613 628532
rect 306933 628212 306973 628532
rect 306573 628172 306973 628212
rect 307292 628532 307692 628572
rect 307292 628212 307332 628532
rect 307652 628212 307692 628532
rect 307292 628172 307692 628212
rect 308011 628532 308411 628572
rect 308011 628212 308051 628532
rect 308371 628212 308411 628532
rect 308011 628172 308411 628212
rect 308730 628532 309130 628572
rect 308730 628212 308770 628532
rect 309090 628212 309130 628532
rect 308730 628172 309130 628212
rect 309449 628532 309849 628572
rect 309449 628212 309489 628532
rect 309809 628212 309849 628532
rect 309449 628172 309849 628212
rect 310168 628532 310568 628572
rect 310168 628212 310208 628532
rect 310528 628212 310568 628532
rect 310168 628172 310568 628212
rect 310887 628532 311287 628572
rect 310887 628212 310927 628532
rect 311247 628212 311287 628532
rect 310887 628172 311287 628212
rect 304416 627832 304816 627872
rect 304416 627512 304456 627832
rect 304776 627512 304816 627832
rect 304416 627472 304816 627512
rect 305135 627832 305535 627872
rect 305135 627512 305175 627832
rect 305495 627512 305535 627832
rect 305135 627472 305535 627512
rect 305854 627832 306254 627872
rect 305854 627512 305894 627832
rect 306214 627512 306254 627832
rect 305854 627472 306254 627512
rect 306573 627832 306973 627872
rect 306573 627512 306613 627832
rect 306933 627512 306973 627832
rect 306573 627472 306973 627512
rect 307292 627832 307692 627872
rect 307292 627512 307332 627832
rect 307652 627512 307692 627832
rect 307292 627472 307692 627512
rect 308011 627832 308411 627872
rect 308011 627512 308051 627832
rect 308371 627512 308411 627832
rect 308011 627472 308411 627512
rect 308730 627832 309130 627872
rect 308730 627512 308770 627832
rect 309090 627512 309130 627832
rect 308730 627472 309130 627512
rect 309449 627832 309849 627872
rect 309449 627512 309489 627832
rect 309809 627512 309849 627832
rect 309449 627472 309849 627512
rect 310168 627832 310568 627872
rect 310168 627512 310208 627832
rect 310528 627512 310568 627832
rect 310168 627472 310568 627512
rect 310887 627832 311287 627872
rect 310887 627512 310927 627832
rect 311247 627512 311287 627832
rect 310887 627472 311287 627512
rect 304416 627132 304816 627172
rect 304416 626812 304456 627132
rect 304776 626812 304816 627132
rect 304416 626772 304816 626812
rect 305135 627132 305535 627172
rect 305135 626812 305175 627132
rect 305495 626812 305535 627132
rect 305135 626772 305535 626812
rect 305854 627132 306254 627172
rect 305854 626812 305894 627132
rect 306214 626812 306254 627132
rect 305854 626772 306254 626812
rect 306573 627132 306973 627172
rect 306573 626812 306613 627132
rect 306933 626812 306973 627132
rect 306573 626772 306973 626812
rect 307292 627132 307692 627172
rect 307292 626812 307332 627132
rect 307652 626812 307692 627132
rect 307292 626772 307692 626812
rect 308011 627132 308411 627172
rect 308011 626812 308051 627132
rect 308371 626812 308411 627132
rect 308011 626772 308411 626812
rect 308730 627132 309130 627172
rect 308730 626812 308770 627132
rect 309090 626812 309130 627132
rect 308730 626772 309130 626812
rect 309449 627132 309849 627172
rect 309449 626812 309489 627132
rect 309809 626812 309849 627132
rect 309449 626772 309849 626812
rect 310168 627132 310568 627172
rect 310168 626812 310208 627132
rect 310528 626812 310568 627132
rect 310168 626772 310568 626812
rect 310887 627132 311287 627172
rect 310887 626812 310927 627132
rect 311247 626812 311287 627132
rect 310887 626772 311287 626812
rect 304416 626432 304816 626472
rect 304416 626112 304456 626432
rect 304776 626112 304816 626432
rect 304416 626072 304816 626112
rect 305135 626432 305535 626472
rect 305135 626112 305175 626432
rect 305495 626112 305535 626432
rect 305135 626072 305535 626112
rect 305854 626432 306254 626472
rect 305854 626112 305894 626432
rect 306214 626112 306254 626432
rect 305854 626072 306254 626112
rect 306573 626432 306973 626472
rect 306573 626112 306613 626432
rect 306933 626112 306973 626432
rect 306573 626072 306973 626112
rect 307292 626432 307692 626472
rect 307292 626112 307332 626432
rect 307652 626112 307692 626432
rect 307292 626072 307692 626112
rect 308011 626432 308411 626472
rect 308011 626112 308051 626432
rect 308371 626112 308411 626432
rect 308011 626072 308411 626112
rect 308730 626432 309130 626472
rect 308730 626112 308770 626432
rect 309090 626112 309130 626432
rect 308730 626072 309130 626112
rect 309449 626432 309849 626472
rect 309449 626112 309489 626432
rect 309809 626112 309849 626432
rect 309449 626072 309849 626112
rect 310168 626432 310568 626472
rect 310168 626112 310208 626432
rect 310528 626112 310568 626432
rect 310168 626072 310568 626112
rect 310887 626432 311287 626472
rect 310887 626112 310927 626432
rect 311247 626112 311287 626432
rect 310887 626072 311287 626112
rect 304416 625732 304816 625772
rect 304416 625412 304456 625732
rect 304776 625412 304816 625732
rect 304416 625372 304816 625412
rect 305135 625732 305535 625772
rect 305135 625412 305175 625732
rect 305495 625412 305535 625732
rect 305135 625372 305535 625412
rect 305854 625732 306254 625772
rect 305854 625412 305894 625732
rect 306214 625412 306254 625732
rect 305854 625372 306254 625412
rect 306573 625732 306973 625772
rect 306573 625412 306613 625732
rect 306933 625412 306973 625732
rect 306573 625372 306973 625412
rect 307292 625732 307692 625772
rect 307292 625412 307332 625732
rect 307652 625412 307692 625732
rect 307292 625372 307692 625412
rect 308011 625732 308411 625772
rect 308011 625412 308051 625732
rect 308371 625412 308411 625732
rect 308011 625372 308411 625412
rect 308730 625732 309130 625772
rect 308730 625412 308770 625732
rect 309090 625412 309130 625732
rect 308730 625372 309130 625412
rect 309449 625732 309849 625772
rect 309449 625412 309489 625732
rect 309809 625412 309849 625732
rect 309449 625372 309849 625412
rect 310168 625732 310568 625772
rect 310168 625412 310208 625732
rect 310528 625412 310568 625732
rect 310168 625372 310568 625412
rect 310887 625732 311287 625772
rect 310887 625412 310927 625732
rect 311247 625412 311287 625732
rect 310887 625372 311287 625412
<< mimcapcontact >>
rect 304456 631712 304776 632032
rect 305175 631712 305495 632032
rect 305894 631712 306214 632032
rect 306613 631712 306933 632032
rect 307332 631712 307652 632032
rect 308051 631712 308371 632032
rect 308770 631712 309090 632032
rect 309489 631712 309809 632032
rect 310208 631712 310528 632032
rect 310927 631712 311247 632032
rect 304456 631012 304776 631332
rect 305175 631012 305495 631332
rect 305894 631012 306214 631332
rect 306613 631012 306933 631332
rect 307332 631012 307652 631332
rect 308051 631012 308371 631332
rect 308770 631012 309090 631332
rect 309489 631012 309809 631332
rect 310208 631012 310528 631332
rect 310927 631012 311247 631332
rect 304456 630312 304776 630632
rect 305175 630312 305495 630632
rect 305894 630312 306214 630632
rect 306613 630312 306933 630632
rect 307332 630312 307652 630632
rect 308051 630312 308371 630632
rect 308770 630312 309090 630632
rect 309489 630312 309809 630632
rect 310208 630312 310528 630632
rect 310927 630312 311247 630632
rect 304456 629612 304776 629932
rect 305175 629612 305495 629932
rect 305894 629612 306214 629932
rect 306613 629612 306933 629932
rect 307332 629612 307652 629932
rect 308051 629612 308371 629932
rect 308770 629612 309090 629932
rect 309489 629612 309809 629932
rect 310208 629612 310528 629932
rect 310927 629612 311247 629932
rect 304456 628912 304776 629232
rect 305175 628912 305495 629232
rect 305894 628912 306214 629232
rect 306613 628912 306933 629232
rect 307332 628912 307652 629232
rect 308051 628912 308371 629232
rect 308770 628912 309090 629232
rect 309489 628912 309809 629232
rect 310208 628912 310528 629232
rect 310927 628912 311247 629232
rect 304456 628212 304776 628532
rect 305175 628212 305495 628532
rect 305894 628212 306214 628532
rect 306613 628212 306933 628532
rect 307332 628212 307652 628532
rect 308051 628212 308371 628532
rect 308770 628212 309090 628532
rect 309489 628212 309809 628532
rect 310208 628212 310528 628532
rect 310927 628212 311247 628532
rect 304456 627512 304776 627832
rect 305175 627512 305495 627832
rect 305894 627512 306214 627832
rect 306613 627512 306933 627832
rect 307332 627512 307652 627832
rect 308051 627512 308371 627832
rect 308770 627512 309090 627832
rect 309489 627512 309809 627832
rect 310208 627512 310528 627832
rect 310927 627512 311247 627832
rect 304456 626812 304776 627132
rect 305175 626812 305495 627132
rect 305894 626812 306214 627132
rect 306613 626812 306933 627132
rect 307332 626812 307652 627132
rect 308051 626812 308371 627132
rect 308770 626812 309090 627132
rect 309489 626812 309809 627132
rect 310208 626812 310528 627132
rect 310927 626812 311247 627132
rect 304456 626112 304776 626432
rect 305175 626112 305495 626432
rect 305894 626112 306214 626432
rect 306613 626112 306933 626432
rect 307332 626112 307652 626432
rect 308051 626112 308371 626432
rect 308770 626112 309090 626432
rect 309489 626112 309809 626432
rect 310208 626112 310528 626432
rect 310927 626112 311247 626432
rect 304456 625412 304776 625732
rect 305175 625412 305495 625732
rect 305894 625412 306214 625732
rect 306613 625412 306933 625732
rect 307332 625412 307652 625732
rect 308051 625412 308371 625732
rect 308770 625412 309090 625732
rect 309489 625412 309809 625732
rect 310208 625412 310528 625732
rect 310927 625412 311247 625732
<< metal4 >>
rect 170628 690610 526162 690737
rect 170628 690577 222622 690610
rect 170628 684353 170922 690577
rect 173066 684353 173422 690577
rect 175566 684386 222622 690577
rect 224766 690593 526162 690610
rect 224766 690084 324322 690593
rect 224766 684386 289800 690084
rect 175566 684353 289800 684386
rect 170628 684340 289800 684353
rect 294584 684369 324322 690084
rect 326466 690560 526162 690593
rect 326466 684369 510602 690560
rect 294584 684340 510602 684369
rect 170628 684336 510602 684340
rect 515386 684336 520602 690560
rect 525386 684336 526162 690560
rect 170628 684183 526162 684336
rect 343420 651400 525804 651406
rect 285800 650961 525804 651400
rect 285800 650904 510602 650961
rect 285800 650584 336480 650904
rect 285800 644840 289920 650584
rect 294704 644840 298920 650584
rect 303704 644840 304920 650584
rect 309704 644840 310920 650584
rect 315704 645160 336480 650584
rect 341264 645217 510602 650904
rect 515386 645217 520602 650961
rect 525386 645217 525804 650961
rect 341264 645160 525804 645217
rect 315704 644840 525804 645160
rect 285800 644744 525804 644840
rect 560425 644576 566979 644980
rect 335560 642719 342216 642724
rect 335560 642714 342217 642719
rect 298820 642699 305476 642704
rect 309290 642699 315946 642704
rect 298820 642694 305477 642699
rect 298820 642594 298876 642694
rect 298976 642594 299100 642694
rect 299200 642594 299324 642694
rect 299424 642594 299548 642694
rect 299648 642594 299772 642694
rect 299872 642594 299996 642694
rect 300096 642594 300220 642694
rect 300320 642594 300444 642694
rect 300544 642594 300668 642694
rect 300768 642594 300892 642694
rect 300992 642594 301116 642694
rect 301216 642594 301340 642694
rect 301440 642594 301564 642694
rect 301664 642594 301788 642694
rect 301888 642594 302012 642694
rect 302112 642594 302236 642694
rect 302336 642594 302460 642694
rect 302560 642594 302684 642694
rect 302784 642594 302908 642694
rect 303008 642594 303132 642694
rect 303232 642594 303356 642694
rect 303456 642594 303580 642694
rect 303680 642594 303804 642694
rect 303904 642594 304028 642694
rect 304128 642594 304252 642694
rect 304352 642594 304476 642694
rect 304576 642594 304700 642694
rect 304800 642594 304924 642694
rect 305024 642594 305148 642694
rect 305248 642594 305372 642694
rect 305472 642594 305477 642694
rect 298820 642589 305477 642594
rect 309290 642694 315947 642699
rect 309290 642594 309346 642694
rect 309446 642594 309570 642694
rect 309670 642594 309794 642694
rect 309894 642594 310018 642694
rect 310118 642594 310242 642694
rect 310342 642594 310466 642694
rect 310566 642594 310690 642694
rect 310790 642594 310914 642694
rect 311014 642594 311138 642694
rect 311238 642594 311362 642694
rect 311462 642594 311586 642694
rect 311686 642594 311810 642694
rect 311910 642594 312034 642694
rect 312134 642594 312258 642694
rect 312358 642594 312482 642694
rect 312582 642594 312706 642694
rect 312806 642594 312930 642694
rect 313030 642594 313154 642694
rect 313254 642594 313378 642694
rect 313478 642594 313602 642694
rect 313702 642594 313826 642694
rect 313926 642594 314050 642694
rect 314150 642594 314274 642694
rect 314374 642594 314498 642694
rect 314598 642594 314722 642694
rect 314822 642594 314946 642694
rect 315046 642594 315170 642694
rect 315270 642594 315394 642694
rect 315494 642594 315618 642694
rect 315718 642594 315842 642694
rect 315942 642594 315947 642694
rect 309290 642589 315947 642594
rect 335560 642614 335616 642714
rect 335716 642614 335840 642714
rect 335940 642614 336064 642714
rect 336164 642614 336288 642714
rect 336388 642614 336512 642714
rect 336612 642614 336736 642714
rect 336836 642614 336960 642714
rect 337060 642614 337184 642714
rect 337284 642614 337408 642714
rect 337508 642614 337632 642714
rect 337732 642614 337856 642714
rect 337956 642614 338080 642714
rect 338180 642614 338304 642714
rect 338404 642614 338528 642714
rect 338628 642614 338752 642714
rect 338852 642614 338976 642714
rect 339076 642614 339200 642714
rect 339300 642614 339424 642714
rect 339524 642614 339648 642714
rect 339748 642614 339872 642714
rect 339972 642614 340096 642714
rect 340196 642614 340320 642714
rect 340420 642614 340544 642714
rect 340644 642614 340768 642714
rect 340868 642614 340992 642714
rect 341092 642614 341216 642714
rect 341316 642614 341440 642714
rect 341540 642614 341664 642714
rect 341764 642614 341888 642714
rect 341988 642614 342112 642714
rect 342212 642614 342217 642714
rect 335560 642609 342217 642614
rect 298820 642475 305476 642589
rect 309290 642475 315946 642589
rect 335560 642495 342216 642609
rect 335560 642490 342217 642495
rect 298820 642470 305477 642475
rect 298820 642370 298876 642470
rect 298976 642370 299100 642470
rect 299200 642370 299324 642470
rect 299424 642370 299548 642470
rect 299648 642370 299772 642470
rect 299872 642370 299996 642470
rect 300096 642370 300220 642470
rect 300320 642370 300444 642470
rect 300544 642370 300668 642470
rect 300768 642370 300892 642470
rect 300992 642370 301116 642470
rect 301216 642370 301340 642470
rect 301440 642370 301564 642470
rect 301664 642370 301788 642470
rect 301888 642370 302012 642470
rect 302112 642370 302236 642470
rect 302336 642370 302460 642470
rect 302560 642370 302684 642470
rect 302784 642370 302908 642470
rect 303008 642370 303132 642470
rect 303232 642370 303356 642470
rect 303456 642370 303580 642470
rect 303680 642370 303804 642470
rect 303904 642370 304028 642470
rect 304128 642370 304252 642470
rect 304352 642370 304476 642470
rect 304576 642370 304700 642470
rect 304800 642370 304924 642470
rect 305024 642370 305148 642470
rect 305248 642370 305372 642470
rect 305472 642370 305477 642470
rect 298820 642365 305477 642370
rect 309290 642470 315947 642475
rect 309290 642370 309346 642470
rect 309446 642370 309570 642470
rect 309670 642370 309794 642470
rect 309894 642370 310018 642470
rect 310118 642370 310242 642470
rect 310342 642370 310466 642470
rect 310566 642370 310690 642470
rect 310790 642370 310914 642470
rect 311014 642370 311138 642470
rect 311238 642370 311362 642470
rect 311462 642370 311586 642470
rect 311686 642370 311810 642470
rect 311910 642370 312034 642470
rect 312134 642370 312258 642470
rect 312358 642370 312482 642470
rect 312582 642370 312706 642470
rect 312806 642370 312930 642470
rect 313030 642370 313154 642470
rect 313254 642370 313378 642470
rect 313478 642370 313602 642470
rect 313702 642370 313826 642470
rect 313926 642370 314050 642470
rect 314150 642370 314274 642470
rect 314374 642370 314498 642470
rect 314598 642370 314722 642470
rect 314822 642370 314946 642470
rect 315046 642370 315170 642470
rect 315270 642370 315394 642470
rect 315494 642370 315618 642470
rect 315718 642370 315842 642470
rect 315942 642370 315947 642470
rect 309290 642365 315947 642370
rect 335560 642390 335616 642490
rect 335716 642390 335840 642490
rect 335940 642390 336064 642490
rect 336164 642390 336288 642490
rect 336388 642390 336512 642490
rect 336612 642390 336736 642490
rect 336836 642390 336960 642490
rect 337060 642390 337184 642490
rect 337284 642390 337408 642490
rect 337508 642390 337632 642490
rect 337732 642390 337856 642490
rect 337956 642390 338080 642490
rect 338180 642390 338304 642490
rect 338404 642390 338528 642490
rect 338628 642390 338752 642490
rect 338852 642390 338976 642490
rect 339076 642390 339200 642490
rect 339300 642390 339424 642490
rect 339524 642390 339648 642490
rect 339748 642390 339872 642490
rect 339972 642390 340096 642490
rect 340196 642390 340320 642490
rect 340420 642390 340544 642490
rect 340644 642390 340768 642490
rect 340868 642390 340992 642490
rect 341092 642390 341216 642490
rect 341316 642390 341440 642490
rect 341540 642390 341664 642490
rect 341764 642390 341888 642490
rect 341988 642390 342112 642490
rect 342212 642390 342217 642490
rect 335560 642385 342217 642390
rect 298820 642251 305476 642365
rect 309290 642251 315946 642365
rect 335560 642271 342216 642385
rect 335560 642266 342217 642271
rect 298820 642246 305477 642251
rect 298820 642146 298876 642246
rect 298976 642146 299100 642246
rect 299200 642146 299324 642246
rect 299424 642146 299548 642246
rect 299648 642146 299772 642246
rect 299872 642146 299996 642246
rect 300096 642146 300220 642246
rect 300320 642146 300444 642246
rect 300544 642146 300668 642246
rect 300768 642146 300892 642246
rect 300992 642146 301116 642246
rect 301216 642146 301340 642246
rect 301440 642146 301564 642246
rect 301664 642146 301788 642246
rect 301888 642146 302012 642246
rect 302112 642146 302236 642246
rect 302336 642146 302460 642246
rect 302560 642146 302684 642246
rect 302784 642146 302908 642246
rect 303008 642146 303132 642246
rect 303232 642146 303356 642246
rect 303456 642146 303580 642246
rect 303680 642146 303804 642246
rect 303904 642146 304028 642246
rect 304128 642146 304252 642246
rect 304352 642146 304476 642246
rect 304576 642146 304700 642246
rect 304800 642146 304924 642246
rect 305024 642146 305148 642246
rect 305248 642146 305372 642246
rect 305472 642146 305477 642246
rect 298820 642141 305477 642146
rect 309290 642246 315947 642251
rect 309290 642146 309346 642246
rect 309446 642146 309570 642246
rect 309670 642146 309794 642246
rect 309894 642146 310018 642246
rect 310118 642146 310242 642246
rect 310342 642146 310466 642246
rect 310566 642146 310690 642246
rect 310790 642146 310914 642246
rect 311014 642146 311138 642246
rect 311238 642146 311362 642246
rect 311462 642146 311586 642246
rect 311686 642146 311810 642246
rect 311910 642146 312034 642246
rect 312134 642146 312258 642246
rect 312358 642146 312482 642246
rect 312582 642146 312706 642246
rect 312806 642146 312930 642246
rect 313030 642146 313154 642246
rect 313254 642146 313378 642246
rect 313478 642146 313602 642246
rect 313702 642146 313826 642246
rect 313926 642146 314050 642246
rect 314150 642146 314274 642246
rect 314374 642146 314498 642246
rect 314598 642146 314722 642246
rect 314822 642146 314946 642246
rect 315046 642146 315170 642246
rect 315270 642146 315394 642246
rect 315494 642146 315618 642246
rect 315718 642146 315842 642246
rect 315942 642146 315947 642246
rect 309290 642141 315947 642146
rect 335560 642166 335616 642266
rect 335716 642166 335840 642266
rect 335940 642166 336064 642266
rect 336164 642166 336288 642266
rect 336388 642166 336512 642266
rect 336612 642166 336736 642266
rect 336836 642166 336960 642266
rect 337060 642166 337184 642266
rect 337284 642166 337408 642266
rect 337508 642166 337632 642266
rect 337732 642166 337856 642266
rect 337956 642166 338080 642266
rect 338180 642166 338304 642266
rect 338404 642166 338528 642266
rect 338628 642166 338752 642266
rect 338852 642166 338976 642266
rect 339076 642166 339200 642266
rect 339300 642166 339424 642266
rect 339524 642166 339648 642266
rect 339748 642166 339872 642266
rect 339972 642166 340096 642266
rect 340196 642166 340320 642266
rect 340420 642166 340544 642266
rect 340644 642166 340768 642266
rect 340868 642166 340992 642266
rect 341092 642166 341216 642266
rect 341316 642166 341440 642266
rect 341540 642166 341664 642266
rect 341764 642166 341888 642266
rect 341988 642166 342112 642266
rect 342212 642166 342217 642266
rect 335560 642161 342217 642166
rect 298820 642027 305476 642141
rect 309290 642027 315946 642141
rect 335560 642047 342216 642161
rect 335560 642042 342217 642047
rect 298820 642022 305477 642027
rect 298820 641922 298876 642022
rect 298976 641922 299100 642022
rect 299200 641922 299324 642022
rect 299424 641922 299548 642022
rect 299648 641922 299772 642022
rect 299872 641922 299996 642022
rect 300096 641922 300220 642022
rect 300320 641922 300444 642022
rect 300544 641922 300668 642022
rect 300768 641922 300892 642022
rect 300992 641922 301116 642022
rect 301216 641922 301340 642022
rect 301440 641922 301564 642022
rect 301664 641922 301788 642022
rect 301888 641922 302012 642022
rect 302112 641922 302236 642022
rect 302336 641922 302460 642022
rect 302560 641922 302684 642022
rect 302784 641922 302908 642022
rect 303008 641922 303132 642022
rect 303232 641922 303356 642022
rect 303456 641922 303580 642022
rect 303680 641922 303804 642022
rect 303904 641922 304028 642022
rect 304128 641922 304252 642022
rect 304352 641922 304476 642022
rect 304576 641922 304700 642022
rect 304800 641922 304924 642022
rect 305024 641922 305148 642022
rect 305248 641922 305372 642022
rect 305472 641922 305477 642022
rect 298820 641917 305477 641922
rect 309290 642022 315947 642027
rect 309290 641922 309346 642022
rect 309446 641922 309570 642022
rect 309670 641922 309794 642022
rect 309894 641922 310018 642022
rect 310118 641922 310242 642022
rect 310342 641922 310466 642022
rect 310566 641922 310690 642022
rect 310790 641922 310914 642022
rect 311014 641922 311138 642022
rect 311238 641922 311362 642022
rect 311462 641922 311586 642022
rect 311686 641922 311810 642022
rect 311910 641922 312034 642022
rect 312134 641922 312258 642022
rect 312358 641922 312482 642022
rect 312582 641922 312706 642022
rect 312806 641922 312930 642022
rect 313030 641922 313154 642022
rect 313254 641922 313378 642022
rect 313478 641922 313602 642022
rect 313702 641922 313826 642022
rect 313926 641922 314050 642022
rect 314150 641922 314274 642022
rect 314374 641922 314498 642022
rect 314598 641922 314722 642022
rect 314822 641922 314946 642022
rect 315046 641922 315170 642022
rect 315270 641922 315394 642022
rect 315494 641922 315618 642022
rect 315718 641922 315842 642022
rect 315942 641922 315947 642022
rect 309290 641917 315947 641922
rect 335560 641942 335616 642042
rect 335716 641942 335840 642042
rect 335940 641942 336064 642042
rect 336164 641942 336288 642042
rect 336388 641942 336512 642042
rect 336612 641942 336736 642042
rect 336836 641942 336960 642042
rect 337060 641942 337184 642042
rect 337284 641942 337408 642042
rect 337508 641942 337632 642042
rect 337732 641942 337856 642042
rect 337956 641942 338080 642042
rect 338180 641942 338304 642042
rect 338404 641942 338528 642042
rect 338628 641942 338752 642042
rect 338852 641942 338976 642042
rect 339076 641942 339200 642042
rect 339300 641942 339424 642042
rect 339524 641942 339648 642042
rect 339748 641942 339872 642042
rect 339972 641942 340096 642042
rect 340196 641942 340320 642042
rect 340420 641942 340544 642042
rect 340644 641942 340768 642042
rect 340868 641942 340992 642042
rect 341092 641942 341216 642042
rect 341316 641942 341440 642042
rect 341540 641942 341664 642042
rect 341764 641942 341888 642042
rect 341988 641942 342112 642042
rect 342212 641942 342217 642042
rect 335560 641937 342217 641942
rect 298820 641803 305476 641917
rect 309290 641803 315946 641917
rect 335560 641823 342216 641937
rect 335560 641818 342217 641823
rect 298820 641798 305477 641803
rect 298820 641698 298876 641798
rect 298976 641698 299100 641798
rect 299200 641698 299324 641798
rect 299424 641698 299548 641798
rect 299648 641698 299772 641798
rect 299872 641698 299996 641798
rect 300096 641698 300220 641798
rect 300320 641698 300444 641798
rect 300544 641698 300668 641798
rect 300768 641698 300892 641798
rect 300992 641698 301116 641798
rect 301216 641698 301340 641798
rect 301440 641698 301564 641798
rect 301664 641698 301788 641798
rect 301888 641698 302012 641798
rect 302112 641698 302236 641798
rect 302336 641698 302460 641798
rect 302560 641698 302684 641798
rect 302784 641698 302908 641798
rect 303008 641698 303132 641798
rect 303232 641698 303356 641798
rect 303456 641698 303580 641798
rect 303680 641698 303804 641798
rect 303904 641698 304028 641798
rect 304128 641698 304252 641798
rect 304352 641698 304476 641798
rect 304576 641698 304700 641798
rect 304800 641698 304924 641798
rect 305024 641698 305148 641798
rect 305248 641698 305372 641798
rect 305472 641698 305477 641798
rect 298820 641693 305477 641698
rect 309290 641798 315947 641803
rect 309290 641698 309346 641798
rect 309446 641698 309570 641798
rect 309670 641698 309794 641798
rect 309894 641698 310018 641798
rect 310118 641698 310242 641798
rect 310342 641698 310466 641798
rect 310566 641698 310690 641798
rect 310790 641698 310914 641798
rect 311014 641698 311138 641798
rect 311238 641698 311362 641798
rect 311462 641698 311586 641798
rect 311686 641698 311810 641798
rect 311910 641698 312034 641798
rect 312134 641698 312258 641798
rect 312358 641698 312482 641798
rect 312582 641698 312706 641798
rect 312806 641698 312930 641798
rect 313030 641698 313154 641798
rect 313254 641698 313378 641798
rect 313478 641698 313602 641798
rect 313702 641698 313826 641798
rect 313926 641698 314050 641798
rect 314150 641698 314274 641798
rect 314374 641698 314498 641798
rect 314598 641698 314722 641798
rect 314822 641698 314946 641798
rect 315046 641698 315170 641798
rect 315270 641698 315394 641798
rect 315494 641698 315618 641798
rect 315718 641698 315842 641798
rect 315942 641698 315947 641798
rect 309290 641693 315947 641698
rect 335560 641718 335616 641818
rect 335716 641718 335840 641818
rect 335940 641718 336064 641818
rect 336164 641718 336288 641818
rect 336388 641718 336512 641818
rect 336612 641718 336736 641818
rect 336836 641718 336960 641818
rect 337060 641718 337184 641818
rect 337284 641718 337408 641818
rect 337508 641718 337632 641818
rect 337732 641718 337856 641818
rect 337956 641718 338080 641818
rect 338180 641718 338304 641818
rect 338404 641718 338528 641818
rect 338628 641718 338752 641818
rect 338852 641718 338976 641818
rect 339076 641718 339200 641818
rect 339300 641718 339424 641818
rect 339524 641718 339648 641818
rect 339748 641718 339872 641818
rect 339972 641718 340096 641818
rect 340196 641718 340320 641818
rect 340420 641718 340544 641818
rect 340644 641718 340768 641818
rect 340868 641718 340992 641818
rect 341092 641718 341216 641818
rect 341316 641718 341440 641818
rect 341540 641718 341664 641818
rect 341764 641718 341888 641818
rect 341988 641718 342112 641818
rect 342212 641718 342217 641818
rect 335560 641713 342217 641718
rect 298820 641664 305476 641693
rect 309290 641664 315946 641693
rect 335560 641684 342216 641713
rect 300626 640587 311952 640624
rect 300626 639731 300643 640587
rect 311917 639731 311952 640587
rect 289020 637996 298880 638020
rect 289020 637896 297850 637996
rect 297950 637896 298074 637996
rect 298174 637896 298298 637996
rect 298398 637896 298522 637996
rect 298622 637896 298746 637996
rect 298846 637896 298880 637996
rect 289020 637772 298880 637896
rect 289020 637672 297850 637772
rect 297950 637672 298074 637772
rect 298174 637672 298298 637772
rect 298398 637672 298522 637772
rect 298622 637672 298746 637772
rect 298846 637672 298880 637772
rect 289020 637548 298880 637672
rect 289020 637448 297850 637548
rect 297950 637448 298074 637548
rect 298174 637448 298298 637548
rect 298398 637448 298522 637548
rect 298622 637448 298746 637548
rect 298846 637448 298880 637548
rect 289020 637324 298880 637448
rect 289020 637224 297850 637324
rect 297950 637224 298074 637324
rect 298174 637224 298298 637324
rect 298398 637224 298522 637324
rect 298622 637224 298746 637324
rect 298846 637224 298880 637324
rect 289020 637184 298880 637224
rect 289020 631440 289920 637184
rect 294704 637100 298880 637184
rect 294704 637000 297850 637100
rect 297950 637000 298074 637100
rect 298174 637000 298298 637100
rect 298398 637000 298522 637100
rect 298622 637000 298746 637100
rect 298846 637000 298880 637100
rect 294704 636876 298880 637000
rect 294704 636776 297850 636876
rect 297950 636776 298074 636876
rect 298174 636776 298298 636876
rect 298398 636776 298522 636876
rect 298622 636776 298746 636876
rect 298846 636776 298880 636876
rect 294704 636652 298880 636776
rect 294704 636552 297850 636652
rect 297950 636552 298074 636652
rect 298174 636552 298298 636652
rect 298398 636552 298522 636652
rect 298622 636552 298746 636652
rect 298846 636552 298880 636652
rect 294704 636428 298880 636552
rect 294704 636328 297850 636428
rect 297950 636328 298074 636428
rect 298174 636328 298298 636428
rect 298398 636328 298522 636428
rect 298622 636328 298746 636428
rect 298846 636328 298880 636428
rect 294704 636204 298880 636328
rect 294704 636104 297850 636204
rect 297950 636104 298074 636204
rect 298174 636104 298298 636204
rect 298398 636104 298522 636204
rect 298622 636104 298746 636204
rect 298846 636104 298880 636204
rect 294704 635980 298880 636104
rect 294704 635880 297850 635980
rect 297950 635880 298074 635980
rect 298174 635880 298298 635980
rect 298398 635880 298522 635980
rect 298622 635880 298746 635980
rect 298846 635880 298880 635980
rect 294704 635756 298880 635880
rect 294704 635656 297850 635756
rect 297950 635656 298074 635756
rect 298174 635656 298298 635756
rect 298398 635656 298522 635756
rect 298622 635656 298746 635756
rect 298846 635656 298880 635756
rect 294704 635532 298880 635656
rect 294704 635432 297850 635532
rect 297950 635432 298074 635532
rect 298174 635432 298298 635532
rect 298398 635432 298522 635532
rect 298622 635432 298746 635532
rect 298846 635432 298880 635532
rect 294704 635308 298880 635432
rect 294704 635208 297850 635308
rect 297950 635208 298074 635308
rect 298174 635208 298298 635308
rect 298398 635208 298522 635308
rect 298622 635208 298746 635308
rect 298846 635208 298880 635308
rect 294704 635084 298880 635208
rect 294704 634984 297850 635084
rect 297950 634984 298074 635084
rect 298174 634984 298298 635084
rect 298398 634984 298522 635084
rect 298622 634984 298746 635084
rect 298846 634984 298880 635084
rect 294704 634860 298880 634984
rect 294704 634760 297850 634860
rect 297950 634760 298074 634860
rect 298174 634760 298298 634860
rect 298398 634760 298522 634860
rect 298622 634760 298746 634860
rect 298846 634760 298880 634860
rect 294704 634636 298880 634760
rect 294704 634536 297850 634636
rect 297950 634536 298074 634636
rect 298174 634536 298298 634636
rect 298398 634536 298522 634636
rect 298622 634536 298746 634636
rect 298846 634536 298880 634636
rect 294704 634412 298880 634536
rect 294704 634312 297850 634412
rect 297950 634312 298074 634412
rect 298174 634312 298298 634412
rect 298398 634312 298522 634412
rect 298622 634312 298746 634412
rect 298846 634312 298880 634412
rect 294704 634188 298880 634312
rect 294704 634088 297850 634188
rect 297950 634088 298074 634188
rect 298174 634088 298298 634188
rect 298398 634088 298522 634188
rect 298622 634088 298746 634188
rect 298846 634088 298880 634188
rect 294704 633964 298880 634088
rect 294704 633864 297850 633964
rect 297950 633864 298074 633964
rect 298174 633864 298298 633964
rect 298398 633864 298522 633964
rect 298622 633864 298746 633964
rect 298846 633864 298880 633964
rect 294704 633740 298880 633864
rect 294704 633640 297850 633740
rect 297950 633640 298074 633740
rect 298174 633640 298298 633740
rect 298398 633640 298522 633740
rect 298622 633640 298746 633740
rect 298846 633640 298880 633740
rect 294704 633516 298880 633640
rect 294704 633416 297850 633516
rect 297950 633416 298074 633516
rect 298174 633416 298298 633516
rect 298398 633416 298522 633516
rect 298622 633416 298746 633516
rect 298846 633416 298880 633516
rect 294704 633292 298880 633416
rect 294704 633192 297850 633292
rect 297950 633192 298074 633292
rect 298174 633192 298298 633292
rect 298398 633192 298522 633292
rect 298622 633192 298746 633292
rect 298846 633192 298880 633292
rect 294704 633068 298880 633192
rect 294704 632968 297850 633068
rect 297950 632968 298074 633068
rect 298174 632968 298298 633068
rect 298398 632968 298522 633068
rect 298622 632968 298746 633068
rect 298846 632968 298880 633068
rect 294704 632844 298880 632968
rect 294704 632744 297850 632844
rect 297950 632744 298074 632844
rect 298174 632744 298298 632844
rect 298398 632744 298522 632844
rect 298622 632744 298746 632844
rect 298846 632744 298880 632844
rect 294704 632620 298880 632744
rect 294704 632520 297850 632620
rect 297950 632520 298074 632620
rect 298174 632520 298298 632620
rect 298398 632520 298522 632620
rect 298622 632520 298746 632620
rect 298846 632520 298880 632620
rect 294704 632396 298880 632520
rect 300626 632462 311952 639731
rect 560425 639792 560582 644576
rect 566726 639792 566979 644576
rect 342125 638000 342235 638001
rect 342349 638000 342459 638001
rect 342573 638000 342683 638001
rect 342797 638000 342907 638001
rect 343021 638000 343131 638001
rect 300672 632456 311952 632462
rect 341994 637996 525800 638000
rect 341994 637896 342130 637996
rect 342230 637896 342354 637996
rect 342454 637896 342578 637996
rect 342678 637896 342802 637996
rect 342902 637896 343026 637996
rect 343126 637896 525800 637996
rect 341994 637772 525800 637896
rect 341994 637672 342130 637772
rect 342230 637672 342354 637772
rect 342454 637672 342578 637772
rect 342678 637672 342802 637772
rect 342902 637672 343026 637772
rect 343126 637672 525800 637772
rect 341994 637561 525800 637672
rect 341994 637548 510602 637561
rect 341994 637448 342130 637548
rect 342230 637448 342354 637548
rect 342454 637448 342578 637548
rect 342678 637448 342802 637548
rect 342902 637448 343026 637548
rect 343126 637448 510602 637548
rect 341994 637324 510602 637448
rect 341994 637224 342130 637324
rect 342230 637224 342354 637324
rect 342454 637224 342578 637324
rect 342678 637224 342802 637324
rect 342902 637224 343026 637324
rect 343126 637224 510602 637324
rect 341994 637100 510602 637224
rect 341994 637000 342130 637100
rect 342230 637000 342354 637100
rect 342454 637000 342578 637100
rect 342678 637000 342802 637100
rect 342902 637000 343026 637100
rect 343126 637000 510602 637100
rect 341994 636876 510602 637000
rect 341994 636776 342130 636876
rect 342230 636776 342354 636876
rect 342454 636776 342578 636876
rect 342678 636776 342802 636876
rect 342902 636776 343026 636876
rect 343126 636776 510602 636876
rect 341994 636652 510602 636776
rect 341994 636552 342130 636652
rect 342230 636552 342354 636652
rect 342454 636552 342578 636652
rect 342678 636552 342802 636652
rect 342902 636552 343026 636652
rect 343126 636552 510602 636652
rect 341994 636428 510602 636552
rect 341994 636328 342130 636428
rect 342230 636328 342354 636428
rect 342454 636328 342578 636428
rect 342678 636328 342802 636428
rect 342902 636328 343026 636428
rect 343126 636328 510602 636428
rect 341994 636204 510602 636328
rect 341994 636104 342130 636204
rect 342230 636104 342354 636204
rect 342454 636104 342578 636204
rect 342678 636104 342802 636204
rect 342902 636104 343026 636204
rect 343126 636104 510602 636204
rect 341994 635980 510602 636104
rect 341994 635880 342130 635980
rect 342230 635880 342354 635980
rect 342454 635880 342578 635980
rect 342678 635880 342802 635980
rect 342902 635880 343026 635980
rect 343126 635880 510602 635980
rect 341994 635756 510602 635880
rect 341994 635656 342130 635756
rect 342230 635656 342354 635756
rect 342454 635656 342578 635756
rect 342678 635656 342802 635756
rect 342902 635656 343026 635756
rect 343126 635656 510602 635756
rect 341994 635532 510602 635656
rect 341994 635432 342130 635532
rect 342230 635432 342354 635532
rect 342454 635432 342578 635532
rect 342678 635432 342802 635532
rect 342902 635432 343026 635532
rect 343126 635432 510602 635532
rect 341994 635308 510602 635432
rect 341994 635208 342130 635308
rect 342230 635208 342354 635308
rect 342454 635208 342578 635308
rect 342678 635208 342802 635308
rect 342902 635208 343026 635308
rect 343126 635208 510602 635308
rect 341994 635084 510602 635208
rect 341994 634984 342130 635084
rect 342230 634984 342354 635084
rect 342454 634984 342578 635084
rect 342678 634984 342802 635084
rect 342902 634984 343026 635084
rect 343126 634984 510602 635084
rect 341994 634860 510602 634984
rect 341994 634760 342130 634860
rect 342230 634760 342354 634860
rect 342454 634760 342578 634860
rect 342678 634760 342802 634860
rect 342902 634760 343026 634860
rect 343126 634760 510602 634860
rect 341994 634636 510602 634760
rect 341994 634536 342130 634636
rect 342230 634536 342354 634636
rect 342454 634536 342578 634636
rect 342678 634536 342802 634636
rect 342902 634536 343026 634636
rect 343126 634536 510602 634636
rect 341994 634412 510602 634536
rect 341994 634312 342130 634412
rect 342230 634312 342354 634412
rect 342454 634312 342578 634412
rect 342678 634312 342802 634412
rect 342902 634312 343026 634412
rect 343126 634312 510602 634412
rect 341994 634188 510602 634312
rect 341994 634088 342130 634188
rect 342230 634088 342354 634188
rect 342454 634088 342578 634188
rect 342678 634088 342802 634188
rect 342902 634088 343026 634188
rect 343126 634088 510602 634188
rect 341994 633964 510602 634088
rect 341994 633864 342130 633964
rect 342230 633864 342354 633964
rect 342454 633864 342578 633964
rect 342678 633864 342802 633964
rect 342902 633864 343026 633964
rect 343126 633864 510602 633964
rect 341994 633740 510602 633864
rect 341994 633640 342130 633740
rect 342230 633640 342354 633740
rect 342454 633640 342578 633740
rect 342678 633640 342802 633740
rect 342902 633640 343026 633740
rect 343126 633640 510602 633740
rect 341994 633516 510602 633640
rect 341994 633416 342130 633516
rect 342230 633416 342354 633516
rect 342454 633416 342578 633516
rect 342678 633416 342802 633516
rect 342902 633416 343026 633516
rect 343126 633416 510602 633516
rect 341994 633292 510602 633416
rect 341994 633192 342130 633292
rect 342230 633192 342354 633292
rect 342454 633192 342578 633292
rect 342678 633192 342802 633292
rect 342902 633192 343026 633292
rect 343126 633192 510602 633292
rect 341994 633068 510602 633192
rect 341994 632968 342130 633068
rect 342230 632968 342354 633068
rect 342454 632968 342578 633068
rect 342678 632968 342802 633068
rect 342902 632968 343026 633068
rect 343126 632968 510602 633068
rect 341994 632844 510602 632968
rect 341994 632744 342130 632844
rect 342230 632744 342354 632844
rect 342454 632744 342578 632844
rect 342678 632744 342802 632844
rect 342902 632744 343026 632844
rect 343126 632744 510602 632844
rect 341994 632620 510602 632744
rect 341994 632520 342130 632620
rect 342230 632520 342354 632620
rect 342454 632520 342578 632620
rect 342678 632520 342802 632620
rect 342902 632520 343026 632620
rect 343126 632520 510602 632620
rect 294704 632296 297850 632396
rect 297950 632296 298074 632396
rect 298174 632296 298298 632396
rect 298398 632296 298522 632396
rect 298622 632296 298746 632396
rect 298846 632296 298880 632396
rect 294704 632172 298880 632296
rect 294704 632072 297850 632172
rect 297950 632072 298074 632172
rect 298174 632072 298298 632172
rect 298398 632072 298522 632172
rect 298622 632072 298746 632172
rect 298846 632072 298880 632172
rect 341994 632396 510602 632520
rect 341994 632296 342130 632396
rect 342230 632296 342354 632396
rect 342454 632296 342578 632396
rect 342678 632296 342802 632396
rect 342902 632296 343026 632396
rect 343126 632296 510602 632396
rect 341994 632172 510602 632296
rect 304915 632144 305011 632160
rect 294704 631948 298880 632072
rect 294704 631848 297850 631948
rect 297950 631848 298074 631948
rect 298174 631848 298298 631948
rect 298398 631848 298522 631948
rect 298622 631848 298746 631948
rect 298846 631848 298880 631948
rect 294704 631724 298880 631848
rect 294704 631624 297850 631724
rect 297950 631624 298074 631724
rect 298174 631624 298298 631724
rect 298398 631624 298522 631724
rect 298622 631624 298746 631724
rect 298846 631624 298880 631724
rect 294704 631500 298880 631624
rect 294704 631440 297850 631500
rect 289020 631400 297850 631440
rect 297950 631400 298074 631500
rect 298174 631400 298298 631500
rect 298398 631400 298522 631500
rect 298622 631400 298746 631500
rect 298846 631400 298880 631500
rect 289020 631340 298880 631400
rect 304416 632032 304816 632072
rect 304416 631712 304456 632032
rect 304776 631712 304816 632032
rect 304416 631332 304816 631712
rect 304915 631600 304931 632144
rect 304995 631600 305011 632144
rect 305634 632144 305730 632160
rect 304915 631584 305011 631600
rect 305136 632032 305536 632072
rect 305136 631712 305175 632032
rect 305495 631712 305536 632032
rect 304416 631012 304456 631332
rect 304776 631012 304816 631332
rect 304416 630632 304816 631012
rect 304915 631444 305011 631460
rect 304915 630900 304931 631444
rect 304995 630900 305011 631444
rect 304915 630884 305011 630900
rect 305136 631332 305536 631712
rect 305634 631600 305650 632144
rect 305714 631600 305730 632144
rect 306353 632144 306449 632160
rect 305634 631584 305730 631600
rect 305856 632032 306256 632072
rect 305856 631712 305894 632032
rect 306214 631712 306256 632032
rect 305136 631012 305175 631332
rect 305495 631012 305536 631332
rect 304416 630312 304456 630632
rect 304776 630312 304816 630632
rect 304416 629932 304816 630312
rect 304915 630744 305011 630760
rect 304915 630200 304931 630744
rect 304995 630200 305011 630744
rect 304915 630184 305011 630200
rect 305136 630632 305536 631012
rect 305634 631444 305730 631460
rect 305634 630900 305650 631444
rect 305714 630900 305730 631444
rect 305634 630884 305730 630900
rect 305856 631332 306256 631712
rect 306353 631600 306369 632144
rect 306433 631600 306449 632144
rect 307072 632144 307168 632160
rect 306353 631584 306449 631600
rect 306576 632032 306976 632072
rect 306576 631712 306613 632032
rect 306933 631712 306976 632032
rect 305856 631012 305894 631332
rect 306214 631012 306256 631332
rect 305136 630312 305175 630632
rect 305495 630312 305536 630632
rect 304416 629612 304456 629932
rect 304776 629612 304816 629932
rect 304416 629232 304816 629612
rect 304915 630044 305011 630060
rect 304915 629500 304931 630044
rect 304995 629500 305011 630044
rect 304915 629484 305011 629500
rect 305136 629932 305536 630312
rect 305634 630744 305730 630760
rect 305634 630200 305650 630744
rect 305714 630200 305730 630744
rect 305634 630184 305730 630200
rect 305856 630632 306256 631012
rect 306353 631444 306449 631460
rect 306353 630900 306369 631444
rect 306433 630900 306449 631444
rect 306353 630884 306449 630900
rect 306576 631332 306976 631712
rect 307072 631600 307088 632144
rect 307152 631600 307168 632144
rect 307791 632144 307887 632160
rect 307072 631584 307168 631600
rect 307296 632032 307696 632072
rect 307296 631712 307332 632032
rect 307652 631712 307696 632032
rect 306576 631012 306613 631332
rect 306933 631012 306976 631332
rect 305856 630312 305894 630632
rect 306214 630312 306256 630632
rect 305136 629612 305175 629932
rect 305495 629612 305536 629932
rect 304416 628912 304456 629232
rect 304776 628912 304816 629232
rect 304416 628532 304816 628912
rect 304915 629344 305011 629360
rect 304915 628800 304931 629344
rect 304995 628800 305011 629344
rect 304915 628784 305011 628800
rect 305136 629232 305536 629612
rect 305634 630044 305730 630060
rect 305634 629500 305650 630044
rect 305714 629500 305730 630044
rect 305634 629484 305730 629500
rect 305856 629932 306256 630312
rect 306353 630744 306449 630760
rect 306353 630200 306369 630744
rect 306433 630200 306449 630744
rect 306353 630184 306449 630200
rect 306576 630632 306976 631012
rect 307072 631444 307168 631460
rect 307072 630900 307088 631444
rect 307152 630900 307168 631444
rect 307072 630884 307168 630900
rect 307296 631332 307696 631712
rect 307791 631600 307807 632144
rect 307871 631600 307887 632144
rect 308510 632144 308606 632160
rect 307791 631584 307887 631600
rect 308016 632032 308416 632072
rect 308016 631712 308051 632032
rect 308371 631712 308416 632032
rect 307296 631012 307332 631332
rect 307652 631012 307696 631332
rect 306576 630312 306613 630632
rect 306933 630312 306976 630632
rect 305856 629612 305894 629932
rect 306214 629612 306256 629932
rect 305136 628912 305175 629232
rect 305495 628912 305536 629232
rect 304416 628212 304456 628532
rect 304776 628212 304816 628532
rect 304416 627832 304816 628212
rect 304915 628644 305011 628660
rect 304915 628100 304931 628644
rect 304995 628100 305011 628644
rect 304915 628084 305011 628100
rect 305136 628532 305536 628912
rect 305634 629344 305730 629360
rect 305634 628800 305650 629344
rect 305714 628800 305730 629344
rect 305634 628784 305730 628800
rect 305856 629232 306256 629612
rect 306353 630044 306449 630060
rect 306353 629500 306369 630044
rect 306433 629500 306449 630044
rect 306353 629484 306449 629500
rect 306576 629932 306976 630312
rect 307072 630744 307168 630760
rect 307072 630200 307088 630744
rect 307152 630200 307168 630744
rect 307072 630184 307168 630200
rect 307296 630632 307696 631012
rect 307791 631444 307887 631460
rect 307791 630900 307807 631444
rect 307871 630900 307887 631444
rect 307791 630884 307887 630900
rect 308016 631332 308416 631712
rect 308510 631600 308526 632144
rect 308590 631600 308606 632144
rect 309229 632144 309325 632160
rect 308510 631584 308606 631600
rect 308736 632032 309136 632072
rect 308736 631712 308770 632032
rect 309090 631712 309136 632032
rect 308016 631012 308051 631332
rect 308371 631012 308416 631332
rect 307296 630312 307332 630632
rect 307652 630312 307696 630632
rect 306576 629612 306613 629932
rect 306933 629612 306976 629932
rect 305856 628912 305894 629232
rect 306214 628912 306256 629232
rect 305136 628212 305175 628532
rect 305495 628212 305536 628532
rect 304416 627512 304456 627832
rect 304776 627512 304816 627832
rect 304416 627132 304816 627512
rect 304915 627944 305011 627960
rect 304915 627400 304931 627944
rect 304995 627400 305011 627944
rect 304915 627384 305011 627400
rect 305136 627832 305536 628212
rect 305634 628644 305730 628660
rect 305634 628100 305650 628644
rect 305714 628100 305730 628644
rect 305634 628084 305730 628100
rect 305856 628532 306256 628912
rect 306353 629344 306449 629360
rect 306353 628800 306369 629344
rect 306433 628800 306449 629344
rect 306353 628784 306449 628800
rect 306576 629232 306976 629612
rect 307072 630044 307168 630060
rect 307072 629500 307088 630044
rect 307152 629500 307168 630044
rect 307072 629484 307168 629500
rect 307296 629932 307696 630312
rect 307791 630744 307887 630760
rect 307791 630200 307807 630744
rect 307871 630200 307887 630744
rect 307791 630184 307887 630200
rect 308016 630632 308416 631012
rect 308510 631444 308606 631460
rect 308510 630900 308526 631444
rect 308590 630900 308606 631444
rect 308510 630884 308606 630900
rect 308736 631332 309136 631712
rect 309229 631600 309245 632144
rect 309309 631600 309325 632144
rect 309948 632144 310044 632160
rect 309229 631584 309325 631600
rect 309456 632032 309856 632072
rect 309456 631712 309489 632032
rect 309809 631712 309856 632032
rect 308736 631012 308770 631332
rect 309090 631012 309136 631332
rect 308016 630312 308051 630632
rect 308371 630312 308416 630632
rect 307296 629612 307332 629932
rect 307652 629612 307696 629932
rect 306576 628912 306613 629232
rect 306933 628912 306976 629232
rect 305856 628212 305894 628532
rect 306214 628212 306256 628532
rect 305136 627512 305175 627832
rect 305495 627512 305536 627832
rect 304416 626812 304456 627132
rect 304776 626812 304816 627132
rect 304416 626432 304816 626812
rect 304915 627244 305011 627260
rect 304915 626700 304931 627244
rect 304995 626700 305011 627244
rect 304915 626684 305011 626700
rect 305136 627132 305536 627512
rect 305634 627944 305730 627960
rect 305634 627400 305650 627944
rect 305714 627400 305730 627944
rect 305634 627384 305730 627400
rect 305856 627832 306256 628212
rect 306353 628644 306449 628660
rect 306353 628100 306369 628644
rect 306433 628100 306449 628644
rect 306353 628084 306449 628100
rect 306576 628532 306976 628912
rect 307072 629344 307168 629360
rect 307072 628800 307088 629344
rect 307152 628800 307168 629344
rect 307072 628784 307168 628800
rect 307296 629232 307696 629612
rect 307791 630044 307887 630060
rect 307791 629500 307807 630044
rect 307871 629500 307887 630044
rect 307791 629484 307887 629500
rect 308016 629932 308416 630312
rect 308510 630744 308606 630760
rect 308510 630200 308526 630744
rect 308590 630200 308606 630744
rect 308510 630184 308606 630200
rect 308736 630632 309136 631012
rect 309229 631444 309325 631460
rect 309229 630900 309245 631444
rect 309309 630900 309325 631444
rect 309229 630884 309325 630900
rect 309456 631332 309856 631712
rect 309948 631600 309964 632144
rect 310028 631600 310044 632144
rect 310667 632144 310763 632160
rect 309948 631584 310044 631600
rect 310176 632032 310576 632072
rect 310176 631712 310208 632032
rect 310528 631712 310576 632032
rect 309456 631012 309489 631332
rect 309809 631012 309856 631332
rect 308736 630312 308770 630632
rect 309090 630312 309136 630632
rect 308016 629612 308051 629932
rect 308371 629612 308416 629932
rect 307296 628912 307332 629232
rect 307652 628912 307696 629232
rect 306576 628212 306613 628532
rect 306933 628212 306976 628532
rect 305856 627512 305894 627832
rect 306214 627512 306256 627832
rect 305136 626812 305175 627132
rect 305495 626812 305536 627132
rect 217216 626176 299008 626240
rect 217216 626112 217344 626176
rect 217408 626112 217472 626176
rect 217536 626112 217600 626176
rect 217664 626112 217728 626176
rect 217792 626112 217856 626176
rect 217920 626112 217984 626176
rect 218048 626112 218112 626176
rect 218176 626112 218240 626176
rect 218304 626112 218368 626176
rect 218432 626112 218496 626176
rect 218560 626112 218624 626176
rect 218688 626112 218752 626176
rect 218816 626112 218880 626176
rect 218944 626112 219008 626176
rect 219072 626112 219136 626176
rect 219200 626112 219264 626176
rect 219328 626112 219392 626176
rect 219456 626112 219520 626176
rect 219584 626112 219648 626176
rect 219712 626112 219776 626176
rect 219840 626112 219904 626176
rect 219968 626112 220032 626176
rect 220096 626112 220160 626176
rect 220224 626112 220288 626176
rect 220352 626112 220416 626176
rect 220480 626112 220544 626176
rect 220608 626112 220672 626176
rect 220736 626112 220800 626176
rect 220864 626112 220928 626176
rect 220992 626112 221056 626176
rect 221120 626112 221184 626176
rect 221248 626112 221312 626176
rect 221376 626112 221440 626176
rect 221504 626112 221568 626176
rect 221632 626112 221696 626176
rect 221760 626112 221824 626176
rect 221888 626112 221952 626176
rect 222016 626112 222080 626176
rect 222144 626112 227640 626176
rect 227704 626112 227768 626176
rect 227832 626112 227896 626176
rect 227960 626112 228024 626176
rect 228088 626112 228152 626176
rect 228216 626112 228280 626176
rect 228344 626112 228408 626176
rect 228472 626112 228536 626176
rect 228600 626112 228664 626176
rect 228728 626112 228792 626176
rect 228856 626112 228920 626176
rect 228984 626112 229048 626176
rect 229112 626112 229176 626176
rect 229240 626112 229304 626176
rect 229368 626112 229432 626176
rect 229496 626112 229560 626176
rect 229624 626112 229688 626176
rect 229752 626112 229816 626176
rect 229880 626112 229944 626176
rect 230008 626112 230072 626176
rect 230136 626112 230200 626176
rect 230264 626112 230328 626176
rect 230392 626112 230456 626176
rect 230520 626112 230584 626176
rect 230648 626112 230712 626176
rect 230776 626112 230840 626176
rect 230904 626112 230968 626176
rect 231032 626112 231096 626176
rect 231160 626112 231224 626176
rect 231288 626112 231352 626176
rect 231416 626112 231480 626176
rect 231544 626112 231608 626176
rect 231672 626112 231736 626176
rect 231800 626112 231864 626176
rect 231928 626112 231992 626176
rect 232056 626112 232120 626176
rect 232184 626112 232248 626176
rect 232312 626112 232376 626176
rect 232440 626112 297856 626176
rect 297920 626112 297984 626176
rect 298048 626112 298112 626176
rect 298176 626112 298240 626176
rect 298304 626112 298368 626176
rect 298432 626112 298496 626176
rect 298560 626112 298624 626176
rect 298688 626112 298752 626176
rect 298816 626112 298880 626176
rect 298944 626112 299008 626176
rect 217216 626048 299008 626112
rect 217216 625984 217344 626048
rect 217408 625984 217472 626048
rect 217536 625984 217600 626048
rect 217664 625984 217728 626048
rect 217792 625984 217856 626048
rect 217920 625984 217984 626048
rect 218048 625984 218112 626048
rect 218176 625984 218240 626048
rect 218304 625984 218368 626048
rect 218432 625984 218496 626048
rect 218560 625984 218624 626048
rect 218688 625984 218752 626048
rect 218816 625984 218880 626048
rect 218944 625984 219008 626048
rect 219072 625984 219136 626048
rect 219200 625984 219264 626048
rect 219328 625984 219392 626048
rect 219456 625984 219520 626048
rect 219584 625984 219648 626048
rect 219712 625984 219776 626048
rect 219840 625984 219904 626048
rect 219968 625984 220032 626048
rect 220096 625984 220160 626048
rect 220224 625984 220288 626048
rect 220352 625984 220416 626048
rect 220480 625984 220544 626048
rect 220608 625984 220672 626048
rect 220736 625984 220800 626048
rect 220864 625984 220928 626048
rect 220992 625984 221056 626048
rect 221120 625984 221184 626048
rect 221248 625984 221312 626048
rect 221376 625984 221440 626048
rect 221504 625984 221568 626048
rect 221632 625984 221696 626048
rect 221760 625984 221824 626048
rect 221888 625984 221952 626048
rect 222016 625984 222080 626048
rect 222144 625984 227640 626048
rect 227704 625984 227768 626048
rect 227832 625984 227896 626048
rect 227960 625984 228024 626048
rect 228088 625984 228152 626048
rect 228216 625984 228280 626048
rect 228344 625984 228408 626048
rect 228472 625984 228536 626048
rect 228600 625984 228664 626048
rect 228728 625984 228792 626048
rect 228856 625984 228920 626048
rect 228984 625984 229048 626048
rect 229112 625984 229176 626048
rect 229240 625984 229304 626048
rect 229368 625984 229432 626048
rect 229496 625984 229560 626048
rect 229624 625984 229688 626048
rect 229752 625984 229816 626048
rect 229880 625984 229944 626048
rect 230008 625984 230072 626048
rect 230136 625984 230200 626048
rect 230264 625984 230328 626048
rect 230392 625984 230456 626048
rect 230520 625984 230584 626048
rect 230648 625984 230712 626048
rect 230776 625984 230840 626048
rect 230904 625984 230968 626048
rect 231032 625984 231096 626048
rect 231160 625984 231224 626048
rect 231288 625984 231352 626048
rect 231416 625984 231480 626048
rect 231544 625984 231608 626048
rect 231672 625984 231736 626048
rect 231800 625984 231864 626048
rect 231928 625984 231992 626048
rect 232056 625984 232120 626048
rect 232184 625984 232248 626048
rect 232312 625984 232376 626048
rect 232440 625984 297856 626048
rect 297920 625984 297984 626048
rect 298048 625984 298112 626048
rect 298176 625984 298240 626048
rect 298304 625984 298368 626048
rect 298432 625984 298496 626048
rect 298560 625984 298624 626048
rect 298688 625984 298752 626048
rect 298816 625984 298880 626048
rect 298944 625984 299008 626048
rect 217216 625920 299008 625984
rect 217216 625856 217344 625920
rect 217408 625856 217472 625920
rect 217536 625856 217600 625920
rect 217664 625856 217728 625920
rect 217792 625856 217856 625920
rect 217920 625856 217984 625920
rect 218048 625856 218112 625920
rect 218176 625856 218240 625920
rect 218304 625856 218368 625920
rect 218432 625856 218496 625920
rect 218560 625856 218624 625920
rect 218688 625856 218752 625920
rect 218816 625856 218880 625920
rect 218944 625856 219008 625920
rect 219072 625856 219136 625920
rect 219200 625856 219264 625920
rect 219328 625856 219392 625920
rect 219456 625856 219520 625920
rect 219584 625856 219648 625920
rect 219712 625856 219776 625920
rect 219840 625856 219904 625920
rect 219968 625856 220032 625920
rect 220096 625856 220160 625920
rect 220224 625856 220288 625920
rect 220352 625856 220416 625920
rect 220480 625856 220544 625920
rect 220608 625856 220672 625920
rect 220736 625856 220800 625920
rect 220864 625856 220928 625920
rect 220992 625856 221056 625920
rect 221120 625856 221184 625920
rect 221248 625856 221312 625920
rect 221376 625856 221440 625920
rect 221504 625856 221568 625920
rect 221632 625856 221696 625920
rect 221760 625856 221824 625920
rect 221888 625856 221952 625920
rect 222016 625856 222080 625920
rect 222144 625856 227640 625920
rect 227704 625856 227768 625920
rect 227832 625856 227896 625920
rect 227960 625856 228024 625920
rect 228088 625856 228152 625920
rect 228216 625856 228280 625920
rect 228344 625856 228408 625920
rect 228472 625856 228536 625920
rect 228600 625856 228664 625920
rect 228728 625856 228792 625920
rect 228856 625856 228920 625920
rect 228984 625856 229048 625920
rect 229112 625856 229176 625920
rect 229240 625856 229304 625920
rect 229368 625856 229432 625920
rect 229496 625856 229560 625920
rect 229624 625856 229688 625920
rect 229752 625856 229816 625920
rect 229880 625856 229944 625920
rect 230008 625856 230072 625920
rect 230136 625856 230200 625920
rect 230264 625856 230328 625920
rect 230392 625856 230456 625920
rect 230520 625856 230584 625920
rect 230648 625856 230712 625920
rect 230776 625856 230840 625920
rect 230904 625856 230968 625920
rect 231032 625856 231096 625920
rect 231160 625856 231224 625920
rect 231288 625856 231352 625920
rect 231416 625856 231480 625920
rect 231544 625856 231608 625920
rect 231672 625856 231736 625920
rect 231800 625856 231864 625920
rect 231928 625856 231992 625920
rect 232056 625856 232120 625920
rect 232184 625856 232248 625920
rect 232312 625856 232376 625920
rect 232440 625856 297856 625920
rect 297920 625856 297984 625920
rect 298048 625856 298112 625920
rect 298176 625856 298240 625920
rect 298304 625856 298368 625920
rect 298432 625856 298496 625920
rect 298560 625856 298624 625920
rect 298688 625856 298752 625920
rect 298816 625856 298880 625920
rect 298944 625856 299008 625920
rect 217216 625792 299008 625856
rect 217216 625728 217344 625792
rect 217408 625728 217472 625792
rect 217536 625728 217600 625792
rect 217664 625728 217728 625792
rect 217792 625728 217856 625792
rect 217920 625728 217984 625792
rect 218048 625728 218112 625792
rect 218176 625728 218240 625792
rect 218304 625728 218368 625792
rect 218432 625728 218496 625792
rect 218560 625728 218624 625792
rect 218688 625728 218752 625792
rect 218816 625728 218880 625792
rect 218944 625728 219008 625792
rect 219072 625728 219136 625792
rect 219200 625728 219264 625792
rect 219328 625728 219392 625792
rect 219456 625728 219520 625792
rect 219584 625728 219648 625792
rect 219712 625728 219776 625792
rect 219840 625728 219904 625792
rect 219968 625728 220032 625792
rect 220096 625728 220160 625792
rect 220224 625728 220288 625792
rect 220352 625728 220416 625792
rect 220480 625728 220544 625792
rect 220608 625728 220672 625792
rect 220736 625728 220800 625792
rect 220864 625728 220928 625792
rect 220992 625728 221056 625792
rect 221120 625728 221184 625792
rect 221248 625728 221312 625792
rect 221376 625728 221440 625792
rect 221504 625728 221568 625792
rect 221632 625728 221696 625792
rect 221760 625728 221824 625792
rect 221888 625728 221952 625792
rect 222016 625728 222080 625792
rect 222144 625728 227640 625792
rect 227704 625728 227768 625792
rect 227832 625728 227896 625792
rect 227960 625728 228024 625792
rect 228088 625728 228152 625792
rect 228216 625728 228280 625792
rect 228344 625728 228408 625792
rect 228472 625728 228536 625792
rect 228600 625728 228664 625792
rect 228728 625728 228792 625792
rect 228856 625728 228920 625792
rect 228984 625728 229048 625792
rect 229112 625728 229176 625792
rect 229240 625728 229304 625792
rect 229368 625728 229432 625792
rect 229496 625728 229560 625792
rect 229624 625728 229688 625792
rect 229752 625728 229816 625792
rect 229880 625728 229944 625792
rect 230008 625728 230072 625792
rect 230136 625728 230200 625792
rect 230264 625728 230328 625792
rect 230392 625728 230456 625792
rect 230520 625728 230584 625792
rect 230648 625728 230712 625792
rect 230776 625728 230840 625792
rect 230904 625728 230968 625792
rect 231032 625728 231096 625792
rect 231160 625728 231224 625792
rect 231288 625728 231352 625792
rect 231416 625728 231480 625792
rect 231544 625728 231608 625792
rect 231672 625728 231736 625792
rect 231800 625728 231864 625792
rect 231928 625728 231992 625792
rect 232056 625728 232120 625792
rect 232184 625728 232248 625792
rect 232312 625728 232376 625792
rect 232440 625728 297856 625792
rect 297920 625728 297984 625792
rect 298048 625728 298112 625792
rect 298176 625728 298240 625792
rect 298304 625728 298368 625792
rect 298432 625728 298496 625792
rect 298560 625728 298624 625792
rect 298688 625728 298752 625792
rect 298816 625728 298880 625792
rect 298944 625728 299008 625792
rect 217216 625664 299008 625728
rect 304416 626112 304456 626432
rect 304776 626112 304816 626432
rect 304416 625732 304816 626112
rect 304915 626544 305011 626560
rect 304915 626000 304931 626544
rect 304995 626000 305011 626544
rect 304915 625984 305011 626000
rect 305136 626432 305536 626812
rect 305634 627244 305730 627260
rect 305634 626700 305650 627244
rect 305714 626700 305730 627244
rect 305634 626684 305730 626700
rect 305856 627132 306256 627512
rect 306353 627944 306449 627960
rect 306353 627400 306369 627944
rect 306433 627400 306449 627944
rect 306353 627384 306449 627400
rect 306576 627832 306976 628212
rect 307072 628644 307168 628660
rect 307072 628100 307088 628644
rect 307152 628100 307168 628644
rect 307072 628084 307168 628100
rect 307296 628532 307696 628912
rect 307791 629344 307887 629360
rect 307791 628800 307807 629344
rect 307871 628800 307887 629344
rect 307791 628784 307887 628800
rect 308016 629232 308416 629612
rect 308510 630044 308606 630060
rect 308510 629500 308526 630044
rect 308590 629500 308606 630044
rect 308510 629484 308606 629500
rect 308736 629932 309136 630312
rect 309229 630744 309325 630760
rect 309229 630200 309245 630744
rect 309309 630200 309325 630744
rect 309229 630184 309325 630200
rect 309456 630632 309856 631012
rect 309948 631444 310044 631460
rect 309948 630900 309964 631444
rect 310028 630900 310044 631444
rect 309948 630884 310044 630900
rect 310176 631332 310576 631712
rect 310667 631600 310683 632144
rect 310747 631600 310763 632144
rect 311386 632144 311482 632160
rect 310887 632032 311296 632072
rect 310887 631712 310927 632032
rect 311247 631712 311296 632032
rect 310887 631672 311296 631712
rect 310667 631584 310763 631600
rect 310176 631012 310208 631332
rect 310528 631012 310576 631332
rect 309456 630312 309489 630632
rect 309809 630312 309856 630632
rect 308736 629612 308770 629932
rect 309090 629612 309136 629932
rect 308016 628912 308051 629232
rect 308371 628912 308416 629232
rect 307296 628212 307332 628532
rect 307652 628212 307696 628532
rect 306576 627512 306613 627832
rect 306933 627512 306976 627832
rect 305856 626812 305894 627132
rect 306214 626812 306256 627132
rect 305136 626112 305175 626432
rect 305495 626112 305536 626432
rect 304416 625412 304456 625732
rect 304776 625412 304816 625732
rect 304416 625204 304816 625412
rect 304915 625844 305011 625860
rect 304915 625300 304931 625844
rect 304995 625300 305011 625844
rect 304915 625284 305011 625300
rect 305136 625732 305536 626112
rect 305634 626544 305730 626560
rect 305634 626000 305650 626544
rect 305714 626000 305730 626544
rect 305634 625984 305730 626000
rect 305856 626432 306256 626812
rect 306353 627244 306449 627260
rect 306353 626700 306369 627244
rect 306433 626700 306449 627244
rect 306353 626684 306449 626700
rect 306576 627132 306976 627512
rect 307072 627944 307168 627960
rect 307072 627400 307088 627944
rect 307152 627400 307168 627944
rect 307072 627384 307168 627400
rect 307296 627832 307696 628212
rect 307791 628644 307887 628660
rect 307791 628100 307807 628644
rect 307871 628100 307887 628644
rect 307791 628084 307887 628100
rect 308016 628532 308416 628912
rect 308510 629344 308606 629360
rect 308510 628800 308526 629344
rect 308590 628800 308606 629344
rect 308510 628784 308606 628800
rect 308736 629232 309136 629612
rect 309229 630044 309325 630060
rect 309229 629500 309245 630044
rect 309309 629500 309325 630044
rect 309229 629484 309325 629500
rect 309456 629932 309856 630312
rect 309948 630744 310044 630760
rect 309948 630200 309964 630744
rect 310028 630200 310044 630744
rect 309948 630184 310044 630200
rect 310176 630632 310576 631012
rect 310667 631444 310763 631460
rect 310667 630900 310683 631444
rect 310747 630900 310763 631444
rect 310667 630884 310763 630900
rect 310896 631332 311296 631672
rect 311386 631600 311402 632144
rect 311466 631600 311482 632144
rect 311386 631584 311482 631600
rect 341994 632072 342130 632172
rect 342230 632072 342354 632172
rect 342454 632072 342578 632172
rect 342678 632072 342802 632172
rect 342902 632072 343026 632172
rect 343126 632072 510602 632172
rect 341994 631948 510602 632072
rect 341994 631848 342130 631948
rect 342230 631848 342354 631948
rect 342454 631848 342578 631948
rect 342678 631848 342802 631948
rect 342902 631848 343026 631948
rect 343126 631848 510602 631948
rect 341994 631817 510602 631848
rect 515386 631817 520602 637561
rect 525386 631817 525800 637561
rect 341994 631724 525800 631817
rect 341994 631624 342130 631724
rect 342230 631624 342354 631724
rect 342454 631624 342578 631724
rect 342678 631624 342802 631724
rect 342902 631624 343026 631724
rect 343126 631624 525800 631724
rect 341994 631500 525800 631624
rect 310896 631012 310927 631332
rect 311247 631012 311296 631332
rect 310176 630312 310208 630632
rect 310528 630312 310576 630632
rect 309456 629612 309489 629932
rect 309809 629612 309856 629932
rect 308736 628912 308770 629232
rect 309090 628912 309136 629232
rect 308016 628212 308051 628532
rect 308371 628212 308416 628532
rect 307296 627512 307332 627832
rect 307652 627512 307696 627832
rect 306576 626812 306613 627132
rect 306933 626812 306976 627132
rect 305856 626112 305894 626432
rect 306214 626112 306256 626432
rect 305136 625412 305175 625732
rect 305495 625412 305536 625732
rect 305136 625204 305536 625412
rect 305634 625844 305730 625860
rect 305634 625300 305650 625844
rect 305714 625300 305730 625844
rect 305634 625284 305730 625300
rect 305856 625732 306256 626112
rect 306353 626544 306449 626560
rect 306353 626000 306369 626544
rect 306433 626000 306449 626544
rect 306353 625984 306449 626000
rect 306576 626432 306976 626812
rect 307072 627244 307168 627260
rect 307072 626700 307088 627244
rect 307152 626700 307168 627244
rect 307072 626684 307168 626700
rect 307296 627132 307696 627512
rect 307791 627944 307887 627960
rect 307791 627400 307807 627944
rect 307871 627400 307887 627944
rect 307791 627384 307887 627400
rect 308016 627832 308416 628212
rect 308510 628644 308606 628660
rect 308510 628100 308526 628644
rect 308590 628100 308606 628644
rect 308510 628084 308606 628100
rect 308736 628532 309136 628912
rect 309229 629344 309325 629360
rect 309229 628800 309245 629344
rect 309309 628800 309325 629344
rect 309229 628784 309325 628800
rect 309456 629232 309856 629612
rect 309948 630044 310044 630060
rect 309948 629500 309964 630044
rect 310028 629500 310044 630044
rect 309948 629484 310044 629500
rect 310176 629932 310576 630312
rect 310667 630744 310763 630760
rect 310667 630200 310683 630744
rect 310747 630200 310763 630744
rect 310667 630184 310763 630200
rect 310896 630632 311296 631012
rect 311386 631444 311482 631460
rect 311386 630900 311402 631444
rect 311466 630900 311482 631444
rect 341994 631400 342130 631500
rect 342230 631400 342354 631500
rect 342454 631400 342578 631500
rect 342678 631400 342802 631500
rect 342902 631400 343026 631500
rect 343126 631400 525800 631500
rect 341994 631344 525800 631400
rect 560425 634576 566979 639792
rect 311386 630884 311482 630900
rect 310896 630312 310927 630632
rect 311247 630312 311296 630632
rect 310176 629612 310208 629932
rect 310528 629612 310576 629932
rect 309456 628912 309489 629232
rect 309809 628912 309856 629232
rect 308736 628212 308770 628532
rect 309090 628212 309136 628532
rect 308016 627512 308051 627832
rect 308371 627512 308416 627832
rect 307296 626812 307332 627132
rect 307652 626812 307696 627132
rect 306576 626112 306613 626432
rect 306933 626112 306976 626432
rect 305856 625412 305894 625732
rect 306214 625412 306256 625732
rect 305856 625204 306256 625412
rect 306353 625844 306449 625860
rect 306353 625300 306369 625844
rect 306433 625300 306449 625844
rect 306353 625284 306449 625300
rect 306576 625732 306976 626112
rect 307072 626544 307168 626560
rect 307072 626000 307088 626544
rect 307152 626000 307168 626544
rect 307072 625984 307168 626000
rect 307296 626432 307696 626812
rect 307791 627244 307887 627260
rect 307791 626700 307807 627244
rect 307871 626700 307887 627244
rect 307791 626684 307887 626700
rect 308016 627132 308416 627512
rect 308510 627944 308606 627960
rect 308510 627400 308526 627944
rect 308590 627400 308606 627944
rect 308510 627384 308606 627400
rect 308736 627832 309136 628212
rect 309229 628644 309325 628660
rect 309229 628100 309245 628644
rect 309309 628100 309325 628644
rect 309229 628084 309325 628100
rect 309456 628532 309856 628912
rect 309948 629344 310044 629360
rect 309948 628800 309964 629344
rect 310028 628800 310044 629344
rect 309948 628784 310044 628800
rect 310176 629232 310576 629612
rect 310667 630044 310763 630060
rect 310667 629500 310683 630044
rect 310747 629500 310763 630044
rect 310667 629484 310763 629500
rect 310896 629932 311296 630312
rect 311386 630744 311482 630760
rect 311386 630200 311402 630744
rect 311466 630200 311482 630744
rect 311386 630184 311482 630200
rect 310896 629612 310927 629932
rect 311247 629612 311296 629932
rect 310176 628912 310208 629232
rect 310528 628912 310576 629232
rect 309456 628212 309489 628532
rect 309809 628212 309856 628532
rect 308736 627512 308770 627832
rect 309090 627512 309136 627832
rect 308016 626812 308051 627132
rect 308371 626812 308416 627132
rect 307296 626112 307332 626432
rect 307652 626112 307696 626432
rect 306576 625412 306613 625732
rect 306933 625412 306976 625732
rect 306576 625204 306976 625412
rect 307072 625844 307168 625860
rect 307072 625300 307088 625844
rect 307152 625300 307168 625844
rect 307072 625284 307168 625300
rect 307296 625732 307696 626112
rect 307791 626544 307887 626560
rect 307791 626000 307807 626544
rect 307871 626000 307887 626544
rect 307791 625984 307887 626000
rect 308016 626432 308416 626812
rect 308510 627244 308606 627260
rect 308510 626700 308526 627244
rect 308590 626700 308606 627244
rect 308510 626684 308606 626700
rect 308736 627132 309136 627512
rect 309229 627944 309325 627960
rect 309229 627400 309245 627944
rect 309309 627400 309325 627944
rect 309229 627384 309325 627400
rect 309456 627832 309856 628212
rect 309948 628644 310044 628660
rect 309948 628100 309964 628644
rect 310028 628100 310044 628644
rect 309948 628084 310044 628100
rect 310176 628532 310576 628912
rect 310667 629344 310763 629360
rect 310667 628800 310683 629344
rect 310747 628800 310763 629344
rect 310667 628784 310763 628800
rect 310896 629232 311296 629612
rect 311386 630044 311482 630060
rect 311386 629500 311402 630044
rect 311466 629500 311482 630044
rect 311386 629484 311482 629500
rect 560425 629792 560582 634576
rect 566726 629792 566979 634576
rect 310896 628912 310927 629232
rect 311247 628912 311296 629232
rect 310176 628212 310208 628532
rect 310528 628212 310576 628532
rect 309456 627512 309489 627832
rect 309809 627512 309856 627832
rect 308736 626812 308770 627132
rect 309090 626812 309136 627132
rect 308016 626112 308051 626432
rect 308371 626112 308416 626432
rect 307296 625412 307332 625732
rect 307652 625412 307696 625732
rect 307296 625204 307696 625412
rect 307791 625844 307887 625860
rect 307791 625300 307807 625844
rect 307871 625300 307887 625844
rect 307791 625284 307887 625300
rect 308016 625732 308416 626112
rect 308510 626544 308606 626560
rect 308510 626000 308526 626544
rect 308590 626000 308606 626544
rect 308510 625984 308606 626000
rect 308736 626432 309136 626812
rect 309229 627244 309325 627260
rect 309229 626700 309245 627244
rect 309309 626700 309325 627244
rect 309229 626684 309325 626700
rect 309456 627132 309856 627512
rect 309948 627944 310044 627960
rect 309948 627400 309964 627944
rect 310028 627400 310044 627944
rect 309948 627384 310044 627400
rect 310176 627832 310576 628212
rect 310667 628644 310763 628660
rect 310667 628100 310683 628644
rect 310747 628100 310763 628644
rect 310667 628084 310763 628100
rect 310896 628532 311296 628912
rect 311386 629344 311482 629360
rect 311386 628800 311402 629344
rect 311466 628800 311482 629344
rect 311386 628784 311482 628800
rect 319399 628868 319601 628869
rect 319399 628668 319400 628868
rect 319600 628668 319601 628868
rect 319399 628667 319601 628668
rect 319833 628868 320035 628869
rect 319833 628668 319834 628868
rect 320034 628668 320035 628868
rect 319833 628667 320035 628668
rect 320267 628868 320469 628869
rect 320267 628668 320268 628868
rect 320468 628668 320469 628868
rect 320267 628667 320469 628668
rect 320701 628868 320903 628869
rect 320701 628668 320702 628868
rect 320902 628668 320903 628868
rect 320701 628667 320903 628668
rect 321135 628868 321337 628869
rect 321135 628668 321136 628868
rect 321336 628668 321337 628868
rect 321135 628667 321337 628668
rect 321569 628868 321771 628869
rect 321569 628668 321570 628868
rect 321770 628668 321771 628868
rect 321569 628667 321771 628668
rect 322003 628868 322205 628869
rect 322003 628668 322004 628868
rect 322204 628668 322205 628868
rect 322003 628667 322205 628668
rect 322437 628868 322639 628869
rect 322437 628668 322438 628868
rect 322638 628668 322639 628868
rect 322437 628667 322639 628668
rect 322871 628868 323073 628869
rect 322871 628668 322872 628868
rect 323072 628668 323073 628868
rect 322871 628667 323073 628668
rect 323305 628868 323507 628869
rect 323305 628668 323306 628868
rect 323506 628668 323507 628868
rect 323305 628667 323507 628668
rect 323739 628868 323941 628869
rect 323739 628668 323740 628868
rect 323940 628668 323941 628868
rect 323739 628667 323941 628668
rect 324139 628868 324341 628869
rect 324139 628668 324140 628868
rect 324340 628668 324341 628868
rect 324139 628667 324341 628668
rect 324539 628868 324741 628869
rect 324539 628668 324540 628868
rect 324740 628668 324741 628868
rect 324539 628667 324741 628668
rect 324939 628868 325141 628869
rect 324939 628668 324940 628868
rect 325140 628668 325141 628868
rect 324939 628667 325141 628668
rect 325339 628868 325541 628869
rect 325339 628668 325340 628868
rect 325540 628668 325541 628868
rect 325339 628667 325541 628668
rect 325739 628868 325941 628869
rect 325739 628668 325740 628868
rect 325940 628668 325941 628868
rect 325739 628667 325941 628668
rect 326139 628868 326341 628869
rect 326139 628668 326140 628868
rect 326340 628668 326341 628868
rect 326139 628667 326341 628668
rect 326539 628868 326741 628869
rect 326539 628668 326540 628868
rect 326740 628668 326741 628868
rect 326539 628667 326741 628668
rect 326939 628868 327141 628869
rect 326939 628668 326940 628868
rect 327140 628668 327141 628868
rect 326939 628667 327141 628668
rect 327339 628868 327541 628869
rect 327339 628668 327340 628868
rect 327540 628668 327541 628868
rect 327339 628667 327541 628668
rect 328939 628868 329141 628869
rect 328939 628668 328940 628868
rect 329140 628668 329141 628868
rect 328939 628667 329141 628668
rect 329339 628868 329541 628869
rect 329339 628668 329340 628868
rect 329540 628668 329541 628868
rect 329339 628667 329541 628668
rect 329739 628868 329941 628869
rect 329739 628668 329740 628868
rect 329940 628668 329941 628868
rect 329739 628667 329941 628668
rect 330139 628868 330341 628869
rect 330139 628668 330140 628868
rect 330340 628668 330341 628868
rect 330139 628667 330341 628668
rect 330539 628868 330741 628869
rect 330539 628668 330540 628868
rect 330740 628668 330741 628868
rect 330539 628667 330741 628668
rect 330939 628868 331141 628869
rect 330939 628668 330940 628868
rect 331140 628668 331141 628868
rect 330939 628667 331141 628668
rect 331339 628868 331541 628869
rect 331339 628668 331340 628868
rect 331540 628668 331541 628868
rect 331339 628667 331541 628668
rect 331739 628868 331941 628869
rect 331739 628668 331740 628868
rect 331940 628668 331941 628868
rect 331739 628667 331941 628668
rect 332139 628868 332341 628869
rect 332139 628668 332140 628868
rect 332340 628668 332341 628868
rect 332139 628667 332341 628668
rect 310896 628212 310927 628532
rect 311247 628212 311296 628532
rect 310176 627512 310208 627832
rect 310528 627512 310576 627832
rect 309456 626812 309489 627132
rect 309809 626812 309856 627132
rect 308736 626112 308770 626432
rect 309090 626112 309136 626432
rect 308016 625412 308051 625732
rect 308371 625412 308416 625732
rect 308016 625204 308416 625412
rect 308510 625844 308606 625860
rect 308510 625300 308526 625844
rect 308590 625300 308606 625844
rect 308510 625284 308606 625300
rect 308736 625732 309136 626112
rect 309229 626544 309325 626560
rect 309229 626000 309245 626544
rect 309309 626000 309325 626544
rect 309229 625984 309325 626000
rect 309456 626432 309856 626812
rect 309948 627244 310044 627260
rect 309948 626700 309964 627244
rect 310028 626700 310044 627244
rect 309948 626684 310044 626700
rect 310176 627132 310576 627512
rect 310667 627944 310763 627960
rect 310667 627400 310683 627944
rect 310747 627400 310763 627944
rect 310667 627384 310763 627400
rect 310896 627832 311296 628212
rect 311386 628644 311482 628660
rect 311386 628100 311402 628644
rect 311466 628100 311482 628644
rect 319399 628434 319601 628435
rect 319399 628234 319400 628434
rect 319600 628234 319601 628434
rect 319399 628233 319601 628234
rect 319833 628434 320035 628435
rect 319833 628234 319834 628434
rect 320034 628234 320035 628434
rect 319833 628233 320035 628234
rect 320267 628434 320469 628435
rect 320267 628234 320268 628434
rect 320468 628234 320469 628434
rect 320267 628233 320469 628234
rect 320701 628434 320903 628435
rect 320701 628234 320702 628434
rect 320902 628234 320903 628434
rect 320701 628233 320903 628234
rect 321135 628434 321337 628435
rect 321135 628234 321136 628434
rect 321336 628234 321337 628434
rect 321135 628233 321337 628234
rect 321569 628434 321771 628435
rect 321569 628234 321570 628434
rect 321770 628234 321771 628434
rect 321569 628233 321771 628234
rect 322003 628434 322205 628435
rect 322003 628234 322004 628434
rect 322204 628234 322205 628434
rect 322003 628233 322205 628234
rect 322437 628434 322639 628435
rect 322437 628234 322438 628434
rect 322638 628234 322639 628434
rect 322437 628233 322639 628234
rect 322871 628434 323073 628435
rect 322871 628234 322872 628434
rect 323072 628234 323073 628434
rect 322871 628233 323073 628234
rect 323305 628434 323507 628435
rect 323305 628234 323306 628434
rect 323506 628234 323507 628434
rect 323305 628233 323507 628234
rect 323739 628434 323941 628435
rect 323739 628234 323740 628434
rect 323940 628234 323941 628434
rect 323739 628233 323941 628234
rect 311386 628084 311482 628100
rect 319399 628000 319601 628001
rect 310896 627512 310927 627832
rect 311247 627512 311296 627832
rect 310176 626812 310208 627132
rect 310528 626812 310576 627132
rect 309456 626112 309489 626432
rect 309809 626112 309856 626432
rect 308736 625412 308770 625732
rect 309090 625412 309136 625732
rect 308736 625204 309136 625412
rect 309229 625844 309325 625860
rect 309229 625300 309245 625844
rect 309309 625300 309325 625844
rect 309229 625284 309325 625300
rect 309456 625732 309856 626112
rect 309948 626544 310044 626560
rect 309948 626000 309964 626544
rect 310028 626000 310044 626544
rect 309948 625984 310044 626000
rect 310176 626432 310576 626812
rect 310667 627244 310763 627260
rect 310667 626700 310683 627244
rect 310747 626700 310763 627244
rect 310667 626684 310763 626700
rect 310896 627132 311296 627512
rect 311386 627944 311482 627960
rect 311386 627400 311402 627944
rect 311466 627400 311482 627944
rect 319399 627800 319400 628000
rect 319600 627800 319601 628000
rect 319399 627799 319601 627800
rect 319833 628000 320035 628001
rect 319833 627800 319834 628000
rect 320034 627800 320035 628000
rect 319833 627799 320035 627800
rect 320267 628000 320469 628001
rect 320267 627800 320268 628000
rect 320468 627800 320469 628000
rect 320267 627799 320469 627800
rect 320701 628000 320903 628001
rect 320701 627800 320702 628000
rect 320902 627800 320903 628000
rect 320701 627799 320903 627800
rect 321135 628000 321337 628001
rect 321135 627800 321136 628000
rect 321336 627800 321337 628000
rect 321135 627799 321337 627800
rect 321569 628000 321771 628001
rect 321569 627800 321570 628000
rect 321770 627800 321771 628000
rect 321569 627799 321771 627800
rect 322003 628000 322205 628001
rect 322003 627800 322004 628000
rect 322204 627800 322205 628000
rect 322003 627799 322205 627800
rect 322437 628000 322639 628001
rect 322437 627800 322438 628000
rect 322638 627800 322639 628000
rect 322437 627799 322639 627800
rect 322871 628000 323073 628001
rect 322871 627800 322872 628000
rect 323072 627800 323073 628000
rect 322871 627799 323073 627800
rect 323305 628000 323507 628001
rect 323305 627800 323306 628000
rect 323506 627800 323507 628000
rect 323305 627799 323507 627800
rect 323739 628000 323941 628001
rect 323739 627800 323740 628000
rect 323940 627800 323941 628000
rect 323739 627799 323941 627800
rect 311386 627384 311482 627400
rect 312957 627286 333269 627287
rect 310896 626812 310927 627132
rect 311247 626812 311296 627132
rect 310176 626112 310208 626432
rect 310528 626112 310576 626432
rect 309456 625412 309489 625732
rect 309809 625412 309856 625732
rect 309456 625204 309856 625412
rect 309948 625844 310044 625860
rect 309948 625300 309964 625844
rect 310028 625300 310044 625844
rect 309948 625284 310044 625300
rect 310176 625732 310576 626112
rect 310667 626544 310763 626560
rect 310667 626000 310683 626544
rect 310747 626000 310763 626544
rect 310667 625984 310763 626000
rect 310896 626432 311296 626812
rect 311386 627244 311482 627260
rect 311386 626700 311402 627244
rect 311466 626700 311482 627244
rect 311386 626684 311482 626700
rect 310896 626112 310927 626432
rect 311247 626112 311296 626432
rect 310176 625412 310208 625732
rect 310528 625412 310576 625732
rect 310176 625204 310576 625412
rect 310667 625844 310763 625860
rect 310667 625300 310683 625844
rect 310747 625300 310763 625844
rect 310667 625284 310763 625300
rect 310896 625732 311296 626112
rect 311386 626544 311482 626560
rect 311386 626000 311402 626544
rect 311466 626000 311482 626544
rect 312957 626314 312958 627286
rect 333268 626314 333269 627286
rect 312957 626313 333269 626314
rect 311386 625984 311482 626000
rect 310896 625412 310927 625732
rect 311247 625412 311296 625732
rect 310896 625212 311296 625412
rect 311386 625844 311482 625860
rect 311386 625300 311402 625844
rect 311466 625300 311482 625844
rect 311386 625284 311482 625300
rect 310896 625204 311316 625212
rect 304416 625197 311316 625204
rect 289020 624596 298880 624620
rect 289020 624496 297850 624596
rect 297950 624496 298074 624596
rect 298174 624496 298298 624596
rect 298398 624496 298522 624596
rect 298622 624496 298746 624596
rect 298846 624496 298880 624596
rect 289020 624372 298880 624496
rect 289020 624272 297850 624372
rect 297950 624272 298074 624372
rect 298174 624272 298298 624372
rect 298398 624272 298522 624372
rect 298622 624272 298746 624372
rect 298846 624272 298880 624372
rect 289020 624148 298880 624272
rect 289020 624048 297850 624148
rect 297950 624048 298074 624148
rect 298174 624048 298298 624148
rect 298398 624048 298522 624148
rect 298622 624048 298746 624148
rect 298846 624048 298880 624148
rect 289020 623924 298880 624048
rect 289020 623824 297850 623924
rect 297950 623824 298074 623924
rect 298174 623824 298298 623924
rect 298398 623824 298522 623924
rect 298622 623824 298746 623924
rect 298846 623824 298880 623924
rect 289020 623784 298880 623824
rect 289020 618040 289920 623784
rect 294704 623700 298880 623784
rect 294704 623600 297850 623700
rect 297950 623600 298074 623700
rect 298174 623600 298298 623700
rect 298398 623600 298522 623700
rect 298622 623600 298746 623700
rect 298846 623600 298880 623700
rect 294704 623476 298880 623600
rect 294704 623376 297850 623476
rect 297950 623376 298074 623476
rect 298174 623376 298298 623476
rect 298398 623376 298522 623476
rect 298622 623376 298746 623476
rect 298846 623376 298880 623476
rect 294704 623252 298880 623376
rect 294704 623152 297850 623252
rect 297950 623152 298074 623252
rect 298174 623152 298298 623252
rect 298398 623152 298522 623252
rect 298622 623152 298746 623252
rect 298846 623152 298880 623252
rect 294704 623028 298880 623152
rect 294704 622928 297850 623028
rect 297950 622928 298074 623028
rect 298174 622928 298298 623028
rect 298398 622928 298522 623028
rect 298622 622928 298746 623028
rect 298846 622928 298880 623028
rect 294704 622804 298880 622928
rect 294704 622704 297850 622804
rect 297950 622704 298074 622804
rect 298174 622704 298298 622804
rect 298398 622704 298522 622804
rect 298622 622704 298746 622804
rect 298846 622704 298880 622804
rect 294704 622580 298880 622704
rect 294704 622480 297850 622580
rect 297950 622480 298074 622580
rect 298174 622480 298298 622580
rect 298398 622480 298522 622580
rect 298622 622480 298746 622580
rect 298846 622480 298880 622580
rect 294704 622356 298880 622480
rect 294704 622256 297850 622356
rect 297950 622256 298074 622356
rect 298174 622256 298298 622356
rect 298398 622256 298522 622356
rect 298622 622256 298746 622356
rect 298846 622256 298880 622356
rect 294704 622132 298880 622256
rect 294704 622032 297850 622132
rect 297950 622032 298074 622132
rect 298174 622032 298298 622132
rect 298398 622032 298522 622132
rect 298622 622032 298746 622132
rect 298846 622032 298880 622132
rect 294704 621908 298880 622032
rect 294704 621808 297850 621908
rect 297950 621808 298074 621908
rect 298174 621808 298298 621908
rect 298398 621808 298522 621908
rect 298622 621808 298746 621908
rect 298846 621808 298880 621908
rect 294704 621684 298880 621808
rect 294704 621584 297850 621684
rect 297950 621584 298074 621684
rect 298174 621584 298298 621684
rect 298398 621584 298522 621684
rect 298622 621584 298746 621684
rect 298846 621584 298880 621684
rect 294704 621460 298880 621584
rect 294704 621360 297850 621460
rect 297950 621360 298074 621460
rect 298174 621360 298298 621460
rect 298398 621360 298522 621460
rect 298622 621360 298746 621460
rect 298846 621360 298880 621460
rect 294704 621236 298880 621360
rect 294704 621136 297850 621236
rect 297950 621136 298074 621236
rect 298174 621136 298298 621236
rect 298398 621136 298522 621236
rect 298622 621136 298746 621236
rect 298846 621136 298880 621236
rect 294704 621012 298880 621136
rect 294704 620912 297850 621012
rect 297950 620912 298074 621012
rect 298174 620912 298298 621012
rect 298398 620912 298522 621012
rect 298622 620912 298746 621012
rect 298846 620912 298880 621012
rect 294704 620788 298880 620912
rect 294704 620688 297850 620788
rect 297950 620688 298074 620788
rect 298174 620688 298298 620788
rect 298398 620688 298522 620788
rect 298622 620688 298746 620788
rect 298846 620688 298880 620788
rect 294704 620564 298880 620688
rect 294704 620464 297850 620564
rect 297950 620464 298074 620564
rect 298174 620464 298298 620564
rect 298398 620464 298522 620564
rect 298622 620464 298746 620564
rect 298846 620464 298880 620564
rect 294704 620340 298880 620464
rect 294704 620240 297850 620340
rect 297950 620240 298074 620340
rect 298174 620240 298298 620340
rect 298398 620240 298522 620340
rect 298622 620240 298746 620340
rect 298846 620240 298880 620340
rect 294704 620116 298880 620240
rect 303590 620151 312722 625197
rect 294704 620016 297850 620116
rect 297950 620016 298074 620116
rect 298174 620016 298298 620116
rect 298398 620016 298522 620116
rect 298622 620016 298746 620116
rect 298846 620016 298880 620116
rect 294704 619892 298880 620016
rect 294704 619792 297850 619892
rect 297950 619792 298074 619892
rect 298174 619792 298298 619892
rect 298398 619792 298522 619892
rect 298622 619792 298746 619892
rect 298846 619792 298880 619892
rect 303588 620149 312722 620151
rect 303588 619869 303590 620149
rect 304218 619869 312081 620149
rect 312709 619869 312722 620149
rect 303588 619867 312722 619869
rect 303590 619866 312722 619867
rect 342000 624596 525804 624606
rect 342000 624496 342130 624596
rect 342230 624496 342354 624596
rect 342454 624496 342578 624596
rect 342678 624496 342802 624596
rect 342902 624496 343026 624596
rect 343126 624496 525804 624596
rect 342000 624372 525804 624496
rect 342000 624272 342130 624372
rect 342230 624272 342354 624372
rect 342454 624272 342578 624372
rect 342678 624272 342802 624372
rect 342902 624272 343026 624372
rect 343126 624272 525804 624372
rect 342000 624161 525804 624272
rect 342000 624148 510602 624161
rect 342000 624048 342130 624148
rect 342230 624048 342354 624148
rect 342454 624048 342578 624148
rect 342678 624048 342802 624148
rect 342902 624048 343026 624148
rect 343126 624048 510602 624148
rect 342000 623924 510602 624048
rect 342000 623824 342130 623924
rect 342230 623824 342354 623924
rect 342454 623824 342578 623924
rect 342678 623824 342802 623924
rect 342902 623824 343026 623924
rect 343126 623824 510602 623924
rect 342000 623700 510602 623824
rect 342000 623600 342130 623700
rect 342230 623600 342354 623700
rect 342454 623600 342578 623700
rect 342678 623600 342802 623700
rect 342902 623600 343026 623700
rect 343126 623600 510602 623700
rect 342000 623476 510602 623600
rect 342000 623376 342130 623476
rect 342230 623376 342354 623476
rect 342454 623376 342578 623476
rect 342678 623376 342802 623476
rect 342902 623376 343026 623476
rect 343126 623376 510602 623476
rect 342000 623252 510602 623376
rect 342000 623152 342130 623252
rect 342230 623152 342354 623252
rect 342454 623152 342578 623252
rect 342678 623152 342802 623252
rect 342902 623152 343026 623252
rect 343126 623152 510602 623252
rect 342000 623028 510602 623152
rect 342000 622928 342130 623028
rect 342230 622928 342354 623028
rect 342454 622928 342578 623028
rect 342678 622928 342802 623028
rect 342902 622928 343026 623028
rect 343126 622928 510602 623028
rect 342000 622804 510602 622928
rect 342000 622704 342130 622804
rect 342230 622704 342354 622804
rect 342454 622704 342578 622804
rect 342678 622704 342802 622804
rect 342902 622704 343026 622804
rect 343126 622704 510602 622804
rect 342000 622580 510602 622704
rect 342000 622480 342130 622580
rect 342230 622480 342354 622580
rect 342454 622480 342578 622580
rect 342678 622480 342802 622580
rect 342902 622480 343026 622580
rect 343126 622480 510602 622580
rect 342000 622356 510602 622480
rect 342000 622256 342130 622356
rect 342230 622256 342354 622356
rect 342454 622256 342578 622356
rect 342678 622256 342802 622356
rect 342902 622256 343026 622356
rect 343126 622256 510602 622356
rect 342000 622132 510602 622256
rect 342000 622032 342130 622132
rect 342230 622032 342354 622132
rect 342454 622032 342578 622132
rect 342678 622032 342802 622132
rect 342902 622032 343026 622132
rect 343126 622032 510602 622132
rect 342000 621908 510602 622032
rect 342000 621808 342130 621908
rect 342230 621808 342354 621908
rect 342454 621808 342578 621908
rect 342678 621808 342802 621908
rect 342902 621808 343026 621908
rect 343126 621808 510602 621908
rect 342000 621684 510602 621808
rect 342000 621584 342130 621684
rect 342230 621584 342354 621684
rect 342454 621584 342578 621684
rect 342678 621584 342802 621684
rect 342902 621584 343026 621684
rect 343126 621584 510602 621684
rect 342000 621460 510602 621584
rect 342000 621360 342130 621460
rect 342230 621360 342354 621460
rect 342454 621360 342578 621460
rect 342678 621360 342802 621460
rect 342902 621360 343026 621460
rect 343126 621360 510602 621460
rect 342000 621236 510602 621360
rect 342000 621136 342130 621236
rect 342230 621136 342354 621236
rect 342454 621136 342578 621236
rect 342678 621136 342802 621236
rect 342902 621136 343026 621236
rect 343126 621136 510602 621236
rect 342000 621012 510602 621136
rect 342000 620912 342130 621012
rect 342230 620912 342354 621012
rect 342454 620912 342578 621012
rect 342678 620912 342802 621012
rect 342902 620912 343026 621012
rect 343126 620912 510602 621012
rect 342000 620788 510602 620912
rect 342000 620688 342130 620788
rect 342230 620688 342354 620788
rect 342454 620688 342578 620788
rect 342678 620688 342802 620788
rect 342902 620688 343026 620788
rect 343126 620688 510602 620788
rect 342000 620564 510602 620688
rect 342000 620464 342130 620564
rect 342230 620464 342354 620564
rect 342454 620464 342578 620564
rect 342678 620464 342802 620564
rect 342902 620464 343026 620564
rect 343126 620464 510602 620564
rect 342000 620340 510602 620464
rect 342000 620240 342130 620340
rect 342230 620240 342354 620340
rect 342454 620240 342578 620340
rect 342678 620240 342802 620340
rect 342902 620240 343026 620340
rect 343126 620240 510602 620340
rect 342000 620116 510602 620240
rect 342000 620016 342130 620116
rect 342230 620016 342354 620116
rect 342454 620016 342578 620116
rect 342678 620016 342802 620116
rect 342902 620016 343026 620116
rect 343126 620016 510602 620116
rect 342000 619892 510602 620016
rect 294704 619668 298880 619792
rect 294704 619568 297850 619668
rect 297950 619568 298074 619668
rect 298174 619568 298298 619668
rect 298398 619568 298522 619668
rect 298622 619568 298746 619668
rect 298846 619568 298880 619668
rect 294704 619444 298880 619568
rect 294704 619344 297850 619444
rect 297950 619344 298074 619444
rect 298174 619344 298298 619444
rect 298398 619344 298522 619444
rect 298622 619344 298746 619444
rect 298846 619344 298880 619444
rect 294704 619220 298880 619344
rect 294704 619120 297850 619220
rect 297950 619120 298074 619220
rect 298174 619120 298298 619220
rect 298398 619120 298522 619220
rect 298622 619120 298746 619220
rect 298846 619120 298880 619220
rect 294704 618996 298880 619120
rect 294704 618896 297850 618996
rect 297950 618896 298074 618996
rect 298174 618896 298298 618996
rect 298398 618896 298522 618996
rect 298622 618896 298746 618996
rect 298846 618896 298880 618996
rect 294704 618772 298880 618896
rect 294704 618672 297850 618772
rect 297950 618672 298074 618772
rect 298174 618672 298298 618772
rect 298398 618672 298522 618772
rect 298622 618672 298746 618772
rect 298846 618672 298880 618772
rect 294704 618548 298880 618672
rect 294704 618448 297850 618548
rect 297950 618448 298074 618548
rect 298174 618448 298298 618548
rect 298398 618448 298522 618548
rect 298622 618448 298746 618548
rect 298846 618448 298880 618548
rect 294704 618324 298880 618448
rect 294704 618224 297850 618324
rect 297950 618224 298074 618324
rect 298174 618224 298298 618324
rect 298398 618224 298522 618324
rect 298622 618224 298746 618324
rect 298846 618224 298880 618324
rect 294704 618100 298880 618224
rect 294704 618040 297850 618100
rect 289020 618000 297850 618040
rect 297950 618000 298074 618100
rect 298174 618000 298298 618100
rect 298398 618000 298522 618100
rect 298622 618000 298746 618100
rect 298846 618000 298880 618100
rect 289020 617940 298880 618000
rect 342000 619792 342130 619892
rect 342230 619792 342354 619892
rect 342454 619792 342578 619892
rect 342678 619792 342802 619892
rect 342902 619792 343026 619892
rect 343126 619792 510602 619892
rect 342000 619668 510602 619792
rect 342000 619568 342130 619668
rect 342230 619568 342354 619668
rect 342454 619568 342578 619668
rect 342678 619568 342802 619668
rect 342902 619568 343026 619668
rect 343126 619568 510602 619668
rect 342000 619444 510602 619568
rect 342000 619344 342130 619444
rect 342230 619344 342354 619444
rect 342454 619344 342578 619444
rect 342678 619344 342802 619444
rect 342902 619344 343026 619444
rect 343126 619344 510602 619444
rect 342000 619220 510602 619344
rect 342000 619120 342130 619220
rect 342230 619120 342354 619220
rect 342454 619120 342578 619220
rect 342678 619120 342802 619220
rect 342902 619120 343026 619220
rect 343126 619120 510602 619220
rect 342000 618996 510602 619120
rect 342000 618896 342130 618996
rect 342230 618896 342354 618996
rect 342454 618896 342578 618996
rect 342678 618896 342802 618996
rect 342902 618896 343026 618996
rect 343126 618896 510602 618996
rect 342000 618772 510602 618896
rect 342000 618672 342130 618772
rect 342230 618672 342354 618772
rect 342454 618672 342578 618772
rect 342678 618672 342802 618772
rect 342902 618672 343026 618772
rect 343126 618672 510602 618772
rect 342000 618548 510602 618672
rect 342000 618448 342130 618548
rect 342230 618448 342354 618548
rect 342454 618448 342578 618548
rect 342678 618448 342802 618548
rect 342902 618448 343026 618548
rect 343126 618448 510602 618548
rect 342000 618417 510602 618448
rect 515386 618417 520602 624161
rect 525386 618417 525804 624161
rect 342000 618324 525804 618417
rect 342000 618224 342130 618324
rect 342230 618224 342354 618324
rect 342454 618224 342578 618324
rect 342678 618224 342802 618324
rect 342902 618224 343026 618324
rect 343126 618224 525804 618324
rect 342000 618100 525804 618224
rect 342000 618000 342130 618100
rect 342230 618000 342354 618100
rect 342454 618000 342578 618100
rect 342678 618000 342802 618100
rect 342902 618000 343026 618100
rect 343126 618000 525804 618100
rect 342000 617944 525804 618000
rect 335560 615499 342216 615504
rect 335560 615494 342217 615499
rect 298820 615479 305476 615484
rect 309290 615479 315946 615484
rect 298820 615474 305477 615479
rect 298820 615374 298876 615474
rect 298976 615374 299100 615474
rect 299200 615374 299324 615474
rect 299424 615374 299548 615474
rect 299648 615374 299772 615474
rect 299872 615374 299996 615474
rect 300096 615374 300220 615474
rect 300320 615374 300444 615474
rect 300544 615374 300668 615474
rect 300768 615374 300892 615474
rect 300992 615374 301116 615474
rect 301216 615374 301340 615474
rect 301440 615374 301564 615474
rect 301664 615374 301788 615474
rect 301888 615374 302012 615474
rect 302112 615374 302236 615474
rect 302336 615374 302460 615474
rect 302560 615374 302684 615474
rect 302784 615374 302908 615474
rect 303008 615374 303132 615474
rect 303232 615374 303356 615474
rect 303456 615374 303580 615474
rect 303680 615374 303804 615474
rect 303904 615374 304028 615474
rect 304128 615374 304252 615474
rect 304352 615374 304476 615474
rect 304576 615374 304700 615474
rect 304800 615374 304924 615474
rect 305024 615374 305148 615474
rect 305248 615374 305372 615474
rect 305472 615374 305477 615474
rect 298820 615369 305477 615374
rect 309290 615474 315947 615479
rect 309290 615374 309346 615474
rect 309446 615374 309570 615474
rect 309670 615374 309794 615474
rect 309894 615374 310018 615474
rect 310118 615374 310242 615474
rect 310342 615374 310466 615474
rect 310566 615374 310690 615474
rect 310790 615374 310914 615474
rect 311014 615374 311138 615474
rect 311238 615374 311362 615474
rect 311462 615374 311586 615474
rect 311686 615374 311810 615474
rect 311910 615374 312034 615474
rect 312134 615374 312258 615474
rect 312358 615374 312482 615474
rect 312582 615374 312706 615474
rect 312806 615374 312930 615474
rect 313030 615374 313154 615474
rect 313254 615374 313378 615474
rect 313478 615374 313602 615474
rect 313702 615374 313826 615474
rect 313926 615374 314050 615474
rect 314150 615374 314274 615474
rect 314374 615374 314498 615474
rect 314598 615374 314722 615474
rect 314822 615374 314946 615474
rect 315046 615374 315170 615474
rect 315270 615374 315394 615474
rect 315494 615374 315618 615474
rect 315718 615374 315842 615474
rect 315942 615374 315947 615474
rect 309290 615369 315947 615374
rect 335560 615394 335616 615494
rect 335716 615394 335840 615494
rect 335940 615394 336064 615494
rect 336164 615394 336288 615494
rect 336388 615394 336512 615494
rect 336612 615394 336736 615494
rect 336836 615394 336960 615494
rect 337060 615394 337184 615494
rect 337284 615394 337408 615494
rect 337508 615394 337632 615494
rect 337732 615394 337856 615494
rect 337956 615394 338080 615494
rect 338180 615394 338304 615494
rect 338404 615394 338528 615494
rect 338628 615394 338752 615494
rect 338852 615394 338976 615494
rect 339076 615394 339200 615494
rect 339300 615394 339424 615494
rect 339524 615394 339648 615494
rect 339748 615394 339872 615494
rect 339972 615394 340096 615494
rect 340196 615394 340320 615494
rect 340420 615394 340544 615494
rect 340644 615394 340768 615494
rect 340868 615394 340992 615494
rect 341092 615394 341216 615494
rect 341316 615394 341440 615494
rect 341540 615394 341664 615494
rect 341764 615394 341888 615494
rect 341988 615394 342112 615494
rect 342212 615394 342217 615494
rect 335560 615389 342217 615394
rect 298820 615255 305476 615369
rect 309290 615255 315946 615369
rect 335560 615275 342216 615389
rect 335560 615270 342217 615275
rect 298820 615250 305477 615255
rect 298820 615150 298876 615250
rect 298976 615150 299100 615250
rect 299200 615150 299324 615250
rect 299424 615150 299548 615250
rect 299648 615150 299772 615250
rect 299872 615150 299996 615250
rect 300096 615150 300220 615250
rect 300320 615150 300444 615250
rect 300544 615150 300668 615250
rect 300768 615150 300892 615250
rect 300992 615150 301116 615250
rect 301216 615150 301340 615250
rect 301440 615150 301564 615250
rect 301664 615150 301788 615250
rect 301888 615150 302012 615250
rect 302112 615150 302236 615250
rect 302336 615150 302460 615250
rect 302560 615150 302684 615250
rect 302784 615150 302908 615250
rect 303008 615150 303132 615250
rect 303232 615150 303356 615250
rect 303456 615150 303580 615250
rect 303680 615150 303804 615250
rect 303904 615150 304028 615250
rect 304128 615150 304252 615250
rect 304352 615150 304476 615250
rect 304576 615150 304700 615250
rect 304800 615150 304924 615250
rect 305024 615150 305148 615250
rect 305248 615150 305372 615250
rect 305472 615150 305477 615250
rect 298820 615145 305477 615150
rect 309290 615250 315947 615255
rect 309290 615150 309346 615250
rect 309446 615150 309570 615250
rect 309670 615150 309794 615250
rect 309894 615150 310018 615250
rect 310118 615150 310242 615250
rect 310342 615150 310466 615250
rect 310566 615150 310690 615250
rect 310790 615150 310914 615250
rect 311014 615150 311138 615250
rect 311238 615150 311362 615250
rect 311462 615150 311586 615250
rect 311686 615150 311810 615250
rect 311910 615150 312034 615250
rect 312134 615150 312258 615250
rect 312358 615150 312482 615250
rect 312582 615150 312706 615250
rect 312806 615150 312930 615250
rect 313030 615150 313154 615250
rect 313254 615150 313378 615250
rect 313478 615150 313602 615250
rect 313702 615150 313826 615250
rect 313926 615150 314050 615250
rect 314150 615150 314274 615250
rect 314374 615150 314498 615250
rect 314598 615150 314722 615250
rect 314822 615150 314946 615250
rect 315046 615150 315170 615250
rect 315270 615150 315394 615250
rect 315494 615150 315618 615250
rect 315718 615150 315842 615250
rect 315942 615150 315947 615250
rect 309290 615145 315947 615150
rect 335560 615170 335616 615270
rect 335716 615170 335840 615270
rect 335940 615170 336064 615270
rect 336164 615170 336288 615270
rect 336388 615170 336512 615270
rect 336612 615170 336736 615270
rect 336836 615170 336960 615270
rect 337060 615170 337184 615270
rect 337284 615170 337408 615270
rect 337508 615170 337632 615270
rect 337732 615170 337856 615270
rect 337956 615170 338080 615270
rect 338180 615170 338304 615270
rect 338404 615170 338528 615270
rect 338628 615170 338752 615270
rect 338852 615170 338976 615270
rect 339076 615170 339200 615270
rect 339300 615170 339424 615270
rect 339524 615170 339648 615270
rect 339748 615170 339872 615270
rect 339972 615170 340096 615270
rect 340196 615170 340320 615270
rect 340420 615170 340544 615270
rect 340644 615170 340768 615270
rect 340868 615170 340992 615270
rect 341092 615170 341216 615270
rect 341316 615170 341440 615270
rect 341540 615170 341664 615270
rect 341764 615170 341888 615270
rect 341988 615170 342112 615270
rect 342212 615170 342217 615270
rect 335560 615165 342217 615170
rect 298820 615031 305476 615145
rect 309290 615031 315946 615145
rect 335560 615051 342216 615165
rect 335560 615046 342217 615051
rect 298820 615026 305477 615031
rect 298820 614926 298876 615026
rect 298976 614926 299100 615026
rect 299200 614926 299324 615026
rect 299424 614926 299548 615026
rect 299648 614926 299772 615026
rect 299872 614926 299996 615026
rect 300096 614926 300220 615026
rect 300320 614926 300444 615026
rect 300544 614926 300668 615026
rect 300768 614926 300892 615026
rect 300992 614926 301116 615026
rect 301216 614926 301340 615026
rect 301440 614926 301564 615026
rect 301664 614926 301788 615026
rect 301888 614926 302012 615026
rect 302112 614926 302236 615026
rect 302336 614926 302460 615026
rect 302560 614926 302684 615026
rect 302784 614926 302908 615026
rect 303008 614926 303132 615026
rect 303232 614926 303356 615026
rect 303456 614926 303580 615026
rect 303680 614926 303804 615026
rect 303904 614926 304028 615026
rect 304128 614926 304252 615026
rect 304352 614926 304476 615026
rect 304576 614926 304700 615026
rect 304800 614926 304924 615026
rect 305024 614926 305148 615026
rect 305248 614926 305372 615026
rect 305472 614926 305477 615026
rect 298820 614921 305477 614926
rect 309290 615026 315947 615031
rect 309290 614926 309346 615026
rect 309446 614926 309570 615026
rect 309670 614926 309794 615026
rect 309894 614926 310018 615026
rect 310118 614926 310242 615026
rect 310342 614926 310466 615026
rect 310566 614926 310690 615026
rect 310790 614926 310914 615026
rect 311014 614926 311138 615026
rect 311238 614926 311362 615026
rect 311462 614926 311586 615026
rect 311686 614926 311810 615026
rect 311910 614926 312034 615026
rect 312134 614926 312258 615026
rect 312358 614926 312482 615026
rect 312582 614926 312706 615026
rect 312806 614926 312930 615026
rect 313030 614926 313154 615026
rect 313254 614926 313378 615026
rect 313478 614926 313602 615026
rect 313702 614926 313826 615026
rect 313926 614926 314050 615026
rect 314150 614926 314274 615026
rect 314374 614926 314498 615026
rect 314598 614926 314722 615026
rect 314822 614926 314946 615026
rect 315046 614926 315170 615026
rect 315270 614926 315394 615026
rect 315494 614926 315618 615026
rect 315718 614926 315842 615026
rect 315942 614926 315947 615026
rect 309290 614921 315947 614926
rect 335560 614946 335616 615046
rect 335716 614946 335840 615046
rect 335940 614946 336064 615046
rect 336164 614946 336288 615046
rect 336388 614946 336512 615046
rect 336612 614946 336736 615046
rect 336836 614946 336960 615046
rect 337060 614946 337184 615046
rect 337284 614946 337408 615046
rect 337508 614946 337632 615046
rect 337732 614946 337856 615046
rect 337956 614946 338080 615046
rect 338180 614946 338304 615046
rect 338404 614946 338528 615046
rect 338628 614946 338752 615046
rect 338852 614946 338976 615046
rect 339076 614946 339200 615046
rect 339300 614946 339424 615046
rect 339524 614946 339648 615046
rect 339748 614946 339872 615046
rect 339972 614946 340096 615046
rect 340196 614946 340320 615046
rect 340420 614946 340544 615046
rect 340644 614946 340768 615046
rect 340868 614946 340992 615046
rect 341092 614946 341216 615046
rect 341316 614946 341440 615046
rect 341540 614946 341664 615046
rect 341764 614946 341888 615046
rect 341988 614946 342112 615046
rect 342212 614946 342217 615046
rect 335560 614941 342217 614946
rect 298820 614807 305476 614921
rect 309290 614807 315946 614921
rect 335560 614827 342216 614941
rect 335560 614822 342217 614827
rect 298820 614802 305477 614807
rect 298820 614702 298876 614802
rect 298976 614702 299100 614802
rect 299200 614702 299324 614802
rect 299424 614702 299548 614802
rect 299648 614702 299772 614802
rect 299872 614702 299996 614802
rect 300096 614702 300220 614802
rect 300320 614702 300444 614802
rect 300544 614702 300668 614802
rect 300768 614702 300892 614802
rect 300992 614702 301116 614802
rect 301216 614702 301340 614802
rect 301440 614702 301564 614802
rect 301664 614702 301788 614802
rect 301888 614702 302012 614802
rect 302112 614702 302236 614802
rect 302336 614702 302460 614802
rect 302560 614702 302684 614802
rect 302784 614702 302908 614802
rect 303008 614702 303132 614802
rect 303232 614702 303356 614802
rect 303456 614702 303580 614802
rect 303680 614702 303804 614802
rect 303904 614702 304028 614802
rect 304128 614702 304252 614802
rect 304352 614702 304476 614802
rect 304576 614702 304700 614802
rect 304800 614702 304924 614802
rect 305024 614702 305148 614802
rect 305248 614702 305372 614802
rect 305472 614702 305477 614802
rect 298820 614697 305477 614702
rect 309290 614802 315947 614807
rect 309290 614702 309346 614802
rect 309446 614702 309570 614802
rect 309670 614702 309794 614802
rect 309894 614702 310018 614802
rect 310118 614702 310242 614802
rect 310342 614702 310466 614802
rect 310566 614702 310690 614802
rect 310790 614702 310914 614802
rect 311014 614702 311138 614802
rect 311238 614702 311362 614802
rect 311462 614702 311586 614802
rect 311686 614702 311810 614802
rect 311910 614702 312034 614802
rect 312134 614702 312258 614802
rect 312358 614702 312482 614802
rect 312582 614702 312706 614802
rect 312806 614702 312930 614802
rect 313030 614702 313154 614802
rect 313254 614702 313378 614802
rect 313478 614702 313602 614802
rect 313702 614702 313826 614802
rect 313926 614702 314050 614802
rect 314150 614702 314274 614802
rect 314374 614702 314498 614802
rect 314598 614702 314722 614802
rect 314822 614702 314946 614802
rect 315046 614702 315170 614802
rect 315270 614702 315394 614802
rect 315494 614702 315618 614802
rect 315718 614702 315842 614802
rect 315942 614702 315947 614802
rect 309290 614697 315947 614702
rect 335560 614722 335616 614822
rect 335716 614722 335840 614822
rect 335940 614722 336064 614822
rect 336164 614722 336288 614822
rect 336388 614722 336512 614822
rect 336612 614722 336736 614822
rect 336836 614722 336960 614822
rect 337060 614722 337184 614822
rect 337284 614722 337408 614822
rect 337508 614722 337632 614822
rect 337732 614722 337856 614822
rect 337956 614722 338080 614822
rect 338180 614722 338304 614822
rect 338404 614722 338528 614822
rect 338628 614722 338752 614822
rect 338852 614722 338976 614822
rect 339076 614722 339200 614822
rect 339300 614722 339424 614822
rect 339524 614722 339648 614822
rect 339748 614722 339872 614822
rect 339972 614722 340096 614822
rect 340196 614722 340320 614822
rect 340420 614722 340544 614822
rect 340644 614722 340768 614822
rect 340868 614722 340992 614822
rect 341092 614722 341216 614822
rect 341316 614722 341440 614822
rect 341540 614722 341664 614822
rect 341764 614722 341888 614822
rect 341988 614722 342112 614822
rect 342212 614722 342217 614822
rect 335560 614717 342217 614722
rect 298820 614583 305476 614697
rect 309290 614583 315946 614697
rect 335560 614603 342216 614717
rect 335560 614598 342217 614603
rect 298820 614578 305477 614583
rect 298820 614478 298876 614578
rect 298976 614478 299100 614578
rect 299200 614478 299324 614578
rect 299424 614478 299548 614578
rect 299648 614478 299772 614578
rect 299872 614478 299996 614578
rect 300096 614478 300220 614578
rect 300320 614478 300444 614578
rect 300544 614478 300668 614578
rect 300768 614478 300892 614578
rect 300992 614478 301116 614578
rect 301216 614478 301340 614578
rect 301440 614478 301564 614578
rect 301664 614478 301788 614578
rect 301888 614478 302012 614578
rect 302112 614478 302236 614578
rect 302336 614478 302460 614578
rect 302560 614478 302684 614578
rect 302784 614478 302908 614578
rect 303008 614478 303132 614578
rect 303232 614478 303356 614578
rect 303456 614478 303580 614578
rect 303680 614478 303804 614578
rect 303904 614478 304028 614578
rect 304128 614478 304252 614578
rect 304352 614478 304476 614578
rect 304576 614478 304700 614578
rect 304800 614478 304924 614578
rect 305024 614478 305148 614578
rect 305248 614478 305372 614578
rect 305472 614478 305477 614578
rect 298820 614473 305477 614478
rect 309290 614578 315947 614583
rect 309290 614478 309346 614578
rect 309446 614478 309570 614578
rect 309670 614478 309794 614578
rect 309894 614478 310018 614578
rect 310118 614478 310242 614578
rect 310342 614478 310466 614578
rect 310566 614478 310690 614578
rect 310790 614478 310914 614578
rect 311014 614478 311138 614578
rect 311238 614478 311362 614578
rect 311462 614478 311586 614578
rect 311686 614478 311810 614578
rect 311910 614478 312034 614578
rect 312134 614478 312258 614578
rect 312358 614478 312482 614578
rect 312582 614478 312706 614578
rect 312806 614478 312930 614578
rect 313030 614478 313154 614578
rect 313254 614478 313378 614578
rect 313478 614478 313602 614578
rect 313702 614478 313826 614578
rect 313926 614478 314050 614578
rect 314150 614478 314274 614578
rect 314374 614478 314498 614578
rect 314598 614478 314722 614578
rect 314822 614478 314946 614578
rect 315046 614478 315170 614578
rect 315270 614478 315394 614578
rect 315494 614478 315618 614578
rect 315718 614478 315842 614578
rect 315942 614478 315947 614578
rect 309290 614473 315947 614478
rect 335560 614498 335616 614598
rect 335716 614498 335840 614598
rect 335940 614498 336064 614598
rect 336164 614498 336288 614598
rect 336388 614498 336512 614598
rect 336612 614498 336736 614598
rect 336836 614498 336960 614598
rect 337060 614498 337184 614598
rect 337284 614498 337408 614598
rect 337508 614498 337632 614598
rect 337732 614498 337856 614598
rect 337956 614498 338080 614598
rect 338180 614498 338304 614598
rect 338404 614498 338528 614598
rect 338628 614498 338752 614598
rect 338852 614498 338976 614598
rect 339076 614498 339200 614598
rect 339300 614498 339424 614598
rect 339524 614498 339648 614598
rect 339748 614498 339872 614598
rect 339972 614498 340096 614598
rect 340196 614498 340320 614598
rect 340420 614498 340544 614598
rect 340644 614498 340768 614598
rect 340868 614498 340992 614598
rect 341092 614498 341216 614598
rect 341316 614498 341440 614598
rect 341540 614498 341664 614598
rect 341764 614498 341888 614598
rect 341988 614498 342112 614598
rect 342212 614498 342217 614598
rect 335560 614493 342217 614498
rect 298820 614444 305476 614473
rect 309290 614444 315946 614473
rect 335560 614464 342216 614493
rect 316300 611176 525804 611206
rect 285800 611084 525804 611176
rect 285800 611080 336480 611084
rect 285800 610764 298920 611080
rect 285800 605020 289920 610764
rect 294704 605336 298920 610764
rect 303704 605336 304920 611080
rect 309704 605336 310920 611080
rect 315704 605340 336480 611080
rect 341264 610761 525804 611084
rect 341264 605340 510602 610761
rect 315704 605336 510602 605340
rect 294704 605020 510602 605336
rect 285800 605017 510602 605020
rect 515386 605017 520602 610761
rect 525386 605017 525804 610761
rect 285800 604544 525804 605017
rect 285800 604520 316300 604544
rect 560425 597806 566979 629792
rect 316064 597324 566979 597806
rect 316064 591580 317480 597324
rect 322264 591580 325480 597324
rect 330264 591580 566979 597324
rect 316064 591240 566979 591580
rect 316060 591140 566980 591240
rect 556059 555354 562613 559520
rect 556059 550570 556255 555354
rect 562319 550570 562613 555354
rect 556059 545354 562613 550570
rect 556059 540570 556255 545354
rect 562319 540570 562613 545354
rect 556059 540155 562613 540570
rect 573464 500138 576816 500473
rect 573464 500074 573553 500138
rect 573617 500074 573633 500138
rect 573697 500074 573713 500138
rect 573777 500074 573793 500138
rect 573857 500074 573873 500138
rect 573937 500074 573953 500138
rect 574017 500074 574033 500138
rect 574097 500074 574113 500138
rect 574177 500074 574193 500138
rect 574257 500074 574273 500138
rect 574337 500074 574353 500138
rect 574417 500074 574433 500138
rect 574497 500074 574513 500138
rect 574577 500074 574593 500138
rect 574657 500074 574673 500138
rect 574737 500074 574753 500138
rect 574817 500074 574833 500138
rect 574897 500074 574913 500138
rect 574977 500074 574993 500138
rect 575057 500074 575073 500138
rect 575137 500074 575153 500138
rect 575217 500074 575233 500138
rect 575297 500074 575313 500138
rect 575377 500074 575393 500138
rect 575457 500074 575473 500138
rect 575537 500074 575553 500138
rect 575617 500074 575633 500138
rect 575697 500074 575713 500138
rect 575777 500074 575793 500138
rect 575857 500074 575873 500138
rect 575937 500074 575953 500138
rect 576017 500074 576033 500138
rect 576097 500074 576113 500138
rect 576177 500074 576193 500138
rect 576257 500074 576273 500138
rect 576337 500074 576353 500138
rect 576417 500074 576433 500138
rect 576497 500074 576513 500138
rect 576577 500074 576593 500138
rect 576657 500074 576673 500138
rect 576737 500074 576816 500138
rect 13814 462486 17684 462771
rect 13814 462422 13897 462486
rect 13961 462422 13977 462486
rect 14041 462422 14057 462486
rect 14121 462422 14137 462486
rect 14201 462422 14217 462486
rect 14281 462422 14297 462486
rect 14361 462422 14377 462486
rect 14441 462422 14457 462486
rect 14521 462422 14537 462486
rect 14601 462422 14617 462486
rect 14681 462422 14697 462486
rect 14761 462422 14777 462486
rect 14841 462422 14857 462486
rect 14921 462422 14937 462486
rect 15001 462422 15017 462486
rect 15081 462422 15097 462486
rect 15161 462422 15177 462486
rect 15241 462422 15257 462486
rect 15321 462422 15337 462486
rect 15401 462422 15417 462486
rect 15481 462422 15497 462486
rect 15561 462422 15577 462486
rect 15641 462422 15657 462486
rect 15721 462422 15737 462486
rect 15801 462422 15817 462486
rect 15881 462422 15897 462486
rect 15961 462422 15977 462486
rect 16041 462422 16057 462486
rect 16121 462422 16137 462486
rect 16201 462422 16217 462486
rect 16281 462422 16297 462486
rect 16361 462422 16377 462486
rect 16441 462422 16457 462486
rect 16521 462422 16537 462486
rect 16601 462422 16617 462486
rect 16681 462422 16697 462486
rect 16761 462422 16777 462486
rect 16841 462422 16857 462486
rect 16921 462422 16937 462486
rect 17001 462422 17017 462486
rect 17081 462422 17097 462486
rect 17161 462422 17177 462486
rect 17241 462422 17257 462486
rect 17321 462422 17337 462486
rect 17401 462422 17417 462486
rect 17481 462422 17497 462486
rect 17561 462422 17684 462486
rect 13814 419264 17684 462422
rect 13814 419200 13911 419264
rect 13975 419200 13991 419264
rect 14055 419200 14071 419264
rect 14135 419200 14151 419264
rect 14215 419200 14231 419264
rect 14295 419200 14311 419264
rect 14375 419200 14391 419264
rect 14455 419200 14471 419264
rect 14535 419200 14551 419264
rect 14615 419200 14631 419264
rect 14695 419200 14711 419264
rect 14775 419200 14791 419264
rect 14855 419200 14871 419264
rect 14935 419200 14951 419264
rect 15015 419200 15031 419264
rect 15095 419200 15111 419264
rect 15175 419200 15191 419264
rect 15255 419200 15271 419264
rect 15335 419200 15351 419264
rect 15415 419200 15431 419264
rect 15495 419200 15511 419264
rect 15575 419200 15591 419264
rect 15655 419200 15671 419264
rect 15735 419200 15751 419264
rect 15815 419200 15831 419264
rect 15895 419200 15911 419264
rect 15975 419200 15991 419264
rect 16055 419200 16071 419264
rect 16135 419200 16151 419264
rect 16215 419200 16231 419264
rect 16295 419200 16311 419264
rect 16375 419200 16391 419264
rect 16455 419200 16471 419264
rect 16535 419200 16551 419264
rect 16615 419200 16631 419264
rect 16695 419200 16711 419264
rect 16775 419200 16791 419264
rect 16855 419200 16871 419264
rect 16935 419200 16951 419264
rect 17015 419200 17031 419264
rect 17095 419200 17111 419264
rect 17175 419200 17191 419264
rect 17255 419200 17271 419264
rect 17335 419200 17351 419264
rect 17415 419200 17431 419264
rect 17495 419200 17511 419264
rect 17575 419200 17684 419264
rect 13814 227257 17684 419200
rect 573464 455716 576816 500074
rect 573464 455652 573591 455716
rect 573655 455652 573671 455716
rect 573735 455652 573751 455716
rect 573815 455652 573831 455716
rect 573895 455652 573911 455716
rect 573975 455652 573991 455716
rect 574055 455652 574071 455716
rect 574135 455652 574151 455716
rect 574215 455652 574231 455716
rect 574295 455652 574311 455716
rect 574375 455652 574391 455716
rect 574455 455652 574471 455716
rect 574535 455652 574551 455716
rect 574615 455652 574631 455716
rect 574695 455652 574711 455716
rect 574775 455652 574791 455716
rect 574855 455652 574871 455716
rect 574935 455652 574951 455716
rect 575015 455652 575031 455716
rect 575095 455652 575111 455716
rect 575175 455652 575191 455716
rect 575255 455652 575271 455716
rect 575335 455652 575351 455716
rect 575415 455652 575431 455716
rect 575495 455652 575511 455716
rect 575575 455652 575591 455716
rect 575655 455652 575671 455716
rect 575735 455652 575751 455716
rect 575815 455652 575831 455716
rect 575895 455652 575911 455716
rect 575975 455652 575991 455716
rect 576055 455652 576071 455716
rect 576135 455652 576151 455716
rect 576215 455652 576231 455716
rect 576295 455652 576311 455716
rect 576375 455652 576391 455716
rect 576455 455652 576471 455716
rect 576535 455652 576551 455716
rect 576615 455652 576631 455716
rect 576695 455652 576816 455716
rect 13811 196222 17688 227257
rect 13811 191438 13997 196222
rect 17421 191438 17688 196222
rect 13811 191098 17688 191438
rect 573464 196222 576816 455652
rect 573464 191438 573605 196222
rect 576629 191438 576816 196222
rect 573464 191191 576816 191438
<< via4 >>
rect 312958 626314 333268 627286
<< mimcap2 >>
rect 300726 639272 301126 639312
rect 300726 638952 300766 639272
rect 301086 638952 301126 639272
rect 300726 638912 301126 638952
rect 301848 639272 302248 639312
rect 301848 638952 301888 639272
rect 302208 638952 302248 639272
rect 301848 638912 302248 638952
rect 302970 639272 303370 639312
rect 302970 638952 303010 639272
rect 303330 638952 303370 639272
rect 302970 638912 303370 638952
rect 304092 639272 304492 639312
rect 304092 638952 304132 639272
rect 304452 638952 304492 639272
rect 304092 638912 304492 638952
rect 305214 639272 305614 639312
rect 305214 638952 305254 639272
rect 305574 638952 305614 639272
rect 305214 638912 305614 638952
rect 306336 639272 306736 639312
rect 306336 638952 306376 639272
rect 306696 638952 306736 639272
rect 306336 638912 306736 638952
rect 307458 639272 307858 639312
rect 307458 638952 307498 639272
rect 307818 638952 307858 639272
rect 307458 638912 307858 638952
rect 308580 639272 308980 639312
rect 308580 638952 308620 639272
rect 308940 638952 308980 639272
rect 308580 638912 308980 638952
rect 309702 639272 310102 639312
rect 309702 638952 309742 639272
rect 310062 638952 310102 639272
rect 309702 638912 310102 638952
rect 310824 639272 311224 639312
rect 310824 638952 310864 639272
rect 311184 638952 311224 639272
rect 310824 638912 311224 638952
rect 300726 638572 301126 638612
rect 300726 638252 300766 638572
rect 301086 638252 301126 638572
rect 300726 638212 301126 638252
rect 301848 638572 302248 638612
rect 301848 638252 301888 638572
rect 302208 638252 302248 638572
rect 301848 638212 302248 638252
rect 302970 638572 303370 638612
rect 302970 638252 303010 638572
rect 303330 638252 303370 638572
rect 302970 638212 303370 638252
rect 304092 638572 304492 638612
rect 304092 638252 304132 638572
rect 304452 638252 304492 638572
rect 304092 638212 304492 638252
rect 305214 638572 305614 638612
rect 305214 638252 305254 638572
rect 305574 638252 305614 638572
rect 305214 638212 305614 638252
rect 306336 638572 306736 638612
rect 306336 638252 306376 638572
rect 306696 638252 306736 638572
rect 306336 638212 306736 638252
rect 307458 638572 307858 638612
rect 307458 638252 307498 638572
rect 307818 638252 307858 638572
rect 307458 638212 307858 638252
rect 308580 638572 308980 638612
rect 308580 638252 308620 638572
rect 308940 638252 308980 638572
rect 308580 638212 308980 638252
rect 309702 638572 310102 638612
rect 309702 638252 309742 638572
rect 310062 638252 310102 638572
rect 309702 638212 310102 638252
rect 310824 638572 311224 638612
rect 310824 638252 310864 638572
rect 311184 638252 311224 638572
rect 310824 638212 311224 638252
rect 300726 637872 301126 637912
rect 300726 637552 300766 637872
rect 301086 637552 301126 637872
rect 300726 637512 301126 637552
rect 301848 637872 302248 637912
rect 301848 637552 301888 637872
rect 302208 637552 302248 637872
rect 301848 637512 302248 637552
rect 302970 637872 303370 637912
rect 302970 637552 303010 637872
rect 303330 637552 303370 637872
rect 302970 637512 303370 637552
rect 304092 637872 304492 637912
rect 304092 637552 304132 637872
rect 304452 637552 304492 637872
rect 304092 637512 304492 637552
rect 305214 637872 305614 637912
rect 305214 637552 305254 637872
rect 305574 637552 305614 637872
rect 305214 637512 305614 637552
rect 306336 637872 306736 637912
rect 306336 637552 306376 637872
rect 306696 637552 306736 637872
rect 306336 637512 306736 637552
rect 307458 637872 307858 637912
rect 307458 637552 307498 637872
rect 307818 637552 307858 637872
rect 307458 637512 307858 637552
rect 308580 637872 308980 637912
rect 308580 637552 308620 637872
rect 308940 637552 308980 637872
rect 308580 637512 308980 637552
rect 309702 637872 310102 637912
rect 309702 637552 309742 637872
rect 310062 637552 310102 637872
rect 309702 637512 310102 637552
rect 310824 637872 311224 637912
rect 310824 637552 310864 637872
rect 311184 637552 311224 637872
rect 310824 637512 311224 637552
rect 300726 637172 301126 637212
rect 300726 636852 300766 637172
rect 301086 636852 301126 637172
rect 300726 636812 301126 636852
rect 301848 637172 302248 637212
rect 301848 636852 301888 637172
rect 302208 636852 302248 637172
rect 301848 636812 302248 636852
rect 302970 637172 303370 637212
rect 302970 636852 303010 637172
rect 303330 636852 303370 637172
rect 302970 636812 303370 636852
rect 304092 637172 304492 637212
rect 304092 636852 304132 637172
rect 304452 636852 304492 637172
rect 304092 636812 304492 636852
rect 305214 637172 305614 637212
rect 305214 636852 305254 637172
rect 305574 636852 305614 637172
rect 305214 636812 305614 636852
rect 306336 637172 306736 637212
rect 306336 636852 306376 637172
rect 306696 636852 306736 637172
rect 306336 636812 306736 636852
rect 307458 637172 307858 637212
rect 307458 636852 307498 637172
rect 307818 636852 307858 637172
rect 307458 636812 307858 636852
rect 308580 637172 308980 637212
rect 308580 636852 308620 637172
rect 308940 636852 308980 637172
rect 308580 636812 308980 636852
rect 309702 637172 310102 637212
rect 309702 636852 309742 637172
rect 310062 636852 310102 637172
rect 309702 636812 310102 636852
rect 310824 637172 311224 637212
rect 310824 636852 310864 637172
rect 311184 636852 311224 637172
rect 310824 636812 311224 636852
rect 300726 636472 301126 636512
rect 300726 636152 300766 636472
rect 301086 636152 301126 636472
rect 300726 636112 301126 636152
rect 301848 636472 302248 636512
rect 301848 636152 301888 636472
rect 302208 636152 302248 636472
rect 301848 636112 302248 636152
rect 302970 636472 303370 636512
rect 302970 636152 303010 636472
rect 303330 636152 303370 636472
rect 302970 636112 303370 636152
rect 304092 636472 304492 636512
rect 304092 636152 304132 636472
rect 304452 636152 304492 636472
rect 304092 636112 304492 636152
rect 305214 636472 305614 636512
rect 305214 636152 305254 636472
rect 305574 636152 305614 636472
rect 305214 636112 305614 636152
rect 306336 636472 306736 636512
rect 306336 636152 306376 636472
rect 306696 636152 306736 636472
rect 306336 636112 306736 636152
rect 307458 636472 307858 636512
rect 307458 636152 307498 636472
rect 307818 636152 307858 636472
rect 307458 636112 307858 636152
rect 308580 636472 308980 636512
rect 308580 636152 308620 636472
rect 308940 636152 308980 636472
rect 308580 636112 308980 636152
rect 309702 636472 310102 636512
rect 309702 636152 309742 636472
rect 310062 636152 310102 636472
rect 309702 636112 310102 636152
rect 310824 636472 311224 636512
rect 310824 636152 310864 636472
rect 311184 636152 311224 636472
rect 310824 636112 311224 636152
rect 300726 635772 301126 635812
rect 300726 635452 300766 635772
rect 301086 635452 301126 635772
rect 300726 635412 301126 635452
rect 301848 635772 302248 635812
rect 301848 635452 301888 635772
rect 302208 635452 302248 635772
rect 301848 635412 302248 635452
rect 302970 635772 303370 635812
rect 302970 635452 303010 635772
rect 303330 635452 303370 635772
rect 302970 635412 303370 635452
rect 304092 635772 304492 635812
rect 304092 635452 304132 635772
rect 304452 635452 304492 635772
rect 304092 635412 304492 635452
rect 305214 635772 305614 635812
rect 305214 635452 305254 635772
rect 305574 635452 305614 635772
rect 305214 635412 305614 635452
rect 306336 635772 306736 635812
rect 306336 635452 306376 635772
rect 306696 635452 306736 635772
rect 306336 635412 306736 635452
rect 307458 635772 307858 635812
rect 307458 635452 307498 635772
rect 307818 635452 307858 635772
rect 307458 635412 307858 635452
rect 308580 635772 308980 635812
rect 308580 635452 308620 635772
rect 308940 635452 308980 635772
rect 308580 635412 308980 635452
rect 309702 635772 310102 635812
rect 309702 635452 309742 635772
rect 310062 635452 310102 635772
rect 309702 635412 310102 635452
rect 310824 635772 311224 635812
rect 310824 635452 310864 635772
rect 311184 635452 311224 635772
rect 310824 635412 311224 635452
rect 300726 635072 301126 635112
rect 300726 634752 300766 635072
rect 301086 634752 301126 635072
rect 300726 634712 301126 634752
rect 301848 635072 302248 635112
rect 301848 634752 301888 635072
rect 302208 634752 302248 635072
rect 301848 634712 302248 634752
rect 302970 635072 303370 635112
rect 302970 634752 303010 635072
rect 303330 634752 303370 635072
rect 302970 634712 303370 634752
rect 304092 635072 304492 635112
rect 304092 634752 304132 635072
rect 304452 634752 304492 635072
rect 304092 634712 304492 634752
rect 305214 635072 305614 635112
rect 305214 634752 305254 635072
rect 305574 634752 305614 635072
rect 305214 634712 305614 634752
rect 306336 635072 306736 635112
rect 306336 634752 306376 635072
rect 306696 634752 306736 635072
rect 306336 634712 306736 634752
rect 307458 635072 307858 635112
rect 307458 634752 307498 635072
rect 307818 634752 307858 635072
rect 307458 634712 307858 634752
rect 308580 635072 308980 635112
rect 308580 634752 308620 635072
rect 308940 634752 308980 635072
rect 308580 634712 308980 634752
rect 309702 635072 310102 635112
rect 309702 634752 309742 635072
rect 310062 634752 310102 635072
rect 309702 634712 310102 634752
rect 310824 635072 311224 635112
rect 310824 634752 310864 635072
rect 311184 634752 311224 635072
rect 310824 634712 311224 634752
rect 300726 634372 301126 634412
rect 300726 634052 300766 634372
rect 301086 634052 301126 634372
rect 300726 634012 301126 634052
rect 301848 634372 302248 634412
rect 301848 634052 301888 634372
rect 302208 634052 302248 634372
rect 301848 634012 302248 634052
rect 302970 634372 303370 634412
rect 302970 634052 303010 634372
rect 303330 634052 303370 634372
rect 302970 634012 303370 634052
rect 304092 634372 304492 634412
rect 304092 634052 304132 634372
rect 304452 634052 304492 634372
rect 304092 634012 304492 634052
rect 305214 634372 305614 634412
rect 305214 634052 305254 634372
rect 305574 634052 305614 634372
rect 305214 634012 305614 634052
rect 306336 634372 306736 634412
rect 306336 634052 306376 634372
rect 306696 634052 306736 634372
rect 306336 634012 306736 634052
rect 307458 634372 307858 634412
rect 307458 634052 307498 634372
rect 307818 634052 307858 634372
rect 307458 634012 307858 634052
rect 308580 634372 308980 634412
rect 308580 634052 308620 634372
rect 308940 634052 308980 634372
rect 308580 634012 308980 634052
rect 309702 634372 310102 634412
rect 309702 634052 309742 634372
rect 310062 634052 310102 634372
rect 309702 634012 310102 634052
rect 310824 634372 311224 634412
rect 310824 634052 310864 634372
rect 311184 634052 311224 634372
rect 310824 634012 311224 634052
rect 300726 633672 301126 633712
rect 300726 633352 300766 633672
rect 301086 633352 301126 633672
rect 300726 633312 301126 633352
rect 301848 633672 302248 633712
rect 301848 633352 301888 633672
rect 302208 633352 302248 633672
rect 301848 633312 302248 633352
rect 302970 633672 303370 633712
rect 302970 633352 303010 633672
rect 303330 633352 303370 633672
rect 302970 633312 303370 633352
rect 304092 633672 304492 633712
rect 304092 633352 304132 633672
rect 304452 633352 304492 633672
rect 304092 633312 304492 633352
rect 305214 633672 305614 633712
rect 305214 633352 305254 633672
rect 305574 633352 305614 633672
rect 305214 633312 305614 633352
rect 306336 633672 306736 633712
rect 306336 633352 306376 633672
rect 306696 633352 306736 633672
rect 306336 633312 306736 633352
rect 307458 633672 307858 633712
rect 307458 633352 307498 633672
rect 307818 633352 307858 633672
rect 307458 633312 307858 633352
rect 308580 633672 308980 633712
rect 308580 633352 308620 633672
rect 308940 633352 308980 633672
rect 308580 633312 308980 633352
rect 309702 633672 310102 633712
rect 309702 633352 309742 633672
rect 310062 633352 310102 633672
rect 309702 633312 310102 633352
rect 310824 633672 311224 633712
rect 310824 633352 310864 633672
rect 311184 633352 311224 633672
rect 310824 633312 311224 633352
rect 300726 632972 301126 633012
rect 300726 632652 300766 632972
rect 301086 632652 301126 632972
rect 300726 632612 301126 632652
rect 301848 632972 302248 633012
rect 301848 632652 301888 632972
rect 302208 632652 302248 632972
rect 301848 632612 302248 632652
rect 302970 632972 303370 633012
rect 302970 632652 303010 632972
rect 303330 632652 303370 632972
rect 302970 632612 303370 632652
rect 304092 632972 304492 633012
rect 304092 632652 304132 632972
rect 304452 632652 304492 632972
rect 304092 632612 304492 632652
rect 305214 632972 305614 633012
rect 305214 632652 305254 632972
rect 305574 632652 305614 632972
rect 305214 632612 305614 632652
rect 306336 632972 306736 633012
rect 306336 632652 306376 632972
rect 306696 632652 306736 632972
rect 306336 632612 306736 632652
rect 307458 632972 307858 633012
rect 307458 632652 307498 632972
rect 307818 632652 307858 632972
rect 307458 632612 307858 632652
rect 308580 632972 308980 633012
rect 308580 632652 308620 632972
rect 308940 632652 308980 632972
rect 308580 632612 308980 632652
rect 309702 632972 310102 633012
rect 309702 632652 309742 632972
rect 310062 632652 310102 632972
rect 309702 632612 310102 632652
rect 310824 632972 311224 633012
rect 310824 632652 310864 632972
rect 311184 632652 311224 632972
rect 310824 632612 311224 632652
<< mimcap2contact >>
rect 300766 638952 301086 639272
rect 301888 638952 302208 639272
rect 303010 638952 303330 639272
rect 304132 638952 304452 639272
rect 305254 638952 305574 639272
rect 306376 638952 306696 639272
rect 307498 638952 307818 639272
rect 308620 638952 308940 639272
rect 309742 638952 310062 639272
rect 310864 638952 311184 639272
rect 300766 638252 301086 638572
rect 301888 638252 302208 638572
rect 303010 638252 303330 638572
rect 304132 638252 304452 638572
rect 305254 638252 305574 638572
rect 306376 638252 306696 638572
rect 307498 638252 307818 638572
rect 308620 638252 308940 638572
rect 309742 638252 310062 638572
rect 310864 638252 311184 638572
rect 300766 637552 301086 637872
rect 301888 637552 302208 637872
rect 303010 637552 303330 637872
rect 304132 637552 304452 637872
rect 305254 637552 305574 637872
rect 306376 637552 306696 637872
rect 307498 637552 307818 637872
rect 308620 637552 308940 637872
rect 309742 637552 310062 637872
rect 310864 637552 311184 637872
rect 300766 636852 301086 637172
rect 301888 636852 302208 637172
rect 303010 636852 303330 637172
rect 304132 636852 304452 637172
rect 305254 636852 305574 637172
rect 306376 636852 306696 637172
rect 307498 636852 307818 637172
rect 308620 636852 308940 637172
rect 309742 636852 310062 637172
rect 310864 636852 311184 637172
rect 300766 636152 301086 636472
rect 301888 636152 302208 636472
rect 303010 636152 303330 636472
rect 304132 636152 304452 636472
rect 305254 636152 305574 636472
rect 306376 636152 306696 636472
rect 307498 636152 307818 636472
rect 308620 636152 308940 636472
rect 309742 636152 310062 636472
rect 310864 636152 311184 636472
rect 300766 635452 301086 635772
rect 301888 635452 302208 635772
rect 303010 635452 303330 635772
rect 304132 635452 304452 635772
rect 305254 635452 305574 635772
rect 306376 635452 306696 635772
rect 307498 635452 307818 635772
rect 308620 635452 308940 635772
rect 309742 635452 310062 635772
rect 310864 635452 311184 635772
rect 300766 634752 301086 635072
rect 301888 634752 302208 635072
rect 303010 634752 303330 635072
rect 304132 634752 304452 635072
rect 305254 634752 305574 635072
rect 306376 634752 306696 635072
rect 307498 634752 307818 635072
rect 308620 634752 308940 635072
rect 309742 634752 310062 635072
rect 310864 634752 311184 635072
rect 300766 634052 301086 634372
rect 301888 634052 302208 634372
rect 303010 634052 303330 634372
rect 304132 634052 304452 634372
rect 305254 634052 305574 634372
rect 306376 634052 306696 634372
rect 307498 634052 307818 634372
rect 308620 634052 308940 634372
rect 309742 634052 310062 634372
rect 310864 634052 311184 634372
rect 300766 633352 301086 633672
rect 301888 633352 302208 633672
rect 303010 633352 303330 633672
rect 304132 633352 304452 633672
rect 305254 633352 305574 633672
rect 306376 633352 306696 633672
rect 307498 633352 307818 633672
rect 308620 633352 308940 633672
rect 309742 633352 310062 633672
rect 310864 633352 311184 633672
rect 300766 632652 301086 632972
rect 301888 632652 302208 632972
rect 303010 632652 303330 632972
rect 304132 632652 304452 632972
rect 305254 632652 305574 632972
rect 306376 632652 306696 632972
rect 307498 632652 307818 632972
rect 308620 632652 308940 632972
rect 309742 632652 310062 632972
rect 310864 632652 311184 632972
<< metal5 >>
rect 300672 639456 333286 639731
rect 300672 639272 333442 639456
rect 300672 638952 300766 639272
rect 301086 638952 301888 639272
rect 302208 638952 303010 639272
rect 303330 638952 304132 639272
rect 304452 638952 305254 639272
rect 305574 638952 306376 639272
rect 306696 638952 307498 639272
rect 307818 638952 308620 639272
rect 308940 638952 309742 639272
rect 310062 638952 310864 639272
rect 311184 638952 333442 639272
rect 300672 638572 333442 638952
rect 300672 638252 300766 638572
rect 301086 638252 301888 638572
rect 302208 638252 303010 638572
rect 303330 638252 304132 638572
rect 304452 638252 305254 638572
rect 305574 638252 306376 638572
rect 306696 638252 307498 638572
rect 307818 638252 308620 638572
rect 308940 638252 309742 638572
rect 310062 638252 310864 638572
rect 311184 638252 333442 638572
rect 300672 637872 333442 638252
rect 300672 637552 300766 637872
rect 301086 637552 301888 637872
rect 302208 637552 303010 637872
rect 303330 637552 304132 637872
rect 304452 637552 305254 637872
rect 305574 637552 306376 637872
rect 306696 637552 307498 637872
rect 307818 637552 308620 637872
rect 308940 637552 309742 637872
rect 310062 637552 310864 637872
rect 311184 637552 333442 637872
rect 300672 637172 333442 637552
rect 300672 636852 300766 637172
rect 301086 636852 301888 637172
rect 302208 636852 303010 637172
rect 303330 636852 304132 637172
rect 304452 636852 305254 637172
rect 305574 636852 306376 637172
rect 306696 636852 307498 637172
rect 307818 636852 308620 637172
rect 308940 636852 309742 637172
rect 310062 636852 310864 637172
rect 311184 636852 333442 637172
rect 300672 636472 333442 636852
rect 300672 636152 300766 636472
rect 301086 636152 301888 636472
rect 302208 636152 303010 636472
rect 303330 636152 304132 636472
rect 304452 636152 305254 636472
rect 305574 636152 306376 636472
rect 306696 636152 307498 636472
rect 307818 636152 308620 636472
rect 308940 636152 309742 636472
rect 310062 636152 310864 636472
rect 311184 636152 333442 636472
rect 300672 635772 333442 636152
rect 300672 635452 300766 635772
rect 301086 635452 301888 635772
rect 302208 635452 303010 635772
rect 303330 635452 304132 635772
rect 304452 635452 305254 635772
rect 305574 635452 306376 635772
rect 306696 635452 307498 635772
rect 307818 635452 308620 635772
rect 308940 635452 309742 635772
rect 310062 635452 310864 635772
rect 311184 635452 333442 635772
rect 300672 635072 333442 635452
rect 300672 634752 300766 635072
rect 301086 634752 301888 635072
rect 302208 634752 303010 635072
rect 303330 634752 304132 635072
rect 304452 634752 305254 635072
rect 305574 634752 306376 635072
rect 306696 634752 307498 635072
rect 307818 634752 308620 635072
rect 308940 634752 309742 635072
rect 310062 634752 310864 635072
rect 311184 634752 333442 635072
rect 300672 634372 333442 634752
rect 300672 634052 300766 634372
rect 301086 634052 301888 634372
rect 302208 634052 303010 634372
rect 303330 634052 304132 634372
rect 304452 634052 305254 634372
rect 305574 634052 306376 634372
rect 306696 634052 307498 634372
rect 307818 634052 308620 634372
rect 308940 634052 309742 634372
rect 310062 634052 310864 634372
rect 311184 634052 333442 634372
rect 300672 633672 333442 634052
rect 300672 633352 300766 633672
rect 301086 633352 301888 633672
rect 302208 633352 303010 633672
rect 303330 633352 304132 633672
rect 304452 633352 305254 633672
rect 305574 633352 306376 633672
rect 306696 633352 307498 633672
rect 307818 633352 308620 633672
rect 308940 633352 309742 633672
rect 310062 633352 310864 633672
rect 311184 633352 333442 633672
rect 300672 632972 333442 633352
rect 300672 632652 300766 632972
rect 301086 632652 301888 632972
rect 302208 632652 303010 632972
rect 303330 632652 304132 632972
rect 304452 632652 305254 632972
rect 305574 632652 306376 632972
rect 306696 632652 307498 632972
rect 307818 632652 308620 632972
rect 308940 632652 309742 632972
rect 310062 632652 310864 632972
rect 311184 632652 333442 632972
rect 300672 627286 333442 632652
rect 300672 626314 312958 627286
rect 333268 626314 333442 627286
rect 300672 626254 333442 626314
rect 312958 626216 333442 626254
<< res2p85 >>
rect 313270 632356 313844 635684
rect 314088 632356 314662 635684
rect 314906 632356 315480 635684
rect 316542 632766 317116 637070
rect 317360 632766 317934 637070
rect 318178 632766 318752 637070
rect 318996 632766 319570 637070
rect 321450 630700 322024 637008
rect 322268 630700 322842 637008
rect 323086 630700 323660 637008
rect 323904 630700 324478 637008
rect 324722 630700 325296 637008
rect 325540 630700 326114 637008
rect 326358 630700 326932 637008
rect 327176 630700 327750 637008
rect 327994 630700 328568 637008
rect 328812 630700 329386 637008
rect 329630 630700 330204 637008
rect 330448 630700 331022 637008
rect 331266 630700 331840 637008
rect 332084 630700 332658 637008
rect 332902 630700 333476 637008
rect 333720 630700 334294 637008
rect 334538 630700 335112 637008
<< pnp3p40 >>
rect 334944 617724 340788 627424
<< labels >>
flabel metal3 s 572152 640142 580220 644150 0 FreeSans 20000 0 0 0 VCCD1
flabel metal3 s 567038 550960 577302 554546 0 FreeSans 20000 0 0 0 VDDA1
flabel metal3 s 511190 664896 514962 676272 0 FreeSans 20000 90 0 0 VSSA1
flabel metal3 s 561703 191929 571721 195859 0 FreeSans 20000 0 0 0 VSSD1
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
flabel metal1 302950 624008 303412 624206 1 FreeSans 1600 0 0 0 bandgaptop_flat_0/porst
flabel metal1 319346 628330 324014 629006 1 FreeSans 1600 0 0 0 bandgaptop_flat_0/Vbg
flabel metal2 300892 620234 302674 620304 1 FreeSans 800 0 0 0 bandgaptop_flat_0/ampcurrentsource_0/Vq
flabel metal2 300892 620444 302674 620514 1 FreeSans 800 0 0 0 bandgaptop_flat_0/ampcurrentsource_0/Vx
flabel locali 301752 621204 301834 621232 1 FreeSans 800 0 0 0 bandgaptop_flat_0/ampcurrentsource_0/GND!
flabel metal2 307644 616944 307660 617068 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/VDD!
flabel metal2 308298 620172 308314 620296 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Vq
flabel metal2 308240 622432 308256 622512 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Va
flabel metal2 307468 622292 307484 622372 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Vb
flabel metal2 308974 619876 309068 620142 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Vgate
flabel metal2 307250 619876 307344 620142 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Vgate
flabel metal1 305892 619890 305926 619982 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/vg
flabel metal2 309992 616744 310014 616868 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/Vx
flabel psubdiffcont 304770 620548 304870 622148 5 FreeSans 800 0 0 0 bandgaptop_flat_0/amplifier_0/GND!
flabel psubdiff 310220 622148 310420 622248 5 FreeSans 800 180 0 0 bandgaptop_flat_0/amplifier_0/GND!
rlabel via1 314086 616924 314132 616968 5 bandgaptop_flat_0/currentmirror_0/Vgate
rlabel metal3 314808 616568 314942 616686 5 bandgaptop_flat_0/currentmirror_0/VDD!
flabel metal1 321614 625108 321914 625208 5 FreeSans 1600 0 0 0 bandgaptop_flat_0/currentmirror_0/Vbg
flabel metal2 321614 625708 321814 625808 5 FreeSans 1600 0 0 0 bandgaptop_flat_0/currentmirror_0/Vb
flabel metal2 321614 626308 321814 626408 5 FreeSans 1600 0 0 0 bandgaptop_flat_0/currentmirror_0/Va
flabel metal2 333810 617726 334946 618674 7 FreeSans 1600 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/Vbneg
flabel metal2 323088 637006 323658 637438 1 FreeSans 800 90 0 0 bandgaptop_flat_0/bandgapcorev3_0/VbEnd
flabel metal2 323906 630270 324476 630702 1 FreeSans 800 90 0 0 bandgaptop_flat_0/bandgapcorev3_0/VbgEnd
flabel metal2 322270 636206 322840 637438 1 FreeSans 800 90 0 0 bandgaptop_flat_0/bandgapcorev3_0/VaEnd
flabel metal2 332014 630004 332706 630696 1 FreeSans 1600 90 0 0 bandgaptop_flat_0/bandgapcorev3_0/Vbg
flabel metal2 333644 629998 334348 630702 1 FreeSans 1600 90 0 0 bandgaptop_flat_0/bandgapcorev3_0/Vb
flabel metal1 332826 629432 333530 630004 3 FreeSans 1600 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/Va
flabel locali 340982 621162 341068 621382 3 FreeSans 1600 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/GND!
flabel locali 340312 627036 340560 627140 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,0]/Emitter
flabel locali 340400 626465 340501 626514 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,0]/Collector
flabel locali 340406 626624 340524 626664 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,0]/Base
flabel locali 339024 627036 339272 627140 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,1]/Emitter
flabel locali 339112 626465 339213 626514 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,1]/Collector
flabel locali 339118 626624 339236 626664 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,1]/Base
flabel locali 337736 627036 337984 627140 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,2]/Emitter
flabel locali 337824 626465 337925 626514 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,2]/Collector
flabel locali 337830 626624 337948 626664 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,2]/Base
flabel locali 336448 627036 336696 627140 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,3]/Emitter
flabel locali 336536 626465 336637 626514 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,3]/Collector
flabel locali 336542 626624 336660 626664 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,3]/Base
flabel locali 335160 627036 335408 627140 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,4]/Emitter
flabel locali 335248 626465 335349 626514 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,4]/Collector
flabel locali 335254 626624 335372 626664 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[0,4]/Base
flabel locali 340312 625748 340560 625852 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,0]/Emitter
flabel locali 340400 625177 340501 625226 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,0]/Collector
flabel locali 340406 625336 340524 625376 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,0]/Base
flabel locali 339024 625748 339272 625852 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,1]/Emitter
flabel locali 339112 625177 339213 625226 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,1]/Collector
flabel locali 339118 625336 339236 625376 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,1]/Base
flabel locali 337736 625748 337984 625852 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,2]/Emitter
flabel locali 337824 625177 337925 625226 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,2]/Collector
flabel locali 337830 625336 337948 625376 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,2]/Base
flabel locali 336448 625748 336696 625852 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,3]/Emitter
flabel locali 336536 625177 336637 625226 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,3]/Collector
flabel locali 336542 625336 336660 625376 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,3]/Base
flabel locali 335160 625748 335408 625852 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,4]/Emitter
flabel locali 335248 625177 335349 625226 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,4]/Collector
flabel locali 335254 625336 335372 625376 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[1,4]/Base
flabel locali 340312 624460 340560 624564 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,0]/Emitter
flabel locali 340400 623889 340501 623938 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,0]/Collector
flabel locali 340406 624048 340524 624088 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,0]/Base
flabel locali 339024 624460 339272 624564 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,1]/Emitter
flabel locali 339112 623889 339213 623938 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,1]/Collector
flabel locali 339118 624048 339236 624088 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,1]/Base
flabel locali 337736 624460 337984 624564 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,2]/Emitter
flabel locali 337824 623889 337925 623938 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,2]/Collector
flabel locali 337830 624048 337948 624088 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,2]/Base
flabel locali 336448 624460 336696 624564 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,3]/Emitter
flabel locali 336536 623889 336637 623938 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,3]/Collector
flabel locali 336542 624048 336660 624088 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,3]/Base
flabel locali 335160 624460 335408 624564 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,4]/Emitter
flabel locali 335248 623889 335349 623938 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,4]/Collector
flabel locali 335254 624048 335372 624088 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[2,4]/Base
flabel locali 340312 623172 340560 623276 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,0]/Emitter
flabel locali 340400 622601 340501 622650 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,0]/Collector
flabel locali 340406 622760 340524 622800 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,0]/Base
flabel locali 339024 623172 339272 623276 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,1]/Emitter
flabel locali 339112 622601 339213 622650 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,1]/Collector
flabel locali 339118 622760 339236 622800 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,1]/Base
flabel locali 337736 623172 337984 623276 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,2]/Emitter
flabel locali 337824 622601 337925 622650 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,2]/Collector
flabel locali 337830 622760 337948 622800 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,2]/Base
flabel locali 336448 623172 336696 623276 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,3]/Emitter
flabel locali 336536 622601 336637 622650 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,3]/Collector
flabel locali 336542 622760 336660 622800 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,3]/Base
flabel locali 335160 623172 335408 623276 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,4]/Emitter
flabel locali 335248 622601 335349 622650 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,4]/Collector
flabel locali 335254 622760 335372 622800 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[3,4]/Base
flabel locali 340312 621884 340560 621988 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,0]/Emitter
flabel locali 340400 621313 340501 621362 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,0]/Collector
flabel locali 340406 621472 340524 621512 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,0]/Base
flabel locali 339024 621884 339272 621988 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,1]/Emitter
flabel locali 339112 621313 339213 621362 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,1]/Collector
flabel locali 339118 621472 339236 621512 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,1]/Base
flabel locali 337736 621884 337984 621988 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,2]/Emitter
flabel locali 337824 621313 337925 621362 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,2]/Collector
flabel locali 337830 621472 337948 621512 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,2]/Base
flabel locali 336448 621884 336696 621988 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,3]/Emitter
flabel locali 336536 621313 336637 621362 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,3]/Collector
flabel locali 336542 621472 336660 621512 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,3]/Base
flabel locali 335160 621884 335408 621988 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,4]/Emitter
flabel locali 335248 621313 335349 621362 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,4]/Collector
flabel locali 335254 621472 335372 621512 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[4,4]/Base
flabel locali 340312 620596 340560 620700 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,0]/Emitter
flabel locali 340400 620025 340501 620074 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,0]/Collector
flabel locali 340406 620184 340524 620224 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,0]/Base
flabel locali 339024 620596 339272 620700 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,1]/Emitter
flabel locali 339112 620025 339213 620074 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,1]/Collector
flabel locali 339118 620184 339236 620224 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,1]/Base
flabel locali 337736 620596 337984 620700 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,2]/Emitter
flabel locali 337824 620025 337925 620074 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,2]/Collector
flabel locali 337830 620184 337948 620224 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,2]/Base
flabel locali 336448 620596 336696 620700 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,3]/Emitter
flabel locali 336536 620025 336637 620074 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,3]/Collector
flabel locali 336542 620184 336660 620224 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,3]/Base
flabel locali 335160 620596 335408 620700 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,4]/Emitter
flabel locali 335248 620025 335349 620074 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,4]/Collector
flabel locali 335254 620184 335372 620224 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[5,4]/Base
flabel locali 340312 619308 340560 619412 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,0]/Emitter
flabel locali 340400 618737 340501 618786 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,0]/Collector
flabel locali 340406 618896 340524 618936 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,0]/Base
flabel locali 339024 619308 339272 619412 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,1]/Emitter
flabel locali 339112 618737 339213 618786 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,1]/Collector
flabel locali 339118 618896 339236 618936 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,1]/Base
flabel locali 337736 619308 337984 619412 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,2]/Emitter
flabel locali 337824 618737 337925 618786 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,2]/Collector
flabel locali 337830 618896 337948 618936 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,2]/Base
flabel locali 336448 619308 336696 619412 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,3]/Emitter
flabel locali 336536 618737 336637 618786 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,3]/Collector
flabel locali 336542 618896 336660 618936 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,3]/Base
flabel locali 335160 619308 335408 619412 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,4]/Emitter
flabel locali 335248 618737 335349 618786 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,4]/Collector
flabel locali 335254 618896 335372 618936 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[6,4]/Base
flabel locali 340312 618020 340560 618124 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,0]/Emitter
flabel locali 340400 617449 340501 617498 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,0]/Collector
flabel locali 340406 617608 340524 617648 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,0]/Base
flabel locali 339024 618020 339272 618124 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,1]/Emitter
flabel locali 339112 617449 339213 617498 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,1]/Collector
flabel locali 339118 617608 339236 617648 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,1]/Base
flabel locali 337736 618020 337984 618124 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,2]/Emitter
flabel locali 337824 617449 337925 617498 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,2]/Collector
flabel locali 337830 617608 337948 617648 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,2]/Base
flabel locali 336448 618020 336696 618124 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,3]/Emitter
flabel locali 336536 617449 336637 617498 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,3]/Collector
flabel locali 336542 617608 336660 617648 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,3]/Base
flabel locali 335160 618020 335408 618124 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,4]/Emitter
flabel locali 335248 617449 335349 617498 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,4]/Collector
flabel locali 335254 617608 335372 617648 0 FreeSans 400 0 0 0 bandgaptop_flat_0/bandgapcorev3_0/sky130_fd_pr__pnp_05v5_W3p40L3p40_0[7,4]/Base
rlabel psubdiffcont 297848 614448 341088 615448 1 bandgaptop_flat_0/GND
rlabel metal3 301938 616506 302648 616928 1 bandgaptop_flat_0/VDD
<< end >>
