magic
tech sky130A
magscale 1 2
timestamp 1620316209
<< nwell >>
rect -396 -13355 396 13355
<< pmoslvt >>
rect -200 4536 200 13136
rect -200 -4300 200 4300
rect -200 -13136 200 -4536
<< pdiff >>
rect -258 13124 -200 13136
rect -258 4548 -246 13124
rect -212 4548 -200 13124
rect -258 4536 -200 4548
rect 200 13124 258 13136
rect 200 4548 212 13124
rect 246 4548 258 13124
rect 200 4536 258 4548
rect -258 4288 -200 4300
rect -258 -4288 -246 4288
rect -212 -4288 -200 4288
rect -258 -4300 -200 -4288
rect 200 4288 258 4300
rect 200 -4288 212 4288
rect 246 -4288 258 4288
rect 200 -4300 258 -4288
rect -258 -4548 -200 -4536
rect -258 -13124 -246 -4548
rect -212 -13124 -200 -4548
rect -258 -13136 -200 -13124
rect 200 -4548 258 -4536
rect 200 -13124 212 -4548
rect 246 -13124 258 -4548
rect 200 -13136 258 -13124
<< pdiffc >>
rect -246 4548 -212 13124
rect 212 4548 246 13124
rect -246 -4288 -212 4288
rect 212 -4288 246 4288
rect -246 -13124 -212 -4548
rect 212 -13124 246 -4548
<< nsubdiff >>
rect -360 13285 360 13319
rect -360 -13285 -326 13285
rect 326 -13285 360 13285
rect -360 -13319 360 -13285
<< poly >>
rect -200 13217 200 13233
rect -200 13183 -184 13217
rect 184 13183 200 13217
rect -200 13136 200 13183
rect -200 4489 200 4536
rect -200 4455 -184 4489
rect 184 4455 200 4489
rect -200 4439 200 4455
rect -200 4381 200 4397
rect -200 4347 -184 4381
rect 184 4347 200 4381
rect -200 4300 200 4347
rect -200 -4347 200 -4300
rect -200 -4381 -184 -4347
rect 184 -4381 200 -4347
rect -200 -4397 200 -4381
rect -200 -4455 200 -4439
rect -200 -4489 -184 -4455
rect 184 -4489 200 -4455
rect -200 -4536 200 -4489
rect -200 -13183 200 -13136
rect -200 -13217 -184 -13183
rect 184 -13217 200 -13183
rect -200 -13233 200 -13217
<< polycont >>
rect -184 13183 184 13217
rect -184 4455 184 4489
rect -184 4347 184 4381
rect -184 -4381 184 -4347
rect -184 -4489 184 -4455
rect -184 -13217 184 -13183
<< locali >>
rect -360 13285 360 13319
rect -360 -13285 -326 13285
rect -200 13183 -184 13217
rect 184 13183 200 13217
rect -246 13124 -212 13140
rect -246 4532 -212 4548
rect 212 13124 246 13140
rect 212 4532 246 4548
rect -200 4455 -184 4489
rect 184 4455 200 4489
rect -200 4347 -184 4381
rect 184 4347 200 4381
rect -246 4288 -212 4304
rect -246 -4304 -212 -4288
rect 212 4288 246 4304
rect 212 -4304 246 -4288
rect -200 -4381 -184 -4347
rect 184 -4381 200 -4347
rect -200 -4489 -184 -4455
rect 184 -4489 200 -4455
rect -246 -4548 -212 -4532
rect -246 -13140 -212 -13124
rect 212 -4548 246 -4532
rect 212 -13140 246 -13124
rect -200 -13217 -184 -13183
rect 184 -13217 200 -13183
rect 326 -13285 360 13285
rect -360 -13319 360 -13285
<< viali >>
rect -184 13183 184 13217
rect -246 4548 -212 13124
rect 212 4548 246 13124
rect -184 4455 184 4489
rect -184 4347 184 4381
rect -246 -4288 -212 4288
rect 212 -4288 246 4288
rect -184 -4381 184 -4347
rect -184 -4489 184 -4455
rect -246 -13124 -212 -4548
rect 212 -13124 246 -4548
rect -184 -13217 184 -13183
<< metal1 >>
rect -196 13217 196 13223
rect -196 13183 -184 13217
rect 184 13183 196 13217
rect -196 13177 196 13183
rect -252 13124 -206 13136
rect -252 4548 -246 13124
rect -212 4548 -206 13124
rect -252 4536 -206 4548
rect 206 13124 252 13136
rect 206 4548 212 13124
rect 246 4548 252 13124
rect 206 4536 252 4548
rect -196 4489 196 4495
rect -196 4455 -184 4489
rect 184 4455 196 4489
rect -196 4449 196 4455
rect -196 4381 196 4387
rect -196 4347 -184 4381
rect 184 4347 196 4381
rect -196 4341 196 4347
rect -252 4288 -206 4300
rect -252 -4288 -246 4288
rect -212 -4288 -206 4288
rect -252 -4300 -206 -4288
rect 206 4288 252 4300
rect 206 -4288 212 4288
rect 246 -4288 252 4288
rect 206 -4300 252 -4288
rect -196 -4347 196 -4341
rect -196 -4381 -184 -4347
rect 184 -4381 196 -4347
rect -196 -4387 196 -4381
rect -196 -4455 196 -4449
rect -196 -4489 -184 -4455
rect 184 -4489 196 -4455
rect -196 -4495 196 -4489
rect -252 -4548 -206 -4536
rect -252 -13124 -246 -4548
rect -212 -13124 -206 -4548
rect -252 -13136 -206 -13124
rect 206 -4548 252 -4536
rect 206 -13124 212 -4548
rect 246 -13124 252 -4548
rect 206 -13136 252 -13124
rect -196 -13183 196 -13177
rect -196 -13217 -184 -13183
rect 184 -13217 196 -13183
rect -196 -13223 196 -13217
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -343 -13302 343 13302
string parameters w 43 l 2 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
