magic
tech sky130A
magscale 1 2
timestamp 1620417585
<< xpolycontact >>
rect -2579 50 -2509 482
rect -2579 -482 -2509 -50
rect -2261 50 -2191 482
rect -2261 -482 -2191 -50
rect -1943 50 -1873 482
rect -1943 -482 -1873 -50
rect -1625 50 -1555 482
rect -1625 -482 -1555 -50
rect -1307 50 -1237 482
rect -1307 -482 -1237 -50
rect -989 50 -919 482
rect -989 -482 -919 -50
rect -671 50 -601 482
rect -671 -482 -601 -50
rect -353 50 -283 482
rect -353 -482 -283 -50
rect -35 50 35 482
rect -35 -482 35 -50
rect 283 50 353 482
rect 283 -482 353 -50
rect 601 50 671 482
rect 601 -482 671 -50
rect 919 50 989 482
rect 919 -482 989 -50
rect 1237 50 1307 482
rect 1237 -482 1307 -50
rect 1555 50 1625 482
rect 1555 -482 1625 -50
rect 1873 50 1943 482
rect 1873 -482 1943 -50
rect 2191 50 2261 482
rect 2191 -482 2261 -50
rect 2509 50 2579 482
rect 2509 -482 2579 -50
<< xpolyres >>
rect -2579 -50 -2509 50
rect -2261 -50 -2191 50
rect -1943 -50 -1873 50
rect -1625 -50 -1555 50
rect -1307 -50 -1237 50
rect -989 -50 -919 50
rect -671 -50 -601 50
rect -353 -50 -283 50
rect -35 -50 35 50
rect 283 -50 353 50
rect 601 -50 671 50
rect 919 -50 989 50
rect 1237 -50 1307 50
rect 1555 -50 1625 50
rect 1873 -50 1943 50
rect 2191 -50 2261 50
rect 2509 -50 2579 50
<< viali >>
rect -2563 67 -2525 464
rect -2245 67 -2207 464
rect -1927 67 -1889 464
rect -1609 67 -1571 464
rect -1291 67 -1253 464
rect -973 67 -935 464
rect -655 67 -617 464
rect -337 67 -299 464
rect -19 67 19 464
rect 299 67 337 464
rect 617 67 655 464
rect 935 67 973 464
rect 1253 67 1291 464
rect 1571 67 1609 464
rect 1889 67 1927 464
rect 2207 67 2245 464
rect 2525 67 2563 464
rect -2563 -464 -2525 -67
rect -2245 -464 -2207 -67
rect -1927 -464 -1889 -67
rect -1609 -464 -1571 -67
rect -1291 -464 -1253 -67
rect -973 -464 -935 -67
rect -655 -464 -617 -67
rect -337 -464 -299 -67
rect -19 -464 19 -67
rect 299 -464 337 -67
rect 617 -464 655 -67
rect 935 -464 973 -67
rect 1253 -464 1291 -67
rect 1571 -464 1609 -67
rect 1889 -464 1927 -67
rect 2207 -464 2245 -67
rect 2525 -464 2563 -67
<< metal1 >>
rect -2569 464 -2519 476
rect -2569 67 -2563 464
rect -2525 67 -2519 464
rect -2569 55 -2519 67
rect -2251 464 -2201 476
rect -2251 67 -2245 464
rect -2207 67 -2201 464
rect -2251 55 -2201 67
rect -1933 464 -1883 476
rect -1933 67 -1927 464
rect -1889 67 -1883 464
rect -1933 55 -1883 67
rect -1615 464 -1565 476
rect -1615 67 -1609 464
rect -1571 67 -1565 464
rect -1615 55 -1565 67
rect -1297 464 -1247 476
rect -1297 67 -1291 464
rect -1253 67 -1247 464
rect -1297 55 -1247 67
rect -979 464 -929 476
rect -979 67 -973 464
rect -935 67 -929 464
rect -979 55 -929 67
rect -661 464 -611 476
rect -661 67 -655 464
rect -617 67 -611 464
rect -661 55 -611 67
rect -343 464 -293 476
rect -343 67 -337 464
rect -299 67 -293 464
rect -343 55 -293 67
rect -25 464 25 476
rect -25 67 -19 464
rect 19 67 25 464
rect -25 55 25 67
rect 293 464 343 476
rect 293 67 299 464
rect 337 67 343 464
rect 293 55 343 67
rect 611 464 661 476
rect 611 67 617 464
rect 655 67 661 464
rect 611 55 661 67
rect 929 464 979 476
rect 929 67 935 464
rect 973 67 979 464
rect 929 55 979 67
rect 1247 464 1297 476
rect 1247 67 1253 464
rect 1291 67 1297 464
rect 1247 55 1297 67
rect 1565 464 1615 476
rect 1565 67 1571 464
rect 1609 67 1615 464
rect 1565 55 1615 67
rect 1883 464 1933 476
rect 1883 67 1889 464
rect 1927 67 1933 464
rect 1883 55 1933 67
rect 2201 464 2251 476
rect 2201 67 2207 464
rect 2245 67 2251 464
rect 2201 55 2251 67
rect 2519 464 2569 476
rect 2519 67 2525 464
rect 2563 67 2569 464
rect 2519 55 2569 67
rect -2569 -67 -2519 -55
rect -2569 -464 -2563 -67
rect -2525 -464 -2519 -67
rect -2569 -476 -2519 -464
rect -2251 -67 -2201 -55
rect -2251 -464 -2245 -67
rect -2207 -464 -2201 -67
rect -2251 -476 -2201 -464
rect -1933 -67 -1883 -55
rect -1933 -464 -1927 -67
rect -1889 -464 -1883 -67
rect -1933 -476 -1883 -464
rect -1615 -67 -1565 -55
rect -1615 -464 -1609 -67
rect -1571 -464 -1565 -67
rect -1615 -476 -1565 -464
rect -1297 -67 -1247 -55
rect -1297 -464 -1291 -67
rect -1253 -464 -1247 -67
rect -1297 -476 -1247 -464
rect -979 -67 -929 -55
rect -979 -464 -973 -67
rect -935 -464 -929 -67
rect -979 -476 -929 -464
rect -661 -67 -611 -55
rect -661 -464 -655 -67
rect -617 -464 -611 -67
rect -661 -476 -611 -464
rect -343 -67 -293 -55
rect -343 -464 -337 -67
rect -299 -464 -293 -67
rect -343 -476 -293 -464
rect -25 -67 25 -55
rect -25 -464 -19 -67
rect 19 -464 25 -67
rect -25 -476 25 -464
rect 293 -67 343 -55
rect 293 -464 299 -67
rect 337 -464 343 -67
rect 293 -476 343 -464
rect 611 -67 661 -55
rect 611 -464 617 -67
rect 655 -464 661 -67
rect 611 -476 661 -464
rect 929 -67 979 -55
rect 929 -464 935 -67
rect 973 -464 979 -67
rect 929 -476 979 -464
rect 1247 -67 1297 -55
rect 1247 -464 1253 -67
rect 1291 -464 1297 -67
rect 1247 -476 1297 -464
rect 1565 -67 1615 -55
rect 1565 -464 1571 -67
rect 1609 -464 1615 -67
rect 1565 -476 1615 -464
rect 1883 -67 1933 -55
rect 1883 -464 1889 -67
rect 1927 -464 1933 -67
rect 1883 -476 1933 -464
rect 2201 -67 2251 -55
rect 2201 -464 2207 -67
rect 2245 -464 2251 -67
rect 2201 -476 2251 -464
rect 2519 -67 2569 -55
rect 2519 -464 2525 -67
rect 2563 -464 2569 -67
rect 2519 -476 2569 -464
<< res0p35 >>
rect -2581 -52 -2507 52
rect -2263 -52 -2189 52
rect -1945 -52 -1871 52
rect -1627 -52 -1553 52
rect -1309 -52 -1235 52
rect -991 -52 -917 52
rect -673 -52 -599 52
rect -355 -52 -281 52
rect -37 -52 37 52
rect 281 -52 355 52
rect 599 -52 673 52
rect 917 -52 991 52
rect 1235 -52 1309 52
rect 1553 -52 1627 52
rect 1871 -52 1945 52
rect 2189 -52 2263 52
rect 2507 -52 2581 52
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 0.50 m 1 nx 17 wmin 0.350 lmin 0.50 rho 2000 val 3.542k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
