magic
tech sky130A
magscale 1 2
timestamp 1620244706
<< error_p >>
rect -801 4464 -729 4498
rect 729 4464 801 4498
rect -801 4426 -767 4464
rect 767 4426 801 4464
rect -671 2704 -601 2848
rect -353 2704 -283 2848
rect -35 2704 35 2848
rect 283 2704 353 2848
rect 601 2704 671 2848
rect -671 936 -601 1080
rect -353 936 -283 1080
rect -35 936 35 1080
rect 283 936 353 1080
rect 601 936 671 1080
rect -671 -832 -601 -688
rect -353 -832 -283 -688
rect -35 -832 35 -688
rect 283 -832 353 -688
rect 601 -832 671 -688
rect -671 -2600 -601 -2456
rect -353 -2600 -283 -2456
rect -35 -2600 35 -2456
rect 283 -2600 353 -2456
rect 601 -2600 671 -2456
rect -801 -4430 -767 -4426
rect 767 -4430 801 -4426
rect -801 -4464 -733 -4430
rect 733 -4464 801 -4430
rect -767 -4498 -729 -4464
rect 729 -4498 767 -4464
<< pwell >>
rect -837 -4534 837 4534
<< psubdiff >>
rect -801 4464 -705 4498
rect 705 4464 801 4498
rect -801 4402 -767 4464
rect 767 4402 801 4464
rect -801 -4464 -767 -4402
rect 767 -4464 801 -4402
rect -801 -4498 -705 -4464
rect 705 -4498 801 -4464
<< psubdiffcont >>
rect -705 4464 705 4498
rect -801 -4402 -767 4402
rect 767 -4402 801 4402
rect -705 -4498 705 -4464
<< xpolycontact >>
rect -671 3936 -601 4368
rect -671 2704 -601 3136
rect -353 3936 -283 4368
rect -353 2704 -283 3136
rect -35 3936 35 4368
rect -35 2704 35 3136
rect 283 3936 353 4368
rect 283 2704 353 3136
rect 601 3936 671 4368
rect 601 2704 671 3136
rect -671 2168 -601 2600
rect -671 936 -601 1368
rect -353 2168 -283 2600
rect -353 936 -283 1368
rect -35 2168 35 2600
rect -35 936 35 1368
rect 283 2168 353 2600
rect 283 936 353 1368
rect 601 2168 671 2600
rect 601 936 671 1368
rect -671 400 -601 832
rect -671 -832 -601 -400
rect -353 400 -283 832
rect -353 -832 -283 -400
rect -35 400 35 832
rect -35 -832 35 -400
rect 283 400 353 832
rect 283 -832 353 -400
rect 601 400 671 832
rect 601 -832 671 -400
rect -671 -1368 -601 -936
rect -671 -2600 -601 -2168
rect -353 -1368 -283 -936
rect -353 -2600 -283 -2168
rect -35 -1368 35 -936
rect -35 -2600 35 -2168
rect 283 -1368 353 -936
rect 283 -2600 353 -2168
rect 601 -1368 671 -936
rect 601 -2600 671 -2168
rect -671 -3136 -601 -2704
rect -671 -4368 -601 -3936
rect -353 -3136 -283 -2704
rect -353 -4368 -283 -3936
rect -35 -3136 35 -2704
rect -35 -4368 35 -3936
rect 283 -3136 353 -2704
rect 283 -4368 353 -3936
rect 601 -3136 671 -2704
rect 601 -4368 671 -3936
<< xpolyres >>
rect -671 3136 -601 3936
rect -353 3136 -283 3936
rect -35 3136 35 3936
rect 283 3136 353 3936
rect 601 3136 671 3936
rect -671 1368 -601 2168
rect -353 1368 -283 2168
rect -35 1368 35 2168
rect 283 1368 353 2168
rect 601 1368 671 2168
rect -671 -400 -601 400
rect -353 -400 -283 400
rect -35 -400 35 400
rect 283 -400 353 400
rect 601 -400 671 400
rect -671 -2168 -601 -1368
rect -353 -2168 -283 -1368
rect -35 -2168 35 -1368
rect 283 -2168 353 -1368
rect 601 -2168 671 -1368
rect -671 -3936 -601 -3136
rect -353 -3936 -283 -3136
rect -35 -3936 35 -3136
rect 283 -3936 353 -3136
rect 601 -3936 671 -3136
<< locali >>
rect -801 4464 -767 4498
rect 767 4464 801 4498
rect -801 -4498 -767 -4464
rect 767 -4498 801 -4464
<< viali >>
rect -767 4464 -705 4498
rect -705 4464 705 4498
rect 705 4464 767 4498
rect -801 4402 -767 4464
rect -801 -4402 -767 4402
rect 767 4402 801 4464
rect -655 3953 -617 4350
rect -337 3953 -299 4350
rect -19 3953 19 4350
rect 299 3953 337 4350
rect 617 3953 655 4350
rect -655 2722 -617 3119
rect -337 2722 -299 3119
rect -19 2722 19 3119
rect 299 2722 337 3119
rect 617 2722 655 3119
rect -655 2185 -617 2582
rect -337 2185 -299 2582
rect -19 2185 19 2582
rect 299 2185 337 2582
rect 617 2185 655 2582
rect -655 954 -617 1351
rect -337 954 -299 1351
rect -19 954 19 1351
rect 299 954 337 1351
rect 617 954 655 1351
rect -655 417 -617 814
rect -337 417 -299 814
rect -19 417 19 814
rect 299 417 337 814
rect 617 417 655 814
rect -655 -814 -617 -417
rect -337 -814 -299 -417
rect -19 -814 19 -417
rect 299 -814 337 -417
rect 617 -814 655 -417
rect -655 -1351 -617 -954
rect -337 -1351 -299 -954
rect -19 -1351 19 -954
rect 299 -1351 337 -954
rect 617 -1351 655 -954
rect -655 -2582 -617 -2185
rect -337 -2582 -299 -2185
rect -19 -2582 19 -2185
rect 299 -2582 337 -2185
rect 617 -2582 655 -2185
rect -655 -3119 -617 -2722
rect -337 -3119 -299 -2722
rect -19 -3119 19 -2722
rect 299 -3119 337 -2722
rect 617 -3119 655 -2722
rect -655 -4350 -617 -3953
rect -337 -4350 -299 -3953
rect -19 -4350 19 -3953
rect 299 -4350 337 -3953
rect 617 -4350 655 -3953
rect -801 -4464 -767 -4402
rect 767 -4402 801 4402
rect 767 -4464 801 -4402
rect -767 -4498 -705 -4464
rect -705 -4498 705 -4464
rect 705 -4498 767 -4464
<< metal1 >>
rect -779 4498 779 4504
rect -779 4476 -767 4498
rect -807 4464 -767 4476
rect 767 4476 779 4498
rect 767 4464 807 4476
rect -807 -4464 -801 4464
rect -767 4458 767 4464
rect -767 -4458 -761 4458
rect -661 4350 -611 4362
rect -661 3953 -655 4350
rect -617 3953 -611 4350
rect -661 3941 -611 3953
rect -343 4350 -293 4362
rect -343 3953 -337 4350
rect -299 3953 -293 4350
rect -343 3941 -293 3953
rect -25 4350 25 4362
rect -25 3953 -19 4350
rect 19 3953 25 4350
rect -25 3941 25 3953
rect 293 4350 343 4362
rect 293 3953 299 4350
rect 337 3953 343 4350
rect 293 3941 343 3953
rect 611 4350 661 4362
rect 611 3953 617 4350
rect 655 3953 661 4350
rect 611 3941 661 3953
rect -661 3119 -611 3131
rect -661 2722 -655 3119
rect -617 2722 -611 3119
rect -661 2710 -611 2722
rect -343 3119 -293 3131
rect -343 2722 -337 3119
rect -299 2722 -293 3119
rect -343 2710 -293 2722
rect -25 3119 25 3131
rect -25 2722 -19 3119
rect 19 2722 25 3119
rect -25 2710 25 2722
rect 293 3119 343 3131
rect 293 2722 299 3119
rect 337 2722 343 3119
rect 293 2710 343 2722
rect 611 3119 661 3131
rect 611 2722 617 3119
rect 655 2722 661 3119
rect 611 2710 661 2722
rect -661 2582 -611 2594
rect -661 2185 -655 2582
rect -617 2185 -611 2582
rect -661 2173 -611 2185
rect -343 2582 -293 2594
rect -343 2185 -337 2582
rect -299 2185 -293 2582
rect -343 2173 -293 2185
rect -25 2582 25 2594
rect -25 2185 -19 2582
rect 19 2185 25 2582
rect -25 2173 25 2185
rect 293 2582 343 2594
rect 293 2185 299 2582
rect 337 2185 343 2582
rect 293 2173 343 2185
rect 611 2582 661 2594
rect 611 2185 617 2582
rect 655 2185 661 2582
rect 611 2173 661 2185
rect -661 1351 -611 1363
rect -661 954 -655 1351
rect -617 954 -611 1351
rect -661 942 -611 954
rect -343 1351 -293 1363
rect -343 954 -337 1351
rect -299 954 -293 1351
rect -343 942 -293 954
rect -25 1351 25 1363
rect -25 954 -19 1351
rect 19 954 25 1351
rect -25 942 25 954
rect 293 1351 343 1363
rect 293 954 299 1351
rect 337 954 343 1351
rect 293 942 343 954
rect 611 1351 661 1363
rect 611 954 617 1351
rect 655 954 661 1351
rect 611 942 661 954
rect -661 814 -611 826
rect -661 417 -655 814
rect -617 417 -611 814
rect -661 405 -611 417
rect -343 814 -293 826
rect -343 417 -337 814
rect -299 417 -293 814
rect -343 405 -293 417
rect -25 814 25 826
rect -25 417 -19 814
rect 19 417 25 814
rect -25 405 25 417
rect 293 814 343 826
rect 293 417 299 814
rect 337 417 343 814
rect 293 405 343 417
rect 611 814 661 826
rect 611 417 617 814
rect 655 417 661 814
rect 611 405 661 417
rect -661 -417 -611 -405
rect -661 -814 -655 -417
rect -617 -814 -611 -417
rect -661 -826 -611 -814
rect -343 -417 -293 -405
rect -343 -814 -337 -417
rect -299 -814 -293 -417
rect -343 -826 -293 -814
rect -25 -417 25 -405
rect -25 -814 -19 -417
rect 19 -814 25 -417
rect -25 -826 25 -814
rect 293 -417 343 -405
rect 293 -814 299 -417
rect 337 -814 343 -417
rect 293 -826 343 -814
rect 611 -417 661 -405
rect 611 -814 617 -417
rect 655 -814 661 -417
rect 611 -826 661 -814
rect -661 -954 -611 -942
rect -661 -1351 -655 -954
rect -617 -1351 -611 -954
rect -661 -1363 -611 -1351
rect -343 -954 -293 -942
rect -343 -1351 -337 -954
rect -299 -1351 -293 -954
rect -343 -1363 -293 -1351
rect -25 -954 25 -942
rect -25 -1351 -19 -954
rect 19 -1351 25 -954
rect -25 -1363 25 -1351
rect 293 -954 343 -942
rect 293 -1351 299 -954
rect 337 -1351 343 -954
rect 293 -1363 343 -1351
rect 611 -954 661 -942
rect 611 -1351 617 -954
rect 655 -1351 661 -954
rect 611 -1363 661 -1351
rect -661 -2185 -611 -2173
rect -661 -2582 -655 -2185
rect -617 -2582 -611 -2185
rect -661 -2594 -611 -2582
rect -343 -2185 -293 -2173
rect -343 -2582 -337 -2185
rect -299 -2582 -293 -2185
rect -343 -2594 -293 -2582
rect -25 -2185 25 -2173
rect -25 -2582 -19 -2185
rect 19 -2582 25 -2185
rect -25 -2594 25 -2582
rect 293 -2185 343 -2173
rect 293 -2582 299 -2185
rect 337 -2582 343 -2185
rect 293 -2594 343 -2582
rect 611 -2185 661 -2173
rect 611 -2582 617 -2185
rect 655 -2582 661 -2185
rect 611 -2594 661 -2582
rect -661 -2722 -611 -2710
rect -661 -3119 -655 -2722
rect -617 -3119 -611 -2722
rect -661 -3131 -611 -3119
rect -343 -2722 -293 -2710
rect -343 -3119 -337 -2722
rect -299 -3119 -293 -2722
rect -343 -3131 -293 -3119
rect -25 -2722 25 -2710
rect -25 -3119 -19 -2722
rect 19 -3119 25 -2722
rect -25 -3131 25 -3119
rect 293 -2722 343 -2710
rect 293 -3119 299 -2722
rect 337 -3119 343 -2722
rect 293 -3131 343 -3119
rect 611 -2722 661 -2710
rect 611 -3119 617 -2722
rect 655 -3119 661 -2722
rect 611 -3131 661 -3119
rect -661 -3953 -611 -3941
rect -661 -4350 -655 -3953
rect -617 -4350 -611 -3953
rect -661 -4362 -611 -4350
rect -343 -3953 -293 -3941
rect -343 -4350 -337 -3953
rect -299 -4350 -293 -3953
rect -343 -4362 -293 -4350
rect -25 -3953 25 -3941
rect -25 -4350 -19 -3953
rect 19 -4350 25 -3953
rect -25 -4362 25 -4350
rect 293 -3953 343 -3941
rect 293 -4350 299 -3953
rect 337 -4350 343 -3953
rect 293 -4362 343 -4350
rect 611 -3953 661 -3941
rect 611 -4350 617 -3953
rect 655 -4350 661 -3953
rect 611 -4362 661 -4350
rect 761 -4458 767 4458
rect -767 -4464 767 -4458
rect 801 -4464 807 4464
rect -807 -4476 -767 -4464
rect -779 -4498 -767 -4476
rect 767 -4476 807 -4464
rect 767 -4498 779 -4476
rect -779 -4504 779 -4498
<< res0p35 >>
rect -673 3134 -599 3938
rect -355 3134 -281 3938
rect -37 3134 37 3938
rect 281 3134 355 3938
rect 599 3134 673 3938
rect -673 1366 -599 2170
rect -355 1366 -281 2170
rect -37 1366 37 2170
rect 281 1366 355 2170
rect 599 1366 673 2170
rect -673 -402 -599 402
rect -355 -402 -281 402
rect -37 -402 37 402
rect 281 -402 355 402
rect 599 -402 673 402
rect -673 -2170 -599 -1366
rect -355 -2170 -281 -1366
rect -37 -2170 37 -1366
rect 281 -2170 355 -1366
rect 599 -2170 673 -1366
rect -673 -3938 -599 -3134
rect -355 -3938 -281 -3134
rect -37 -3938 37 -3134
rect 281 -3938 355 -3134
rect 599 -3938 673 -3134
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string FIXED_BBOX -784 -4481 784 4481
string parameters w 0.350 l 4 m 5 nx 5 wmin 0.350 lmin 0.50 rho 2000 val 23.542k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 vias 1 viagb 100 viagt 100 viagl 100 viagr 100
string library sky130
<< end >>
