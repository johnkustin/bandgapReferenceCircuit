magic
tech sky130A
magscale 1 2
timestamp 1620244706
<< error_p >>
rect -512 52 -442 196
rect -194 52 -124 196
rect 124 52 194 196
rect 442 52 512 196
<< xpolycontact >>
rect -512 1236 -442 1668
rect -512 52 -442 484
rect -194 1236 -124 1668
rect -194 52 -124 484
rect 124 1236 194 1668
rect 124 52 194 484
rect 442 1236 512 1668
rect 442 52 512 484
rect -512 -484 -442 -52
rect -512 -1668 -442 -1236
rect -194 -484 -124 -52
rect -194 -1668 -124 -1236
rect 124 -484 194 -52
rect 124 -1668 194 -1236
rect 442 -484 512 -52
rect 442 -1668 512 -1236
<< xpolyres >>
rect -512 484 -442 1236
rect -194 484 -124 1236
rect 124 484 194 1236
rect 442 484 512 1236
rect -512 -1236 -442 -484
rect -194 -1236 -124 -484
rect 124 -1236 194 -484
rect 442 -1236 512 -484
<< viali >>
rect -496 1253 -458 1650
rect -178 1253 -140 1650
rect 140 1253 178 1650
rect 458 1253 496 1650
rect -496 70 -458 467
rect -178 70 -140 467
rect 140 70 178 467
rect 458 70 496 467
rect -496 -467 -458 -70
rect -178 -467 -140 -70
rect 140 -467 178 -70
rect 458 -467 496 -70
rect -496 -1650 -458 -1253
rect -178 -1650 -140 -1253
rect 140 -1650 178 -1253
rect 458 -1650 496 -1253
<< metal1 >>
rect -502 1650 -452 1662
rect -502 1253 -496 1650
rect -458 1253 -452 1650
rect -502 1241 -452 1253
rect -184 1650 -134 1662
rect -184 1253 -178 1650
rect -140 1253 -134 1650
rect -184 1241 -134 1253
rect 134 1650 184 1662
rect 134 1253 140 1650
rect 178 1253 184 1650
rect 134 1241 184 1253
rect 452 1650 502 1662
rect 452 1253 458 1650
rect 496 1253 502 1650
rect 452 1241 502 1253
rect -502 467 -452 479
rect -502 70 -496 467
rect -458 70 -452 467
rect -502 58 -452 70
rect -184 467 -134 479
rect -184 70 -178 467
rect -140 70 -134 467
rect -184 58 -134 70
rect 134 467 184 479
rect 134 70 140 467
rect 178 70 184 467
rect 134 58 184 70
rect 452 467 502 479
rect 452 70 458 467
rect 496 70 502 467
rect 452 58 502 70
rect -502 -70 -452 -58
rect -502 -467 -496 -70
rect -458 -467 -452 -70
rect -502 -479 -452 -467
rect -184 -70 -134 -58
rect -184 -467 -178 -70
rect -140 -467 -134 -70
rect -184 -479 -134 -467
rect 134 -70 184 -58
rect 134 -467 140 -70
rect 178 -467 184 -70
rect 134 -479 184 -467
rect 452 -70 502 -58
rect 452 -467 458 -70
rect 496 -467 502 -70
rect 452 -479 502 -467
rect -502 -1253 -452 -1241
rect -502 -1650 -496 -1253
rect -458 -1650 -452 -1253
rect -502 -1662 -452 -1650
rect -184 -1253 -134 -1241
rect -184 -1650 -178 -1253
rect -140 -1650 -134 -1253
rect -184 -1662 -134 -1650
rect 134 -1253 184 -1241
rect 134 -1650 140 -1253
rect 178 -1650 184 -1253
rect 134 -1662 184 -1650
rect 452 -1253 502 -1241
rect 452 -1650 458 -1253
rect 496 -1650 502 -1253
rect 452 -1662 502 -1650
<< res0p35 >>
rect -514 482 -440 1238
rect -196 482 -122 1238
rect 122 482 196 1238
rect 440 482 514 1238
rect -514 -1238 -440 -482
rect -196 -1238 -122 -482
rect 122 -1238 196 -482
rect 440 -1238 514 -482
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string parameters w 0.350 l 3.763 m 2 nx 4 wmin 0.350 lmin 0.50 rho 2000 val 22.188k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
