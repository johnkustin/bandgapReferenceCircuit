magic
tech sky130A
magscale 1 2
timestamp 1620886664
<< xpolycontact >>
rect -69 487 69 919
rect -69 -919 69 -487
<< xpolyres >>
rect -69 -487 69 487
<< viali >>
rect -53 504 53 901
rect -53 -901 53 -504
<< metal1 >>
rect -59 901 59 913
rect -59 504 -53 901
rect 53 504 59 901
rect -59 492 59 504
rect -59 -504 59 -492
rect -59 -901 -53 -504
rect 53 -901 59 -504
rect -59 -913 59 -901
<< res0p69 >>
rect -71 -489 71 489
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p69
string parameters w 0.690 l 4.87 m 1 nx 1 wmin 0.690 lmin 0.50 rho 2000 val 14.171k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 wmax 0.690 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
