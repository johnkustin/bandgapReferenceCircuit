magic
tech sky130A
magscale 1 2
timestamp 1620244706
<< error_p >>
rect -35 11232 35 11376
rect -35 9512 35 9656
rect -35 7792 35 7936
rect -35 6072 35 6216
rect -35 4352 35 4496
rect -35 2632 35 2776
rect -35 912 35 1056
rect -35 -808 35 -664
rect -35 -2528 35 -2384
rect -35 -4248 35 -4104
rect -35 -5968 35 -5824
rect -35 -7688 35 -7544
rect -35 -9408 35 -9264
rect -35 -11128 35 -10984
<< pwell >>
rect -201 -13014 201 13014
<< psubdiff >>
rect -165 12944 -69 12978
rect 69 12944 165 12978
rect -165 12882 -131 12944
rect 131 12882 165 12944
rect -165 -12944 -131 -12882
rect 131 -12944 165 -12882
rect -165 -12978 -69 -12944
rect 69 -12978 165 -12944
<< psubdiffcont >>
rect -69 12944 69 12978
rect -165 -12882 -131 12882
rect 131 -12882 165 12882
rect -69 -12978 69 -12944
<< xpolycontact >>
rect -35 12416 35 12848
rect -35 11232 35 11664
rect -35 10696 35 11128
rect -35 9512 35 9944
rect -35 8976 35 9408
rect -35 7792 35 8224
rect -35 7256 35 7688
rect -35 6072 35 6504
rect -35 5536 35 5968
rect -35 4352 35 4784
rect -35 3816 35 4248
rect -35 2632 35 3064
rect -35 2096 35 2528
rect -35 912 35 1344
rect -35 376 35 808
rect -35 -808 35 -376
rect -35 -1344 35 -912
rect -35 -2528 35 -2096
rect -35 -3064 35 -2632
rect -35 -4248 35 -3816
rect -35 -4784 35 -4352
rect -35 -5968 35 -5536
rect -35 -6504 35 -6072
rect -35 -7688 35 -7256
rect -35 -8224 35 -7792
rect -35 -9408 35 -8976
rect -35 -9944 35 -9512
rect -35 -11128 35 -10696
rect -35 -11664 35 -11232
rect -35 -12848 35 -12416
<< xpolyres >>
rect -35 11664 35 12416
rect -35 9944 35 10696
rect -35 8224 35 8976
rect -35 6504 35 7256
rect -35 4784 35 5536
rect -35 3064 35 3816
rect -35 1344 35 2096
rect -35 -376 35 376
rect -35 -2096 35 -1344
rect -35 -3816 35 -3064
rect -35 -5536 35 -4784
rect -35 -7256 35 -6504
rect -35 -8976 35 -8224
rect -35 -10696 35 -9944
rect -35 -12416 35 -11664
<< locali >>
rect -165 12944 -69 12978
rect 69 12944 165 12978
rect -165 12882 -131 12944
rect 131 12882 165 12944
rect -165 -12944 -131 -12882
rect 131 -12944 165 -12882
rect -165 -12978 -69 -12944
rect 69 -12978 165 -12944
<< viali >>
rect -19 12433 19 12830
rect -19 11250 19 11647
rect -19 10713 19 11110
rect -19 9530 19 9927
rect -19 8993 19 9390
rect -19 7810 19 8207
rect -19 7273 19 7670
rect -19 6090 19 6487
rect -19 5553 19 5950
rect -19 4370 19 4767
rect -19 3833 19 4230
rect -19 2650 19 3047
rect -19 2113 19 2510
rect -19 930 19 1327
rect -19 393 19 790
rect -19 -790 19 -393
rect -19 -1327 19 -930
rect -19 -2510 19 -2113
rect -19 -3047 19 -2650
rect -19 -4230 19 -3833
rect -19 -4767 19 -4370
rect -19 -5950 19 -5553
rect -19 -6487 19 -6090
rect -19 -7670 19 -7273
rect -19 -8207 19 -7810
rect -19 -9390 19 -8993
rect -19 -9927 19 -9530
rect -19 -11110 19 -10713
rect -19 -11647 19 -11250
rect -19 -12830 19 -12433
<< metal1 >>
rect -25 12830 25 12842
rect -25 12433 -19 12830
rect 19 12433 25 12830
rect -25 12421 25 12433
rect -25 11647 25 11659
rect -25 11250 -19 11647
rect 19 11250 25 11647
rect -25 11238 25 11250
rect -25 11110 25 11122
rect -25 10713 -19 11110
rect 19 10713 25 11110
rect -25 10701 25 10713
rect -25 9927 25 9939
rect -25 9530 -19 9927
rect 19 9530 25 9927
rect -25 9518 25 9530
rect -25 9390 25 9402
rect -25 8993 -19 9390
rect 19 8993 25 9390
rect -25 8981 25 8993
rect -25 8207 25 8219
rect -25 7810 -19 8207
rect 19 7810 25 8207
rect -25 7798 25 7810
rect -25 7670 25 7682
rect -25 7273 -19 7670
rect 19 7273 25 7670
rect -25 7261 25 7273
rect -25 6487 25 6499
rect -25 6090 -19 6487
rect 19 6090 25 6487
rect -25 6078 25 6090
rect -25 5950 25 5962
rect -25 5553 -19 5950
rect 19 5553 25 5950
rect -25 5541 25 5553
rect -25 4767 25 4779
rect -25 4370 -19 4767
rect 19 4370 25 4767
rect -25 4358 25 4370
rect -25 4230 25 4242
rect -25 3833 -19 4230
rect 19 3833 25 4230
rect -25 3821 25 3833
rect -25 3047 25 3059
rect -25 2650 -19 3047
rect 19 2650 25 3047
rect -25 2638 25 2650
rect -25 2510 25 2522
rect -25 2113 -19 2510
rect 19 2113 25 2510
rect -25 2101 25 2113
rect -25 1327 25 1339
rect -25 930 -19 1327
rect 19 930 25 1327
rect -25 918 25 930
rect -25 790 25 802
rect -25 393 -19 790
rect 19 393 25 790
rect -25 381 25 393
rect -25 -393 25 -381
rect -25 -790 -19 -393
rect 19 -790 25 -393
rect -25 -802 25 -790
rect -25 -930 25 -918
rect -25 -1327 -19 -930
rect 19 -1327 25 -930
rect -25 -1339 25 -1327
rect -25 -2113 25 -2101
rect -25 -2510 -19 -2113
rect 19 -2510 25 -2113
rect -25 -2522 25 -2510
rect -25 -2650 25 -2638
rect -25 -3047 -19 -2650
rect 19 -3047 25 -2650
rect -25 -3059 25 -3047
rect -25 -3833 25 -3821
rect -25 -4230 -19 -3833
rect 19 -4230 25 -3833
rect -25 -4242 25 -4230
rect -25 -4370 25 -4358
rect -25 -4767 -19 -4370
rect 19 -4767 25 -4370
rect -25 -4779 25 -4767
rect -25 -5553 25 -5541
rect -25 -5950 -19 -5553
rect 19 -5950 25 -5553
rect -25 -5962 25 -5950
rect -25 -6090 25 -6078
rect -25 -6487 -19 -6090
rect 19 -6487 25 -6090
rect -25 -6499 25 -6487
rect -25 -7273 25 -7261
rect -25 -7670 -19 -7273
rect 19 -7670 25 -7273
rect -25 -7682 25 -7670
rect -25 -7810 25 -7798
rect -25 -8207 -19 -7810
rect 19 -8207 25 -7810
rect -25 -8219 25 -8207
rect -25 -8993 25 -8981
rect -25 -9390 -19 -8993
rect 19 -9390 25 -8993
rect -25 -9402 25 -9390
rect -25 -9530 25 -9518
rect -25 -9927 -19 -9530
rect 19 -9927 25 -9530
rect -25 -9939 25 -9927
rect -25 -10713 25 -10701
rect -25 -11110 -19 -10713
rect 19 -11110 25 -10713
rect -25 -11122 25 -11110
rect -25 -11250 25 -11238
rect -25 -11647 -19 -11250
rect 19 -11647 25 -11250
rect -25 -11659 25 -11647
rect -25 -12433 25 -12421
rect -25 -12830 -19 -12433
rect 19 -12830 25 -12433
rect -25 -12842 25 -12830
<< res0p35 >>
rect -37 11662 37 12418
rect -37 9942 37 10698
rect -37 8222 37 8978
rect -37 6502 37 7258
rect -37 4782 37 5538
rect -37 3062 37 3818
rect -37 1342 37 2098
rect -37 -378 37 378
rect -37 -2098 37 -1342
rect -37 -3818 37 -3062
rect -37 -5538 37 -4782
rect -37 -7258 37 -6502
rect -37 -8978 37 -8222
rect -37 -10698 37 -9942
rect -37 -12418 37 -11662
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string FIXED_BBOX -148 -12961 148 12961
string parameters w 0.350 l 3.763 m 15 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 22.188k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
